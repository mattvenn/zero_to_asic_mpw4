magic
tech sky130A
magscale 1 2
timestamp 1640364529
<< metal1 >>
rect 331214 702992 331220 703044
rect 331272 703032 331278 703044
rect 332502 703032 332508 703044
rect 331272 703004 332508 703032
rect 331272 702992 331278 703004
rect 332502 702992 332508 703004
rect 332560 702992 332566 703044
rect 170306 702924 170312 702976
rect 170364 702964 170370 702976
rect 281534 702964 281540 702976
rect 170364 702936 281540 702964
rect 170364 702924 170370 702936
rect 281534 702924 281540 702936
rect 281592 702924 281598 702976
rect 62022 702856 62028 702908
rect 62080 702896 62086 702908
rect 267642 702896 267648 702908
rect 62080 702868 267648 702896
rect 62080 702856 62086 702868
rect 267642 702856 267648 702868
rect 267700 702856 267706 702908
rect 276014 702856 276020 702908
rect 276072 702896 276078 702908
rect 478506 702896 478512 702908
rect 276072 702868 478512 702896
rect 276072 702856 276078 702868
rect 478506 702856 478512 702868
rect 478564 702856 478570 702908
rect 202782 702788 202788 702840
rect 202840 702828 202846 702840
rect 273254 702828 273260 702840
rect 202840 702800 273260 702828
rect 202840 702788 202846 702800
rect 273254 702788 273260 702800
rect 273312 702788 273318 702840
rect 349798 702788 349804 702840
rect 349856 702828 349862 702840
rect 494790 702828 494796 702840
rect 349856 702800 494796 702828
rect 349856 702788 349862 702800
rect 494790 702788 494796 702800
rect 494848 702788 494854 702840
rect 233878 702720 233884 702772
rect 233936 702760 233942 702772
rect 397362 702760 397368 702772
rect 233936 702732 397368 702760
rect 233936 702720 233942 702732
rect 397362 702720 397368 702732
rect 397420 702720 397426 702772
rect 197262 702652 197268 702704
rect 197320 702692 197326 702704
rect 364978 702692 364984 702704
rect 197320 702664 364984 702692
rect 197320 702652 197326 702664
rect 364978 702652 364984 702664
rect 365036 702652 365042 702704
rect 382918 702652 382924 702704
rect 382976 702692 382982 702704
rect 462314 702692 462320 702704
rect 382976 702664 462320 702692
rect 382976 702652 382982 702664
rect 462314 702652 462320 702664
rect 462372 702652 462378 702704
rect 95142 702584 95148 702636
rect 95200 702624 95206 702636
rect 300118 702624 300124 702636
rect 95200 702596 300124 702624
rect 95200 702584 95206 702596
rect 300118 702584 300124 702596
rect 300176 702624 300182 702636
rect 300762 702624 300768 702636
rect 300176 702596 300768 702624
rect 300176 702584 300182 702596
rect 300762 702584 300768 702596
rect 300820 702584 300826 702636
rect 363598 702584 363604 702636
rect 363656 702624 363662 702636
rect 543458 702624 543464 702636
rect 363656 702596 543464 702624
rect 363656 702584 363662 702596
rect 543458 702584 543464 702596
rect 543516 702584 543522 702636
rect 86862 702516 86868 702568
rect 86920 702556 86926 702568
rect 235166 702556 235172 702568
rect 86920 702528 235172 702556
rect 86920 702516 86926 702528
rect 235166 702516 235172 702528
rect 235224 702516 235230 702568
rect 264238 702516 264244 702568
rect 264296 702556 264302 702568
rect 559650 702556 559656 702568
rect 264296 702528 559656 702556
rect 264296 702516 264302 702528
rect 559650 702516 559656 702528
rect 559708 702516 559714 702568
rect 8110 702448 8116 702500
rect 8168 702488 8174 702500
rect 88794 702488 88800 702500
rect 8168 702460 88800 702488
rect 8168 702448 8174 702460
rect 88794 702448 88800 702460
rect 88852 702448 88858 702500
rect 99282 702448 99288 702500
rect 99340 702488 99346 702500
rect 527174 702488 527180 702500
rect 99340 702460 527180 702488
rect 99340 702448 99346 702460
rect 527174 702448 527180 702460
rect 527232 702448 527238 702500
rect 129642 700340 129648 700392
rect 129700 700380 129706 700392
rect 137830 700380 137836 700392
rect 129700 700352 137836 700380
rect 129700 700340 129706 700352
rect 137830 700340 137836 700352
rect 137888 700340 137894 700392
rect 68278 700272 68284 700324
rect 68336 700312 68342 700324
rect 105446 700312 105452 700324
rect 68336 700284 105452 700312
rect 68336 700272 68342 700284
rect 105446 700272 105452 700284
rect 105504 700272 105510 700324
rect 130378 700272 130384 700324
rect 130436 700312 130442 700324
rect 218974 700312 218980 700324
rect 130436 700284 218980 700312
rect 130436 700272 130442 700284
rect 218974 700272 218980 700284
rect 219032 700272 219038 700324
rect 283834 700272 283840 700324
rect 283892 700312 283898 700324
rect 295334 700312 295340 700324
rect 283892 700284 295340 700312
rect 283892 700272 283898 700284
rect 295334 700272 295340 700284
rect 295392 700272 295398 700324
rect 300762 700272 300768 700324
rect 300820 700312 300826 700324
rect 360194 700312 360200 700324
rect 300820 700284 360200 700312
rect 300820 700272 300826 700284
rect 360194 700272 360200 700284
rect 360252 700272 360258 700324
rect 374638 700272 374644 700324
rect 374696 700312 374702 700324
rect 429838 700312 429844 700324
rect 374696 700284 429844 700312
rect 374696 700272 374702 700284
rect 429838 700272 429844 700284
rect 429896 700272 429902 700324
rect 24302 699660 24308 699712
rect 24360 699700 24366 699712
rect 25498 699700 25504 699712
rect 24360 699672 25504 699700
rect 24360 699660 24366 699672
rect 25498 699660 25504 699672
rect 25556 699660 25562 699712
rect 65794 699660 65800 699712
rect 65852 699700 65858 699712
rect 72970 699700 72976 699712
rect 65852 699672 72976 699700
rect 65852 699660 65858 699672
rect 72970 699660 72976 699672
rect 73028 699660 73034 699712
rect 87598 699660 87604 699712
rect 87656 699700 87662 699712
rect 89162 699700 89168 699712
rect 87656 699672 89168 699700
rect 87656 699660 87662 699672
rect 89162 699660 89168 699672
rect 89220 699660 89226 699712
rect 327718 698912 327724 698964
rect 327776 698952 327782 698964
rect 348786 698952 348792 698964
rect 327776 698924 348792 698952
rect 327776 698912 327782 698924
rect 348786 698912 348792 698924
rect 348844 698912 348850 698964
rect 3418 683136 3424 683188
rect 3476 683176 3482 683188
rect 11698 683176 11704 683188
rect 3476 683148 11704 683176
rect 3476 683136 3482 683148
rect 11698 683136 11704 683148
rect 11756 683136 11762 683188
rect 3510 670692 3516 670744
rect 3568 670732 3574 670744
rect 14458 670732 14464 670744
rect 3568 670704 14464 670732
rect 3568 670692 3574 670704
rect 14458 670692 14464 670704
rect 14516 670692 14522 670744
rect 3418 658112 3424 658164
rect 3476 658152 3482 658164
rect 7558 658152 7564 658164
rect 3476 658124 7564 658152
rect 3476 658112 3482 658124
rect 7558 658112 7564 658124
rect 7616 658112 7622 658164
rect 3418 632068 3424 632120
rect 3476 632108 3482 632120
rect 17218 632108 17224 632120
rect 3476 632080 17224 632108
rect 3476 632068 3482 632080
rect 17218 632068 17224 632080
rect 17276 632068 17282 632120
rect 3142 618264 3148 618316
rect 3200 618304 3206 618316
rect 15838 618304 15844 618316
rect 3200 618276 15844 618304
rect 3200 618264 3206 618276
rect 15838 618264 15844 618276
rect 15896 618264 15902 618316
rect 3234 605820 3240 605872
rect 3292 605860 3298 605872
rect 90358 605860 90364 605872
rect 3292 605832 90364 605860
rect 3292 605820 3298 605832
rect 90358 605820 90364 605832
rect 90416 605820 90422 605872
rect 74626 598952 74632 599004
rect 74684 598992 74690 599004
rect 98638 598992 98644 599004
rect 74684 598964 98644 598992
rect 74684 598952 74690 598964
rect 98638 598952 98644 598964
rect 98696 598952 98702 599004
rect 349154 598884 349160 598936
rect 349212 598924 349218 598936
rect 349798 598924 349804 598936
rect 349212 598896 349804 598924
rect 349212 598884 349218 598896
rect 349798 598884 349804 598896
rect 349856 598884 349862 598936
rect 70302 597524 70308 597576
rect 70360 597564 70366 597576
rect 349154 597564 349160 597576
rect 70360 597536 349160 597564
rect 70360 597524 70366 597536
rect 349154 597524 349160 597536
rect 349212 597524 349218 597576
rect 67450 596776 67456 596828
rect 67508 596816 67514 596828
rect 170398 596816 170404 596828
rect 67508 596788 170404 596816
rect 67508 596776 67514 596788
rect 170398 596776 170404 596788
rect 170456 596776 170462 596828
rect 86862 594872 86868 594924
rect 86920 594912 86926 594924
rect 113174 594912 113180 594924
rect 86920 594884 113180 594912
rect 86920 594872 86926 594884
rect 113174 594872 113180 594884
rect 113232 594872 113238 594924
rect 65978 594804 65984 594856
rect 66036 594844 66042 594856
rect 295334 594844 295340 594856
rect 66036 594816 295340 594844
rect 66036 594804 66042 594816
rect 295334 594804 295340 594816
rect 295392 594844 295398 594856
rect 295978 594844 295984 594856
rect 295392 594816 295984 594844
rect 295392 594804 295398 594816
rect 295978 594804 295984 594816
rect 296036 594804 296042 594856
rect 90358 594396 90364 594448
rect 90416 594436 90422 594448
rect 91094 594436 91100 594448
rect 90416 594408 91100 594436
rect 90416 594396 90422 594408
rect 91094 594396 91100 594408
rect 91152 594396 91158 594448
rect 40034 594056 40040 594108
rect 40092 594096 40098 594108
rect 89806 594096 89812 594108
rect 40092 594068 89812 594096
rect 40092 594056 40098 594068
rect 89806 594056 89812 594068
rect 89864 594056 89870 594108
rect 73982 593376 73988 593428
rect 74040 593416 74046 593428
rect 116578 593416 116584 593428
rect 74040 593388 116584 593416
rect 74040 593376 74046 593388
rect 116578 593376 116584 593388
rect 116636 593376 116642 593428
rect 25498 592628 25504 592680
rect 25556 592668 25562 592680
rect 80330 592668 80336 592680
rect 25556 592640 80336 592668
rect 25556 592628 25562 592640
rect 80330 592628 80336 592640
rect 80388 592628 80394 592680
rect 75638 592084 75644 592136
rect 75696 592124 75702 592136
rect 96614 592124 96620 592136
rect 75696 592096 96620 592124
rect 75696 592084 75702 592096
rect 96614 592084 96620 592096
rect 96672 592084 96678 592136
rect 84102 592016 84108 592068
rect 84160 592056 84166 592068
rect 112530 592056 112536 592068
rect 84160 592028 112536 592056
rect 84160 592016 84166 592028
rect 112530 592016 112536 592028
rect 112588 592016 112594 592068
rect 7558 591268 7564 591320
rect 7616 591308 7622 591320
rect 69106 591308 69112 591320
rect 7616 591280 69112 591308
rect 7616 591268 7622 591280
rect 69106 591268 69112 591280
rect 69164 591268 69170 591320
rect 70118 590724 70124 590776
rect 70176 590764 70182 590776
rect 73154 590764 73160 590776
rect 70176 590736 73160 590764
rect 70176 590724 70182 590736
rect 73154 590724 73160 590736
rect 73212 590724 73218 590776
rect 86770 590724 86776 590776
rect 86828 590764 86834 590776
rect 115290 590764 115296 590776
rect 86828 590736 115296 590764
rect 86828 590724 86834 590736
rect 115290 590724 115296 590736
rect 115348 590724 115354 590776
rect 69106 590656 69112 590708
rect 69164 590696 69170 590708
rect 70394 590696 70400 590708
rect 69164 590668 70400 590696
rect 69164 590656 69170 590668
rect 70394 590656 70400 590668
rect 70452 590656 70458 590708
rect 73062 590656 73068 590708
rect 73120 590696 73126 590708
rect 81710 590696 81716 590708
rect 73120 590668 81716 590696
rect 73120 590656 73126 590668
rect 81710 590656 81716 590668
rect 81768 590656 81774 590708
rect 85022 590656 85028 590708
rect 85080 590696 85086 590708
rect 86862 590696 86868 590708
rect 85080 590668 86868 590696
rect 85080 590656 85086 590668
rect 86862 590656 86868 590668
rect 86920 590656 86926 590708
rect 204254 590696 204260 590708
rect 86972 590668 204260 590696
rect 86218 590588 86224 590640
rect 86276 590628 86282 590640
rect 86972 590628 87000 590668
rect 204254 590656 204260 590668
rect 204312 590656 204318 590708
rect 86276 590600 87000 590628
rect 86276 590588 86282 590600
rect 70394 589908 70400 589960
rect 70452 589948 70458 589960
rect 89070 589948 89076 589960
rect 70452 589920 89076 589948
rect 70452 589908 70458 589920
rect 89070 589908 89076 589920
rect 89128 589908 89134 589960
rect 100754 589908 100760 589960
rect 100812 589948 100818 589960
rect 111058 589948 111064 589960
rect 100812 589920 111064 589948
rect 100812 589908 100818 589920
rect 111058 589908 111064 589920
rect 111116 589908 111122 589960
rect 3418 589296 3424 589348
rect 3476 589336 3482 589348
rect 74902 589336 74908 589348
rect 3476 589308 74908 589336
rect 3476 589296 3482 589308
rect 74902 589296 74908 589308
rect 74960 589336 74966 589348
rect 75638 589336 75644 589348
rect 74960 589308 75644 589336
rect 74960 589296 74966 589308
rect 75638 589296 75644 589308
rect 75696 589296 75702 589348
rect 76742 589296 76748 589348
rect 76800 589336 76806 589348
rect 100754 589336 100760 589348
rect 76800 589308 100760 589336
rect 76800 589296 76806 589308
rect 100754 589296 100760 589308
rect 100812 589296 100818 589348
rect 187602 589296 187608 589348
rect 187660 589336 187666 589348
rect 255958 589336 255964 589348
rect 187660 589308 255964 589336
rect 187660 589296 187666 589308
rect 255958 589296 255964 589308
rect 256016 589296 256022 589348
rect 79778 588480 79784 588532
rect 79836 588520 79842 588532
rect 79836 588492 93854 588520
rect 79836 588480 79842 588492
rect 72418 588412 72424 588464
rect 72476 588452 72482 588464
rect 72878 588452 72884 588464
rect 72476 588424 72884 588452
rect 72476 588412 72482 588424
rect 72878 588412 72884 588424
rect 72936 588452 72942 588464
rect 72936 588424 74534 588452
rect 72936 588412 72942 588424
rect 74506 587976 74534 588424
rect 80698 588412 80704 588464
rect 80756 588452 80762 588464
rect 89162 588452 89168 588464
rect 80756 588424 89168 588452
rect 80756 588412 80762 588424
rect 89162 588412 89168 588424
rect 89220 588412 89226 588464
rect 77266 588084 84194 588112
rect 77266 587976 77294 588084
rect 74506 587948 77294 587976
rect 55030 587868 55036 587920
rect 55088 587908 55094 587920
rect 66806 587908 66812 587920
rect 55088 587880 66812 587908
rect 55088 587868 55094 587880
rect 66806 587868 66812 587880
rect 66864 587868 66870 587920
rect 84166 587704 84194 588084
rect 93826 587908 93854 588492
rect 105538 587908 105544 587920
rect 93826 587880 105544 587908
rect 105538 587868 105544 587880
rect 105596 587868 105602 587920
rect 93118 587704 93124 587716
rect 84166 587676 93124 587704
rect 93118 587664 93124 587676
rect 93176 587664 93182 587716
rect 88886 587392 88892 587444
rect 88944 587392 88950 587444
rect 88904 587172 88932 587392
rect 88886 587120 88892 587172
rect 88944 587120 88950 587172
rect 89162 586576 89168 586628
rect 89220 586616 89226 586628
rect 106918 586616 106924 586628
rect 89220 586588 106924 586616
rect 89220 586576 89226 586588
rect 106918 586576 106924 586588
rect 106976 586576 106982 586628
rect 59078 586508 59084 586560
rect 59136 586548 59142 586560
rect 66254 586548 66260 586560
rect 59136 586520 66260 586548
rect 59136 586508 59142 586520
rect 66254 586508 66260 586520
rect 66312 586508 66318 586560
rect 91738 586508 91744 586560
rect 91796 586548 91802 586560
rect 95234 586548 95240 586560
rect 91796 586520 95240 586548
rect 91796 586508 91802 586520
rect 95234 586508 95240 586520
rect 95292 586508 95298 586560
rect 57882 585148 57888 585200
rect 57940 585188 57946 585200
rect 66806 585188 66812 585200
rect 57940 585160 66812 585188
rect 57940 585148 57946 585160
rect 66806 585148 66812 585160
rect 66864 585148 66870 585200
rect 67542 585148 67548 585200
rect 67600 585188 67606 585200
rect 68278 585188 68284 585200
rect 67600 585160 68284 585188
rect 67600 585148 67606 585160
rect 68278 585148 68284 585160
rect 68336 585148 68342 585200
rect 91370 584400 91376 584452
rect 91428 584440 91434 584452
rect 95142 584440 95148 584452
rect 91428 584412 95148 584440
rect 91428 584400 91434 584412
rect 95142 584400 95148 584412
rect 95200 584440 95206 584452
rect 132494 584440 132500 584452
rect 95200 584412 132500 584440
rect 95200 584400 95206 584412
rect 132494 584400 132500 584412
rect 132552 584400 132558 584452
rect 91186 583652 91192 583704
rect 91244 583692 91250 583704
rect 99282 583692 99288 583704
rect 91244 583664 99288 583692
rect 91244 583652 91250 583664
rect 99282 583652 99288 583664
rect 99340 583692 99346 583704
rect 104158 583692 104164 583704
rect 99340 583664 104164 583692
rect 99340 583652 99346 583664
rect 104158 583652 104164 583664
rect 104216 583652 104222 583704
rect 48130 582360 48136 582412
rect 48188 582400 48194 582412
rect 66806 582400 66812 582412
rect 48188 582372 66812 582400
rect 48188 582360 48194 582372
rect 66806 582360 66812 582372
rect 66864 582360 66870 582412
rect 64690 581000 64696 581052
rect 64748 581040 64754 581052
rect 66438 581040 66444 581052
rect 64748 581012 66444 581040
rect 64748 581000 64754 581012
rect 66438 581000 66444 581012
rect 66496 581000 66502 581052
rect 91738 581000 91744 581052
rect 91796 581040 91802 581052
rect 142798 581040 142804 581052
rect 91796 581012 142804 581040
rect 91796 581000 91802 581012
rect 142798 581000 142804 581012
rect 142856 581000 142862 581052
rect 52270 579640 52276 579692
rect 52328 579680 52334 579692
rect 66806 579680 66812 579692
rect 52328 579652 66812 579680
rect 52328 579640 52334 579652
rect 66806 579640 66812 579652
rect 66864 579640 66870 579692
rect 91738 579640 91744 579692
rect 91796 579680 91802 579692
rect 108298 579680 108304 579692
rect 91796 579652 108304 579680
rect 91796 579640 91802 579652
rect 108298 579640 108304 579652
rect 108356 579640 108362 579692
rect 91738 578212 91744 578264
rect 91796 578252 91802 578264
rect 120718 578252 120724 578264
rect 91796 578224 120724 578252
rect 91796 578212 91802 578224
rect 120718 578212 120724 578224
rect 120776 578212 120782 578264
rect 17218 576104 17224 576156
rect 17276 576144 17282 576156
rect 67358 576144 67364 576156
rect 17276 576116 67364 576144
rect 17276 576104 17282 576116
rect 67358 576104 67364 576116
rect 67416 576104 67422 576156
rect 91094 576104 91100 576156
rect 91152 576144 91158 576156
rect 123018 576144 123024 576156
rect 91152 576116 123024 576144
rect 91152 576104 91158 576116
rect 123018 576104 123024 576116
rect 123076 576104 123082 576156
rect 61838 574064 61844 574116
rect 61896 574104 61902 574116
rect 67082 574104 67088 574116
rect 61896 574076 67088 574104
rect 61896 574064 61902 574076
rect 67082 574064 67088 574076
rect 67140 574064 67146 574116
rect 91094 574064 91100 574116
rect 91152 574104 91158 574116
rect 97258 574104 97264 574116
rect 91152 574076 97264 574104
rect 91152 574064 91158 574076
rect 97258 574064 97264 574076
rect 97316 574064 97322 574116
rect 60642 571344 60648 571396
rect 60700 571384 60706 571396
rect 66806 571384 66812 571396
rect 60700 571356 66812 571384
rect 60700 571344 60706 571356
rect 66806 571344 66812 571356
rect 66864 571344 66870 571396
rect 91094 571344 91100 571396
rect 91152 571384 91158 571396
rect 115198 571384 115204 571396
rect 91152 571356 115204 571384
rect 91152 571344 91158 571356
rect 115198 571344 115204 571356
rect 115256 571344 115262 571396
rect 149698 571344 149704 571396
rect 149756 571384 149762 571396
rect 266354 571384 266360 571396
rect 149756 571356 266360 571384
rect 149756 571344 149762 571356
rect 266354 571344 266360 571356
rect 266412 571344 266418 571396
rect 91094 569984 91100 570036
rect 91152 570024 91158 570036
rect 94498 570024 94504 570036
rect 91152 569996 94504 570024
rect 91152 569984 91158 569996
rect 94498 569984 94504 569996
rect 94556 569984 94562 570036
rect 93118 569916 93124 569968
rect 93176 569956 93182 569968
rect 353294 569956 353300 569968
rect 93176 569928 353300 569956
rect 93176 569916 93182 569928
rect 353294 569916 353300 569928
rect 353352 569916 353358 569968
rect 67358 569848 67364 569900
rect 67416 569888 67422 569900
rect 68278 569888 68284 569900
rect 67416 569860 68284 569888
rect 67416 569848 67422 569860
rect 68278 569848 68284 569860
rect 68336 569848 68342 569900
rect 91186 569168 91192 569220
rect 91244 569208 91250 569220
rect 126974 569208 126980 569220
rect 91244 569180 126980 569208
rect 91244 569168 91250 569180
rect 126974 569168 126980 569180
rect 127032 569168 127038 569220
rect 63310 568556 63316 568608
rect 63368 568596 63374 568608
rect 66806 568596 66812 568608
rect 63368 568568 66812 568596
rect 63368 568556 63374 568568
rect 66806 568556 66812 568568
rect 66864 568556 66870 568608
rect 91094 568556 91100 568608
rect 91152 568596 91158 568608
rect 100018 568596 100024 568608
rect 91152 568568 100024 568596
rect 91152 568556 91158 568568
rect 100018 568556 100024 568568
rect 100076 568556 100082 568608
rect 126974 568556 126980 568608
rect 127032 568596 127038 568608
rect 213914 568596 213920 568608
rect 127032 568568 213920 568596
rect 127032 568556 127038 568568
rect 213914 568556 213920 568568
rect 213972 568556 213978 568608
rect 273254 567672 273260 567724
rect 273312 567712 273318 567724
rect 273898 567712 273904 567724
rect 273312 567684 273904 567712
rect 273312 567672 273318 567684
rect 273898 567672 273904 567684
rect 273956 567672 273962 567724
rect 133874 567304 133880 567316
rect 122806 567276 133880 567304
rect 64782 567196 64788 567248
rect 64840 567236 64846 567248
rect 66714 567236 66720 567248
rect 64840 567208 66720 567236
rect 64840 567196 64846 567208
rect 66714 567196 66720 567208
rect 66772 567196 66778 567248
rect 89806 567196 89812 567248
rect 89864 567236 89870 567248
rect 122806 567236 122834 567276
rect 133874 567264 133880 567276
rect 133932 567304 133938 567316
rect 209038 567304 209044 567316
rect 133932 567276 209044 567304
rect 133932 567264 133938 567276
rect 209038 567264 209044 567276
rect 209096 567264 209102 567316
rect 89864 567208 122834 567236
rect 89864 567196 89870 567208
rect 197170 567196 197176 567248
rect 197228 567236 197234 567248
rect 273254 567236 273260 567248
rect 197228 567208 273260 567236
rect 197228 567196 197234 567208
rect 273254 567196 273260 567208
rect 273312 567196 273318 567248
rect 53098 566448 53104 566500
rect 53156 566488 53162 566500
rect 67450 566488 67456 566500
rect 53156 566460 67456 566488
rect 53156 566448 53162 566460
rect 67450 566448 67456 566460
rect 67508 566448 67514 566500
rect 94498 566448 94504 566500
rect 94556 566488 94562 566500
rect 137094 566488 137100 566500
rect 94556 566460 137100 566488
rect 94556 566448 94562 566460
rect 137094 566448 137100 566460
rect 137152 566448 137158 566500
rect 3418 565836 3424 565888
rect 3476 565876 3482 565888
rect 43438 565876 43444 565888
rect 3476 565848 43444 565876
rect 3476 565836 3482 565848
rect 43438 565836 43444 565848
rect 43496 565836 43502 565888
rect 91370 565836 91376 565888
rect 91428 565876 91434 565888
rect 102778 565876 102784 565888
rect 91428 565848 102784 565876
rect 91428 565836 91434 565848
rect 102778 565836 102784 565848
rect 102836 565836 102842 565888
rect 136634 565836 136640 565888
rect 136692 565876 136698 565888
rect 137094 565876 137100 565888
rect 136692 565848 137100 565876
rect 136692 565836 136698 565848
rect 137094 565836 137100 565848
rect 137152 565876 137158 565888
rect 291194 565876 291200 565888
rect 137152 565848 291200 565876
rect 137152 565836 137158 565848
rect 291194 565836 291200 565848
rect 291252 565836 291258 565888
rect 177298 564476 177304 564528
rect 177356 564516 177362 564528
rect 259454 564516 259460 564528
rect 177356 564488 259460 564516
rect 177356 564476 177362 564488
rect 259454 564476 259460 564488
rect 259512 564476 259518 564528
rect 50890 564408 50896 564460
rect 50948 564448 50954 564460
rect 66806 564448 66812 564460
rect 50948 564420 66812 564448
rect 50948 564408 50954 564420
rect 66806 564408 66812 564420
rect 66864 564408 66870 564460
rect 91370 564408 91376 564460
rect 91428 564448 91434 564460
rect 107010 564448 107016 564460
rect 91428 564420 107016 564448
rect 91428 564408 91434 564420
rect 107010 564408 107016 564420
rect 107068 564408 107074 564460
rect 115290 564408 115296 564460
rect 115348 564448 115354 564460
rect 117958 564448 117964 564460
rect 115348 564420 117964 564448
rect 115348 564408 115354 564420
rect 117958 564408 117964 564420
rect 118016 564408 118022 564460
rect 166810 564408 166816 564460
rect 166868 564448 166874 564460
rect 298094 564448 298100 564460
rect 166868 564420 298100 564448
rect 166868 564408 166874 564420
rect 298094 564408 298100 564420
rect 298152 564408 298158 564460
rect 195882 563116 195888 563168
rect 195940 563156 195946 563168
rect 271874 563156 271880 563168
rect 195940 563128 271880 563156
rect 195940 563116 195946 563128
rect 271874 563116 271880 563128
rect 271932 563116 271938 563168
rect 50982 563048 50988 563100
rect 51040 563088 51046 563100
rect 66806 563088 66812 563100
rect 51040 563060 66812 563088
rect 51040 563048 51046 563060
rect 66806 563048 66812 563060
rect 66864 563048 66870 563100
rect 91370 563048 91376 563100
rect 91428 563088 91434 563100
rect 134702 563088 134708 563100
rect 91428 563060 134708 563088
rect 91428 563048 91434 563060
rect 134702 563048 134708 563060
rect 134760 563048 134766 563100
rect 206278 563048 206284 563100
rect 206336 563088 206342 563100
rect 582834 563088 582840 563100
rect 206336 563060 582840 563088
rect 206336 563048 206342 563060
rect 582834 563048 582840 563060
rect 582892 563048 582898 563100
rect 52362 561688 52368 561740
rect 52420 561728 52426 561740
rect 66806 561728 66812 561740
rect 52420 561700 66812 561728
rect 52420 561688 52426 561700
rect 66806 561688 66812 561700
rect 66864 561688 66870 561740
rect 111058 561688 111064 561740
rect 111116 561728 111122 561740
rect 111702 561728 111708 561740
rect 111116 561700 111708 561728
rect 111116 561688 111122 561700
rect 111702 561688 111708 561700
rect 111760 561728 111766 561740
rect 358906 561728 358912 561740
rect 111760 561700 358912 561728
rect 111760 561688 111766 561700
rect 358906 561688 358912 561700
rect 358964 561688 358970 561740
rect 263594 561620 263600 561672
rect 263652 561660 263658 561672
rect 264238 561660 264244 561672
rect 263652 561632 264244 561660
rect 263652 561620 263658 561632
rect 264238 561620 264244 561632
rect 264296 561620 264302 561672
rect 197078 560328 197084 560380
rect 197136 560368 197142 560380
rect 288434 560368 288440 560380
rect 197136 560340 288440 560368
rect 197136 560328 197142 560340
rect 288434 560328 288440 560340
rect 288492 560328 288498 560380
rect 41322 560260 41328 560312
rect 41380 560300 41386 560312
rect 66806 560300 66812 560312
rect 41380 560272 66812 560300
rect 41380 560260 41386 560272
rect 66806 560260 66812 560272
rect 66864 560260 66870 560312
rect 146938 560260 146944 560312
rect 146996 560300 147002 560312
rect 263594 560300 263600 560312
rect 146996 560272 263600 560300
rect 146996 560260 147002 560272
rect 263594 560260 263600 560272
rect 263652 560260 263658 560312
rect 192478 558968 192484 559020
rect 192536 559008 192542 559020
rect 287054 559008 287060 559020
rect 192536 558980 287060 559008
rect 192536 558968 192542 558980
rect 287054 558968 287060 558980
rect 287112 558968 287118 559020
rect 63402 558900 63408 558952
rect 63460 558940 63466 558952
rect 66806 558940 66812 558952
rect 63460 558912 66812 558940
rect 63460 558900 63466 558912
rect 66806 558900 66812 558912
rect 66864 558900 66870 558952
rect 89622 558900 89628 558952
rect 89680 558940 89686 558952
rect 122098 558940 122104 558952
rect 89680 558912 122104 558940
rect 89680 558900 89686 558912
rect 122098 558900 122104 558912
rect 122156 558900 122162 558952
rect 160002 558900 160008 558952
rect 160060 558940 160066 558952
rect 309134 558940 309140 558952
rect 160060 558912 309140 558940
rect 160060 558900 160066 558912
rect 309134 558900 309140 558912
rect 309192 558900 309198 558952
rect 59170 558424 59176 558476
rect 59228 558464 59234 558476
rect 62022 558464 62028 558476
rect 59228 558436 62028 558464
rect 59228 558424 59234 558436
rect 62022 558424 62028 558436
rect 62080 558424 62086 558476
rect 97258 558152 97264 558204
rect 97316 558192 97322 558204
rect 122926 558192 122932 558204
rect 97316 558164 122932 558192
rect 97316 558152 97322 558164
rect 122926 558152 122932 558164
rect 122984 558152 122990 558204
rect 198826 558152 198832 558204
rect 198884 558192 198890 558204
rect 331214 558192 331220 558204
rect 198884 558164 331220 558192
rect 198884 558152 198890 558164
rect 331214 558152 331220 558164
rect 331272 558152 331278 558204
rect 62022 557540 62028 557592
rect 62080 557580 62086 557592
rect 66806 557580 66812 557592
rect 62080 557552 66812 557580
rect 62080 557540 62086 557552
rect 66806 557540 66812 557552
rect 66864 557540 66870 557592
rect 195422 557540 195428 557592
rect 195480 557580 195486 557592
rect 357434 557580 357440 557592
rect 195480 557552 357440 557580
rect 195480 557540 195486 557552
rect 357434 557540 357440 557552
rect 357492 557540 357498 557592
rect 92382 556792 92388 556844
rect 92440 556832 92446 556844
rect 152458 556832 152464 556844
rect 92440 556804 152464 556832
rect 92440 556792 92446 556804
rect 152458 556792 152464 556804
rect 152516 556792 152522 556844
rect 204254 556792 204260 556844
rect 204312 556832 204318 556844
rect 582374 556832 582380 556844
rect 204312 556804 582380 556832
rect 204312 556792 204318 556804
rect 582374 556792 582380 556804
rect 582432 556792 582438 556844
rect 91186 556180 91192 556232
rect 91244 556220 91250 556232
rect 121454 556220 121460 556232
rect 91244 556192 121460 556220
rect 91244 556180 91250 556192
rect 121454 556180 121460 556192
rect 121512 556180 121518 556232
rect 181530 556180 181536 556232
rect 181588 556220 181594 556232
rect 251818 556220 251824 556232
rect 181588 556192 251824 556220
rect 181588 556180 181594 556192
rect 251818 556180 251824 556192
rect 251876 556180 251882 556232
rect 324314 555228 324320 555280
rect 324372 555268 324378 555280
rect 324866 555268 324872 555280
rect 324372 555240 324872 555268
rect 324372 555228 324378 555240
rect 324866 555228 324872 555240
rect 324924 555268 324930 555280
rect 327718 555268 327724 555280
rect 324924 555240 327724 555268
rect 324924 555228 324930 555240
rect 327718 555228 327724 555240
rect 327776 555228 327782 555280
rect 187050 554820 187056 554872
rect 187108 554860 187114 554872
rect 324314 554860 324320 554872
rect 187108 554832 324320 554860
rect 187108 554820 187114 554832
rect 324314 554820 324320 554832
rect 324372 554820 324378 554872
rect 53650 554752 53656 554804
rect 53708 554792 53714 554804
rect 66806 554792 66812 554804
rect 53708 554764 66812 554792
rect 53708 554752 53714 554764
rect 66806 554752 66812 554764
rect 66864 554752 66870 554804
rect 91738 554752 91744 554804
rect 91796 554792 91802 554804
rect 106182 554792 106188 554804
rect 91796 554764 106188 554792
rect 91796 554752 91802 554764
rect 106182 554752 106188 554764
rect 106240 554792 106246 554804
rect 244918 554792 244924 554804
rect 106240 554764 244924 554792
rect 106240 554752 106246 554764
rect 244918 554752 244924 554764
rect 244976 554752 244982 554804
rect 49602 554004 49608 554056
rect 49660 554044 49666 554056
rect 65978 554044 65984 554056
rect 49660 554016 65984 554044
rect 49660 554004 49666 554016
rect 65978 554004 65984 554016
rect 66036 554044 66042 554056
rect 66530 554044 66536 554056
rect 66036 554016 66536 554044
rect 66036 554004 66042 554016
rect 66530 554004 66536 554016
rect 66588 554004 66594 554056
rect 198550 554004 198556 554056
rect 198608 554044 198614 554056
rect 583018 554044 583024 554056
rect 198608 554016 583024 554044
rect 198608 554004 198614 554016
rect 583018 554004 583024 554016
rect 583076 554004 583082 554056
rect 91738 553392 91744 553444
rect 91796 553432 91802 553444
rect 112438 553432 112444 553444
rect 91796 553404 112444 553432
rect 91796 553392 91802 553404
rect 112438 553392 112444 553404
rect 112496 553392 112502 553444
rect 188338 553392 188344 553444
rect 188396 553432 188402 553444
rect 270494 553432 270500 553444
rect 188396 553404 270500 553432
rect 188396 553392 188402 553404
rect 270494 553392 270500 553404
rect 270552 553392 270558 553444
rect 91738 552100 91744 552152
rect 91796 552140 91802 552152
rect 97350 552140 97356 552152
rect 91796 552112 97356 552140
rect 91796 552100 91802 552112
rect 97350 552100 97356 552112
rect 97408 552100 97414 552152
rect 193858 552100 193864 552152
rect 193916 552140 193922 552152
rect 296714 552140 296720 552152
rect 193916 552112 296720 552140
rect 193916 552100 193922 552112
rect 296714 552100 296720 552112
rect 296772 552100 296778 552152
rect 91186 552032 91192 552084
rect 91244 552072 91250 552084
rect 100110 552072 100116 552084
rect 91244 552044 100116 552072
rect 91244 552032 91250 552044
rect 100110 552032 100116 552044
rect 100168 552032 100174 552084
rect 112530 552032 112536 552084
rect 112588 552072 112594 552084
rect 226978 552072 226984 552084
rect 112588 552044 226984 552072
rect 112588 552032 112594 552044
rect 226978 552032 226984 552044
rect 227036 552032 227042 552084
rect 198642 551284 198648 551336
rect 198700 551324 198706 551336
rect 582742 551324 582748 551336
rect 198700 551296 582748 551324
rect 198700 551284 198706 551296
rect 582742 551284 582748 551296
rect 582800 551284 582806 551336
rect 91186 550604 91192 550656
rect 91244 550644 91250 550656
rect 108942 550644 108948 550656
rect 91244 550616 108948 550644
rect 91244 550604 91250 550616
rect 108942 550604 108948 550616
rect 109000 550644 109006 550656
rect 124858 550644 124864 550656
rect 109000 550616 124864 550644
rect 109000 550604 109006 550616
rect 124858 550604 124864 550616
rect 124916 550604 124922 550656
rect 180150 550604 180156 550656
rect 180208 550644 180214 550656
rect 229094 550644 229100 550656
rect 180208 550616 229100 550644
rect 180208 550604 180214 550616
rect 229094 550604 229100 550616
rect 229152 550604 229158 550656
rect 295978 549856 295984 549908
rect 296036 549896 296042 549908
rect 351914 549896 351920 549908
rect 296036 549868 351920 549896
rect 296036 549856 296042 549868
rect 351914 549856 351920 549868
rect 351972 549856 351978 549908
rect 161382 549312 161388 549364
rect 161440 549352 161446 549364
rect 215386 549352 215392 549364
rect 161440 549324 215392 549352
rect 161440 549312 161446 549324
rect 215386 549312 215392 549324
rect 215444 549312 215450 549364
rect 56502 549244 56508 549296
rect 56560 549284 56566 549296
rect 66438 549284 66444 549296
rect 56560 549256 66444 549284
rect 56560 549244 56566 549256
rect 66438 549244 66444 549256
rect 66496 549244 66502 549296
rect 189810 549244 189816 549296
rect 189868 549284 189874 549296
rect 304994 549284 305000 549296
rect 189868 549256 305000 549284
rect 189868 549244 189874 549256
rect 304994 549244 305000 549256
rect 305052 549244 305058 549296
rect 180058 547952 180064 548004
rect 180116 547992 180122 548004
rect 285122 547992 285128 548004
rect 180116 547964 285128 547992
rect 180116 547952 180122 547964
rect 285122 547952 285128 547964
rect 285180 547952 285186 548004
rect 59262 547884 59268 547936
rect 59320 547924 59326 547936
rect 66438 547924 66444 547936
rect 59320 547896 66444 547924
rect 59320 547884 59326 547896
rect 66438 547884 66444 547896
rect 66496 547884 66502 547936
rect 91462 547884 91468 547936
rect 91520 547924 91526 547936
rect 95326 547924 95332 547936
rect 91520 547896 95332 547924
rect 91520 547884 91526 547896
rect 95326 547884 95332 547896
rect 95384 547884 95390 547936
rect 184198 547884 184204 547936
rect 184256 547924 184262 547936
rect 343634 547924 343640 547936
rect 184256 547896 343640 547924
rect 184256 547884 184262 547896
rect 343634 547884 343640 547896
rect 343692 547884 343698 547936
rect 95326 547136 95332 547188
rect 95384 547176 95390 547188
rect 245654 547176 245660 547188
rect 95384 547148 245660 547176
rect 95384 547136 95390 547148
rect 245654 547136 245660 547148
rect 245712 547136 245718 547188
rect 91186 546456 91192 546508
rect 91244 546496 91250 546508
rect 97258 546496 97264 546508
rect 91244 546468 97264 546496
rect 91244 546456 91250 546468
rect 97258 546456 97264 546468
rect 97316 546456 97322 546508
rect 126882 546456 126888 546508
rect 126940 546496 126946 546508
rect 339954 546496 339960 546508
rect 126940 546468 339960 546496
rect 126940 546456 126946 546468
rect 339954 546456 339960 546468
rect 340012 546456 340018 546508
rect 185578 545164 185584 545216
rect 185636 545204 185642 545216
rect 220814 545204 220820 545216
rect 185636 545176 220820 545204
rect 185636 545164 185642 545176
rect 220814 545164 220820 545176
rect 220872 545164 220878 545216
rect 48222 545096 48228 545148
rect 48280 545136 48286 545148
rect 66806 545136 66812 545148
rect 48280 545108 66812 545136
rect 48280 545096 48286 545108
rect 66806 545096 66812 545108
rect 66864 545096 66870 545148
rect 91186 545096 91192 545148
rect 91244 545136 91250 545148
rect 94498 545136 94504 545148
rect 91244 545108 94504 545136
rect 91244 545096 91250 545108
rect 94498 545096 94504 545108
rect 94556 545096 94562 545148
rect 188430 545096 188436 545148
rect 188488 545136 188494 545148
rect 290090 545136 290096 545148
rect 188488 545108 290096 545136
rect 188488 545096 188494 545108
rect 290090 545096 290096 545108
rect 290148 545096 290154 545148
rect 328454 545096 328460 545148
rect 328512 545136 328518 545148
rect 375466 545136 375472 545148
rect 328512 545108 375472 545136
rect 328512 545096 328518 545108
rect 375466 545096 375472 545108
rect 375524 545096 375530 545148
rect 194134 543804 194140 543856
rect 194192 543844 194198 543856
rect 223666 543844 223672 543856
rect 194192 543816 223672 543844
rect 194192 543804 194198 543816
rect 223666 543804 223672 543816
rect 223724 543804 223730 543856
rect 330018 543804 330024 543856
rect 330076 543844 330082 543856
rect 364426 543844 364432 543856
rect 330076 543816 364432 543844
rect 330076 543804 330082 543816
rect 364426 543804 364432 543816
rect 364484 543804 364490 543856
rect 55122 543736 55128 543788
rect 55180 543776 55186 543788
rect 66806 543776 66812 543788
rect 55180 543748 66812 543776
rect 55180 543736 55186 543748
rect 66806 543736 66812 543748
rect 66864 543736 66870 543788
rect 91830 543736 91836 543788
rect 91888 543776 91894 543788
rect 93670 543776 93676 543788
rect 91888 543748 93676 543776
rect 91888 543736 91894 543748
rect 93670 543736 93676 543748
rect 93728 543776 93734 543788
rect 284294 543776 284300 543788
rect 93728 543748 284300 543776
rect 93728 543736 93734 543748
rect 284294 543736 284300 543748
rect 284352 543736 284358 543788
rect 311894 543736 311900 543788
rect 311952 543776 311958 543788
rect 356238 543776 356244 543788
rect 311952 543748 356244 543776
rect 311952 543736 311958 543748
rect 356238 543736 356244 543748
rect 356296 543736 356302 543788
rect 11698 542988 11704 543040
rect 11756 543028 11762 543040
rect 36538 543028 36544 543040
rect 11756 543000 36544 543028
rect 11756 542988 11762 543000
rect 36538 542988 36544 543000
rect 36596 542988 36602 543040
rect 166902 542444 166908 542496
rect 166960 542484 166966 542496
rect 306650 542484 306656 542496
rect 166960 542456 306656 542484
rect 166960 542444 166966 542456
rect 306650 542444 306656 542456
rect 306708 542444 306714 542496
rect 338298 542444 338304 542496
rect 338356 542484 338362 542496
rect 363046 542484 363052 542496
rect 338356 542456 363052 542484
rect 338356 542444 338362 542456
rect 363046 542444 363052 542456
rect 363104 542444 363110 542496
rect 36538 542376 36544 542428
rect 36596 542416 36602 542428
rect 37182 542416 37188 542428
rect 36596 542388 37188 542416
rect 36596 542376 36602 542388
rect 37182 542376 37188 542388
rect 37240 542416 37246 542428
rect 66806 542416 66812 542428
rect 37240 542388 66812 542416
rect 37240 542376 37246 542388
rect 66806 542376 66812 542388
rect 66864 542376 66870 542428
rect 91186 542376 91192 542428
rect 91244 542416 91250 542428
rect 98730 542416 98736 542428
rect 91244 542388 98736 542416
rect 91244 542376 91250 542388
rect 98730 542376 98736 542388
rect 98788 542376 98794 542428
rect 195238 542376 195244 542428
rect 195296 542416 195302 542428
rect 356146 542416 356152 542428
rect 195296 542388 356152 542416
rect 195296 542376 195302 542388
rect 356146 542376 356152 542388
rect 356204 542376 356210 542428
rect 209038 542308 209044 542360
rect 209096 542348 209102 542360
rect 210418 542348 210424 542360
rect 209096 542320 210424 542348
rect 209096 542308 209102 542320
rect 210418 542308 210424 542320
rect 210476 542308 210482 542360
rect 244918 542308 244924 542360
rect 244976 542348 244982 542360
rect 247034 542348 247040 542360
rect 244976 542320 247040 542348
rect 244976 542308 244982 542320
rect 247034 542308 247040 542320
rect 247092 542308 247098 542360
rect 14458 541628 14464 541680
rect 14516 541668 14522 541680
rect 67082 541668 67088 541680
rect 14516 541640 67088 541668
rect 14516 541628 14522 541640
rect 67082 541628 67088 541640
rect 67140 541668 67146 541680
rect 67358 541668 67364 541680
rect 67140 541640 67364 541668
rect 67140 541628 67146 541640
rect 67358 541628 67364 541640
rect 67416 541628 67422 541680
rect 91186 541628 91192 541680
rect 91244 541668 91250 541680
rect 128354 541668 128360 541680
rect 91244 541640 128360 541668
rect 91244 541628 91250 541640
rect 128354 541628 128360 541640
rect 128412 541628 128418 541680
rect 199470 541628 199476 541680
rect 199528 541668 199534 541680
rect 204254 541668 204260 541680
rect 199528 541640 204260 541668
rect 199528 541628 199534 541640
rect 204254 541628 204260 541640
rect 204312 541668 204318 541680
rect 207014 541668 207020 541680
rect 204312 541640 207020 541668
rect 204312 541628 204318 541640
rect 207014 541628 207020 541640
rect 207072 541628 207078 541680
rect 331674 541016 331680 541068
rect 331732 541056 331738 541068
rect 360286 541056 360292 541068
rect 331732 541028 360292 541056
rect 331732 541016 331738 541028
rect 360286 541016 360292 541028
rect 360344 541016 360350 541068
rect 128354 540948 128360 541000
rect 128412 540988 128418 541000
rect 129642 540988 129648 541000
rect 128412 540960 129648 540988
rect 128412 540948 128418 540960
rect 129642 540948 129648 540960
rect 129700 540988 129706 541000
rect 258442 540988 258448 541000
rect 129700 540960 258448 540988
rect 129700 540948 129706 540960
rect 258442 540948 258448 540960
rect 258500 540948 258506 541000
rect 316586 540948 316592 541000
rect 316644 540988 316650 541000
rect 364518 540988 364524 541000
rect 316644 540960 364524 540988
rect 316644 540948 316650 540960
rect 364518 540948 364524 540960
rect 364576 540948 364582 541000
rect 3418 540200 3424 540252
rect 3476 540240 3482 540252
rect 3476 540212 64874 540240
rect 3476 540200 3482 540212
rect 64846 539696 64874 540212
rect 67266 539724 67272 539776
rect 67324 539764 67330 539776
rect 67324 539736 71912 539764
rect 67324 539724 67330 539736
rect 64846 539668 70440 539696
rect 70412 539640 70440 539668
rect 71884 539640 71912 539736
rect 88168 539668 93854 539696
rect 88168 539640 88196 539668
rect 61930 539588 61936 539640
rect 61988 539628 61994 539640
rect 67542 539628 67548 539640
rect 61988 539600 67548 539628
rect 61988 539588 61994 539600
rect 67542 539588 67548 539600
rect 67600 539588 67606 539640
rect 70394 539588 70400 539640
rect 70452 539588 70458 539640
rect 71866 539588 71872 539640
rect 71924 539588 71930 539640
rect 88150 539588 88156 539640
rect 88208 539588 88214 539640
rect 92382 539588 92388 539640
rect 92440 539628 92446 539640
rect 93210 539628 93216 539640
rect 92440 539600 93216 539628
rect 92440 539588 92446 539600
rect 93210 539588 93216 539600
rect 93268 539588 93274 539640
rect 93826 539628 93854 539668
rect 129642 539656 129648 539708
rect 129700 539696 129706 539708
rect 357526 539696 357532 539708
rect 129700 539668 357532 539696
rect 129700 539656 129706 539668
rect 357526 539656 357532 539668
rect 357584 539656 357590 539708
rect 250622 539628 250628 539640
rect 93826 539600 250628 539628
rect 250622 539588 250628 539600
rect 250680 539588 250686 539640
rect 347682 539588 347688 539640
rect 347740 539628 347746 539640
rect 580258 539628 580264 539640
rect 347740 539600 580264 539628
rect 347740 539588 347746 539600
rect 580258 539588 580264 539600
rect 580316 539588 580322 539640
rect 67450 539520 67456 539572
rect 67508 539520 67514 539572
rect 273898 539520 273904 539572
rect 273956 539560 273962 539572
rect 275646 539560 275652 539572
rect 273956 539532 275652 539560
rect 273956 539520 273962 539532
rect 275646 539520 275652 539532
rect 275704 539520 275710 539572
rect 278038 539520 278044 539572
rect 278096 539560 278102 539572
rect 278958 539560 278964 539572
rect 278096 539532 278964 539560
rect 278096 539520 278102 539532
rect 278958 539520 278964 539532
rect 279016 539520 279022 539572
rect 67468 539368 67496 539520
rect 270862 539452 270868 539504
rect 270920 539492 270926 539504
rect 273990 539492 273996 539504
rect 270920 539464 273996 539492
rect 270920 539452 270926 539464
rect 273990 539452 273996 539464
rect 274048 539452 274054 539504
rect 67450 539316 67456 539368
rect 67508 539316 67514 539368
rect 57790 538908 57796 538960
rect 57848 538948 57854 538960
rect 65794 538948 65800 538960
rect 57848 538920 65800 538948
rect 57848 538908 57854 538920
rect 65794 538908 65800 538920
rect 65852 538948 65858 538960
rect 65978 538948 65984 538960
rect 65852 538920 65984 538948
rect 65852 538908 65858 538920
rect 65978 538908 65984 538920
rect 66036 538908 66042 538960
rect 175918 538908 175924 538960
rect 175976 538948 175982 538960
rect 194134 538948 194140 538960
rect 175976 538920 194140 538948
rect 175976 538908 175982 538920
rect 194134 538908 194140 538920
rect 194192 538908 194198 538960
rect 3418 538840 3424 538892
rect 3476 538880 3482 538892
rect 89714 538880 89720 538892
rect 3476 538852 89720 538880
rect 3476 538840 3482 538852
rect 89714 538840 89720 538852
rect 89772 538840 89778 538892
rect 157978 538840 157984 538892
rect 158036 538880 158042 538892
rect 195238 538880 195244 538892
rect 158036 538852 195244 538880
rect 158036 538840 158042 538852
rect 195238 538840 195244 538852
rect 195296 538840 195302 538892
rect 199378 538296 199384 538348
rect 199436 538336 199442 538348
rect 255590 538336 255596 538348
rect 199436 538308 255596 538336
rect 199436 538296 199442 538308
rect 255590 538296 255596 538308
rect 255648 538296 255654 538348
rect 347038 538296 347044 538348
rect 347096 538336 347102 538348
rect 359090 538336 359096 538348
rect 347096 538308 359096 538336
rect 347096 538296 347102 538308
rect 359090 538296 359096 538308
rect 359148 538296 359154 538348
rect 65978 538228 65984 538280
rect 66036 538268 66042 538280
rect 76742 538268 76748 538280
rect 66036 538240 76748 538268
rect 66036 538228 66042 538240
rect 76742 538228 76748 538240
rect 76800 538228 76806 538280
rect 195238 538228 195244 538280
rect 195296 538268 195302 538280
rect 216674 538268 216680 538280
rect 195296 538240 216680 538268
rect 195296 538228 195302 538240
rect 216674 538228 216680 538240
rect 216732 538228 216738 538280
rect 220906 538228 220912 538280
rect 220964 538268 220970 538280
rect 356330 538268 356336 538280
rect 220964 538240 356336 538268
rect 220964 538228 220970 538240
rect 356330 538228 356336 538240
rect 356388 538228 356394 538280
rect 88610 538160 88616 538212
rect 88668 538200 88674 538212
rect 89622 538200 89628 538212
rect 88668 538172 89628 538200
rect 88668 538160 88674 538172
rect 89622 538160 89628 538172
rect 89680 538160 89686 538212
rect 130378 538200 130384 538212
rect 93826 538172 130384 538200
rect 86862 538092 86868 538144
rect 86920 538132 86926 538144
rect 93826 538132 93854 538172
rect 130378 538160 130384 538172
rect 130436 538160 130442 538212
rect 86920 538104 93854 538132
rect 86920 538092 86926 538104
rect 8202 537480 8208 537532
rect 8260 537520 8266 537532
rect 91278 537520 91284 537532
rect 8260 537492 91284 537520
rect 8260 537480 8266 537492
rect 91278 537480 91284 537492
rect 91336 537480 91342 537532
rect 198090 537480 198096 537532
rect 198148 537520 198154 537532
rect 220906 537520 220912 537532
rect 198148 537492 220912 537520
rect 198148 537480 198154 537492
rect 220906 537480 220912 537492
rect 220964 537480 220970 537532
rect 323670 537480 323676 537532
rect 323728 537520 323734 537532
rect 580166 537520 580172 537532
rect 323728 537492 580172 537520
rect 323728 537480 323734 537492
rect 580166 537480 580172 537492
rect 580224 537480 580230 537532
rect 178770 536800 178776 536852
rect 178828 536840 178834 536852
rect 233878 536840 233884 536852
rect 178828 536812 233884 536840
rect 178828 536800 178834 536812
rect 233878 536800 233884 536812
rect 233936 536840 233942 536852
rect 234062 536840 234068 536852
rect 233936 536812 234068 536840
rect 233936 536800 233942 536812
rect 234062 536800 234068 536812
rect 234120 536800 234126 536852
rect 337102 536800 337108 536852
rect 337160 536840 337166 536852
rect 371326 536840 371332 536852
rect 337160 536812 371332 536840
rect 337160 536800 337166 536812
rect 371326 536800 371332 536812
rect 371384 536800 371390 536852
rect 43438 536732 43444 536784
rect 43496 536772 43502 536784
rect 69566 536772 69572 536784
rect 43496 536744 69572 536772
rect 43496 536732 43502 536744
rect 69566 536732 69572 536744
rect 69624 536732 69630 536784
rect 75178 536732 75184 536784
rect 75236 536772 75242 536784
rect 129642 536772 129648 536784
rect 75236 536744 129648 536772
rect 75236 536732 75242 536744
rect 129642 536732 129648 536744
rect 129700 536732 129706 536784
rect 84286 536460 84292 536512
rect 84344 536500 84350 536512
rect 89070 536500 89076 536512
rect 84344 536472 89076 536500
rect 84344 536460 84350 536472
rect 89070 536460 89076 536472
rect 89128 536460 89134 536512
rect 15838 536052 15844 536104
rect 15896 536092 15902 536104
rect 43990 536092 43996 536104
rect 15896 536064 43996 536092
rect 15896 536052 15902 536064
rect 43990 536052 43996 536064
rect 44048 536092 44054 536104
rect 73154 536092 73160 536104
rect 44048 536064 73160 536092
rect 44048 536052 44054 536064
rect 73154 536052 73160 536064
rect 73212 536052 73218 536104
rect 81526 535576 81532 535628
rect 81584 535616 81590 535628
rect 83458 535616 83464 535628
rect 81584 535588 83464 535616
rect 81584 535576 81590 535588
rect 83458 535576 83464 535588
rect 83516 535576 83522 535628
rect 198734 535576 198740 535628
rect 198792 535616 198798 535628
rect 200390 535616 200396 535628
rect 198792 535588 200396 535616
rect 198792 535576 198798 535588
rect 200390 535576 200396 535588
rect 200448 535576 200454 535628
rect 130470 535508 130476 535560
rect 130528 535548 130534 535560
rect 308398 535548 308404 535560
rect 130528 535520 308404 535548
rect 130528 535508 130534 535520
rect 308398 535508 308404 535520
rect 308456 535508 308462 535560
rect 327442 535508 327448 535560
rect 327500 535548 327506 535560
rect 361666 535548 361672 535560
rect 327500 535520 361672 535548
rect 327500 535508 327506 535520
rect 361666 535508 361672 535520
rect 361724 535508 361730 535560
rect 89622 535440 89628 535492
rect 89680 535480 89686 535492
rect 90450 535480 90456 535492
rect 89680 535452 90456 535480
rect 89680 535440 89686 535452
rect 90450 535440 90456 535452
rect 90508 535440 90514 535492
rect 201402 535440 201408 535492
rect 201460 535480 201466 535492
rect 208670 535480 208676 535492
rect 201460 535452 208676 535480
rect 201460 535440 201466 535452
rect 208670 535440 208676 535452
rect 208728 535440 208734 535492
rect 247586 535440 247592 535492
rect 247644 535480 247650 535492
rect 582374 535480 582380 535492
rect 247644 535452 582380 535480
rect 247644 535440 247650 535452
rect 582374 535440 582380 535452
rect 582432 535440 582438 535492
rect 202046 535276 202052 535288
rect 200086 535248 202052 535276
rect 175182 534760 175188 534812
rect 175240 534800 175246 534812
rect 200086 534800 200114 535248
rect 202046 535236 202052 535248
rect 202104 535236 202110 535288
rect 175240 534772 200114 534800
rect 175240 534760 175246 534772
rect 11698 534692 11704 534744
rect 11756 534732 11762 534744
rect 91186 534732 91192 534744
rect 11756 534704 91192 534732
rect 11756 534692 11762 534704
rect 91186 534692 91192 534704
rect 91244 534692 91250 534744
rect 67726 534012 67732 534064
rect 67784 534052 67790 534064
rect 76558 534052 76564 534064
rect 67784 534024 76564 534052
rect 67784 534012 67790 534024
rect 76558 534012 76564 534024
rect 76616 534012 76622 534064
rect 164142 533332 164148 533384
rect 164200 533372 164206 533384
rect 191190 533372 191196 533384
rect 164200 533344 191196 533372
rect 164200 533332 164206 533344
rect 191190 533332 191196 533344
rect 191248 533332 191254 533384
rect 77846 532788 77852 532840
rect 77904 532828 77910 532840
rect 100938 532828 100944 532840
rect 77904 532800 100944 532828
rect 77904 532788 77910 532800
rect 100938 532788 100944 532800
rect 100996 532788 101002 532840
rect 48130 532720 48136 532772
rect 48188 532760 48194 532772
rect 162854 532760 162860 532772
rect 48188 532732 162860 532760
rect 48188 532720 48194 532732
rect 162854 532720 162860 532732
rect 162912 532760 162918 532772
rect 164142 532760 164148 532772
rect 162912 532732 164148 532760
rect 162912 532720 162918 532732
rect 164142 532720 164148 532732
rect 164200 532720 164206 532772
rect 100938 532652 100944 532704
rect 100996 532692 101002 532704
rect 197354 532692 197360 532704
rect 100996 532664 197360 532692
rect 100996 532652 101002 532664
rect 197354 532652 197360 532664
rect 197412 532652 197418 532704
rect 17862 531972 17868 532024
rect 17920 532012 17926 532024
rect 91094 532012 91100 532024
rect 17920 531984 91100 532012
rect 17920 531972 17926 531984
rect 91094 531972 91100 531984
rect 91152 531972 91158 532024
rect 358722 531972 358728 532024
rect 358780 532012 358786 532024
rect 358906 532012 358912 532024
rect 358780 531984 358912 532012
rect 358780 531972 358786 531984
rect 358906 531972 358912 531984
rect 358964 532012 358970 532024
rect 582742 532012 582748 532024
rect 358964 531984 582748 532012
rect 358964 531972 358970 531984
rect 582742 531972 582748 531984
rect 582800 531972 582806 532024
rect 41322 531224 41328 531276
rect 41380 531264 41386 531276
rect 195422 531264 195428 531276
rect 41380 531236 195428 531264
rect 41380 531224 41386 531236
rect 195422 531224 195428 531236
rect 195480 531224 195486 531276
rect 64690 530544 64696 530596
rect 64748 530584 64754 530596
rect 79318 530584 79324 530596
rect 64748 530556 79324 530584
rect 64748 530544 64754 530556
rect 79318 530544 79324 530556
rect 79376 530544 79382 530596
rect 177390 529864 177396 529916
rect 177448 529904 177454 529916
rect 197354 529904 197360 529916
rect 177448 529876 197360 529904
rect 177448 529864 177454 529876
rect 197354 529864 197360 529876
rect 197412 529864 197418 529916
rect 59078 529252 59084 529304
rect 59136 529292 59142 529304
rect 85574 529292 85580 529304
rect 59136 529264 85580 529292
rect 59136 529252 59142 529264
rect 85574 529252 85580 529264
rect 85632 529252 85638 529304
rect 80054 529184 80060 529236
rect 80112 529224 80118 529236
rect 129734 529224 129740 529236
rect 80112 529196 129740 529224
rect 80112 529184 80118 529196
rect 129734 529184 129740 529196
rect 129792 529184 129798 529236
rect 129734 528572 129740 528624
rect 129792 528612 129798 528624
rect 177298 528612 177304 528624
rect 129792 528584 177304 528612
rect 129792 528572 129798 528584
rect 177298 528572 177304 528584
rect 177356 528572 177362 528624
rect 124858 528504 124864 528556
rect 124916 528544 124922 528556
rect 197354 528544 197360 528556
rect 124916 528516 197360 528544
rect 124916 528504 124922 528516
rect 197354 528504 197360 528516
rect 197412 528504 197418 528556
rect 70486 527484 70492 527536
rect 70544 527524 70550 527536
rect 71038 527524 71044 527536
rect 70544 527496 71044 527524
rect 70544 527484 70550 527496
rect 71038 527484 71044 527496
rect 71096 527484 71102 527536
rect 71038 527144 71044 527196
rect 71096 527184 71102 527196
rect 124950 527184 124956 527196
rect 71096 527156 124956 527184
rect 71096 527144 71102 527156
rect 124950 527144 124956 527156
rect 125008 527144 125014 527196
rect 358722 527144 358728 527196
rect 358780 527184 358786 527196
rect 367094 527184 367100 527196
rect 358780 527156 367100 527184
rect 358780 527144 358786 527156
rect 367094 527144 367100 527156
rect 367152 527144 367158 527196
rect 34422 525036 34428 525088
rect 34480 525076 34486 525088
rect 197998 525076 198004 525088
rect 34480 525048 198004 525076
rect 34480 525036 34486 525048
rect 197998 525036 198004 525048
rect 198056 525036 198062 525088
rect 358722 524424 358728 524476
rect 358780 524464 358786 524476
rect 378226 524464 378232 524476
rect 358780 524436 378232 524464
rect 358780 524424 358786 524436
rect 378226 524424 378232 524436
rect 378284 524424 378290 524476
rect 66898 523676 66904 523728
rect 66956 523716 66962 523728
rect 188430 523716 188436 523728
rect 66956 523688 188436 523716
rect 66956 523676 66962 523688
rect 188430 523676 188436 523688
rect 188488 523676 188494 523728
rect 189718 522248 189724 522300
rect 189776 522288 189782 522300
rect 197446 522288 197452 522300
rect 189776 522260 197452 522288
rect 189776 522248 189782 522260
rect 197446 522248 197452 522260
rect 197504 522248 197510 522300
rect 358722 522248 358728 522300
rect 358780 522288 358786 522300
rect 582374 522288 582380 522300
rect 358780 522260 582380 522288
rect 358780 522248 358786 522260
rect 582374 522248 582380 522260
rect 582432 522248 582438 522300
rect 147582 521636 147588 521688
rect 147640 521676 147646 521688
rect 197354 521676 197360 521688
rect 147640 521648 197360 521676
rect 147640 521636 147646 521648
rect 197354 521636 197360 521648
rect 197412 521636 197418 521688
rect 46842 520888 46848 520940
rect 46900 520928 46906 520940
rect 195330 520928 195336 520940
rect 46900 520900 195336 520928
rect 46900 520888 46906 520900
rect 195330 520888 195336 520900
rect 195388 520888 195394 520940
rect 56502 520208 56508 520260
rect 56560 520248 56566 520260
rect 189810 520248 189816 520260
rect 56560 520220 189816 520248
rect 56560 520208 56566 520220
rect 189810 520208 189816 520220
rect 189868 520208 189874 520260
rect 357894 520004 357900 520056
rect 357952 520044 357958 520056
rect 360194 520044 360200 520056
rect 357952 520016 360200 520044
rect 357952 520004 357958 520016
rect 360194 520004 360200 520016
rect 360252 520004 360258 520056
rect 162118 518916 162124 518968
rect 162176 518956 162182 518968
rect 197354 518956 197360 518968
rect 162176 518928 197360 518956
rect 162176 518916 162182 518928
rect 197354 518916 197360 518928
rect 197412 518916 197418 518968
rect 39942 518168 39948 518220
rect 40000 518208 40006 518220
rect 184382 518208 184388 518220
rect 40000 518180 184388 518208
rect 40000 518168 40006 518180
rect 184382 518168 184388 518180
rect 184440 518168 184446 518220
rect 66162 517420 66168 517472
rect 66220 517460 66226 517472
rect 187050 517460 187056 517472
rect 66220 517432 187056 517460
rect 66220 517420 66226 517432
rect 187050 517420 187056 517432
rect 187108 517420 187114 517472
rect 176010 516128 176016 516180
rect 176068 516168 176074 516180
rect 197354 516168 197360 516180
rect 176068 516140 197360 516168
rect 176068 516128 176074 516140
rect 197354 516128 197360 516140
rect 197412 516128 197418 516180
rect 358722 516128 358728 516180
rect 358780 516168 358786 516180
rect 375374 516168 375380 516180
rect 358780 516140 375380 516168
rect 358780 516128 358786 516140
rect 375374 516128 375380 516140
rect 375432 516128 375438 516180
rect 2774 514768 2780 514820
rect 2832 514808 2838 514820
rect 4798 514808 4804 514820
rect 2832 514780 4804 514808
rect 2832 514768 2838 514780
rect 4798 514768 4804 514780
rect 4856 514768 4862 514820
rect 358630 514768 358636 514820
rect 358688 514808 358694 514820
rect 360194 514808 360200 514820
rect 358688 514780 360200 514808
rect 358688 514768 358694 514780
rect 360194 514768 360200 514780
rect 360252 514768 360258 514820
rect 45462 514020 45468 514072
rect 45520 514060 45526 514072
rect 191098 514060 191104 514072
rect 45520 514032 191104 514060
rect 45520 514020 45526 514032
rect 191098 514020 191104 514032
rect 191156 514020 191162 514072
rect 156598 512592 156604 512644
rect 156656 512632 156662 512644
rect 199470 512632 199476 512644
rect 156656 512604 199476 512632
rect 156656 512592 156662 512604
rect 199470 512592 199476 512604
rect 199528 512592 199534 512644
rect 124950 510552 124956 510604
rect 125008 510592 125014 510604
rect 197354 510592 197360 510604
rect 125008 510564 197360 510592
rect 125008 510552 125014 510564
rect 197354 510552 197360 510564
rect 197412 510552 197418 510604
rect 169018 506472 169024 506524
rect 169076 506512 169082 506524
rect 197354 506512 197360 506524
rect 169076 506484 197360 506512
rect 169076 506472 169082 506484
rect 197354 506472 197360 506484
rect 197412 506472 197418 506524
rect 357618 505724 357624 505776
rect 357676 505764 357682 505776
rect 367186 505764 367192 505776
rect 357676 505736 367192 505764
rect 357676 505724 357682 505736
rect 367186 505724 367192 505736
rect 367244 505724 367250 505776
rect 358722 505112 358728 505164
rect 358780 505152 358786 505164
rect 385034 505152 385040 505164
rect 358780 505124 385040 505152
rect 358780 505112 358786 505124
rect 385034 505112 385040 505124
rect 385092 505112 385098 505164
rect 358722 502324 358728 502376
rect 358780 502364 358786 502376
rect 369946 502364 369952 502376
rect 358780 502336 369952 502364
rect 358780 502324 358786 502336
rect 369946 502324 369952 502336
rect 370004 502324 370010 502376
rect 3510 502256 3516 502308
rect 3568 502296 3574 502308
rect 11698 502296 11704 502308
rect 3568 502268 11704 502296
rect 3568 502256 3574 502268
rect 11698 502256 11704 502268
rect 11756 502256 11762 502308
rect 177298 500896 177304 500948
rect 177356 500936 177362 500948
rect 197354 500936 197360 500948
rect 177356 500908 197360 500936
rect 177356 500896 177362 500908
rect 197354 500896 197360 500908
rect 197412 500896 197418 500948
rect 358722 499536 358728 499588
rect 358780 499576 358786 499588
rect 371418 499576 371424 499588
rect 358780 499548 371424 499576
rect 358780 499536 358786 499548
rect 371418 499536 371424 499548
rect 371476 499536 371482 499588
rect 356330 496748 356336 496800
rect 356388 496788 356394 496800
rect 357158 496788 357164 496800
rect 356388 496760 357164 496788
rect 356388 496748 356394 496760
rect 357158 496748 357164 496760
rect 357216 496788 357222 496800
rect 582926 496788 582932 496800
rect 357216 496760 582932 496788
rect 357216 496748 357222 496760
rect 582926 496748 582932 496760
rect 582984 496748 582990 496800
rect 188430 495456 188436 495508
rect 188488 495496 188494 495508
rect 197354 495496 197360 495508
rect 188488 495468 197360 495496
rect 188488 495456 188494 495468
rect 197354 495456 197360 495468
rect 197412 495456 197418 495508
rect 358630 493960 358636 494012
rect 358688 494000 358694 494012
rect 412634 494000 412640 494012
rect 358688 493972 412640 494000
rect 358688 493960 358694 493972
rect 412634 493960 412640 493972
rect 412692 493960 412698 494012
rect 130378 492668 130384 492720
rect 130436 492708 130442 492720
rect 197354 492708 197360 492720
rect 130436 492680 197360 492708
rect 130436 492668 130442 492680
rect 197354 492668 197360 492680
rect 197412 492668 197418 492720
rect 152550 489880 152556 489932
rect 152608 489920 152614 489932
rect 197354 489920 197360 489932
rect 152608 489892 197360 489920
rect 152608 489880 152614 489892
rect 197354 489880 197360 489892
rect 197412 489880 197418 489932
rect 152458 487772 152464 487824
rect 152516 487812 152522 487824
rect 180794 487812 180800 487824
rect 152516 487784 180800 487812
rect 152516 487772 152522 487784
rect 180794 487772 180800 487784
rect 180852 487812 180858 487824
rect 182082 487812 182088 487824
rect 180852 487784 182088 487812
rect 180852 487772 180858 487784
rect 182082 487772 182088 487784
rect 182140 487772 182146 487824
rect 182082 487160 182088 487212
rect 182140 487200 182146 487212
rect 197354 487200 197360 487212
rect 182140 487172 197360 487200
rect 182140 487160 182146 487172
rect 197354 487160 197360 487172
rect 197412 487160 197418 487212
rect 358722 487160 358728 487212
rect 358780 487200 358786 487212
rect 372614 487200 372620 487212
rect 358780 487172 372620 487200
rect 358780 487160 358786 487172
rect 372614 487160 372620 487172
rect 372672 487160 372678 487212
rect 358722 484372 358728 484424
rect 358780 484412 358786 484424
rect 369854 484412 369860 484424
rect 358780 484384 369860 484412
rect 358780 484372 358786 484384
rect 369854 484372 369860 484384
rect 369912 484372 369918 484424
rect 191098 480428 191104 480480
rect 191156 480468 191162 480480
rect 197354 480468 197360 480480
rect 191156 480440 197360 480468
rect 191156 480428 191162 480440
rect 197354 480428 197360 480440
rect 197412 480428 197418 480480
rect 116578 478116 116584 478168
rect 116636 478156 116642 478168
rect 128446 478156 128452 478168
rect 116636 478128 128452 478156
rect 116636 478116 116642 478128
rect 128446 478116 128452 478128
rect 128504 478116 128510 478168
rect 128446 477504 128452 477556
rect 128504 477544 128510 477556
rect 176654 477544 176660 477556
rect 128504 477516 176660 477544
rect 128504 477504 128510 477516
rect 176654 477504 176660 477516
rect 176712 477544 176718 477556
rect 197354 477544 197360 477556
rect 176712 477516 197360 477544
rect 176712 477504 176718 477516
rect 197354 477504 197360 477516
rect 197412 477504 197418 477556
rect 358722 477504 358728 477556
rect 358780 477544 358786 477556
rect 362954 477544 362960 477556
rect 358780 477516 362960 477544
rect 358780 477504 358786 477516
rect 362954 477504 362960 477516
rect 363012 477504 363018 477556
rect 147122 476756 147128 476808
rect 147180 476796 147186 476808
rect 198090 476796 198096 476808
rect 147180 476768 198096 476796
rect 147180 476756 147186 476768
rect 198090 476756 198096 476768
rect 198148 476756 198154 476808
rect 68278 476076 68284 476128
rect 68336 476116 68342 476128
rect 68922 476116 68928 476128
rect 68336 476088 68928 476116
rect 68336 476076 68342 476088
rect 68922 476076 68928 476088
rect 68980 476116 68986 476128
rect 147122 476116 147128 476128
rect 68980 476088 147128 476116
rect 68980 476076 68986 476088
rect 147122 476076 147128 476088
rect 147180 476116 147186 476128
rect 147490 476116 147496 476128
rect 147180 476088 147496 476116
rect 147180 476076 147186 476088
rect 147490 476076 147496 476088
rect 147548 476076 147554 476128
rect 3326 475328 3332 475380
rect 3384 475368 3390 475380
rect 8202 475368 8208 475380
rect 3384 475340 8208 475368
rect 3384 475328 3390 475340
rect 8202 475328 8208 475340
rect 8260 475368 8266 475380
rect 25498 475368 25504 475380
rect 8260 475340 25504 475368
rect 8260 475328 8266 475340
rect 25498 475328 25504 475340
rect 25556 475328 25562 475380
rect 144178 474716 144184 474768
rect 144236 474756 144242 474768
rect 197354 474756 197360 474768
rect 144236 474728 197360 474756
rect 144236 474716 144242 474728
rect 197354 474716 197360 474728
rect 197412 474716 197418 474768
rect 358722 474716 358728 474768
rect 358780 474756 358786 474768
rect 375558 474756 375564 474768
rect 358780 474728 375564 474756
rect 358780 474716 358786 474728
rect 375558 474716 375564 474728
rect 375616 474716 375622 474768
rect 140038 473356 140044 473408
rect 140096 473396 140102 473408
rect 197354 473396 197360 473408
rect 140096 473368 197360 473396
rect 140096 473356 140102 473368
rect 197354 473356 197360 473368
rect 197412 473356 197418 473408
rect 358722 471996 358728 472048
rect 358780 472036 358786 472048
rect 368566 472036 368572 472048
rect 358780 472008 368572 472036
rect 358780 471996 358786 472008
rect 368566 471996 368572 472008
rect 368624 471996 368630 472048
rect 195790 470704 195796 470756
rect 195848 470744 195854 470756
rect 197630 470744 197636 470756
rect 195848 470716 197636 470744
rect 195848 470704 195854 470716
rect 197630 470704 197636 470716
rect 197688 470704 197694 470756
rect 358722 470568 358728 470620
rect 358780 470608 358786 470620
rect 380894 470608 380900 470620
rect 358780 470580 380900 470608
rect 358780 470568 358786 470580
rect 380894 470568 380900 470580
rect 380952 470568 380958 470620
rect 165522 467848 165528 467900
rect 165580 467888 165586 467900
rect 197354 467888 197360 467900
rect 165580 467860 197360 467888
rect 165580 467848 165586 467860
rect 197354 467848 197360 467860
rect 197412 467848 197418 467900
rect 358722 467848 358728 467900
rect 358780 467888 358786 467900
rect 363138 467888 363144 467900
rect 358780 467860 363144 467888
rect 358780 467848 358786 467860
rect 363138 467848 363144 467860
rect 363196 467848 363202 467900
rect 105538 467780 105544 467832
rect 105596 467820 105602 467832
rect 187510 467820 187516 467832
rect 105596 467792 187516 467820
rect 105596 467780 105602 467792
rect 187510 467780 187516 467792
rect 187568 467820 187574 467832
rect 191190 467820 191196 467832
rect 187568 467792 191196 467820
rect 187568 467780 187574 467792
rect 191190 467780 191196 467792
rect 191248 467780 191254 467832
rect 62022 467100 62028 467152
rect 62080 467140 62086 467152
rect 95234 467140 95240 467152
rect 62080 467112 95240 467140
rect 62080 467100 62086 467112
rect 95234 467100 95240 467112
rect 95292 467100 95298 467152
rect 104894 466420 104900 466472
rect 104952 466460 104958 466472
rect 105538 466460 105544 466472
rect 104952 466432 105544 466460
rect 104952 466420 104958 466432
rect 105538 466420 105544 466432
rect 105596 466420 105602 466472
rect 60458 465672 60464 465724
rect 60516 465712 60522 465724
rect 78766 465712 78772 465724
rect 60516 465684 78772 465712
rect 60516 465672 60522 465684
rect 78766 465672 78772 465684
rect 78824 465672 78830 465724
rect 124950 465060 124956 465112
rect 125008 465100 125014 465112
rect 171042 465100 171048 465112
rect 125008 465072 171048 465100
rect 125008 465060 125014 465072
rect 171042 465060 171048 465072
rect 171100 465100 171106 465112
rect 197354 465100 197360 465112
rect 171100 465072 197360 465100
rect 171100 465060 171106 465072
rect 197354 465060 197360 465072
rect 197412 465060 197418 465112
rect 356330 465060 356336 465112
rect 356388 465100 356394 465112
rect 356790 465100 356796 465112
rect 356388 465072 356796 465100
rect 356388 465060 356394 465072
rect 356790 465060 356796 465072
rect 356848 465100 356854 465112
rect 582374 465100 582380 465112
rect 356848 465072 582380 465100
rect 356848 465060 356854 465072
rect 582374 465060 582380 465072
rect 582432 465060 582438 465112
rect 358078 464992 358084 465044
rect 358136 465032 358142 465044
rect 365714 465032 365720 465044
rect 358136 465004 365720 465032
rect 358136 464992 358142 465004
rect 365714 464992 365720 465004
rect 365772 464992 365778 465044
rect 106182 464312 106188 464364
rect 106240 464352 106246 464364
rect 120810 464352 120816 464364
rect 106240 464324 120816 464352
rect 106240 464312 106246 464324
rect 120810 464312 120816 464324
rect 120868 464312 120874 464364
rect 64782 463700 64788 463752
rect 64840 463740 64846 463752
rect 180242 463740 180248 463752
rect 64840 463712 180248 463740
rect 64840 463700 64846 463712
rect 180242 463700 180248 463712
rect 180300 463700 180306 463752
rect 93762 462952 93768 463004
rect 93820 462992 93826 463004
rect 107654 462992 107660 463004
rect 93820 462964 107660 462992
rect 93820 462952 93826 462964
rect 107654 462952 107660 462964
rect 107712 462952 107718 463004
rect 3510 462340 3516 462392
rect 3568 462380 3574 462392
rect 14550 462380 14556 462392
rect 3568 462352 14556 462380
rect 3568 462340 3574 462352
rect 14550 462340 14556 462352
rect 14608 462340 14614 462392
rect 127618 462340 127624 462392
rect 127676 462380 127682 462392
rect 197354 462380 197360 462392
rect 127676 462352 197360 462380
rect 127676 462340 127682 462352
rect 197354 462340 197360 462352
rect 197412 462340 197418 462392
rect 358722 462340 358728 462392
rect 358780 462380 358786 462392
rect 385126 462380 385132 462392
rect 358780 462352 385132 462380
rect 358780 462340 358786 462352
rect 385126 462340 385132 462352
rect 385184 462340 385190 462392
rect 59078 461660 59084 461712
rect 59136 461700 59142 461712
rect 72418 461700 72424 461712
rect 59136 461672 72424 461700
rect 59136 461660 59142 461672
rect 72418 461660 72424 461672
rect 72476 461660 72482 461712
rect 52270 461592 52276 461644
rect 52328 461632 52334 461644
rect 78030 461632 78036 461644
rect 52328 461604 78036 461632
rect 52328 461592 52334 461604
rect 78030 461592 78036 461604
rect 78088 461592 78094 461644
rect 76006 461456 76012 461508
rect 76064 461496 76070 461508
rect 76558 461496 76564 461508
rect 76064 461468 76564 461496
rect 76064 461456 76070 461468
rect 76558 461456 76564 461468
rect 76616 461456 76622 461508
rect 76558 460912 76564 460964
rect 76616 460952 76622 460964
rect 173894 460952 173900 460964
rect 76616 460924 173900 460952
rect 76616 460912 76622 460924
rect 173894 460912 173900 460924
rect 173952 460912 173958 460964
rect 65978 460164 65984 460216
rect 66036 460204 66042 460216
rect 77938 460204 77944 460216
rect 66036 460176 77944 460204
rect 66036 460164 66042 460176
rect 77938 460164 77944 460176
rect 77996 460164 78002 460216
rect 143442 460164 143448 460216
rect 143500 460204 143506 460216
rect 197354 460204 197360 460216
rect 143500 460176 197360 460204
rect 143500 460164 143506 460176
rect 197354 460164 197360 460176
rect 197412 460164 197418 460216
rect 370038 460164 370044 460216
rect 370096 460204 370102 460216
rect 582558 460204 582564 460216
rect 370096 460176 582564 460204
rect 370096 460164 370102 460176
rect 582558 460164 582564 460176
rect 582616 460164 582622 460216
rect 142798 459552 142804 459604
rect 142856 459592 142862 459604
rect 143442 459592 143448 459604
rect 142856 459564 143448 459592
rect 142856 459552 142862 459564
rect 143442 459552 143448 459564
rect 143500 459552 143506 459604
rect 358446 459552 358452 459604
rect 358504 459592 358510 459604
rect 370038 459592 370044 459604
rect 358504 459564 370044 459592
rect 358504 459552 358510 459564
rect 370038 459552 370044 459564
rect 370096 459552 370102 459604
rect 4798 459484 4804 459536
rect 4856 459524 4862 459536
rect 112530 459524 112536 459536
rect 4856 459496 112536 459524
rect 4856 459484 4862 459496
rect 112530 459484 112536 459496
rect 112588 459484 112594 459536
rect 64782 458804 64788 458856
rect 64840 458844 64846 458856
rect 73246 458844 73252 458856
rect 64840 458816 73252 458844
rect 64840 458804 64846 458816
rect 73246 458804 73252 458816
rect 73304 458804 73310 458856
rect 131758 458192 131764 458244
rect 131816 458232 131822 458244
rect 197354 458232 197360 458244
rect 131816 458204 197360 458232
rect 131816 458192 131822 458204
rect 197354 458192 197360 458204
rect 197412 458192 197418 458244
rect 108298 458124 108304 458176
rect 108356 458164 108362 458176
rect 115290 458164 115296 458176
rect 108356 458136 115296 458164
rect 108356 458124 108362 458136
rect 115290 458124 115296 458136
rect 115348 458124 115354 458176
rect 52270 456764 52276 456816
rect 52328 456804 52334 456816
rect 67634 456804 67640 456816
rect 52328 456776 67640 456804
rect 52328 456764 52334 456776
rect 67634 456764 67640 456776
rect 67692 456804 67698 456816
rect 68830 456804 68836 456816
rect 67692 456776 68836 456804
rect 67692 456764 67698 456776
rect 68830 456764 68836 456776
rect 68888 456764 68894 456816
rect 63310 456016 63316 456068
rect 63368 456056 63374 456068
rect 67634 456056 67640 456068
rect 63368 456028 67640 456056
rect 63368 456016 63374 456028
rect 67634 456016 67640 456028
rect 67692 456056 67698 456068
rect 68646 456056 68652 456068
rect 67692 456028 68652 456056
rect 67692 456016 67698 456028
rect 68646 456016 68652 456028
rect 68704 456016 68710 456068
rect 68830 456016 68836 456068
rect 68888 456056 68894 456068
rect 81434 456056 81440 456068
rect 68888 456028 81440 456056
rect 68888 456016 68894 456028
rect 81434 456016 81440 456028
rect 81492 456016 81498 456068
rect 68646 455404 68652 455456
rect 68704 455444 68710 455456
rect 185670 455444 185676 455456
rect 68704 455416 185676 455444
rect 68704 455404 68710 455416
rect 185670 455404 185676 455416
rect 185728 455404 185734 455456
rect 358722 455404 358728 455456
rect 358780 455444 358786 455456
rect 387794 455444 387800 455456
rect 358780 455416 387800 455444
rect 358780 455404 358786 455416
rect 387794 455404 387800 455416
rect 387852 455444 387858 455456
rect 582834 455444 582840 455456
rect 387852 455416 582840 455444
rect 387852 455404 387858 455416
rect 582834 455404 582840 455416
rect 582892 455404 582898 455456
rect 55030 455336 55036 455388
rect 55088 455376 55094 455388
rect 56410 455376 56416 455388
rect 55088 455348 56416 455376
rect 55088 455336 55094 455348
rect 56410 455336 56416 455348
rect 56468 455336 56474 455388
rect 63310 454656 63316 454708
rect 63368 454696 63374 454708
rect 75914 454696 75920 454708
rect 63368 454668 75920 454696
rect 63368 454656 63374 454668
rect 75914 454656 75920 454668
rect 75972 454656 75978 454708
rect 102778 454656 102784 454708
rect 102836 454696 102842 454708
rect 125594 454696 125600 454708
rect 102836 454668 125600 454696
rect 102836 454656 102842 454668
rect 125594 454656 125600 454668
rect 125652 454656 125658 454708
rect 56410 454044 56416 454096
rect 56468 454084 56474 454096
rect 87046 454084 87052 454096
rect 56468 454056 87052 454084
rect 56468 454044 56474 454056
rect 87046 454044 87052 454056
rect 87104 454044 87110 454096
rect 17218 453976 17224 454028
rect 17276 454016 17282 454028
rect 17862 454016 17868 454028
rect 17276 453988 17868 454016
rect 17276 453976 17282 453988
rect 17862 453976 17868 453988
rect 17920 453976 17926 454028
rect 65610 453296 65616 453348
rect 65668 453336 65674 453348
rect 75178 453336 75184 453348
rect 65668 453308 75184 453336
rect 65668 453296 65674 453308
rect 75178 453296 75184 453308
rect 75236 453296 75242 453348
rect 17218 452616 17224 452668
rect 17276 452656 17282 452668
rect 124214 452656 124220 452668
rect 17276 452628 124220 452656
rect 17276 452616 17282 452628
rect 124214 452616 124220 452628
rect 124272 452616 124278 452668
rect 358722 452616 358728 452668
rect 358780 452656 358786 452668
rect 376754 452656 376760 452668
rect 358780 452628 376760 452656
rect 358780 452616 358786 452628
rect 376754 452616 376760 452628
rect 376812 452616 376818 452668
rect 3418 451868 3424 451920
rect 3476 451908 3482 451920
rect 121546 451908 121552 451920
rect 3476 451880 121552 451908
rect 3476 451868 3482 451880
rect 121546 451868 121552 451880
rect 121604 451908 121610 451920
rect 124950 451908 124956 451920
rect 121604 451880 124956 451908
rect 121604 451868 121610 451880
rect 124950 451868 124956 451880
rect 125008 451868 125014 451920
rect 116118 451256 116124 451308
rect 116176 451296 116182 451308
rect 156598 451296 156604 451308
rect 116176 451268 156604 451296
rect 116176 451256 116182 451268
rect 156598 451256 156604 451268
rect 156656 451256 156662 451308
rect 66070 450576 66076 450628
rect 66128 450616 66134 450628
rect 91094 450616 91100 450628
rect 66128 450588 91100 450616
rect 66128 450576 66134 450588
rect 91094 450576 91100 450588
rect 91152 450576 91158 450628
rect 48130 450508 48136 450560
rect 48188 450548 48194 450560
rect 80882 450548 80888 450560
rect 48188 450520 80888 450548
rect 48188 450508 48194 450520
rect 80882 450508 80888 450520
rect 80940 450508 80946 450560
rect 96246 450508 96252 450560
rect 96304 450548 96310 450560
rect 128446 450548 128452 450560
rect 96304 450520 128452 450548
rect 96304 450508 96310 450520
rect 128446 450508 128452 450520
rect 128504 450508 128510 450560
rect 91094 449896 91100 449948
rect 91152 449936 91158 449948
rect 91554 449936 91560 449948
rect 91152 449908 91560 449936
rect 91152 449896 91158 449908
rect 91554 449896 91560 449908
rect 91612 449936 91618 449948
rect 159450 449936 159456 449948
rect 91612 449908 159456 449936
rect 91612 449896 91618 449908
rect 159450 449896 159456 449908
rect 159508 449896 159514 449948
rect 358722 449896 358728 449948
rect 358780 449936 358786 449948
rect 364334 449936 364340 449948
rect 358780 449908 364340 449936
rect 358780 449896 358786 449908
rect 364334 449896 364340 449908
rect 364392 449896 364398 449948
rect 106918 449828 106924 449880
rect 106976 449868 106982 449880
rect 131758 449868 131764 449880
rect 106976 449840 131764 449868
rect 106976 449828 106982 449840
rect 131758 449828 131764 449840
rect 131816 449828 131822 449880
rect 115198 449352 115204 449404
rect 115256 449392 115262 449404
rect 120626 449392 120632 449404
rect 115256 449364 120632 449392
rect 115256 449352 115262 449364
rect 120626 449352 120632 449364
rect 120684 449352 120690 449404
rect 57698 449216 57704 449268
rect 57756 449256 57762 449268
rect 78674 449256 78680 449268
rect 57756 449228 78680 449256
rect 57756 449216 57762 449228
rect 78674 449216 78680 449228
rect 78732 449216 78738 449268
rect 14550 449148 14556 449200
rect 14608 449188 14614 449200
rect 68830 449188 68836 449200
rect 14608 449160 68836 449188
rect 14608 449148 14614 449160
rect 68830 449148 68836 449160
rect 68888 449148 68894 449200
rect 368382 449148 368388 449200
rect 368440 449188 368446 449200
rect 582466 449188 582472 449200
rect 368440 449160 582472 449188
rect 368440 449148 368446 449160
rect 582466 449148 582472 449160
rect 582524 449148 582530 449200
rect 3142 448536 3148 448588
rect 3200 448576 3206 448588
rect 14458 448576 14464 448588
rect 3200 448548 14464 448576
rect 3200 448536 3206 448548
rect 14458 448536 14464 448548
rect 14516 448536 14522 448588
rect 68830 448536 68836 448588
rect 68888 448576 68894 448588
rect 103514 448576 103520 448588
rect 68888 448548 103520 448576
rect 68888 448536 68894 448548
rect 103514 448536 103520 448548
rect 103572 448576 103578 448588
rect 103698 448576 103704 448588
rect 103572 448548 103704 448576
rect 103572 448536 103578 448548
rect 103698 448536 103704 448548
rect 103756 448536 103762 448588
rect 168282 448536 168288 448588
rect 168340 448576 168346 448588
rect 197354 448576 197360 448588
rect 168340 448548 197360 448576
rect 168340 448536 168346 448548
rect 197354 448536 197360 448548
rect 197412 448536 197418 448588
rect 358722 448536 358728 448588
rect 358780 448576 358786 448588
rect 367278 448576 367284 448588
rect 358780 448548 367284 448576
rect 358780 448536 358786 448548
rect 367278 448536 367284 448548
rect 367336 448576 367342 448588
rect 368382 448576 368388 448588
rect 367336 448548 368388 448576
rect 367336 448536 367342 448548
rect 368382 448536 368388 448548
rect 368440 448536 368446 448588
rect 57882 447788 57888 447840
rect 57940 447828 57946 447840
rect 83826 447828 83832 447840
rect 57940 447800 83832 447828
rect 57940 447788 57946 447800
rect 83826 447788 83832 447800
rect 83884 447788 83890 447840
rect 94774 447788 94780 447840
rect 94832 447828 94838 447840
rect 127618 447828 127624 447840
rect 94832 447800 127624 447828
rect 94832 447788 94838 447800
rect 127618 447788 127624 447800
rect 127676 447788 127682 447840
rect 164878 447788 164884 447840
rect 164936 447828 164942 447840
rect 192570 447828 192576 447840
rect 164936 447800 192576 447828
rect 164936 447788 164942 447800
rect 192570 447788 192576 447800
rect 192628 447788 192634 447840
rect 65886 447108 65892 447160
rect 65944 447148 65950 447160
rect 71038 447148 71044 447160
rect 65944 447120 71044 447148
rect 65944 447108 65950 447120
rect 71038 447108 71044 447120
rect 71096 447108 71102 447160
rect 88886 447108 88892 447160
rect 88944 447148 88950 447160
rect 132586 447148 132592 447160
rect 88944 447120 132592 447148
rect 88944 447108 88950 447120
rect 132586 447108 132592 447120
rect 132644 447108 132650 447160
rect 68922 447040 68928 447092
rect 68980 447080 68986 447092
rect 73154 447080 73160 447092
rect 68980 447052 73160 447080
rect 68980 447040 68986 447052
rect 73154 447040 73160 447052
rect 73212 447040 73218 447092
rect 79318 447040 79324 447092
rect 79376 447080 79382 447092
rect 130470 447080 130476 447092
rect 79376 447052 130476 447080
rect 79376 447040 79382 447052
rect 130470 447040 130476 447052
rect 130528 447040 130534 447092
rect 48038 446360 48044 446412
rect 48096 446400 48102 446412
rect 71866 446400 71872 446412
rect 48096 446372 71872 446400
rect 48096 446360 48102 446372
rect 71866 446360 71872 446372
rect 71924 446400 71930 446412
rect 74810 446400 74816 446412
rect 71924 446372 74816 446400
rect 71924 446360 71930 446372
rect 74810 446360 74816 446372
rect 74868 446360 74874 446412
rect 90358 445748 90364 445800
rect 90416 445788 90422 445800
rect 96522 445788 96528 445800
rect 90416 445760 96528 445788
rect 90416 445748 90422 445760
rect 96522 445748 96528 445760
rect 96580 445748 96586 445800
rect 100846 445748 100852 445800
rect 100904 445788 100910 445800
rect 102226 445788 102232 445800
rect 100904 445760 102232 445788
rect 100904 445748 100910 445760
rect 102226 445748 102232 445760
rect 102284 445748 102290 445800
rect 112530 445748 112536 445800
rect 112588 445788 112594 445800
rect 112898 445788 112904 445800
rect 112588 445760 112904 445788
rect 112588 445748 112594 445760
rect 112898 445748 112904 445760
rect 112956 445788 112962 445800
rect 142890 445788 142896 445800
rect 112956 445760 142896 445788
rect 112956 445748 112962 445760
rect 142890 445748 142896 445760
rect 142948 445748 142954 445800
rect 144270 445748 144276 445800
rect 144328 445788 144334 445800
rect 197354 445788 197360 445800
rect 144328 445760 197360 445788
rect 144328 445748 144334 445760
rect 197354 445748 197360 445760
rect 197412 445748 197418 445800
rect 60550 444456 60556 444508
rect 60608 444496 60614 444508
rect 93026 444496 93032 444508
rect 60608 444468 93032 444496
rect 60608 444456 60614 444468
rect 93026 444456 93032 444468
rect 93084 444456 93090 444508
rect 100754 444456 100760 444508
rect 100812 444496 100818 444508
rect 127618 444496 127624 444508
rect 100812 444468 127624 444496
rect 100812 444456 100818 444468
rect 127618 444456 127624 444468
rect 127676 444456 127682 444508
rect 4798 444388 4804 444440
rect 4856 444428 4862 444440
rect 118694 444428 118700 444440
rect 4856 444400 118700 444428
rect 4856 444388 4862 444400
rect 118694 444388 118700 444400
rect 118752 444428 118758 444440
rect 119154 444428 119160 444440
rect 118752 444400 119160 444428
rect 118752 444388 118758 444400
rect 119154 444388 119160 444400
rect 119212 444428 119218 444440
rect 121638 444428 121644 444440
rect 119212 444400 121644 444428
rect 119212 444388 119218 444400
rect 121638 444388 121644 444400
rect 121696 444388 121702 444440
rect 147490 444320 147496 444372
rect 147548 444360 147554 444372
rect 148318 444360 148324 444372
rect 147548 444332 148324 444360
rect 147548 444320 147554 444332
rect 148318 444320 148324 444332
rect 148376 444320 148382 444372
rect 168374 443640 168380 443692
rect 168432 443680 168438 443692
rect 184290 443680 184296 443692
rect 168432 443652 184296 443680
rect 168432 443640 168438 443652
rect 184290 443640 184296 443652
rect 184348 443640 184354 443692
rect 184382 443640 184388 443692
rect 184440 443680 184446 443692
rect 197354 443680 197360 443692
rect 184440 443652 197360 443680
rect 184440 443640 184446 443652
rect 197354 443640 197360 443652
rect 197412 443640 197418 443692
rect 125502 442960 125508 443012
rect 125560 443000 125566 443012
rect 168374 443000 168380 443012
rect 125560 442972 168380 443000
rect 125560 442960 125566 442972
rect 168374 442960 168380 442972
rect 168432 442960 168438 443012
rect 358722 442960 358728 443012
rect 358780 443000 358786 443012
rect 383654 443000 383660 443012
rect 358780 442972 383660 443000
rect 358780 442960 358786 442972
rect 383654 442960 383660 442972
rect 383712 442960 383718 443012
rect 67358 442892 67364 442944
rect 67416 442932 67422 442944
rect 67818 442932 67824 442944
rect 67416 442904 67824 442932
rect 67416 442892 67422 442904
rect 67818 442892 67824 442904
rect 67876 442892 67882 442944
rect 124122 442008 124128 442060
rect 124180 442048 124186 442060
rect 131758 442048 131764 442060
rect 124180 442020 131764 442048
rect 124180 442008 124186 442020
rect 131758 442008 131764 442020
rect 131816 442008 131822 442060
rect 185670 441532 185676 441584
rect 185728 441572 185734 441584
rect 197354 441572 197360 441584
rect 185728 441544 197360 441572
rect 185728 441532 185734 441544
rect 197354 441532 197360 441544
rect 197412 441532 197418 441584
rect 358722 440240 358728 440292
rect 358780 440280 358786 440292
rect 368474 440280 368480 440292
rect 358780 440252 368480 440280
rect 358780 440240 358786 440252
rect 368474 440240 368480 440252
rect 368532 440240 368538 440292
rect 67358 438880 67364 438932
rect 67416 438920 67422 438932
rect 67634 438920 67640 438932
rect 67416 438892 67640 438920
rect 67416 438880 67422 438892
rect 67634 438880 67640 438892
rect 67692 438880 67698 438932
rect 358722 438880 358728 438932
rect 358780 438920 358786 438932
rect 361758 438920 361764 438932
rect 358780 438892 361764 438920
rect 358780 438880 358786 438892
rect 361758 438880 361764 438892
rect 361816 438880 361822 438932
rect 64690 438812 64696 438864
rect 64748 438852 64754 438864
rect 66806 438852 66812 438864
rect 64748 438824 66812 438852
rect 64748 438812 64754 438824
rect 66806 438812 66812 438824
rect 66864 438812 66870 438864
rect 124122 438200 124128 438252
rect 124180 438240 124186 438252
rect 132494 438240 132500 438252
rect 124180 438212 132500 438240
rect 124180 438200 124186 438212
rect 132494 438200 132500 438212
rect 132552 438240 132558 438252
rect 133138 438240 133144 438252
rect 132552 438212 133144 438240
rect 132552 438200 132558 438212
rect 133138 438200 133144 438212
rect 133196 438200 133202 438252
rect 126238 438132 126244 438184
rect 126296 438172 126302 438184
rect 152550 438172 152556 438184
rect 126296 438144 152556 438172
rect 126296 438132 126302 438144
rect 152550 438132 152556 438144
rect 152608 438132 152614 438184
rect 50798 436092 50804 436144
rect 50856 436132 50862 436144
rect 50856 436104 53052 436132
rect 50856 436092 50862 436104
rect 53024 436064 53052 436104
rect 358722 436092 358728 436144
rect 358780 436132 358786 436144
rect 379514 436132 379520 436144
rect 358780 436104 379520 436132
rect 358780 436092 358786 436104
rect 379514 436092 379520 436104
rect 379572 436092 379578 436144
rect 53098 436064 53104 436076
rect 53011 436036 53104 436064
rect 53098 436024 53104 436036
rect 53156 436064 53162 436076
rect 66714 436064 66720 436076
rect 53156 436036 66720 436064
rect 53156 436024 53162 436036
rect 66714 436024 66720 436036
rect 66772 436024 66778 436076
rect 192570 433304 192576 433356
rect 192628 433344 192634 433356
rect 197354 433344 197360 433356
rect 192628 433316 197360 433344
rect 192628 433304 192634 433316
rect 197354 433304 197360 433316
rect 197412 433304 197418 433356
rect 358722 433304 358728 433356
rect 358780 433344 358786 433356
rect 380986 433344 380992 433356
rect 358780 433316 380992 433344
rect 358780 433304 358786 433316
rect 380986 433304 380992 433316
rect 381044 433304 381050 433356
rect 50890 433236 50896 433288
rect 50948 433276 50954 433288
rect 54938 433276 54944 433288
rect 50948 433248 54944 433276
rect 50948 433236 50954 433248
rect 54938 433236 54944 433248
rect 54996 433236 55002 433288
rect 124122 432556 124128 432608
rect 124180 432596 124186 432608
rect 142798 432596 142804 432608
rect 124180 432568 142804 432596
rect 124180 432556 124186 432568
rect 142798 432556 142804 432568
rect 142856 432556 142862 432608
rect 54938 431944 54944 431996
rect 54996 431984 55002 431996
rect 66806 431984 66812 431996
rect 54996 431956 66812 431984
rect 54996 431944 55002 431956
rect 66806 431944 66812 431956
rect 66864 431944 66870 431996
rect 124122 431876 124128 431928
rect 124180 431916 124186 431928
rect 124306 431916 124312 431928
rect 124180 431888 124312 431916
rect 124180 431876 124186 431888
rect 124306 431876 124312 431888
rect 124364 431916 124370 431928
rect 169110 431916 169116 431928
rect 124364 431888 169116 431916
rect 124364 431876 124370 431888
rect 169110 431876 169116 431888
rect 169168 431876 169174 431928
rect 50982 431196 50988 431248
rect 51040 431236 51046 431248
rect 64690 431236 64696 431248
rect 51040 431208 64696 431236
rect 51040 431196 51046 431208
rect 64690 431196 64696 431208
rect 64748 431236 64754 431248
rect 66806 431236 66812 431248
rect 64748 431208 66812 431236
rect 64748 431196 64754 431208
rect 66806 431196 66812 431208
rect 66864 431196 66870 431248
rect 358722 430584 358728 430636
rect 358780 430624 358786 430636
rect 376846 430624 376852 430636
rect 358780 430596 376852 430624
rect 358780 430584 358786 430596
rect 376846 430584 376852 430596
rect 376904 430584 376910 430636
rect 51074 429088 51080 429140
rect 51132 429128 51138 429140
rect 52362 429128 52368 429140
rect 51132 429100 52368 429128
rect 51132 429088 51138 429100
rect 52362 429088 52368 429100
rect 52420 429128 52426 429140
rect 66806 429128 66812 429140
rect 52420 429100 66812 429128
rect 52420 429088 52426 429100
rect 66806 429088 66812 429100
rect 66864 429088 66870 429140
rect 122742 429088 122748 429140
rect 122800 429128 122806 429140
rect 173158 429128 173164 429140
rect 122800 429100 173164 429128
rect 122800 429088 122806 429100
rect 173158 429088 173164 429100
rect 173216 429088 173222 429140
rect 22738 428408 22744 428460
rect 22796 428448 22802 428460
rect 51074 428448 51080 428460
rect 22796 428420 51080 428448
rect 22796 428408 22802 428420
rect 51074 428408 51080 428420
rect 51132 428408 51138 428460
rect 178678 427796 178684 427848
rect 178736 427836 178742 427848
rect 197354 427836 197360 427848
rect 178736 427808 197360 427836
rect 178736 427796 178742 427808
rect 197354 427796 197360 427808
rect 197412 427796 197418 427848
rect 358722 427796 358728 427848
rect 358780 427836 358786 427848
rect 372706 427836 372712 427848
rect 358780 427808 372712 427836
rect 358780 427796 358786 427808
rect 372706 427796 372712 427808
rect 372764 427796 372770 427848
rect 356698 426776 356704 426828
rect 356756 426816 356762 426828
rect 357526 426816 357532 426828
rect 356756 426788 357532 426816
rect 356756 426776 356762 426788
rect 357526 426776 357532 426788
rect 357584 426776 357590 426828
rect 152458 426436 152464 426488
rect 152516 426476 152522 426488
rect 197354 426476 197360 426488
rect 152516 426448 197360 426476
rect 152516 426436 152522 426448
rect 197354 426436 197360 426448
rect 197412 426436 197418 426488
rect 41322 425688 41328 425740
rect 41380 425728 41386 425740
rect 60734 425728 60740 425740
rect 41380 425700 60740 425728
rect 41380 425688 41386 425700
rect 60734 425688 60740 425700
rect 60792 425688 60798 425740
rect 60734 425076 60740 425128
rect 60792 425116 60798 425128
rect 61838 425116 61844 425128
rect 60792 425088 61844 425116
rect 60792 425076 60798 425088
rect 61838 425076 61844 425088
rect 61896 425116 61902 425128
rect 66714 425116 66720 425128
rect 61896 425088 66720 425116
rect 61896 425076 61902 425088
rect 66714 425076 66720 425088
rect 66772 425076 66778 425128
rect 58894 423648 58900 423700
rect 58952 423688 58958 423700
rect 63402 423688 63408 423700
rect 58952 423660 63408 423688
rect 58952 423648 58958 423660
rect 63402 423648 63408 423660
rect 63460 423688 63466 423700
rect 66806 423688 66812 423700
rect 63460 423660 66812 423688
rect 63460 423648 63466 423660
rect 66806 423648 66812 423660
rect 66864 423648 66870 423700
rect 178862 423648 178868 423700
rect 178920 423688 178926 423700
rect 197354 423688 197360 423700
rect 178920 423660 197360 423688
rect 178920 423648 178926 423660
rect 197354 423648 197360 423660
rect 197412 423648 197418 423700
rect 358722 423648 358728 423700
rect 358780 423688 358786 423700
rect 364610 423688 364616 423700
rect 358780 423660 364616 423688
rect 358780 423648 358786 423660
rect 364610 423648 364616 423660
rect 364668 423688 364674 423700
rect 373994 423688 374000 423700
rect 364668 423660 374000 423688
rect 364668 423648 364674 423660
rect 373994 423648 374000 423660
rect 374052 423648 374058 423700
rect 3418 423580 3424 423632
rect 3476 423620 3482 423632
rect 17218 423620 17224 423632
rect 3476 423592 17224 423620
rect 3476 423580 3482 423592
rect 17218 423580 17224 423592
rect 17276 423580 17282 423632
rect 50982 421540 50988 421592
rect 51040 421580 51046 421592
rect 59170 421580 59176 421592
rect 51040 421552 59176 421580
rect 51040 421540 51046 421552
rect 59170 421540 59176 421552
rect 59228 421580 59234 421592
rect 66254 421580 66260 421592
rect 59228 421552 66260 421580
rect 59228 421540 59234 421552
rect 66254 421540 66260 421552
rect 66312 421540 66318 421592
rect 122926 421540 122932 421592
rect 122984 421580 122990 421592
rect 148962 421580 148968 421592
rect 122984 421552 148968 421580
rect 122984 421540 122990 421552
rect 148962 421540 148968 421552
rect 149020 421580 149026 421592
rect 178770 421580 178776 421592
rect 149020 421552 178776 421580
rect 149020 421540 149026 421552
rect 178770 421540 178776 421552
rect 178828 421540 178834 421592
rect 358722 420928 358728 420980
rect 358780 420968 358786 420980
rect 370130 420968 370136 420980
rect 358780 420940 370136 420968
rect 358780 420928 358786 420940
rect 370130 420928 370136 420940
rect 370188 420928 370194 420980
rect 124122 420860 124128 420912
rect 124180 420900 124186 420912
rect 159358 420900 159364 420912
rect 124180 420872 159364 420900
rect 124180 420860 124186 420872
rect 159358 420860 159364 420872
rect 159416 420860 159422 420912
rect 358722 418208 358728 418260
rect 358780 418248 358786 418260
rect 365806 418248 365812 418260
rect 358780 418220 365812 418248
rect 358780 418208 358786 418220
rect 365806 418208 365812 418220
rect 365864 418208 365870 418260
rect 177298 418140 177304 418192
rect 177356 418180 177362 418192
rect 197354 418180 197360 418192
rect 177356 418152 197360 418180
rect 177356 418140 177362 418152
rect 197354 418140 197360 418152
rect 197412 418140 197418 418192
rect 121178 415352 121184 415404
rect 121236 415392 121242 415404
rect 126974 415392 126980 415404
rect 121236 415364 126980 415392
rect 121236 415352 121242 415364
rect 126974 415352 126980 415364
rect 127032 415352 127038 415404
rect 49602 415284 49608 415336
rect 49660 415324 49666 415336
rect 53650 415324 53656 415336
rect 49660 415296 53656 415324
rect 49660 415284 49666 415296
rect 53650 415284 53656 415296
rect 53708 415284 53714 415336
rect 53650 413992 53656 414044
rect 53708 414032 53714 414044
rect 66806 414032 66812 414044
rect 53708 414004 66812 414032
rect 53708 413992 53714 414004
rect 66806 413992 66812 414004
rect 66864 413992 66870 414044
rect 185670 413992 185676 414044
rect 185728 414032 185734 414044
rect 197354 414032 197360 414044
rect 185728 414004 197360 414032
rect 185728 413992 185734 414004
rect 197354 413992 197360 414004
rect 197412 413992 197418 414044
rect 358722 413992 358728 414044
rect 358780 414032 358786 414044
rect 367370 414032 367376 414044
rect 358780 414004 367376 414032
rect 358780 413992 358786 414004
rect 367370 413992 367376 414004
rect 367428 413992 367434 414044
rect 123846 413244 123852 413296
rect 123904 413284 123910 413296
rect 136634 413284 136640 413296
rect 123904 413256 136640 413284
rect 123904 413244 123910 413256
rect 136634 413244 136640 413256
rect 136692 413244 136698 413296
rect 58986 411272 58992 411324
rect 59044 411312 59050 411324
rect 66898 411312 66904 411324
rect 59044 411284 66904 411312
rect 59044 411272 59050 411284
rect 66898 411272 66904 411284
rect 66956 411272 66962 411324
rect 123570 411272 123576 411324
rect 123628 411312 123634 411324
rect 151078 411312 151084 411324
rect 123628 411284 151084 411312
rect 123628 411272 123634 411284
rect 151078 411272 151084 411284
rect 151136 411272 151142 411324
rect 164142 411272 164148 411324
rect 164200 411312 164206 411324
rect 197354 411312 197360 411324
rect 164200 411284 197360 411312
rect 164200 411272 164206 411284
rect 197354 411272 197360 411284
rect 197412 411272 197418 411324
rect 358722 411272 358728 411324
rect 358780 411312 358786 411324
rect 389174 411312 389180 411324
rect 358780 411284 389180 411312
rect 358780 411272 358786 411284
rect 389174 411272 389180 411284
rect 389232 411272 389238 411324
rect 124858 409776 124864 409828
rect 124916 409816 124922 409828
rect 197354 409816 197360 409828
rect 124916 409788 197360 409816
rect 124916 409776 124922 409788
rect 197354 409776 197360 409788
rect 197412 409776 197418 409828
rect 358722 408552 358728 408604
rect 358780 408592 358786 408604
rect 365898 408592 365904 408604
rect 358780 408564 365904 408592
rect 358780 408552 358786 408564
rect 365898 408552 365904 408564
rect 365956 408552 365962 408604
rect 124122 407872 124128 407924
rect 124180 407912 124186 407924
rect 133874 407912 133880 407924
rect 124180 407884 133880 407912
rect 124180 407872 124186 407884
rect 133874 407872 133880 407884
rect 133932 407912 133938 407924
rect 134610 407912 134616 407924
rect 133932 407884 134616 407912
rect 133932 407872 133938 407884
rect 134610 407872 134616 407884
rect 134668 407872 134674 407924
rect 122098 407056 122104 407108
rect 122156 407096 122162 407108
rect 123018 407096 123024 407108
rect 122156 407068 123024 407096
rect 122156 407056 122162 407068
rect 123018 407056 123024 407068
rect 123076 407056 123082 407108
rect 124122 406172 124128 406224
rect 124180 406212 124186 406224
rect 125502 406212 125508 406224
rect 124180 406184 125508 406212
rect 124180 406172 124186 406184
rect 125502 406172 125508 406184
rect 125560 406172 125566 406224
rect 59262 405764 59268 405816
rect 59320 405804 59326 405816
rect 64598 405804 64604 405816
rect 59320 405776 64604 405804
rect 59320 405764 59326 405776
rect 64598 405764 64604 405776
rect 64656 405804 64662 405816
rect 66254 405804 66260 405816
rect 64656 405776 66260 405804
rect 64656 405764 64662 405776
rect 66254 405764 66260 405776
rect 66312 405764 66318 405816
rect 133230 405696 133236 405748
rect 133288 405736 133294 405748
rect 197354 405736 197360 405748
rect 133288 405708 197360 405736
rect 133288 405696 133294 405708
rect 197354 405696 197360 405708
rect 197412 405696 197418 405748
rect 57882 403588 57888 403640
rect 57940 403628 57946 403640
rect 66254 403628 66260 403640
rect 57940 403600 66260 403628
rect 57940 403588 57946 403600
rect 66254 403588 66260 403600
rect 66312 403588 66318 403640
rect 142890 403588 142896 403640
rect 142948 403628 142954 403640
rect 166994 403628 167000 403640
rect 142948 403600 167000 403628
rect 142948 403588 142954 403600
rect 166994 403588 167000 403600
rect 167052 403588 167058 403640
rect 358722 403520 358728 403572
rect 358780 403560 358786 403572
rect 363230 403560 363236 403572
rect 358780 403532 363236 403560
rect 358780 403520 358786 403532
rect 363230 403520 363236 403532
rect 363288 403520 363294 403572
rect 123754 403384 123760 403436
rect 123812 403424 123818 403436
rect 124858 403424 124864 403436
rect 123812 403396 124864 403424
rect 123812 403384 123818 403396
rect 124858 403384 124864 403396
rect 124916 403384 124922 403436
rect 194042 401616 194048 401668
rect 194100 401656 194106 401668
rect 197354 401656 197360 401668
rect 194100 401628 197360 401656
rect 194100 401616 194106 401628
rect 197354 401616 197360 401628
rect 197412 401616 197418 401668
rect 358722 401616 358728 401668
rect 358780 401656 358786 401668
rect 378134 401656 378140 401668
rect 358780 401628 378140 401656
rect 358780 401616 358786 401628
rect 378134 401616 378140 401628
rect 378192 401616 378198 401668
rect 44082 401548 44088 401600
rect 44140 401588 44146 401600
rect 48222 401588 48228 401600
rect 44140 401560 48228 401588
rect 44140 401548 44146 401560
rect 48222 401548 48228 401560
rect 48280 401588 48286 401600
rect 66254 401588 66260 401600
rect 48280 401560 66260 401588
rect 48280 401548 48286 401560
rect 66254 401548 66260 401560
rect 66312 401548 66318 401600
rect 124122 400868 124128 400920
rect 124180 400908 124186 400920
rect 193214 400908 193220 400920
rect 124180 400880 193220 400908
rect 124180 400868 124186 400880
rect 193214 400868 193220 400880
rect 193272 400868 193278 400920
rect 193214 400188 193220 400240
rect 193272 400228 193278 400240
rect 194134 400228 194140 400240
rect 193272 400200 194140 400228
rect 193272 400188 193278 400200
rect 194134 400188 194140 400200
rect 194192 400188 194198 400240
rect 59998 399440 60004 399492
rect 60056 399480 60062 399492
rect 66254 399480 66260 399492
rect 60056 399452 66260 399480
rect 60056 399440 60062 399452
rect 66254 399440 66260 399452
rect 66312 399440 66318 399492
rect 124122 399440 124128 399492
rect 124180 399480 124186 399492
rect 189902 399480 189908 399492
rect 124180 399452 189908 399480
rect 124180 399440 124186 399452
rect 189902 399440 189908 399452
rect 189960 399440 189966 399492
rect 187050 398828 187056 398880
rect 187108 398868 187114 398880
rect 197354 398868 197360 398880
rect 187108 398840 197360 398868
rect 187108 398828 187114 398840
rect 197354 398828 197360 398840
rect 197412 398828 197418 398880
rect 357986 398828 357992 398880
rect 358044 398868 358050 398880
rect 360470 398868 360476 398880
rect 358044 398840 360476 398868
rect 358044 398828 358050 398840
rect 360470 398828 360476 398840
rect 360528 398828 360534 398880
rect 2774 398692 2780 398744
rect 2832 398732 2838 398744
rect 4798 398732 4804 398744
rect 2832 398704 4804 398732
rect 2832 398692 2838 398704
rect 4798 398692 4804 398704
rect 4856 398692 4862 398744
rect 48222 398080 48228 398132
rect 48280 398120 48286 398132
rect 55122 398120 55128 398132
rect 48280 398092 55128 398120
rect 48280 398080 48286 398092
rect 55122 398080 55128 398092
rect 55180 398120 55186 398132
rect 59998 398120 60004 398132
rect 55180 398092 60004 398120
rect 55180 398080 55186 398092
rect 59998 398080 60004 398092
rect 60056 398080 60062 398132
rect 130470 397468 130476 397520
rect 130528 397508 130534 397520
rect 187050 397508 187056 397520
rect 130528 397480 187056 397508
rect 130528 397468 130534 397480
rect 187050 397468 187056 397480
rect 187108 397468 187114 397520
rect 37182 396720 37188 396772
rect 37240 396760 37246 396772
rect 66990 396760 66996 396772
rect 37240 396732 66996 396760
rect 37240 396720 37246 396732
rect 66990 396720 66996 396732
rect 67048 396760 67054 396772
rect 67266 396760 67272 396772
rect 67048 396732 67272 396760
rect 67048 396720 67054 396732
rect 67266 396720 67272 396732
rect 67324 396720 67330 396772
rect 133138 396720 133144 396772
rect 133196 396760 133202 396772
rect 171134 396760 171140 396772
rect 133196 396732 171140 396760
rect 133196 396720 133202 396732
rect 171134 396720 171140 396732
rect 171192 396720 171198 396772
rect 169662 396040 169668 396092
rect 169720 396080 169726 396092
rect 197354 396080 197360 396092
rect 169720 396052 197360 396080
rect 169720 396040 169726 396052
rect 197354 396040 197360 396052
rect 197412 396040 197418 396092
rect 358722 396040 358728 396092
rect 358780 396080 358786 396092
rect 361850 396080 361856 396092
rect 358780 396052 361856 396080
rect 358780 396040 358786 396052
rect 361850 396040 361856 396052
rect 361908 396040 361914 396092
rect 124122 395292 124128 395344
rect 124180 395332 124186 395344
rect 188522 395332 188528 395344
rect 124180 395304 188528 395332
rect 124180 395292 124186 395304
rect 188522 395292 188528 395304
rect 188580 395292 188586 395344
rect 191650 394680 191656 394732
rect 191708 394720 191714 394732
rect 197354 394720 197360 394732
rect 191708 394692 197360 394720
rect 191708 394680 191714 394692
rect 197354 394680 197360 394692
rect 197412 394680 197418 394732
rect 134518 393320 134524 393372
rect 134576 393360 134582 393372
rect 198458 393360 198464 393372
rect 134576 393332 198464 393360
rect 134576 393320 134582 393332
rect 198458 393320 198464 393332
rect 198516 393320 198522 393372
rect 61930 392028 61936 392080
rect 61988 392068 61994 392080
rect 66162 392068 66168 392080
rect 61988 392040 66168 392068
rect 61988 392028 61994 392040
rect 66162 392028 66168 392040
rect 66220 392068 66226 392080
rect 66622 392068 66628 392080
rect 66220 392040 66628 392068
rect 66220 392028 66226 392040
rect 66622 392028 66628 392040
rect 66680 392028 66686 392080
rect 121454 392028 121460 392080
rect 121512 392068 121518 392080
rect 153194 392068 153200 392080
rect 121512 392040 153200 392068
rect 121512 392028 121518 392040
rect 153194 392028 153200 392040
rect 153252 392028 153258 392080
rect 140130 391960 140136 392012
rect 140188 392000 140194 392012
rect 197354 392000 197360 392012
rect 140188 391972 197360 392000
rect 140188 391960 140194 391972
rect 197354 391960 197360 391972
rect 197412 391960 197418 392012
rect 3418 391212 3424 391264
rect 3476 391252 3482 391264
rect 140038 391252 140044 391264
rect 3476 391224 64874 391252
rect 3476 391212 3482 391224
rect 64846 391048 64874 391224
rect 93826 391224 140044 391252
rect 81434 391048 81440 391060
rect 64846 391020 81440 391048
rect 81434 391008 81440 391020
rect 81492 391008 81498 391060
rect 85850 391008 85856 391060
rect 85908 391048 85914 391060
rect 93826 391048 93854 391224
rect 140038 391212 140044 391224
rect 140096 391212 140102 391264
rect 157978 391212 157984 391264
rect 158036 391252 158042 391264
rect 175274 391252 175280 391264
rect 158036 391224 175280 391252
rect 158036 391212 158042 391224
rect 175274 391212 175280 391224
rect 175332 391212 175338 391264
rect 85908 391020 93854 391048
rect 85908 391008 85914 391020
rect 120442 390260 120448 390312
rect 120500 390300 120506 390312
rect 120810 390300 120816 390312
rect 120500 390272 120816 390300
rect 120500 390260 120506 390272
rect 120810 390260 120816 390272
rect 120868 390260 120874 390312
rect 113082 389784 113088 389836
rect 113140 389824 113146 389836
rect 120718 389824 120724 389836
rect 113140 389796 120724 389824
rect 113140 389784 113146 389796
rect 120718 389784 120724 389796
rect 120776 389784 120782 389836
rect 57698 389240 57704 389292
rect 57756 389280 57762 389292
rect 85574 389280 85580 389292
rect 57756 389252 85580 389280
rect 57756 389240 57762 389252
rect 85574 389240 85580 389252
rect 85632 389240 85638 389292
rect 25498 389172 25504 389224
rect 25556 389212 25562 389224
rect 110414 389212 110420 389224
rect 25556 389184 110420 389212
rect 25556 389172 25562 389184
rect 110414 389172 110420 389184
rect 110472 389212 110478 389224
rect 111426 389212 111432 389224
rect 110472 389184 111432 389212
rect 110472 389172 110478 389184
rect 111426 389172 111432 389184
rect 111484 389172 111490 389224
rect 43990 389104 43996 389156
rect 44048 389144 44054 389156
rect 44048 389116 64874 389144
rect 44048 389104 44054 389116
rect 64846 389076 64874 389116
rect 70302 389104 70308 389156
rect 70360 389144 70366 389156
rect 76650 389144 76656 389156
rect 70360 389116 76656 389144
rect 70360 389104 70366 389116
rect 76650 389104 76656 389116
rect 76708 389104 76714 389156
rect 91646 389104 91652 389156
rect 91704 389144 91710 389156
rect 93210 389144 93216 389156
rect 91704 389116 93216 389144
rect 91704 389104 91710 389116
rect 93210 389104 93216 389116
rect 93268 389104 93274 389156
rect 96246 389104 96252 389156
rect 96304 389144 96310 389156
rect 130470 389144 130476 389156
rect 96304 389116 130476 389144
rect 96304 389104 96310 389116
rect 130470 389104 130476 389116
rect 130528 389104 130534 389156
rect 76374 389076 76380 389088
rect 64846 389048 76380 389076
rect 76374 389036 76380 389048
rect 76432 389036 76438 389088
rect 79502 388492 79508 388544
rect 79560 388532 79566 388544
rect 86218 388532 86224 388544
rect 79560 388504 86224 388532
rect 79560 388492 79566 388504
rect 86218 388492 86224 388504
rect 86276 388492 86282 388544
rect 77846 388424 77852 388476
rect 77904 388464 77910 388476
rect 171778 388464 171784 388476
rect 77904 388436 171784 388464
rect 77904 388424 77910 388436
rect 171778 388424 171784 388436
rect 171836 388464 171842 388476
rect 191098 388464 191104 388476
rect 171836 388436 191104 388464
rect 171836 388424 171842 388436
rect 191098 388424 191104 388436
rect 191156 388424 191162 388476
rect 88518 387812 88524 387864
rect 88576 387852 88582 387864
rect 90358 387852 90364 387864
rect 88576 387824 90364 387852
rect 88576 387812 88582 387824
rect 90358 387812 90364 387824
rect 90416 387812 90422 387864
rect 57790 387744 57796 387796
rect 57848 387784 57854 387796
rect 82078 387784 82084 387796
rect 57848 387756 82084 387784
rect 57848 387744 57854 387756
rect 82078 387744 82084 387756
rect 82136 387744 82142 387796
rect 104158 387744 104164 387796
rect 104216 387784 104222 387796
rect 128354 387784 128360 387796
rect 104216 387756 128360 387784
rect 104216 387744 104222 387756
rect 128354 387744 128360 387756
rect 128412 387744 128418 387796
rect 11698 387064 11704 387116
rect 11756 387104 11762 387116
rect 123662 387104 123668 387116
rect 11756 387076 123668 387104
rect 11756 387064 11762 387076
rect 123662 387064 123668 387076
rect 123720 387104 123726 387116
rect 185762 387104 185768 387116
rect 123720 387076 185768 387104
rect 123720 387064 123726 387076
rect 185762 387064 185768 387076
rect 185820 387064 185826 387116
rect 187234 386384 187240 386436
rect 187292 386424 187298 386436
rect 197354 386424 197360 386436
rect 187292 386396 197360 386424
rect 187292 386384 187298 386396
rect 197354 386384 197360 386396
rect 197412 386384 197418 386436
rect 60458 386316 60464 386368
rect 60516 386356 60522 386368
rect 86954 386356 86960 386368
rect 60516 386328 86960 386356
rect 60516 386316 60522 386328
rect 86954 386316 86960 386328
rect 87012 386316 87018 386368
rect 3418 385636 3424 385688
rect 3476 385676 3482 385688
rect 95234 385676 95240 385688
rect 3476 385648 95240 385676
rect 3476 385636 3482 385648
rect 95234 385636 95240 385648
rect 95292 385636 95298 385688
rect 107194 385636 107200 385688
rect 107252 385676 107258 385688
rect 167086 385676 167092 385688
rect 107252 385648 167092 385676
rect 107252 385636 107258 385648
rect 167086 385636 167092 385648
rect 167144 385636 167150 385688
rect 171042 385636 171048 385688
rect 171100 385676 171106 385688
rect 191098 385676 191104 385688
rect 171100 385648 191104 385676
rect 171100 385636 171106 385648
rect 191098 385636 191104 385648
rect 191156 385636 191162 385688
rect 117590 384276 117596 384328
rect 117648 384316 117654 384328
rect 196618 384316 196624 384328
rect 117648 384288 196624 384316
rect 117648 384276 117654 384288
rect 196618 384276 196624 384288
rect 196676 384276 196682 384328
rect 111794 383664 111800 383716
rect 111852 383704 111858 383716
rect 113082 383704 113088 383716
rect 111852 383676 113088 383704
rect 111852 383664 111858 383676
rect 113082 383664 113088 383676
rect 113140 383704 113146 383716
rect 184290 383704 184296 383716
rect 113140 383676 184296 383704
rect 113140 383664 113146 383676
rect 184290 383664 184296 383676
rect 184348 383664 184354 383716
rect 65978 383596 65984 383648
rect 66036 383636 66042 383648
rect 82814 383636 82820 383648
rect 66036 383608 82820 383636
rect 66036 383596 66042 383608
rect 82814 383596 82820 383608
rect 82872 383596 82878 383648
rect 61838 382916 61844 382968
rect 61896 382956 61902 382968
rect 165614 382956 165620 382968
rect 61896 382928 165620 382956
rect 61896 382916 61902 382928
rect 165614 382916 165620 382928
rect 165672 382916 165678 382968
rect 123478 382236 123484 382288
rect 123536 382276 123542 382288
rect 192662 382276 192668 382288
rect 123536 382248 192668 382276
rect 123536 382236 123542 382248
rect 192662 382236 192668 382248
rect 192720 382236 192726 382288
rect 79962 381488 79968 381540
rect 80020 381528 80026 381540
rect 169846 381528 169852 381540
rect 80020 381500 169852 381528
rect 80020 381488 80026 381500
rect 169846 381488 169852 381500
rect 169904 381488 169910 381540
rect 50890 380876 50896 380928
rect 50948 380916 50954 380928
rect 173158 380916 173164 380928
rect 50948 380888 173164 380916
rect 50948 380876 50954 380888
rect 173158 380876 173164 380888
rect 173216 380876 173222 380928
rect 59078 380808 59084 380860
rect 59136 380848 59142 380860
rect 74534 380848 74540 380860
rect 59136 380820 74540 380848
rect 59136 380808 59142 380820
rect 74534 380808 74540 380820
rect 74592 380808 74598 380860
rect 49602 380128 49608 380180
rect 49660 380168 49666 380180
rect 59078 380168 59084 380180
rect 49660 380140 59084 380168
rect 49660 380128 49666 380140
rect 59078 380128 59084 380140
rect 59136 380128 59142 380180
rect 73154 380128 73160 380180
rect 73212 380168 73218 380180
rect 140130 380168 140136 380180
rect 73212 380140 140136 380168
rect 73212 380128 73218 380140
rect 140130 380128 140136 380140
rect 140188 380128 140194 380180
rect 188522 379516 188528 379568
rect 188580 379556 188586 379568
rect 189810 379556 189816 379568
rect 188580 379528 189816 379556
rect 188580 379516 188586 379528
rect 189810 379516 189816 379528
rect 189868 379556 189874 379568
rect 197354 379556 197360 379568
rect 189868 379528 197360 379556
rect 189868 379516 189874 379528
rect 197354 379516 197360 379528
rect 197412 379516 197418 379568
rect 357894 379516 357900 379568
rect 357952 379556 357958 379568
rect 382274 379556 382280 379568
rect 357952 379528 382280 379556
rect 357952 379516 357958 379528
rect 382274 379516 382280 379528
rect 382332 379516 382338 379568
rect 101398 378768 101404 378820
rect 101456 378808 101462 378820
rect 152550 378808 152556 378820
rect 101456 378780 152556 378808
rect 101456 378768 101462 378780
rect 152550 378768 152556 378780
rect 152608 378768 152614 378820
rect 67266 378156 67272 378208
rect 67324 378196 67330 378208
rect 195238 378196 195244 378208
rect 67324 378168 195244 378196
rect 67324 378156 67330 378168
rect 195238 378156 195244 378168
rect 195296 378156 195302 378208
rect 358354 378088 358360 378140
rect 358412 378128 358418 378140
rect 360378 378128 360384 378140
rect 358412 378100 360384 378128
rect 358412 378088 358418 378100
rect 360378 378088 360384 378100
rect 360436 378088 360442 378140
rect 361482 377952 361488 378004
rect 361540 377992 361546 378004
rect 364518 377992 364524 378004
rect 361540 377964 364524 377992
rect 361540 377952 361546 377964
rect 364518 377952 364524 377964
rect 364576 377952 364582 378004
rect 355318 377544 355324 377596
rect 355376 377584 355382 377596
rect 356238 377584 356244 377596
rect 355376 377556 356244 377584
rect 355376 377544 355382 377556
rect 356238 377544 356244 377556
rect 356296 377544 356302 377596
rect 197078 377476 197084 377528
rect 197136 377516 197142 377528
rect 201586 377516 201592 377528
rect 197136 377488 201592 377516
rect 197136 377476 197142 377488
rect 201586 377476 201592 377488
rect 201644 377476 201650 377528
rect 140682 376796 140688 376848
rect 140740 376836 140746 376848
rect 198734 376836 198740 376848
rect 140740 376808 198740 376836
rect 140740 376796 140746 376808
rect 198734 376796 198740 376808
rect 198792 376836 198798 376848
rect 199102 376836 199108 376848
rect 198792 376808 199108 376836
rect 198792 376796 198798 376808
rect 199102 376796 199108 376808
rect 199160 376796 199166 376848
rect 72418 376728 72424 376780
rect 72476 376768 72482 376780
rect 73062 376768 73068 376780
rect 72476 376740 73068 376768
rect 72476 376728 72482 376740
rect 73062 376728 73068 376740
rect 73120 376768 73126 376780
rect 187050 376768 187056 376780
rect 73120 376740 187056 376768
rect 73120 376728 73126 376740
rect 187050 376728 187056 376740
rect 187108 376728 187114 376780
rect 189902 376660 189908 376712
rect 189960 376700 189966 376712
rect 218054 376700 218060 376712
rect 189960 376672 218060 376700
rect 189960 376660 189966 376672
rect 218054 376660 218060 376672
rect 218112 376700 218118 376712
rect 218238 376700 218244 376712
rect 218112 376672 218244 376700
rect 218112 376660 218118 376672
rect 218238 376660 218244 376672
rect 218296 376660 218302 376712
rect 92382 376048 92388 376100
rect 92440 376088 92446 376100
rect 115658 376088 115664 376100
rect 92440 376060 115664 376088
rect 92440 376048 92446 376060
rect 115658 376048 115664 376060
rect 115716 376048 115722 376100
rect 352650 376048 352656 376100
rect 352708 376088 352714 376100
rect 358814 376088 358820 376100
rect 352708 376060 358820 376088
rect 352708 376048 352714 376060
rect 358814 376048 358820 376060
rect 358872 376048 358878 376100
rect 48222 375980 48228 376032
rect 48280 376020 48286 376032
rect 184382 376020 184388 376032
rect 48280 375992 184388 376020
rect 48280 375980 48286 375992
rect 184382 375980 184388 375992
rect 184440 375980 184446 376032
rect 198734 375980 198740 376032
rect 198792 376020 198798 376032
rect 242158 376020 242164 376032
rect 198792 375992 242164 376020
rect 198792 375980 198798 375992
rect 242158 375980 242164 375992
rect 242216 375980 242222 376032
rect 353938 375980 353944 376032
rect 353996 376020 354002 376032
rect 363230 376020 363236 376032
rect 353996 375992 363236 376020
rect 353996 375980 354002 375992
rect 363230 375980 363236 375992
rect 363288 375980 363294 376032
rect 50982 375300 50988 375352
rect 51040 375340 51046 375352
rect 202230 375340 202236 375352
rect 51040 375312 202236 375340
rect 51040 375300 51046 375312
rect 202230 375300 202236 375312
rect 202288 375300 202294 375352
rect 203518 375300 203524 375352
rect 203576 375340 203582 375352
rect 204990 375340 204996 375352
rect 203576 375312 204996 375340
rect 203576 375300 203582 375312
rect 204990 375300 204996 375312
rect 205048 375300 205054 375352
rect 236638 375300 236644 375352
rect 236696 375340 236702 375352
rect 238110 375340 238116 375352
rect 236696 375312 238116 375340
rect 236696 375300 236702 375312
rect 238110 375300 238116 375312
rect 238168 375300 238174 375352
rect 260098 375300 260104 375352
rect 260156 375340 260162 375352
rect 261478 375340 261484 375352
rect 260156 375312 261484 375340
rect 260156 375300 260162 375312
rect 261478 375300 261484 375312
rect 261536 375300 261542 375352
rect 262490 375300 262496 375352
rect 262548 375340 262554 375352
rect 273070 375340 273076 375352
rect 262548 375312 273076 375340
rect 262548 375300 262554 375312
rect 273070 375300 273076 375312
rect 273128 375300 273134 375352
rect 273990 375300 273996 375352
rect 274048 375340 274054 375352
rect 274726 375340 274732 375352
rect 274048 375312 274732 375340
rect 274048 375300 274054 375312
rect 274726 375300 274732 375312
rect 274784 375300 274790 375352
rect 278038 375300 278044 375352
rect 278096 375340 278102 375352
rect 279694 375340 279700 375352
rect 278096 375312 279700 375340
rect 278096 375300 278102 375312
rect 279694 375300 279700 375312
rect 279752 375300 279758 375352
rect 320174 375300 320180 375352
rect 320232 375340 320238 375352
rect 321278 375340 321284 375352
rect 320232 375312 321284 375340
rect 320232 375300 320238 375312
rect 321278 375300 321284 375312
rect 321336 375300 321342 375352
rect 339494 375300 339500 375352
rect 339552 375340 339558 375352
rect 342346 375340 342352 375352
rect 339552 375312 342352 375340
rect 339552 375300 339558 375312
rect 342346 375300 342352 375312
rect 342404 375300 342410 375352
rect 344462 375300 344468 375352
rect 344520 375340 344526 375352
rect 582374 375340 582380 375352
rect 344520 375312 582380 375340
rect 344520 375300 344526 375312
rect 582374 375300 582380 375312
rect 582432 375300 582438 375352
rect 194594 375232 194600 375284
rect 194652 375272 194658 375284
rect 196802 375272 196808 375284
rect 194652 375244 196808 375272
rect 194652 375232 194658 375244
rect 196802 375232 196808 375244
rect 196860 375232 196866 375284
rect 233878 375232 233884 375284
rect 233936 375272 233942 375284
rect 236454 375272 236460 375284
rect 233936 375244 236460 375272
rect 233936 375232 233942 375244
rect 236454 375232 236460 375244
rect 236512 375232 236518 375284
rect 348418 375232 348424 375284
rect 348476 375272 348482 375284
rect 352742 375272 352748 375284
rect 348476 375244 352748 375272
rect 348476 375232 348482 375244
rect 352742 375232 352748 375244
rect 352800 375232 352806 375284
rect 50798 375096 50804 375148
rect 50856 375136 50862 375148
rect 50982 375136 50988 375148
rect 50856 375108 50988 375136
rect 50856 375096 50862 375108
rect 50982 375096 50988 375108
rect 51040 375096 51046 375148
rect 304258 374824 304264 374876
rect 304316 374864 304322 374876
rect 306190 374864 306196 374876
rect 304316 374836 306196 374864
rect 304316 374824 304322 374836
rect 306190 374824 306196 374836
rect 306248 374824 306254 374876
rect 327718 374824 327724 374876
rect 327776 374864 327782 374876
rect 331214 374864 331220 374876
rect 327776 374836 331220 374864
rect 327776 374824 327782 374836
rect 331214 374824 331220 374836
rect 331272 374824 331278 374876
rect 198918 374620 198924 374672
rect 198976 374660 198982 374672
rect 204346 374660 204352 374672
rect 198976 374632 204352 374660
rect 198976 374620 198982 374632
rect 204346 374620 204352 374632
rect 204404 374620 204410 374672
rect 246390 374620 246396 374672
rect 246448 374660 246454 374672
rect 253198 374660 253204 374672
rect 246448 374632 253204 374660
rect 246448 374620 246454 374632
rect 253198 374620 253204 374632
rect 253256 374620 253262 374672
rect 258718 374620 258724 374672
rect 258776 374660 258782 374672
rect 281350 374660 281356 374672
rect 258776 374632 281356 374660
rect 258776 374620 258782 374632
rect 281350 374620 281356 374632
rect 281408 374620 281414 374672
rect 282178 374620 282184 374672
rect 282236 374660 282242 374672
rect 296254 374660 296260 374672
rect 282236 374632 296260 374660
rect 282236 374620 282242 374632
rect 296254 374620 296260 374632
rect 296312 374620 296318 374672
rect 309870 374620 309876 374672
rect 309928 374660 309934 374672
rect 327902 374660 327908 374672
rect 309928 374632 327908 374660
rect 309928 374620 309934 374632
rect 327902 374620 327908 374632
rect 327960 374620 327966 374672
rect 198734 374280 198740 374332
rect 198792 374320 198798 374332
rect 200022 374320 200028 374332
rect 198792 374292 200028 374320
rect 198792 374280 198798 374292
rect 200022 374280 200028 374292
rect 200080 374280 200086 374332
rect 206462 374280 206468 374332
rect 206520 374320 206526 374332
rect 208302 374320 208308 374332
rect 206520 374292 208308 374320
rect 206520 374280 206526 374292
rect 208302 374280 208308 374292
rect 208360 374280 208366 374332
rect 119982 374008 119988 374060
rect 120040 374048 120046 374060
rect 195330 374048 195336 374060
rect 120040 374020 195336 374048
rect 120040 374008 120046 374020
rect 195330 374008 195336 374020
rect 195388 374008 195394 374060
rect 226978 374008 226984 374060
rect 227036 374048 227042 374060
rect 229830 374048 229836 374060
rect 227036 374020 229836 374048
rect 227036 374008 227042 374020
rect 229830 374008 229836 374020
rect 229888 374008 229894 374060
rect 250438 374008 250444 374060
rect 250496 374048 250502 374060
rect 255958 374048 255964 374060
rect 250496 374020 255964 374048
rect 250496 374008 250502 374020
rect 255958 374008 255964 374020
rect 256016 374008 256022 374060
rect 276658 374008 276664 374060
rect 276716 374048 276722 374060
rect 277670 374048 277676 374060
rect 276716 374020 277676 374048
rect 276716 374008 276722 374020
rect 277670 374008 277676 374020
rect 277728 374008 277734 374060
rect 294598 374008 294604 374060
rect 294656 374048 294662 374060
rect 297910 374048 297916 374060
rect 294656 374020 297916 374048
rect 294656 374008 294662 374020
rect 297910 374008 297916 374020
rect 297968 374008 297974 374060
rect 308398 374008 308404 374060
rect 308456 374048 308462 374060
rect 313918 374048 313924 374060
rect 308456 374020 313924 374048
rect 308456 374008 308462 374020
rect 313918 374008 313924 374020
rect 313976 374008 313982 374060
rect 354030 374008 354036 374060
rect 354088 374048 354094 374060
rect 356054 374048 356060 374060
rect 354088 374020 356060 374048
rect 354088 374008 354094 374020
rect 356054 374008 356060 374020
rect 356112 374008 356118 374060
rect 199010 373328 199016 373380
rect 199068 373368 199074 373380
rect 207014 373368 207020 373380
rect 199068 373340 207020 373368
rect 199068 373328 199074 373340
rect 207014 373328 207020 373340
rect 207072 373328 207078 373380
rect 355410 373328 355416 373380
rect 355468 373368 355474 373380
rect 364426 373368 364432 373380
rect 355468 373340 364432 373368
rect 355468 373328 355474 373340
rect 364426 373328 364432 373340
rect 364484 373328 364490 373380
rect 101398 373260 101404 373312
rect 101456 373300 101462 373312
rect 133230 373300 133236 373312
rect 101456 373272 133236 373300
rect 101456 373260 101462 373272
rect 133230 373260 133236 373272
rect 133288 373260 133294 373312
rect 184290 373260 184296 373312
rect 184348 373300 184354 373312
rect 251818 373300 251824 373312
rect 184348 373272 251824 373300
rect 184348 373260 184354 373272
rect 251818 373260 251824 373272
rect 251876 373260 251882 373312
rect 286318 373260 286324 373312
rect 286376 373300 286382 373312
rect 293954 373300 293960 373312
rect 286376 373272 293960 373300
rect 286376 373260 286382 373272
rect 293954 373260 293960 373272
rect 294012 373260 294018 373312
rect 340138 373260 340144 373312
rect 340196 373300 340202 373312
rect 357618 373300 357624 373312
rect 340196 373272 357624 373300
rect 340196 373260 340202 373272
rect 357618 373260 357624 373272
rect 357676 373260 357682 373312
rect 136818 372648 136824 372700
rect 136876 372688 136882 372700
rect 175918 372688 175924 372700
rect 136876 372660 175924 372688
rect 136876 372648 136882 372660
rect 175918 372648 175924 372660
rect 175976 372648 175982 372700
rect 67542 372580 67548 372632
rect 67600 372620 67606 372632
rect 191190 372620 191196 372632
rect 67600 372592 191196 372620
rect 67600 372580 67606 372592
rect 191190 372580 191196 372592
rect 191248 372580 191254 372632
rect 334618 372580 334624 372632
rect 334676 372620 334682 372632
rect 336734 372620 336740 372632
rect 334676 372592 336740 372620
rect 334676 372580 334682 372592
rect 336734 372580 336740 372592
rect 336792 372580 336798 372632
rect 180242 372512 180248 372564
rect 180300 372552 180306 372564
rect 197262 372552 197268 372564
rect 180300 372524 197268 372552
rect 180300 372512 180306 372524
rect 197262 372512 197268 372524
rect 197320 372552 197326 372564
rect 582926 372552 582932 372564
rect 197320 372524 582932 372552
rect 197320 372512 197326 372524
rect 582926 372512 582932 372524
rect 582984 372512 582990 372564
rect 56410 371832 56416 371884
rect 56468 371872 56474 371884
rect 76558 371872 76564 371884
rect 56468 371844 76564 371872
rect 56468 371832 56474 371844
rect 76558 371832 76564 371844
rect 76616 371832 76622 371884
rect 341518 371832 341524 371884
rect 341576 371872 341582 371884
rect 357526 371872 357532 371884
rect 341576 371844 357532 371872
rect 341576 371832 341582 371844
rect 357526 371832 357532 371844
rect 357584 371832 357590 371884
rect 358078 371832 358084 371884
rect 358136 371872 358142 371884
rect 365898 371872 365904 371884
rect 358136 371844 365904 371872
rect 358136 371832 358142 371844
rect 365898 371832 365904 371844
rect 365956 371832 365962 371884
rect 66898 371220 66904 371272
rect 66956 371260 66962 371272
rect 67358 371260 67364 371272
rect 66956 371232 67364 371260
rect 66956 371220 66962 371232
rect 67358 371220 67364 371232
rect 67416 371260 67422 371272
rect 213178 371260 213184 371272
rect 67416 371232 213184 371260
rect 67416 371220 67422 371232
rect 213178 371220 213184 371232
rect 213236 371220 213242 371272
rect 195330 371152 195336 371204
rect 195388 371192 195394 371204
rect 234614 371192 234620 371204
rect 195388 371164 234620 371192
rect 195388 371152 195394 371164
rect 234614 371152 234620 371164
rect 234672 371152 234678 371204
rect 267642 370540 267648 370592
rect 267700 370580 267706 370592
rect 357710 370580 357716 370592
rect 267700 370552 357716 370580
rect 267700 370540 267706 370552
rect 357710 370540 357716 370552
rect 357768 370540 357774 370592
rect 84838 370472 84844 370524
rect 84896 370512 84902 370524
rect 120718 370512 120724 370524
rect 84896 370484 120724 370512
rect 84896 370472 84902 370484
rect 120718 370472 120724 370484
rect 120776 370472 120782 370524
rect 124858 370472 124864 370524
rect 124916 370512 124922 370524
rect 162762 370512 162768 370524
rect 124916 370484 162768 370512
rect 124916 370472 124922 370484
rect 162762 370472 162768 370484
rect 162820 370512 162826 370524
rect 387794 370512 387800 370524
rect 162820 370484 387800 370512
rect 162820 370472 162826 370484
rect 387794 370472 387800 370484
rect 387852 370472 387858 370524
rect 234614 369860 234620 369912
rect 234672 369900 234678 369912
rect 235258 369900 235264 369912
rect 234672 369872 235264 369900
rect 234672 369860 234678 369872
rect 235258 369860 235264 369872
rect 235316 369860 235322 369912
rect 345658 369180 345664 369232
rect 345716 369220 345722 369232
rect 361666 369220 361672 369232
rect 345716 369192 361672 369220
rect 345716 369180 345722 369192
rect 361666 369180 361672 369192
rect 361724 369180 361730 369232
rect 56502 369112 56508 369164
rect 56560 369152 56566 369164
rect 144270 369152 144276 369164
rect 56560 369124 144276 369152
rect 56560 369112 56566 369124
rect 144270 369112 144276 369124
rect 144328 369112 144334 369164
rect 190362 369112 190368 369164
rect 190420 369152 190426 369164
rect 211798 369152 211804 369164
rect 190420 369124 211804 369152
rect 190420 369112 190426 369124
rect 211798 369112 211804 369124
rect 211856 369112 211862 369164
rect 347038 369112 347044 369164
rect 347096 369152 347102 369164
rect 365806 369152 365812 369164
rect 347096 369124 365812 369152
rect 347096 369112 347102 369124
rect 365806 369112 365812 369124
rect 365864 369112 365870 369164
rect 134610 368908 134616 368960
rect 134668 368948 134674 368960
rect 135162 368948 135168 368960
rect 134668 368920 135168 368948
rect 134668 368908 134674 368920
rect 135162 368908 135168 368920
rect 135220 368908 135226 368960
rect 147674 368568 147680 368620
rect 147732 368608 147738 368620
rect 148318 368608 148324 368620
rect 147732 368580 148324 368608
rect 147732 368568 147738 368580
rect 148318 368568 148324 368580
rect 148376 368608 148382 368620
rect 184290 368608 184296 368620
rect 148376 368580 184296 368608
rect 148376 368568 148382 368580
rect 184290 368568 184296 368580
rect 184348 368568 184354 368620
rect 135162 368500 135168 368552
rect 135220 368540 135226 368552
rect 195238 368540 195244 368552
rect 135220 368512 195244 368540
rect 135220 368500 135226 368512
rect 195238 368500 195244 368512
rect 195296 368500 195302 368552
rect 125410 368432 125416 368484
rect 125468 368472 125474 368484
rect 127710 368472 127716 368484
rect 125468 368444 127716 368472
rect 125468 368432 125474 368444
rect 127710 368432 127716 368444
rect 127768 368432 127774 368484
rect 86218 367820 86224 367872
rect 86276 367860 86282 367872
rect 124766 367860 124772 367872
rect 86276 367832 124772 367860
rect 86276 367820 86282 367832
rect 124766 367820 124772 367832
rect 124824 367820 124830 367872
rect 67726 367752 67732 367804
rect 67784 367792 67790 367804
rect 124858 367792 124864 367804
rect 67784 367764 124864 367792
rect 67784 367752 67790 367764
rect 124858 367752 124864 367764
rect 124916 367752 124922 367804
rect 144822 367752 144828 367804
rect 144880 367792 144886 367804
rect 202874 367792 202880 367804
rect 144880 367764 202880 367792
rect 144880 367752 144886 367764
rect 202874 367752 202880 367764
rect 202932 367792 202938 367804
rect 209130 367792 209136 367804
rect 202932 367764 209136 367792
rect 202932 367752 202938 367764
rect 209130 367752 209136 367764
rect 209188 367752 209194 367804
rect 242250 367752 242256 367804
rect 242308 367792 242314 367804
rect 359090 367792 359096 367804
rect 242308 367764 359096 367792
rect 242308 367752 242314 367764
rect 359090 367752 359096 367764
rect 359148 367752 359154 367804
rect 124214 367072 124220 367124
rect 124272 367112 124278 367124
rect 124766 367112 124772 367124
rect 124272 367084 124772 367112
rect 124272 367072 124278 367084
rect 124766 367072 124772 367084
rect 124824 367112 124830 367124
rect 196618 367112 196624 367124
rect 124824 367084 196624 367112
rect 124824 367072 124830 367084
rect 196618 367072 196624 367084
rect 196676 367072 196682 367124
rect 71682 366936 71688 366988
rect 71740 366976 71746 366988
rect 73798 366976 73804 366988
rect 71740 366948 73804 366976
rect 71740 366936 71746 366948
rect 73798 366936 73804 366948
rect 73856 366936 73862 366988
rect 231854 366800 231860 366852
rect 231912 366840 231918 366852
rect 232590 366840 232596 366852
rect 231912 366812 232596 366840
rect 231912 366800 231918 366812
rect 232590 366800 232596 366812
rect 232648 366800 232654 366852
rect 77938 366392 77944 366444
rect 77996 366432 78002 366444
rect 130378 366432 130384 366444
rect 77996 366404 130384 366432
rect 77996 366392 78002 366404
rect 130378 366392 130384 366404
rect 130436 366392 130442 366444
rect 331950 366392 331956 366444
rect 332008 366432 332014 366444
rect 360286 366432 360292 366444
rect 332008 366404 360292 366432
rect 332008 366392 332014 366404
rect 360286 366392 360292 366404
rect 360344 366392 360350 366444
rect 99006 366324 99012 366376
rect 99064 366364 99070 366376
rect 157426 366364 157432 366376
rect 99064 366336 157432 366364
rect 99064 366324 99070 366336
rect 157426 366324 157432 366336
rect 157484 366324 157490 366376
rect 159358 366324 159364 366376
rect 159416 366364 159422 366376
rect 166810 366364 166816 366376
rect 159416 366336 166816 366364
rect 159416 366324 159422 366336
rect 166810 366324 166816 366336
rect 166868 366364 166874 366376
rect 203610 366364 203616 366376
rect 166868 366336 203616 366364
rect 166868 366324 166874 366336
rect 203610 366324 203616 366336
rect 203668 366324 203674 366376
rect 209038 366324 209044 366376
rect 209096 366364 209102 366376
rect 218054 366364 218060 366376
rect 209096 366336 218060 366364
rect 209096 366324 209102 366336
rect 218054 366324 218060 366336
rect 218112 366324 218118 366376
rect 273254 366324 273260 366376
rect 273312 366364 273318 366376
rect 349246 366364 349252 366376
rect 273312 366336 349252 366364
rect 273312 366324 273318 366336
rect 349246 366324 349252 366336
rect 349304 366324 349310 366376
rect 349798 366324 349804 366376
rect 349856 366364 349862 366376
rect 368566 366364 368572 366376
rect 349856 366336 368572 366364
rect 349856 366324 349862 366336
rect 368566 366324 368572 366336
rect 368624 366324 368630 366376
rect 139486 365712 139492 365764
rect 139544 365752 139550 365764
rect 232590 365752 232596 365764
rect 139544 365724 232596 365752
rect 139544 365712 139550 365724
rect 232590 365712 232596 365724
rect 232648 365712 232654 365764
rect 197170 365644 197176 365696
rect 197228 365684 197234 365696
rect 198826 365684 198832 365696
rect 197228 365656 198832 365684
rect 197228 365644 197234 365656
rect 198826 365644 198832 365656
rect 198884 365644 198890 365696
rect 338942 365032 338948 365084
rect 339000 365072 339006 365084
rect 363046 365072 363052 365084
rect 339000 365044 363052 365072
rect 339000 365032 339006 365044
rect 363046 365032 363052 365044
rect 363104 365032 363110 365084
rect 71590 364964 71596 365016
rect 71648 365004 71654 365016
rect 136818 365004 136824 365016
rect 71648 364976 136824 365004
rect 71648 364964 71654 364976
rect 136818 364964 136824 364976
rect 136876 364964 136882 365016
rect 137278 364964 137284 365016
rect 137336 365004 137342 365016
rect 185394 365004 185400 365016
rect 137336 364976 185400 365004
rect 137336 364964 137342 364976
rect 185394 364964 185400 364976
rect 185452 364964 185458 365016
rect 206370 364964 206376 365016
rect 206428 365004 206434 365016
rect 212534 365004 212540 365016
rect 206428 364976 212540 365004
rect 206428 364964 206434 364976
rect 212534 364964 212540 364976
rect 212592 364964 212598 365016
rect 213270 364964 213276 365016
rect 213328 365004 213334 365016
rect 356330 365004 356336 365016
rect 213328 364976 356336 365004
rect 213328 364964 213334 364976
rect 356330 364964 356336 364976
rect 356388 364964 356394 365016
rect 134702 364352 134708 364404
rect 134760 364392 134766 364404
rect 200114 364392 200120 364404
rect 134760 364364 200120 364392
rect 134760 364352 134766 364364
rect 200114 364352 200120 364364
rect 200172 364392 200178 364404
rect 206278 364392 206284 364404
rect 200172 364364 206284 364392
rect 200172 364352 200178 364364
rect 206278 364352 206284 364364
rect 206336 364352 206342 364404
rect 206462 364352 206468 364404
rect 206520 364392 206526 364404
rect 209222 364392 209228 364404
rect 206520 364364 209228 364392
rect 206520 364352 206526 364364
rect 209222 364352 209228 364364
rect 209280 364352 209286 364404
rect 58894 363604 58900 363656
rect 58952 363644 58958 363656
rect 130378 363644 130384 363656
rect 58952 363616 130384 363644
rect 58952 363604 58958 363616
rect 130378 363604 130384 363616
rect 130436 363604 130442 363656
rect 325602 363604 325608 363656
rect 325660 363644 325666 363656
rect 363138 363644 363144 363656
rect 325660 363616 363144 363644
rect 325660 363604 325666 363616
rect 363138 363604 363144 363616
rect 363196 363604 363202 363656
rect 137278 362992 137284 363044
rect 137336 363032 137342 363044
rect 188338 363032 188344 363044
rect 137336 363004 188344 363032
rect 137336 362992 137342 363004
rect 188338 362992 188344 363004
rect 188396 363032 188402 363044
rect 188706 363032 188712 363044
rect 188396 363004 188712 363032
rect 188396 362992 188402 363004
rect 188706 362992 188712 363004
rect 188764 362992 188770 363044
rect 103422 362924 103428 362976
rect 103480 362964 103486 362976
rect 149698 362964 149704 362976
rect 103480 362936 149704 362964
rect 103480 362924 103486 362936
rect 149698 362924 149704 362936
rect 149756 362924 149762 362976
rect 151722 362924 151728 362976
rect 151780 362964 151786 362976
rect 325602 362964 325608 362976
rect 151780 362936 325608 362964
rect 151780 362924 151786 362936
rect 325602 362924 325608 362936
rect 325660 362924 325666 362976
rect 322290 362244 322296 362296
rect 322348 362284 322354 362296
rect 347774 362284 347780 362296
rect 322348 362256 347780 362284
rect 322348 362244 322354 362256
rect 347774 362244 347780 362256
rect 347832 362244 347838 362296
rect 82078 362176 82084 362228
rect 82136 362216 82142 362228
rect 259546 362216 259552 362228
rect 82136 362188 259552 362216
rect 82136 362176 82142 362188
rect 259546 362176 259552 362188
rect 259604 362216 259610 362228
rect 260098 362216 260104 362228
rect 259604 362188 260104 362216
rect 259604 362176 259610 362188
rect 260098 362176 260104 362188
rect 260156 362176 260162 362228
rect 338850 362176 338856 362228
rect 338908 362216 338914 362228
rect 374086 362216 374092 362228
rect 338908 362188 374092 362216
rect 338908 362176 338914 362188
rect 374086 362176 374092 362188
rect 374144 362176 374150 362228
rect 81618 361564 81624 361616
rect 81676 361604 81682 361616
rect 82078 361604 82084 361616
rect 81676 361576 82084 361604
rect 81676 361564 81682 361576
rect 82078 361564 82084 361576
rect 82136 361564 82142 361616
rect 90542 361564 90548 361616
rect 90600 361604 90606 361616
rect 90600 361576 173940 361604
rect 90600 361564 90606 361576
rect 173912 361468 173940 361576
rect 186130 361496 186136 361548
rect 186188 361536 186194 361548
rect 367278 361536 367284 361548
rect 186188 361508 367284 361536
rect 186188 361496 186194 361508
rect 367278 361496 367284 361508
rect 367336 361496 367342 361548
rect 175090 361468 175096 361480
rect 173912 361440 175096 361468
rect 175090 361428 175096 361440
rect 175148 361468 175154 361480
rect 211154 361468 211160 361480
rect 175148 361440 211160 361468
rect 175148 361428 175154 361440
rect 211154 361428 211160 361440
rect 211212 361428 211218 361480
rect 103330 360816 103336 360868
rect 103388 360856 103394 360868
rect 155310 360856 155316 360868
rect 103388 360828 155316 360856
rect 103388 360816 103394 360828
rect 155310 360816 155316 360828
rect 155368 360816 155374 360868
rect 173342 360272 173348 360324
rect 173400 360312 173406 360324
rect 173894 360312 173900 360324
rect 173400 360284 173900 360312
rect 173400 360272 173406 360284
rect 173894 360272 173900 360284
rect 173952 360272 173958 360324
rect 90450 360204 90456 360256
rect 90508 360244 90514 360256
rect 181530 360244 181536 360256
rect 90508 360216 181536 360244
rect 90508 360204 90514 360216
rect 181530 360204 181536 360216
rect 181588 360204 181594 360256
rect 202138 359524 202144 359576
rect 202196 359564 202202 359576
rect 228358 359564 228364 359576
rect 202196 359536 228364 359564
rect 202196 359524 202202 359536
rect 228358 359524 228364 359536
rect 228416 359524 228422 359576
rect 80146 359456 80152 359508
rect 80204 359496 80210 359508
rect 81342 359496 81348 359508
rect 80204 359468 81348 359496
rect 80204 359456 80210 359468
rect 81342 359456 81348 359468
rect 81400 359496 81406 359508
rect 273254 359496 273260 359508
rect 81400 359468 273260 359496
rect 81400 359456 81406 359468
rect 273254 359456 273260 359468
rect 273312 359456 273318 359508
rect 99098 358776 99104 358828
rect 99156 358816 99162 358828
rect 192478 358816 192484 358828
rect 99156 358788 192484 358816
rect 99156 358776 99162 358788
rect 192478 358776 192484 358788
rect 192536 358776 192542 358828
rect 3326 358708 3332 358760
rect 3384 358748 3390 358760
rect 15838 358748 15844 358760
rect 3384 358720 15844 358748
rect 3384 358708 3390 358720
rect 15838 358708 15844 358720
rect 15896 358708 15902 358760
rect 47578 358708 47584 358760
rect 47636 358748 47642 358760
rect 48038 358748 48044 358760
rect 47636 358720 48044 358748
rect 47636 358708 47642 358720
rect 48038 358708 48044 358720
rect 48096 358708 48102 358760
rect 79318 358096 79324 358148
rect 79376 358136 79382 358148
rect 93854 358136 93860 358148
rect 79376 358108 93860 358136
rect 79376 358096 79382 358108
rect 93854 358096 93860 358108
rect 93912 358096 93918 358148
rect 206462 358096 206468 358148
rect 206520 358136 206526 358148
rect 253934 358136 253940 358148
rect 206520 358108 253940 358136
rect 206520 358096 206526 358108
rect 253934 358096 253940 358108
rect 253992 358096 253998 358148
rect 273898 358096 273904 358148
rect 273956 358136 273962 358148
rect 285674 358136 285680 358148
rect 273956 358108 285680 358136
rect 273956 358096 273962 358108
rect 285674 358096 285680 358108
rect 285732 358096 285738 358148
rect 47578 358028 47584 358080
rect 47636 358068 47642 358080
rect 139486 358068 139492 358080
rect 47636 358040 139492 358068
rect 47636 358028 47642 358040
rect 139486 358028 139492 358040
rect 139544 358028 139550 358080
rect 235534 358028 235540 358080
rect 235592 358068 235598 358080
rect 356146 358068 356152 358080
rect 235592 358040 356152 358068
rect 235592 358028 235598 358040
rect 356146 358028 356152 358040
rect 356204 358028 356210 358080
rect 142982 357484 142988 357536
rect 143040 357524 143046 357536
rect 190086 357524 190092 357536
rect 143040 357496 190092 357524
rect 143040 357484 143046 357496
rect 190086 357484 190092 357496
rect 190144 357484 190150 357536
rect 103514 357416 103520 357468
rect 103572 357456 103578 357468
rect 170398 357456 170404 357468
rect 103572 357428 170404 357456
rect 103572 357416 103578 357428
rect 170398 357416 170404 357428
rect 170456 357416 170462 357468
rect 180058 357348 180064 357400
rect 180116 357388 180122 357400
rect 180334 357388 180340 357400
rect 180116 357360 180340 357388
rect 180116 357348 180122 357360
rect 180334 357348 180340 357360
rect 180392 357348 180398 357400
rect 75730 356736 75736 356788
rect 75788 356776 75794 356788
rect 98822 356776 98828 356788
rect 75788 356748 98828 356776
rect 75788 356736 75794 356748
rect 98822 356736 98828 356748
rect 98880 356736 98886 356788
rect 129826 356736 129832 356788
rect 129884 356776 129890 356788
rect 160002 356776 160008 356788
rect 129884 356748 160008 356776
rect 129884 356736 129890 356748
rect 160002 356736 160008 356748
rect 160060 356776 160066 356788
rect 202138 356776 202144 356788
rect 160060 356748 202144 356776
rect 160060 356736 160066 356748
rect 202138 356736 202144 356748
rect 202196 356736 202202 356788
rect 64598 356668 64604 356720
rect 64656 356708 64662 356720
rect 107746 356708 107752 356720
rect 64656 356680 107752 356708
rect 64656 356668 64662 356680
rect 107746 356668 107752 356680
rect 107804 356668 107810 356720
rect 110322 356668 110328 356720
rect 110380 356708 110386 356720
rect 164234 356708 164240 356720
rect 110380 356680 164240 356708
rect 110380 356668 110386 356680
rect 164234 356668 164240 356680
rect 164292 356668 164298 356720
rect 164694 356668 164700 356720
rect 164752 356708 164758 356720
rect 180334 356708 180340 356720
rect 164752 356680 180340 356708
rect 164752 356668 164758 356680
rect 180334 356668 180340 356680
rect 180392 356668 180398 356720
rect 201402 356668 201408 356720
rect 201460 356708 201466 356720
rect 240226 356708 240232 356720
rect 201460 356680 240232 356708
rect 201460 356668 201466 356680
rect 240226 356668 240232 356680
rect 240284 356668 240290 356720
rect 132586 355988 132592 356040
rect 132644 356028 132650 356040
rect 244274 356028 244280 356040
rect 132644 356000 244280 356028
rect 132644 355988 132650 356000
rect 244274 355988 244280 356000
rect 244332 356028 244338 356040
rect 244918 356028 244924 356040
rect 244332 356000 244924 356028
rect 244332 355988 244338 356000
rect 244918 355988 244924 356000
rect 244976 355988 244982 356040
rect 81342 355308 81348 355360
rect 81400 355348 81406 355360
rect 132586 355348 132592 355360
rect 81400 355320 132592 355348
rect 81400 355308 81406 355320
rect 132586 355308 132592 355320
rect 132644 355308 132650 355360
rect 195882 355308 195888 355360
rect 195940 355348 195946 355360
rect 230474 355348 230480 355360
rect 195940 355320 230480 355348
rect 195940 355308 195946 355320
rect 230474 355308 230480 355320
rect 230532 355308 230538 355360
rect 94498 354696 94504 354748
rect 94556 354736 94562 354748
rect 195882 354736 195888 354748
rect 94556 354708 195888 354736
rect 94556 354696 94562 354708
rect 195882 354696 195888 354708
rect 195940 354696 195946 354748
rect 93210 353948 93216 354000
rect 93268 353988 93274 354000
rect 120718 353988 120724 354000
rect 93268 353960 120724 353988
rect 93268 353948 93274 353960
rect 120718 353948 120724 353960
rect 120776 353948 120782 354000
rect 305638 353948 305644 354000
rect 305696 353988 305702 354000
rect 340874 353988 340880 354000
rect 305696 353960 340880 353988
rect 305696 353948 305702 353960
rect 340874 353948 340880 353960
rect 340932 353948 340938 354000
rect 104894 353336 104900 353388
rect 104952 353376 104958 353388
rect 199378 353376 199384 353388
rect 104952 353348 199384 353376
rect 104952 353336 104958 353348
rect 199378 353336 199384 353348
rect 199436 353336 199442 353388
rect 120626 353268 120632 353320
rect 120684 353308 120690 353320
rect 220078 353308 220084 353320
rect 120684 353280 220084 353308
rect 120684 353268 120690 353280
rect 220078 353268 220084 353280
rect 220136 353268 220142 353320
rect 235258 352588 235264 352640
rect 235316 352628 235322 352640
rect 249794 352628 249800 352640
rect 235316 352600 249800 352628
rect 235316 352588 235322 352600
rect 249794 352588 249800 352600
rect 249852 352588 249858 352640
rect 76650 352520 76656 352572
rect 76708 352560 76714 352572
rect 158714 352560 158720 352572
rect 76708 352532 158720 352560
rect 76708 352520 76714 352532
rect 158714 352520 158720 352532
rect 158772 352520 158778 352572
rect 161290 352520 161296 352572
rect 161348 352560 161354 352572
rect 222194 352560 222200 352572
rect 161348 352532 222200 352560
rect 161348 352520 161354 352532
rect 222194 352520 222200 352532
rect 222252 352520 222258 352572
rect 240778 352520 240784 352572
rect 240836 352560 240842 352572
rect 580166 352560 580172 352572
rect 240836 352532 580172 352560
rect 240836 352520 240842 352532
rect 580166 352520 580172 352532
rect 580224 352520 580230 352572
rect 240226 352180 240232 352232
rect 240284 352220 240290 352232
rect 240778 352220 240784 352232
rect 240284 352192 240784 352220
rect 240284 352180 240290 352192
rect 240778 352180 240784 352192
rect 240836 352180 240842 352232
rect 101490 351908 101496 351960
rect 101548 351948 101554 351960
rect 180058 351948 180064 351960
rect 101548 351920 180064 351948
rect 101548 351908 101554 351920
rect 180058 351908 180064 351920
rect 180116 351908 180122 351960
rect 96430 351228 96436 351280
rect 96488 351268 96494 351280
rect 120626 351268 120632 351280
rect 96488 351240 120632 351268
rect 96488 351228 96494 351240
rect 120626 351228 120632 351240
rect 120684 351228 120690 351280
rect 64690 351160 64696 351212
rect 64748 351200 64754 351212
rect 66990 351200 66996 351212
rect 64748 351172 66996 351200
rect 64748 351160 64754 351172
rect 66990 351160 66996 351172
rect 67048 351200 67054 351212
rect 195238 351200 195244 351212
rect 67048 351172 195244 351200
rect 67048 351160 67054 351172
rect 195238 351160 195244 351172
rect 195296 351160 195302 351212
rect 255314 351160 255320 351212
rect 255372 351200 255378 351212
rect 273990 351200 273996 351212
rect 255372 351172 273996 351200
rect 255372 351160 255378 351172
rect 273990 351160 273996 351172
rect 274048 351160 274054 351212
rect 124122 350548 124128 350600
rect 124180 350588 124186 350600
rect 255314 350588 255320 350600
rect 124180 350560 255320 350588
rect 124180 350548 124186 350560
rect 255314 350548 255320 350560
rect 255372 350548 255378 350600
rect 233142 350480 233148 350532
rect 233200 350520 233206 350532
rect 240134 350520 240140 350532
rect 233200 350492 240140 350520
rect 233200 350480 233206 350492
rect 240134 350480 240140 350492
rect 240192 350480 240198 350532
rect 86862 349868 86868 349920
rect 86920 349908 86926 349920
rect 100018 349908 100024 349920
rect 86920 349880 100024 349908
rect 86920 349868 86926 349880
rect 100018 349868 100024 349880
rect 100076 349868 100082 349920
rect 110414 349868 110420 349920
rect 110472 349908 110478 349920
rect 158898 349908 158904 349920
rect 110472 349880 158904 349908
rect 110472 349868 110478 349880
rect 158898 349868 158904 349880
rect 158956 349868 158962 349920
rect 25498 349800 25504 349852
rect 25556 349840 25562 349852
rect 67818 349840 67824 349852
rect 25556 349812 67824 349840
rect 25556 349800 25562 349812
rect 67818 349800 67824 349812
rect 67876 349840 67882 349852
rect 125686 349840 125692 349852
rect 67876 349812 125692 349840
rect 67876 349800 67882 349812
rect 125686 349800 125692 349812
rect 125744 349840 125750 349852
rect 142982 349840 142988 349852
rect 125744 349812 142988 349840
rect 125744 349800 125750 349812
rect 142982 349800 142988 349812
rect 143040 349800 143046 349852
rect 169202 349800 169208 349852
rect 169260 349840 169266 349852
rect 309134 349840 309140 349852
rect 169260 349812 309140 349840
rect 169260 349800 169266 349812
rect 309134 349800 309140 349812
rect 309192 349800 309198 349852
rect 155310 349596 155316 349648
rect 155368 349636 155374 349648
rect 155862 349636 155868 349648
rect 155368 349608 155868 349636
rect 155368 349596 155374 349608
rect 155862 349596 155868 349608
rect 155920 349596 155926 349648
rect 155862 349120 155868 349172
rect 155920 349160 155926 349172
rect 233142 349160 233148 349172
rect 155920 349132 233148 349160
rect 155920 349120 155926 349132
rect 233142 349120 233148 349132
rect 233200 349120 233206 349172
rect 105538 348372 105544 348424
rect 105596 348412 105602 348424
rect 157978 348412 157984 348424
rect 105596 348384 157984 348412
rect 105596 348372 105602 348384
rect 157978 348372 157984 348384
rect 158036 348372 158042 348424
rect 196802 348372 196808 348424
rect 196860 348412 196866 348424
rect 231118 348412 231124 348424
rect 196860 348384 231124 348412
rect 196860 348372 196866 348384
rect 231118 348372 231124 348384
rect 231176 348372 231182 348424
rect 130378 347828 130384 347880
rect 130436 347868 130442 347880
rect 133874 347868 133880 347880
rect 130436 347840 133880 347868
rect 130436 347828 130442 347840
rect 133874 347828 133880 347840
rect 133932 347828 133938 347880
rect 129090 347760 129096 347812
rect 129148 347800 129154 347812
rect 201586 347800 201592 347812
rect 129148 347772 201592 347800
rect 129148 347760 129154 347772
rect 201586 347760 201592 347772
rect 201644 347800 201650 347812
rect 202230 347800 202236 347812
rect 201644 347772 202236 347800
rect 201644 347760 201650 347772
rect 202230 347760 202236 347772
rect 202288 347760 202294 347812
rect 93762 347012 93768 347064
rect 93820 347052 93826 347064
rect 137278 347052 137284 347064
rect 93820 347024 137284 347052
rect 93820 347012 93826 347024
rect 137278 347012 137284 347024
rect 137336 347012 137342 347064
rect 139302 347012 139308 347064
rect 139360 347052 139366 347064
rect 191650 347052 191656 347064
rect 139360 347024 191656 347052
rect 139360 347012 139366 347024
rect 191650 347012 191656 347024
rect 191708 347012 191714 347064
rect 121546 346400 121552 346452
rect 121604 346440 121610 346452
rect 122742 346440 122748 346452
rect 121604 346412 122748 346440
rect 121604 346400 121610 346412
rect 122742 346400 122748 346412
rect 122800 346440 122806 346452
rect 221458 346440 221464 346452
rect 122800 346412 221464 346440
rect 122800 346400 122806 346412
rect 221458 346400 221464 346412
rect 221516 346400 221522 346452
rect 135162 346332 135168 346384
rect 135220 346372 135226 346384
rect 139394 346372 139400 346384
rect 135220 346344 139400 346372
rect 135220 346332 135226 346344
rect 139394 346332 139400 346344
rect 139452 346332 139458 346384
rect 2774 346264 2780 346316
rect 2832 346304 2838 346316
rect 4798 346304 4804 346316
rect 2832 346276 4804 346304
rect 2832 346264 2838 346276
rect 4798 346264 4804 346276
rect 4856 346264 4862 346316
rect 84102 345720 84108 345772
rect 84160 345760 84166 345772
rect 108482 345760 108488 345772
rect 84160 345732 108488 345760
rect 84160 345720 84166 345732
rect 108482 345720 108488 345732
rect 108540 345720 108546 345772
rect 119338 345720 119344 345772
rect 119396 345760 119402 345772
rect 157334 345760 157340 345772
rect 119396 345732 157340 345760
rect 119396 345720 119402 345732
rect 157334 345720 157340 345732
rect 157392 345720 157398 345772
rect 58894 345652 58900 345704
rect 58952 345692 58958 345704
rect 134518 345692 134524 345704
rect 58952 345664 134524 345692
rect 58952 345652 58958 345664
rect 134518 345652 134524 345664
rect 134576 345652 134582 345704
rect 146110 345040 146116 345092
rect 146168 345080 146174 345092
rect 242250 345080 242256 345092
rect 146168 345052 242256 345080
rect 146168 345040 146174 345052
rect 242250 345040 242256 345052
rect 242308 345040 242314 345092
rect 156598 344496 156604 344548
rect 156656 344536 156662 344548
rect 162946 344536 162952 344548
rect 156656 344508 162952 344536
rect 156656 344496 156662 344508
rect 162946 344496 162952 344508
rect 163004 344496 163010 344548
rect 110322 344360 110328 344412
rect 110380 344400 110386 344412
rect 116670 344400 116676 344412
rect 110380 344372 116676 344400
rect 110380 344360 110386 344372
rect 116670 344360 116676 344372
rect 116728 344360 116734 344412
rect 79686 344292 79692 344344
rect 79744 344332 79750 344344
rect 111058 344332 111064 344344
rect 79744 344304 111064 344332
rect 79744 344292 79750 344304
rect 111058 344292 111064 344304
rect 111116 344292 111122 344344
rect 120718 344292 120724 344344
rect 120776 344332 120782 344344
rect 235534 344332 235540 344344
rect 120776 344304 235540 344332
rect 120776 344292 120782 344304
rect 235534 344292 235540 344304
rect 235592 344292 235598 344344
rect 114462 343680 114468 343732
rect 114520 343720 114526 343732
rect 124030 343720 124036 343732
rect 114520 343692 124036 343720
rect 114520 343680 114526 343692
rect 124030 343680 124036 343692
rect 124088 343680 124094 343732
rect 63402 343612 63408 343664
rect 63460 343652 63466 343664
rect 66898 343652 66904 343664
rect 63460 343624 66904 343652
rect 63460 343612 63466 343624
rect 66898 343612 66904 343624
rect 66956 343612 66962 343664
rect 120074 343612 120080 343664
rect 120132 343652 120138 343664
rect 120718 343652 120724 343664
rect 120132 343624 120724 343652
rect 120132 343612 120138 343624
rect 120718 343612 120724 343624
rect 120776 343612 120782 343664
rect 144638 343612 144644 343664
rect 144696 343652 144702 343664
rect 156598 343652 156604 343664
rect 144696 343624 156604 343652
rect 144696 343612 144702 343624
rect 156598 343612 156604 343624
rect 156656 343612 156662 343664
rect 155770 343544 155776 343596
rect 155828 343584 155834 343596
rect 207106 343584 207112 343596
rect 155828 343556 207112 343584
rect 155828 343544 155834 343556
rect 207106 343544 207112 343556
rect 207164 343544 207170 343596
rect 97902 342932 97908 342984
rect 97960 342972 97966 342984
rect 128998 342972 129004 342984
rect 97960 342944 129004 342972
rect 97960 342932 97966 342944
rect 128998 342932 129004 342944
rect 129056 342932 129062 342984
rect 73798 342864 73804 342916
rect 73856 342904 73862 342916
rect 144638 342904 144644 342916
rect 73856 342876 144644 342904
rect 73856 342864 73862 342876
rect 144638 342864 144644 342876
rect 144696 342864 144702 342916
rect 148962 342864 148968 342916
rect 149020 342904 149026 342916
rect 158898 342904 158904 342916
rect 149020 342876 158904 342904
rect 149020 342864 149026 342876
rect 158898 342864 158904 342876
rect 158956 342864 158962 342916
rect 207106 342320 207112 342372
rect 207164 342360 207170 342372
rect 207658 342360 207664 342372
rect 207164 342332 207664 342360
rect 207164 342320 207170 342332
rect 207658 342320 207664 342332
rect 207716 342320 207722 342372
rect 85390 342252 85396 342304
rect 85448 342292 85454 342304
rect 90542 342292 90548 342304
rect 85448 342264 90548 342292
rect 85448 342252 85454 342264
rect 90542 342252 90548 342264
rect 90600 342252 90606 342304
rect 141418 342252 141424 342304
rect 141476 342292 141482 342304
rect 142062 342292 142068 342304
rect 141476 342264 142068 342292
rect 141476 342252 141482 342264
rect 142062 342252 142068 342264
rect 142120 342292 142126 342304
rect 155126 342292 155132 342304
rect 142120 342264 155132 342292
rect 142120 342252 142126 342264
rect 155126 342252 155132 342264
rect 155184 342252 155190 342304
rect 158806 342252 158812 342304
rect 158864 342292 158870 342304
rect 227070 342292 227076 342304
rect 158864 342264 227076 342292
rect 158864 342252 158870 342264
rect 227070 342252 227076 342264
rect 227128 342252 227134 342304
rect 55030 341504 55036 341556
rect 55088 341544 55094 341556
rect 86954 341544 86960 341556
rect 55088 341516 86960 341544
rect 55088 341504 55094 341516
rect 86954 341504 86960 341516
rect 87012 341504 87018 341556
rect 155218 341504 155224 341556
rect 155276 341544 155282 341556
rect 195238 341544 195244 341556
rect 155276 341516 195244 341544
rect 155276 341504 155282 341516
rect 195238 341504 195244 341516
rect 195296 341504 195302 341556
rect 304258 341504 304264 341556
rect 304316 341544 304322 341556
rect 372706 341544 372712 341556
rect 304316 341516 372712 341544
rect 304316 341504 304322 341516
rect 372706 341504 372712 341516
rect 372764 341504 372770 341556
rect 125042 340960 125048 341012
rect 125100 341000 125106 341012
rect 140774 341000 140780 341012
rect 125100 340972 140780 341000
rect 125100 340960 125106 340972
rect 140774 340960 140780 340972
rect 140832 340960 140838 341012
rect 95142 340892 95148 340944
rect 95200 340932 95206 340944
rect 254026 340932 254032 340944
rect 95200 340904 254032 340932
rect 95200 340892 95206 340904
rect 254026 340892 254032 340904
rect 254084 340892 254090 340944
rect 140774 340824 140780 340876
rect 140832 340864 140838 340876
rect 153194 340864 153200 340876
rect 140832 340836 153200 340864
rect 140832 340824 140838 340836
rect 153194 340824 153200 340836
rect 153252 340864 153258 340876
rect 153838 340864 153844 340876
rect 153252 340836 153844 340864
rect 153252 340824 153258 340836
rect 153838 340824 153844 340836
rect 153896 340824 153902 340876
rect 229738 340212 229744 340264
rect 229796 340252 229802 340264
rect 309778 340252 309784 340264
rect 229796 340224 309784 340252
rect 229796 340212 229802 340224
rect 309778 340212 309784 340224
rect 309836 340212 309842 340264
rect 52362 340144 52368 340196
rect 52420 340184 52426 340196
rect 125042 340184 125048 340196
rect 52420 340156 125048 340184
rect 52420 340144 52426 340156
rect 125042 340144 125048 340156
rect 125100 340144 125106 340196
rect 156690 340144 156696 340196
rect 156748 340184 156754 340196
rect 337378 340184 337384 340196
rect 156748 340156 337384 340184
rect 156748 340144 156754 340156
rect 337378 340144 337384 340156
rect 337436 340144 337442 340196
rect 61838 339464 61844 339516
rect 61896 339504 61902 339516
rect 162302 339504 162308 339516
rect 61896 339476 162308 339504
rect 61896 339464 61902 339476
rect 162302 339464 162308 339476
rect 162360 339464 162366 339516
rect 156598 338784 156604 338836
rect 156656 338824 156662 338836
rect 207750 338824 207756 338836
rect 156656 338796 207756 338824
rect 156656 338784 156662 338796
rect 207750 338784 207756 338796
rect 207808 338784 207814 338836
rect 64782 338716 64788 338768
rect 64840 338756 64846 338768
rect 116578 338756 116584 338768
rect 64840 338728 116584 338756
rect 64840 338716 64846 338728
rect 116578 338716 116584 338728
rect 116636 338716 116642 338768
rect 201402 338716 201408 338768
rect 201460 338756 201466 338768
rect 335354 338756 335360 338768
rect 201460 338728 335360 338756
rect 201460 338716 201466 338728
rect 335354 338716 335360 338728
rect 335412 338716 335418 338768
rect 118510 338172 118516 338224
rect 118568 338212 118574 338224
rect 131114 338212 131120 338224
rect 118568 338184 131120 338212
rect 118568 338172 118574 338184
rect 131114 338172 131120 338184
rect 131172 338172 131178 338224
rect 147674 338172 147680 338224
rect 147732 338212 147738 338224
rect 156874 338212 156880 338224
rect 147732 338184 156880 338212
rect 147732 338172 147738 338184
rect 156874 338172 156880 338184
rect 156932 338172 156938 338224
rect 117222 338104 117228 338156
rect 117280 338144 117286 338156
rect 196802 338144 196808 338156
rect 117280 338116 196808 338144
rect 117280 338104 117286 338116
rect 196802 338104 196808 338116
rect 196860 338104 196866 338156
rect 77294 337424 77300 337476
rect 77352 337464 77358 337476
rect 85574 337464 85580 337476
rect 77352 337436 85580 337464
rect 77352 337424 77358 337436
rect 85574 337424 85580 337436
rect 85632 337424 85638 337476
rect 52178 337356 52184 337408
rect 52236 337396 52242 337408
rect 82814 337396 82820 337408
rect 52236 337368 82820 337396
rect 52236 337356 52242 337368
rect 82814 337356 82820 337368
rect 82872 337356 82878 337408
rect 107378 337356 107384 337408
rect 107436 337396 107442 337408
rect 129090 337396 129096 337408
rect 107436 337368 129096 337396
rect 107436 337356 107442 337368
rect 129090 337356 129096 337368
rect 129148 337356 129154 337408
rect 139210 337356 139216 337408
rect 139268 337396 139274 337408
rect 147674 337396 147680 337408
rect 139268 337368 147680 337396
rect 139268 337356 139274 337368
rect 147674 337356 147680 337368
rect 147732 337356 147738 337408
rect 170398 337356 170404 337408
rect 170456 337396 170462 337408
rect 249058 337396 249064 337408
rect 170456 337368 249064 337396
rect 170456 337356 170462 337368
rect 249058 337356 249064 337368
rect 249116 337356 249122 337408
rect 275278 337356 275284 337408
rect 275336 337396 275342 337408
rect 371326 337396 371332 337408
rect 275336 337368 371332 337396
rect 275336 337356 275342 337368
rect 371326 337356 371332 337368
rect 371384 337356 371390 337408
rect 149606 336812 149612 336864
rect 149664 336852 149670 336864
rect 174538 336852 174544 336864
rect 149664 336824 174544 336852
rect 149664 336812 149670 336824
rect 174538 336812 174544 336824
rect 174596 336812 174602 336864
rect 136542 336744 136548 336796
rect 136600 336784 136606 336796
rect 169846 336784 169852 336796
rect 136600 336756 169852 336784
rect 136600 336744 136606 336756
rect 169846 336744 169852 336756
rect 169904 336744 169910 336796
rect 155770 335996 155776 336048
rect 155828 336036 155834 336048
rect 224402 336036 224408 336048
rect 155828 336008 224408 336036
rect 155828 335996 155834 336008
rect 224402 335996 224408 336008
rect 224460 335996 224466 336048
rect 148134 335384 148140 335436
rect 148192 335424 148198 335436
rect 155126 335424 155132 335436
rect 148192 335396 155132 335424
rect 148192 335384 148198 335396
rect 155126 335384 155132 335396
rect 155184 335384 155190 335436
rect 60642 335316 60648 335368
rect 60700 335356 60706 335368
rect 84654 335356 84660 335368
rect 60700 335328 84660 335356
rect 60700 335316 60706 335328
rect 84654 335316 84660 335328
rect 84712 335316 84718 335368
rect 134886 335316 134892 335368
rect 134944 335356 134950 335368
rect 163498 335356 163504 335368
rect 134944 335328 163504 335356
rect 134944 335316 134950 335328
rect 163498 335316 163504 335328
rect 163556 335316 163562 335368
rect 155126 334772 155132 334824
rect 155184 334812 155190 334824
rect 160738 334812 160744 334824
rect 155184 334784 160744 334812
rect 155184 334772 155190 334784
rect 160738 334772 160744 334784
rect 160796 334772 160802 334824
rect 129274 334636 129280 334688
rect 129332 334676 129338 334688
rect 136542 334676 136548 334688
rect 129332 334648 136548 334676
rect 129332 334636 129338 334648
rect 136542 334636 136548 334648
rect 136600 334636 136606 334688
rect 149054 334636 149060 334688
rect 149112 334676 149118 334688
rect 155862 334676 155868 334688
rect 149112 334648 155868 334676
rect 149112 334636 149118 334648
rect 155862 334636 155868 334648
rect 155920 334636 155926 334688
rect 189902 334636 189908 334688
rect 189960 334676 189966 334688
rect 243630 334676 243636 334688
rect 189960 334648 243636 334676
rect 189960 334636 189966 334648
rect 243630 334636 243636 334648
rect 243688 334636 243694 334688
rect 135162 334568 135168 334620
rect 135220 334608 135226 334620
rect 149606 334608 149612 334620
rect 135220 334580 149612 334608
rect 135220 334568 135226 334580
rect 149606 334568 149612 334580
rect 149664 334568 149670 334620
rect 173158 334568 173164 334620
rect 173216 334608 173222 334620
rect 192662 334608 192668 334620
rect 173216 334580 192668 334608
rect 173216 334568 173222 334580
rect 192662 334568 192668 334580
rect 192720 334568 192726 334620
rect 223022 334568 223028 334620
rect 223080 334608 223086 334620
rect 582374 334608 582380 334620
rect 223080 334580 582380 334608
rect 223080 334568 223086 334580
rect 582374 334568 582380 334580
rect 582432 334568 582438 334620
rect 3418 333956 3424 334008
rect 3476 333996 3482 334008
rect 124214 333996 124220 334008
rect 3476 333968 124220 333996
rect 3476 333956 3482 333968
rect 124214 333956 124220 333968
rect 124272 333996 124278 334008
rect 124950 333996 124956 334008
rect 124272 333968 124956 333996
rect 124272 333956 124278 333968
rect 124950 333956 124956 333968
rect 125008 333956 125014 334008
rect 137094 333956 137100 334008
rect 137152 333996 137158 334008
rect 139486 333996 139492 334008
rect 137152 333968 139492 333996
rect 137152 333956 137158 333968
rect 139486 333956 139492 333968
rect 139544 333956 139550 334008
rect 140774 333956 140780 334008
rect 140832 333996 140838 334008
rect 172698 333996 172704 334008
rect 140832 333968 172704 333996
rect 140832 333956 140838 333968
rect 172698 333956 172704 333968
rect 172756 333956 172762 334008
rect 52270 333888 52276 333940
rect 52328 333928 52334 333940
rect 94314 333928 94320 333940
rect 52328 333900 94320 333928
rect 52328 333888 52334 333900
rect 94314 333888 94320 333900
rect 94372 333888 94378 333940
rect 14 333208 20 333260
rect 72 333248 78 333260
rect 52270 333248 52276 333260
rect 72 333220 52276 333248
rect 72 333208 78 333220
rect 52270 333208 52276 333220
rect 52328 333208 52334 333260
rect 83366 333208 83372 333260
rect 83424 333248 83430 333260
rect 106918 333248 106924 333260
rect 83424 333220 106924 333248
rect 83424 333208 83430 333220
rect 106918 333208 106924 333220
rect 106976 333208 106982 333260
rect 132126 333208 132132 333260
rect 132184 333248 132190 333260
rect 140774 333248 140780 333260
rect 132184 333220 140780 333248
rect 132184 333208 132190 333220
rect 140774 333208 140780 333220
rect 140832 333208 140838 333260
rect 240870 333208 240876 333260
rect 240928 333248 240934 333260
rect 349798 333248 349804 333260
rect 240928 333220 349804 333248
rect 240928 333208 240934 333220
rect 349798 333208 349804 333220
rect 349856 333208 349862 333260
rect 143074 332664 143080 332716
rect 143132 332704 143138 332716
rect 252554 332704 252560 332716
rect 143132 332676 252560 332704
rect 143132 332664 143138 332676
rect 252554 332664 252560 332676
rect 252612 332664 252618 332716
rect 67818 332596 67824 332648
rect 67876 332636 67882 332648
rect 72418 332636 72424 332648
rect 67876 332608 72424 332636
rect 67876 332596 67882 332608
rect 72418 332596 72424 332608
rect 72476 332596 72482 332648
rect 106642 332596 106648 332648
rect 106700 332636 106706 332648
rect 229186 332636 229192 332648
rect 106700 332608 229192 332636
rect 106700 332596 106706 332608
rect 229186 332596 229192 332608
rect 229244 332596 229250 332648
rect 59078 332528 59084 332580
rect 59136 332568 59142 332580
rect 101490 332568 101496 332580
rect 59136 332540 101496 332568
rect 59136 332528 59142 332540
rect 101490 332528 101496 332540
rect 101548 332528 101554 332580
rect 142890 332528 142896 332580
rect 142948 332568 142954 332580
rect 146938 332568 146944 332580
rect 142948 332540 146944 332568
rect 142948 332528 142954 332540
rect 146938 332528 146944 332540
rect 146996 332528 147002 332580
rect 74258 332460 74264 332512
rect 74316 332500 74322 332512
rect 76742 332500 76748 332512
rect 74316 332472 76748 332500
rect 74316 332460 74322 332472
rect 76742 332460 76748 332472
rect 76800 332460 76806 332512
rect 70762 332120 70768 332172
rect 70820 332160 70826 332172
rect 71498 332160 71504 332172
rect 70820 332132 71504 332160
rect 70820 332120 70826 332132
rect 71498 332120 71504 332132
rect 71556 332120 71562 332172
rect 78582 332120 78588 332172
rect 78640 332160 78646 332172
rect 79318 332160 79324 332172
rect 78640 332132 79324 332160
rect 78640 332120 78646 332132
rect 79318 332120 79324 332132
rect 79376 332120 79382 332172
rect 88242 332120 88248 332172
rect 88300 332160 88306 332172
rect 90450 332160 90456 332172
rect 88300 332132 90456 332160
rect 88300 332120 88306 332132
rect 90450 332120 90456 332132
rect 90508 332120 90514 332172
rect 110874 332120 110880 332172
rect 110932 332160 110938 332172
rect 111610 332160 111616 332172
rect 110932 332132 111616 332160
rect 110932 332120 110938 332132
rect 111610 332120 111616 332132
rect 111668 332120 111674 332172
rect 113818 332120 113824 332172
rect 113876 332160 113882 332172
rect 114462 332160 114468 332172
rect 113876 332132 114468 332160
rect 113876 332120 113882 332132
rect 114462 332120 114468 332132
rect 114520 332120 114526 332172
rect 115290 332120 115296 332172
rect 115348 332160 115354 332172
rect 115842 332160 115848 332172
rect 115348 332132 115848 332160
rect 115348 332120 115354 332132
rect 115842 332120 115848 332132
rect 115900 332120 115906 332172
rect 116762 332120 116768 332172
rect 116820 332160 116826 332172
rect 117222 332160 117228 332172
rect 116820 332132 117228 332160
rect 116820 332120 116826 332132
rect 117222 332120 117228 332132
rect 117280 332120 117286 332172
rect 118510 332120 118516 332172
rect 118568 332160 118574 332172
rect 119062 332160 119068 332172
rect 118568 332132 119068 332160
rect 118568 332120 118574 332132
rect 119062 332120 119068 332132
rect 119120 332120 119126 332172
rect 123294 332120 123300 332172
rect 123352 332160 123358 332172
rect 124122 332160 124128 332172
rect 123352 332132 124128 332160
rect 123352 332120 123358 332132
rect 124122 332120 124128 332132
rect 124180 332120 124186 332172
rect 125594 332120 125600 332172
rect 125652 332160 125658 332172
rect 126422 332160 126428 332172
rect 125652 332132 126428 332160
rect 125652 332120 125658 332132
rect 126422 332120 126428 332132
rect 126480 332120 126486 332172
rect 129918 332120 129924 332172
rect 129976 332160 129982 332172
rect 130378 332160 130384 332172
rect 129976 332132 130384 332160
rect 129976 332120 129982 332132
rect 130378 332120 130384 332132
rect 130436 332120 130442 332172
rect 138658 332120 138664 332172
rect 138716 332160 138722 332172
rect 139302 332160 139308 332172
rect 138716 332132 139308 332160
rect 138716 332120 138722 332132
rect 139302 332120 139308 332132
rect 139360 332120 139366 332172
rect 143810 332120 143816 332172
rect 143868 332160 143874 332172
rect 144730 332160 144736 332172
rect 143868 332132 144736 332160
rect 143868 332120 143874 332132
rect 144730 332120 144736 332132
rect 144788 332120 144794 332172
rect 145282 332120 145288 332172
rect 145340 332160 145346 332172
rect 146018 332160 146024 332172
rect 145340 332132 146024 332160
rect 145340 332120 145346 332132
rect 146018 332120 146024 332132
rect 146076 332120 146082 332172
rect 149698 332120 149704 332172
rect 149756 332160 149762 332172
rect 150342 332160 150348 332172
rect 149756 332132 150348 332160
rect 149756 332120 149762 332132
rect 150342 332120 150348 332132
rect 150400 332120 150406 332172
rect 98546 331984 98552 332036
rect 98604 332024 98610 332036
rect 99282 332024 99288 332036
rect 98604 331996 99288 332024
rect 98604 331984 98610 331996
rect 99282 331984 99288 331996
rect 99340 331984 99346 332036
rect 162210 331984 162216 332036
rect 162268 332024 162274 332036
rect 164970 332024 164976 332036
rect 162268 331996 164976 332024
rect 162268 331984 162274 331996
rect 164970 331984 164976 331996
rect 165028 331984 165034 332036
rect 232590 331916 232596 331968
rect 232648 331956 232654 331968
rect 244274 331956 244280 331968
rect 232648 331928 244280 331956
rect 232648 331916 232654 331928
rect 244274 331916 244280 331928
rect 244332 331916 244338 331968
rect 33778 331848 33784 331900
rect 33836 331888 33842 331900
rect 59078 331888 59084 331900
rect 33836 331860 59084 331888
rect 33836 331848 33842 331860
rect 59078 331848 59084 331860
rect 59136 331848 59142 331900
rect 107838 331848 107844 331900
rect 107896 331888 107902 331900
rect 135162 331888 135168 331900
rect 107896 331860 135168 331888
rect 107896 331848 107902 331860
rect 135162 331848 135168 331860
rect 135220 331848 135226 331900
rect 188614 331848 188620 331900
rect 188672 331888 188678 331900
rect 202874 331888 202880 331900
rect 188672 331860 202880 331888
rect 188672 331848 188678 331860
rect 202874 331848 202880 331860
rect 202932 331848 202938 331900
rect 215386 331848 215392 331900
rect 215444 331888 215450 331900
rect 292574 331888 292580 331900
rect 215444 331860 292580 331888
rect 215444 331848 215450 331860
rect 292574 331848 292580 331860
rect 292632 331848 292638 331900
rect 80238 331576 80244 331628
rect 80296 331616 80302 331628
rect 81342 331616 81348 331628
rect 80296 331588 81348 331616
rect 80296 331576 80302 331588
rect 81342 331576 81348 331588
rect 81400 331576 81406 331628
rect 135714 331576 135720 331628
rect 135772 331616 135778 331628
rect 141418 331616 141424 331628
rect 135772 331588 141424 331616
rect 135772 331576 135778 331588
rect 141418 331576 141424 331588
rect 141476 331576 141482 331628
rect 95602 331508 95608 331560
rect 95660 331548 95666 331560
rect 96522 331548 96528 331560
rect 95660 331520 96528 331548
rect 95660 331508 95666 331520
rect 96522 331508 96528 331520
rect 96580 331508 96586 331560
rect 109402 331508 109408 331560
rect 109460 331548 109466 331560
rect 110322 331548 110328 331560
rect 109460 331520 110328 331548
rect 109460 331508 109466 331520
rect 110322 331508 110328 331520
rect 110380 331508 110386 331560
rect 90450 331440 90456 331492
rect 90508 331480 90514 331492
rect 93118 331480 93124 331492
rect 90508 331452 93124 331480
rect 90508 331440 90514 331452
rect 93118 331440 93124 331452
rect 93176 331440 93182 331492
rect 94130 331440 94136 331492
rect 94188 331480 94194 331492
rect 95142 331480 95148 331492
rect 94188 331452 95148 331480
rect 94188 331440 94194 331452
rect 95142 331440 95148 331452
rect 95200 331440 95206 331492
rect 100018 331440 100024 331492
rect 100076 331480 100082 331492
rect 100662 331480 100668 331492
rect 100076 331452 100668 331480
rect 100076 331440 100082 331452
rect 100662 331440 100668 331452
rect 100720 331440 100726 331492
rect 134242 331440 134248 331492
rect 134300 331480 134306 331492
rect 139210 331480 139216 331492
rect 134300 331452 139216 331480
rect 134300 331440 134306 331452
rect 139210 331440 139216 331452
rect 139268 331440 139274 331492
rect 83090 331304 83096 331356
rect 83148 331344 83154 331356
rect 84102 331344 84108 331356
rect 83148 331316 84108 331344
rect 83148 331304 83154 331316
rect 84102 331304 84108 331316
rect 84160 331304 84166 331356
rect 88978 331304 88984 331356
rect 89036 331344 89042 331356
rect 89622 331344 89628 331356
rect 89036 331316 89628 331344
rect 89036 331304 89042 331316
rect 89622 331304 89628 331316
rect 89680 331304 89686 331356
rect 97074 331304 97080 331356
rect 97132 331344 97138 331356
rect 97902 331344 97908 331356
rect 97132 331316 97908 331344
rect 97132 331304 97138 331316
rect 97902 331304 97908 331316
rect 97960 331304 97966 331356
rect 118970 331304 118976 331356
rect 119028 331344 119034 331356
rect 119890 331344 119896 331356
rect 119028 331316 119896 331344
rect 119028 331304 119034 331316
rect 119890 331304 119896 331316
rect 119948 331304 119954 331356
rect 119982 331304 119988 331356
rect 120040 331344 120046 331356
rect 120534 331344 120540 331356
rect 120040 331316 120540 331344
rect 120040 331304 120046 331316
rect 120534 331304 120540 331316
rect 120592 331304 120598 331356
rect 132770 331304 132776 331356
rect 132828 331344 132834 331356
rect 133782 331344 133788 331356
rect 132828 331316 133788 331344
rect 132828 331304 132834 331316
rect 133782 331304 133788 331316
rect 133840 331304 133846 331356
rect 150342 331304 150348 331356
rect 150400 331344 150406 331356
rect 158070 331344 158076 331356
rect 150400 331316 158076 331344
rect 150400 331304 150406 331316
rect 158070 331304 158076 331316
rect 158128 331304 158134 331356
rect 50982 331236 50988 331288
rect 51040 331276 51046 331288
rect 69382 331276 69388 331288
rect 51040 331248 69388 331276
rect 51040 331236 51046 331248
rect 69382 331236 69388 331248
rect 69440 331236 69446 331288
rect 151170 331236 151176 331288
rect 151228 331276 151234 331288
rect 187142 331276 187148 331288
rect 151228 331248 187148 331276
rect 151228 331236 151234 331248
rect 187142 331236 187148 331248
rect 187200 331236 187206 331288
rect 184290 331100 184296 331152
rect 184348 331140 184354 331152
rect 188338 331140 188344 331152
rect 184348 331112 188344 331140
rect 184348 331100 184354 331112
rect 188338 331100 188344 331112
rect 188396 331100 188402 331152
rect 204898 330624 204904 330676
rect 204956 330664 204962 330676
rect 224218 330664 224224 330676
rect 204956 330636 224224 330664
rect 204956 330624 204962 330636
rect 224218 330624 224224 330636
rect 224276 330624 224282 330676
rect 175918 330556 175924 330608
rect 175976 330596 175982 330608
rect 209314 330596 209320 330608
rect 175976 330568 209320 330596
rect 175976 330556 175982 330568
rect 209314 330556 209320 330568
rect 209372 330556 209378 330608
rect 289078 330556 289084 330608
rect 289136 330596 289142 330608
rect 355410 330596 355416 330608
rect 289136 330568 355416 330596
rect 289136 330556 289142 330568
rect 355410 330556 355416 330568
rect 355468 330556 355474 330608
rect 67266 330488 67272 330540
rect 67324 330528 67330 330540
rect 73798 330528 73804 330540
rect 67324 330500 73804 330528
rect 67324 330488 67330 330500
rect 73798 330488 73804 330500
rect 73856 330488 73862 330540
rect 131758 330488 131764 330540
rect 131816 330528 131822 330540
rect 184474 330528 184480 330540
rect 131816 330500 184480 330528
rect 131816 330488 131822 330500
rect 184474 330488 184480 330500
rect 184532 330488 184538 330540
rect 209222 330488 209228 330540
rect 209280 330528 209286 330540
rect 306374 330528 306380 330540
rect 209280 330500 306380 330528
rect 209280 330488 209286 330500
rect 306374 330488 306380 330500
rect 306432 330488 306438 330540
rect 67726 329808 67732 329860
rect 67784 329848 67790 329860
rect 77294 329848 77300 329860
rect 67784 329820 77300 329848
rect 67784 329808 67790 329820
rect 77294 329808 77300 329820
rect 77352 329848 77358 329860
rect 162210 329848 162216 329860
rect 77352 329820 113174 329848
rect 77352 329808 77358 329820
rect 113146 329780 113174 329820
rect 126072 329820 162216 329848
rect 126072 329780 126100 329820
rect 162210 329808 162216 329820
rect 162268 329808 162274 329860
rect 113146 329752 126100 329780
rect 174538 329740 174544 329792
rect 174596 329780 174602 329792
rect 180334 329780 180340 329792
rect 174596 329752 180340 329780
rect 174596 329740 174602 329752
rect 180334 329740 180340 329752
rect 180392 329740 180398 329792
rect 114554 329672 114560 329724
rect 114612 329712 114618 329724
rect 115704 329712 115710 329724
rect 114612 329684 115710 329712
rect 114612 329672 114618 329684
rect 115704 329672 115710 329684
rect 115762 329672 115768 329724
rect 154114 329128 154120 329180
rect 154172 329168 154178 329180
rect 157242 329168 157248 329180
rect 154172 329140 157248 329168
rect 154172 329128 154178 329140
rect 157242 329128 157248 329140
rect 157300 329128 157306 329180
rect 169846 329128 169852 329180
rect 169904 329168 169910 329180
rect 174538 329168 174544 329180
rect 169904 329140 174544 329168
rect 169904 329128 169910 329140
rect 174538 329128 174544 329140
rect 174596 329128 174602 329180
rect 32398 329060 32404 329112
rect 32456 329100 32462 329112
rect 47578 329100 47584 329112
rect 32456 329072 47584 329100
rect 32456 329060 32462 329072
rect 47578 329060 47584 329072
rect 47636 329060 47642 329112
rect 114554 329100 114560 329112
rect 103486 329072 114560 329100
rect 59078 328516 59084 328568
rect 59136 328556 59142 328568
rect 66622 328556 66628 328568
rect 59136 328528 66628 328556
rect 59136 328516 59142 328528
rect 66622 328516 66628 328528
rect 66680 328516 66686 328568
rect 7558 328448 7564 328500
rect 7616 328488 7622 328500
rect 103486 328488 103514 329072
rect 114554 329060 114560 329072
rect 114612 329060 114618 329112
rect 136450 329060 136456 329112
rect 136508 329060 136514 329112
rect 139302 329060 139308 329112
rect 139360 329100 139366 329112
rect 139360 329072 142154 329100
rect 139360 329060 139366 329072
rect 7616 328460 103514 328488
rect 7616 328448 7622 328460
rect 136468 328420 136496 329060
rect 142126 328624 142154 329072
rect 156322 329060 156328 329112
rect 156380 329100 156386 329112
rect 156380 329072 156736 329100
rect 156380 329060 156386 329072
rect 156708 328840 156736 329072
rect 172698 329060 172704 329112
rect 172756 329100 172762 329112
rect 231210 329100 231216 329112
rect 172756 329072 231216 329100
rect 172756 329060 172762 329072
rect 231210 329060 231216 329072
rect 231268 329060 231274 329112
rect 253290 329060 253296 329112
rect 253348 329100 253354 329112
rect 317414 329100 317420 329112
rect 253348 329072 317420 329100
rect 253348 329060 253354 329072
rect 317414 329060 317420 329072
rect 317472 329060 317478 329112
rect 186222 328924 186228 328976
rect 186280 328964 186286 328976
rect 192570 328964 192576 328976
rect 186280 328936 192576 328964
rect 186280 328924 186286 328936
rect 192570 328924 192576 328936
rect 192628 328924 192634 328976
rect 156690 328788 156696 328840
rect 156748 328788 156754 328840
rect 158162 328624 158168 328636
rect 142126 328596 158168 328624
rect 158162 328584 158168 328596
rect 158220 328584 158226 328636
rect 158898 328516 158904 328568
rect 158956 328556 158962 328568
rect 172514 328556 172520 328568
rect 158956 328528 172520 328556
rect 158956 328516 158962 328528
rect 172514 328516 172520 328528
rect 172572 328516 172578 328568
rect 156782 328448 156788 328500
rect 156840 328488 156846 328500
rect 170398 328488 170404 328500
rect 156840 328460 170404 328488
rect 156840 328448 156846 328460
rect 170398 328448 170404 328460
rect 170456 328448 170462 328500
rect 136468 328392 142154 328420
rect 142126 327740 142154 328392
rect 180150 327768 180156 327820
rect 180208 327808 180214 327820
rect 209222 327808 209228 327820
rect 180208 327780 209228 327808
rect 180208 327768 180214 327780
rect 209222 327768 209228 327780
rect 209280 327768 209286 327820
rect 222930 327768 222936 327820
rect 222988 327808 222994 327820
rect 263594 327808 263600 327820
rect 222988 327780 263600 327808
rect 222988 327768 222994 327780
rect 263594 327768 263600 327780
rect 263652 327768 263658 327820
rect 236730 327740 236736 327752
rect 142126 327712 236736 327740
rect 236730 327700 236736 327712
rect 236788 327700 236794 327752
rect 57790 327088 57796 327140
rect 57848 327128 57854 327140
rect 169846 327128 169852 327140
rect 57848 327100 169852 327128
rect 57848 327088 57854 327100
rect 169846 327088 169852 327100
rect 169904 327088 169910 327140
rect 162302 327020 162308 327072
rect 162360 327060 162366 327072
rect 170490 327060 170496 327072
rect 162360 327032 170496 327060
rect 162360 327020 162366 327032
rect 170490 327020 170496 327032
rect 170548 327020 170554 327072
rect 178034 326408 178040 326460
rect 178092 326448 178098 326460
rect 245010 326448 245016 326460
rect 178092 326420 245016 326448
rect 178092 326408 178098 326420
rect 245010 326408 245016 326420
rect 245068 326408 245074 326460
rect 185578 326340 185584 326392
rect 185636 326380 185642 326392
rect 204898 326380 204904 326392
rect 185636 326352 204904 326380
rect 185636 326340 185642 326352
rect 204898 326340 204904 326352
rect 204956 326340 204962 326392
rect 215938 326340 215944 326392
rect 215996 326380 216002 326392
rect 348418 326380 348424 326392
rect 215996 326352 348424 326380
rect 215996 326340 216002 326352
rect 348418 326340 348424 326352
rect 348476 326340 348482 326392
rect 158990 325660 158996 325712
rect 159048 325700 159054 325712
rect 181622 325700 181628 325712
rect 159048 325672 181628 325700
rect 159048 325660 159054 325672
rect 181622 325660 181628 325672
rect 181680 325660 181686 325712
rect 159082 325592 159088 325644
rect 159140 325632 159146 325644
rect 167086 325632 167092 325644
rect 159140 325604 167092 325632
rect 159140 325592 159146 325604
rect 167086 325592 167092 325604
rect 167144 325592 167150 325644
rect 177390 324980 177396 325032
rect 177448 325020 177454 325032
rect 187234 325020 187240 325032
rect 177448 324992 187240 325020
rect 177448 324980 177454 324992
rect 187234 324980 187240 324992
rect 187292 324980 187298 325032
rect 195238 324980 195244 325032
rect 195296 325020 195302 325032
rect 235902 325020 235908 325032
rect 195296 324992 235908 325020
rect 195296 324980 195302 324992
rect 235902 324980 235908 324992
rect 235960 325020 235966 325032
rect 295978 325020 295984 325032
rect 235960 324992 295984 325020
rect 235960 324980 235966 324992
rect 295978 324980 295984 324992
rect 296036 324980 296042 325032
rect 170398 324912 170404 324964
rect 170456 324952 170462 324964
rect 236638 324952 236644 324964
rect 170456 324924 236644 324952
rect 170456 324912 170462 324924
rect 236638 324912 236644 324924
rect 236696 324912 236702 324964
rect 158714 324368 158720 324420
rect 158772 324408 158778 324420
rect 159082 324408 159088 324420
rect 158772 324380 159088 324408
rect 158772 324368 158778 324380
rect 159082 324368 159088 324380
rect 159140 324368 159146 324420
rect 167086 324300 167092 324352
rect 167144 324340 167150 324352
rect 171870 324340 171876 324352
rect 167144 324312 171876 324340
rect 167144 324300 167150 324312
rect 171870 324300 171876 324312
rect 171928 324300 171934 324352
rect 158714 324232 158720 324284
rect 158772 324272 158778 324284
rect 178770 324272 178776 324284
rect 158772 324244 178776 324272
rect 158772 324232 158778 324244
rect 178770 324232 178776 324244
rect 178828 324232 178834 324284
rect 220078 323552 220084 323604
rect 220136 323592 220142 323604
rect 251358 323592 251364 323604
rect 220136 323564 251364 323592
rect 220136 323552 220142 323564
rect 251358 323552 251364 323564
rect 251416 323552 251422 323604
rect 305730 323552 305736 323604
rect 305788 323592 305794 323604
rect 335998 323592 336004 323604
rect 305788 323564 336004 323592
rect 305788 323552 305794 323564
rect 335998 323552 336004 323564
rect 336056 323552 336062 323604
rect 158898 322940 158904 322992
rect 158956 322980 158962 322992
rect 243722 322980 243728 322992
rect 158956 322952 243728 322980
rect 158956 322940 158962 322952
rect 243722 322940 243728 322952
rect 243780 322940 243786 322992
rect 158990 322328 158996 322380
rect 159048 322368 159054 322380
rect 258166 322368 258172 322380
rect 159048 322340 258172 322368
rect 159048 322328 159054 322340
rect 258166 322328 258172 322340
rect 258224 322328 258230 322380
rect 158714 322260 158720 322312
rect 158772 322300 158778 322312
rect 162946 322300 162952 322312
rect 158772 322272 162952 322300
rect 158772 322260 158778 322272
rect 162946 322260 162952 322272
rect 163004 322300 163010 322312
rect 185578 322300 185584 322312
rect 163004 322272 185584 322300
rect 163004 322260 163010 322272
rect 185578 322260 185584 322272
rect 185636 322260 185642 322312
rect 251818 322192 251824 322244
rect 251876 322232 251882 322244
rect 260926 322232 260932 322244
rect 251876 322204 260932 322232
rect 251876 322192 251882 322204
rect 260926 322192 260932 322204
rect 260984 322232 260990 322244
rect 344278 322232 344284 322244
rect 260984 322204 344284 322232
rect 260984 322192 260990 322204
rect 344278 322192 344284 322204
rect 344336 322192 344342 322244
rect 3510 321512 3516 321564
rect 3568 321552 3574 321564
rect 66898 321552 66904 321564
rect 3568 321524 66904 321552
rect 3568 321512 3574 321524
rect 66898 321512 66904 321524
rect 66956 321512 66962 321564
rect 176102 320900 176108 320952
rect 176160 320940 176166 320952
rect 193858 320940 193864 320952
rect 176160 320912 193864 320940
rect 176160 320900 176166 320912
rect 193858 320900 193864 320912
rect 193916 320900 193922 320952
rect 156690 320832 156696 320884
rect 156748 320872 156754 320884
rect 169294 320872 169300 320884
rect 156748 320844 169300 320872
rect 156748 320832 156754 320844
rect 169294 320832 169300 320844
rect 169352 320832 169358 320884
rect 178034 320832 178040 320884
rect 178092 320872 178098 320884
rect 237374 320872 237380 320884
rect 178092 320844 237380 320872
rect 178092 320832 178098 320844
rect 237374 320832 237380 320844
rect 237432 320832 237438 320884
rect 281442 320832 281448 320884
rect 281500 320872 281506 320884
rect 331950 320872 331956 320884
rect 281500 320844 331956 320872
rect 281500 320832 281506 320844
rect 331950 320832 331956 320844
rect 332008 320832 332014 320884
rect 55122 320152 55128 320204
rect 55180 320192 55186 320204
rect 66806 320192 66812 320204
rect 55180 320164 66812 320192
rect 55180 320152 55186 320164
rect 66806 320152 66812 320164
rect 66864 320152 66870 320204
rect 237374 320152 237380 320204
rect 237432 320192 237438 320204
rect 238018 320192 238024 320204
rect 237432 320164 238024 320192
rect 237432 320152 237438 320164
rect 238018 320152 238024 320164
rect 238076 320192 238082 320204
rect 281442 320192 281448 320204
rect 238076 320164 281448 320192
rect 238076 320152 238082 320164
rect 281442 320152 281448 320164
rect 281500 320152 281506 320204
rect 159266 319472 159272 319524
rect 159324 319512 159330 319524
rect 159910 319512 159916 319524
rect 159324 319484 159916 319512
rect 159324 319472 159330 319484
rect 159910 319472 159916 319484
rect 159968 319512 159974 319524
rect 169110 319512 169116 319524
rect 159968 319484 169116 319512
rect 159968 319472 159974 319484
rect 169110 319472 169116 319484
rect 169168 319472 169174 319524
rect 174538 319472 174544 319524
rect 174596 319512 174602 319524
rect 195238 319512 195244 319524
rect 174596 319484 195244 319512
rect 174596 319472 174602 319484
rect 195238 319472 195244 319484
rect 195296 319472 195302 319524
rect 231118 319472 231124 319524
rect 231176 319512 231182 319524
rect 267826 319512 267832 319524
rect 231176 319484 267832 319512
rect 231176 319472 231182 319484
rect 267826 319472 267832 319484
rect 267884 319472 267890 319524
rect 4062 319404 4068 319456
rect 4120 319444 4126 319456
rect 11698 319444 11704 319456
rect 4120 319416 11704 319444
rect 4120 319404 4126 319416
rect 11698 319404 11704 319416
rect 11756 319404 11762 319456
rect 163498 319404 163504 319456
rect 163556 319444 163562 319456
rect 247126 319444 247132 319456
rect 163556 319416 247132 319444
rect 163556 319404 163562 319416
rect 247126 319404 247132 319416
rect 247184 319404 247190 319456
rect 281350 319404 281356 319456
rect 281408 319444 281414 319456
rect 355318 319444 355324 319456
rect 281408 319416 355324 319444
rect 281408 319404 281414 319416
rect 355318 319404 355324 319416
rect 355376 319404 355382 319456
rect 55858 318832 55864 318844
rect 55186 318804 55864 318832
rect 34422 318724 34428 318776
rect 34480 318764 34486 318776
rect 55186 318764 55214 318804
rect 55858 318792 55864 318804
rect 55916 318832 55922 318844
rect 66898 318832 66904 318844
rect 55916 318804 66904 318832
rect 55916 318792 55922 318804
rect 66898 318792 66904 318804
rect 66956 318792 66962 318844
rect 34480 318736 55214 318764
rect 34480 318724 34486 318736
rect 236730 318724 236736 318776
rect 236788 318764 236794 318776
rect 237282 318764 237288 318776
rect 236788 318736 237288 318764
rect 236788 318724 236794 318736
rect 237282 318724 237288 318736
rect 237340 318724 237346 318776
rect 64690 318112 64696 318164
rect 64748 318152 64754 318164
rect 66806 318152 66812 318164
rect 64748 318124 66812 318152
rect 64748 318112 64754 318124
rect 66806 318112 66812 318124
rect 66864 318112 66870 318164
rect 189074 318112 189080 318164
rect 189132 318152 189138 318164
rect 246114 318152 246120 318164
rect 189132 318124 246120 318152
rect 189132 318112 189138 318124
rect 246114 318112 246120 318124
rect 246172 318112 246178 318164
rect 156874 318044 156880 318096
rect 156932 318084 156938 318096
rect 233878 318084 233884 318096
rect 156932 318056 233884 318084
rect 156932 318044 156938 318056
rect 233878 318044 233884 318056
rect 233936 318044 233942 318096
rect 298002 318044 298008 318096
rect 298060 318084 298066 318096
rect 345658 318084 345664 318096
rect 298060 318056 345664 318084
rect 298060 318044 298066 318056
rect 345658 318044 345664 318056
rect 345716 318044 345722 318096
rect 158714 317568 158720 317620
rect 158772 317608 158778 317620
rect 163590 317608 163596 317620
rect 158772 317580 163596 317608
rect 158772 317568 158778 317580
rect 163590 317568 163596 317580
rect 163648 317568 163654 317620
rect 50798 317432 50804 317484
rect 50856 317472 50862 317484
rect 52270 317472 52276 317484
rect 50856 317444 52276 317472
rect 50856 317432 50862 317444
rect 52270 317432 52276 317444
rect 52328 317432 52334 317484
rect 237282 317432 237288 317484
rect 237340 317472 237346 317484
rect 296898 317472 296904 317484
rect 237340 317444 296904 317472
rect 237340 317432 237346 317444
rect 296898 317432 296904 317444
rect 296956 317472 296962 317484
rect 298002 317472 298008 317484
rect 296956 317444 298008 317472
rect 296956 317432 296962 317444
rect 298002 317432 298008 317444
rect 298060 317432 298066 317484
rect 158714 317364 158720 317416
rect 158772 317404 158778 317416
rect 159082 317404 159088 317416
rect 158772 317376 159088 317404
rect 158772 317364 158778 317376
rect 159082 317364 159088 317376
rect 159140 317404 159146 317416
rect 169202 317404 169208 317416
rect 159140 317376 169208 317404
rect 159140 317364 159146 317376
rect 169202 317364 169208 317376
rect 169260 317364 169266 317416
rect 177482 316752 177488 316804
rect 177540 316792 177546 316804
rect 258258 316792 258264 316804
rect 177540 316764 258264 316792
rect 177540 316752 177546 316764
rect 258258 316752 258264 316764
rect 258316 316752 258322 316804
rect 15838 316684 15844 316736
rect 15896 316724 15902 316736
rect 67358 316724 67364 316736
rect 15896 316696 67364 316724
rect 15896 316684 15902 316696
rect 67358 316684 67364 316696
rect 67416 316684 67422 316736
rect 199470 316684 199476 316736
rect 199528 316724 199534 316736
rect 352650 316724 352656 316736
rect 199528 316696 352656 316724
rect 199528 316684 199534 316696
rect 352650 316684 352656 316696
rect 352708 316684 352714 316736
rect 199378 315324 199384 315376
rect 199436 315364 199442 315376
rect 220078 315364 220084 315376
rect 199436 315336 220084 315364
rect 199436 315324 199442 315336
rect 220078 315324 220084 315336
rect 220136 315324 220142 315376
rect 181622 315256 181628 315308
rect 181680 315296 181686 315308
rect 210418 315296 210424 315308
rect 181680 315268 210424 315296
rect 181680 315256 181686 315268
rect 210418 315256 210424 315268
rect 210476 315256 210482 315308
rect 210510 315256 210516 315308
rect 210568 315296 210574 315308
rect 240778 315296 240784 315308
rect 210568 315268 240784 315296
rect 210568 315256 210574 315268
rect 240778 315256 240784 315268
rect 240836 315256 240842 315308
rect 321554 315256 321560 315308
rect 321612 315296 321618 315308
rect 357434 315296 357440 315308
rect 321612 315268 357440 315296
rect 321612 315256 321618 315268
rect 357434 315256 357440 315268
rect 357492 315256 357498 315308
rect 251818 314644 251824 314696
rect 251876 314684 251882 314696
rect 321554 314684 321560 314696
rect 251876 314656 321560 314684
rect 251876 314644 251882 314656
rect 321554 314644 321560 314656
rect 321612 314644 321618 314696
rect 58894 314576 58900 314628
rect 58952 314616 58958 314628
rect 66806 314616 66812 314628
rect 58952 314588 66812 314616
rect 58952 314576 58958 314588
rect 66806 314576 66812 314588
rect 66864 314576 66870 314628
rect 184382 313964 184388 314016
rect 184440 314004 184446 314016
rect 238110 314004 238116 314016
rect 184440 313976 238116 314004
rect 184440 313964 184446 313976
rect 238110 313964 238116 313976
rect 238168 313964 238174 314016
rect 228450 313896 228456 313948
rect 228508 313936 228514 313948
rect 380986 313936 380992 313948
rect 228508 313908 380992 313936
rect 228508 313896 228514 313908
rect 380986 313896 380992 313908
rect 381044 313896 381050 313948
rect 158714 313352 158720 313404
rect 158772 313392 158778 313404
rect 163498 313392 163504 313404
rect 158772 313364 163504 313392
rect 158772 313352 158778 313364
rect 163498 313352 163504 313364
rect 163556 313352 163562 313404
rect 61838 313216 61844 313268
rect 61896 313256 61902 313268
rect 66438 313256 66444 313268
rect 61896 313228 66444 313256
rect 61896 313216 61902 313228
rect 66438 313216 66444 313228
rect 66496 313216 66502 313268
rect 206462 313216 206468 313268
rect 206520 313256 206526 313268
rect 209866 313256 209872 313268
rect 206520 313228 209872 313256
rect 206520 313216 206526 313228
rect 209866 313216 209872 313228
rect 209924 313216 209930 313268
rect 166442 312604 166448 312656
rect 166500 312644 166506 312656
rect 200758 312644 200764 312656
rect 166500 312616 200764 312644
rect 166500 312604 166506 312616
rect 200758 312604 200764 312616
rect 200816 312604 200822 312656
rect 185578 312536 185584 312588
rect 185636 312576 185642 312588
rect 225966 312576 225972 312588
rect 185636 312548 225972 312576
rect 185636 312536 185642 312548
rect 225966 312536 225972 312548
rect 226024 312536 226030 312588
rect 227070 312536 227076 312588
rect 227128 312576 227134 312588
rect 253934 312576 253940 312588
rect 227128 312548 253940 312576
rect 227128 312536 227134 312548
rect 253934 312536 253940 312548
rect 253992 312536 253998 312588
rect 160830 311856 160836 311908
rect 160888 311896 160894 311908
rect 166258 311896 166264 311908
rect 160888 311868 166264 311896
rect 160888 311856 160894 311868
rect 166258 311856 166264 311868
rect 166316 311856 166322 311908
rect 224402 311856 224408 311908
rect 224460 311896 224466 311908
rect 224862 311896 224868 311908
rect 224460 311868 224868 311896
rect 224460 311856 224466 311868
rect 224862 311856 224868 311868
rect 224920 311896 224926 311908
rect 260834 311896 260840 311908
rect 224920 311868 260840 311896
rect 224920 311856 224926 311868
rect 260834 311856 260840 311868
rect 260892 311856 260898 311908
rect 161382 311788 161388 311840
rect 161440 311828 161446 311840
rect 162854 311828 162860 311840
rect 161440 311800 162860 311828
rect 161440 311788 161446 311800
rect 162854 311788 162860 311800
rect 162912 311788 162918 311840
rect 244918 311788 244924 311840
rect 244976 311828 244982 311840
rect 248414 311828 248420 311840
rect 244976 311800 248420 311828
rect 244976 311788 244982 311800
rect 248414 311788 248420 311800
rect 248472 311788 248478 311840
rect 170490 311176 170496 311228
rect 170548 311216 170554 311228
rect 222930 311216 222936 311228
rect 170548 311188 222936 311216
rect 170548 311176 170554 311188
rect 222930 311176 222936 311188
rect 222988 311176 222994 311228
rect 18598 311108 18604 311160
rect 18656 311148 18662 311160
rect 67450 311148 67456 311160
rect 18656 311120 67456 311148
rect 18656 311108 18662 311120
rect 67450 311108 67456 311120
rect 67508 311108 67514 311160
rect 169294 311108 169300 311160
rect 169352 311148 169358 311160
rect 192478 311148 192484 311160
rect 169352 311120 192484 311148
rect 169352 311108 169358 311120
rect 192478 311108 192484 311120
rect 192536 311108 192542 311160
rect 202230 311108 202236 311160
rect 202288 311148 202294 311160
rect 207014 311148 207020 311160
rect 202288 311120 207020 311148
rect 202288 311108 202294 311120
rect 207014 311108 207020 311120
rect 207072 311148 207078 311160
rect 287054 311148 287060 311160
rect 207072 311120 287060 311148
rect 207072 311108 207078 311120
rect 287054 311108 287060 311120
rect 287112 311108 287118 311160
rect 158714 310496 158720 310548
rect 158772 310536 158778 310548
rect 170398 310536 170404 310548
rect 158772 310508 170404 310536
rect 158772 310496 158778 310508
rect 170398 310496 170404 310508
rect 170456 310496 170462 310548
rect 184474 310428 184480 310480
rect 184532 310468 184538 310480
rect 226426 310468 226432 310480
rect 184532 310440 226432 310468
rect 184532 310428 184538 310440
rect 226426 310428 226432 310440
rect 226484 310428 226490 310480
rect 36538 309748 36544 309800
rect 36596 309788 36602 309800
rect 63402 309788 63408 309800
rect 36596 309760 63408 309788
rect 36596 309748 36602 309760
rect 63402 309748 63408 309760
rect 63460 309788 63466 309800
rect 66806 309788 66812 309800
rect 63460 309760 66812 309788
rect 63460 309748 63466 309760
rect 66806 309748 66812 309760
rect 66864 309748 66870 309800
rect 158806 309748 158812 309800
rect 158864 309788 158870 309800
rect 174630 309788 174636 309800
rect 158864 309760 174636 309788
rect 158864 309748 158870 309760
rect 174630 309748 174636 309760
rect 174688 309748 174694 309800
rect 317322 309748 317328 309800
rect 317380 309788 317386 309800
rect 338942 309788 338948 309800
rect 317380 309760 338948 309788
rect 317380 309748 317386 309760
rect 338942 309748 338948 309760
rect 339000 309748 339006 309800
rect 177482 309136 177488 309188
rect 177540 309176 177546 309188
rect 218146 309176 218152 309188
rect 177540 309148 218152 309176
rect 177540 309136 177546 309148
rect 218146 309136 218152 309148
rect 218204 309136 218210 309188
rect 239490 309136 239496 309188
rect 239548 309176 239554 309188
rect 316126 309176 316132 309188
rect 239548 309148 316132 309176
rect 239548 309136 239554 309148
rect 316126 309136 316132 309148
rect 316184 309176 316190 309188
rect 317322 309176 317328 309188
rect 316184 309148 317328 309176
rect 316184 309136 316190 309148
rect 317322 309136 317328 309148
rect 317380 309136 317386 309188
rect 158714 308456 158720 308508
rect 158772 308496 158778 308508
rect 165614 308496 165620 308508
rect 158772 308468 165620 308496
rect 158772 308456 158778 308468
rect 165614 308456 165620 308468
rect 165672 308456 165678 308508
rect 202138 308456 202144 308508
rect 202196 308496 202202 308508
rect 231118 308496 231124 308508
rect 202196 308468 231124 308496
rect 202196 308456 202202 308468
rect 231118 308456 231124 308468
rect 231176 308456 231182 308508
rect 232498 308456 232504 308508
rect 232556 308496 232562 308508
rect 259638 308496 259644 308508
rect 232556 308468 259644 308496
rect 232556 308456 232562 308468
rect 259638 308456 259644 308468
rect 259696 308456 259702 308508
rect 157978 308388 157984 308440
rect 158036 308428 158042 308440
rect 240870 308428 240876 308440
rect 158036 308400 240876 308428
rect 158036 308388 158042 308400
rect 240870 308388 240876 308400
rect 240928 308388 240934 308440
rect 57606 307708 57612 307760
rect 57664 307748 57670 307760
rect 66898 307748 66904 307760
rect 57664 307720 66904 307748
rect 57664 307708 57670 307720
rect 66898 307708 66904 307720
rect 66956 307708 66962 307760
rect 231210 307708 231216 307760
rect 231268 307748 231274 307760
rect 232222 307748 232228 307760
rect 231268 307720 232228 307748
rect 231268 307708 231274 307720
rect 232222 307708 232228 307720
rect 232280 307708 232286 307760
rect 232222 307096 232228 307148
rect 232280 307136 232286 307148
rect 281350 307136 281356 307148
rect 232280 307108 281356 307136
rect 232280 307096 232286 307108
rect 281350 307096 281356 307108
rect 281408 307096 281414 307148
rect 189718 307028 189724 307080
rect 189776 307068 189782 307080
rect 197170 307068 197176 307080
rect 189776 307040 197176 307068
rect 189776 307028 189782 307040
rect 197170 307028 197176 307040
rect 197228 307028 197234 307080
rect 262858 307028 262864 307080
rect 262916 307068 262922 307080
rect 322290 307068 322296 307080
rect 262916 307040 322296 307068
rect 262916 307028 262922 307040
rect 322290 307028 322296 307040
rect 322348 307028 322354 307080
rect 158714 306348 158720 306400
rect 158772 306388 158778 306400
rect 167638 306388 167644 306400
rect 158772 306360 167644 306388
rect 158772 306348 158778 306360
rect 167638 306348 167644 306360
rect 167696 306348 167702 306400
rect 169110 306348 169116 306400
rect 169168 306388 169174 306400
rect 252738 306388 252744 306400
rect 169168 306360 252744 306388
rect 169168 306348 169174 306360
rect 252738 306348 252744 306360
rect 252796 306348 252802 306400
rect 3510 306280 3516 306332
rect 3568 306320 3574 306332
rect 32398 306320 32404 306332
rect 3568 306292 32404 306320
rect 3568 306280 3574 306292
rect 32398 306280 32404 306292
rect 32456 306280 32462 306332
rect 61930 306280 61936 306332
rect 61988 306320 61994 306332
rect 66806 306320 66812 306332
rect 61988 306292 66812 306320
rect 61988 306280 61994 306292
rect 66806 306280 66812 306292
rect 66864 306280 66870 306332
rect 233878 305940 233884 305992
rect 233936 305980 233942 305992
rect 234246 305980 234252 305992
rect 233936 305952 234252 305980
rect 233936 305940 233942 305952
rect 234246 305940 234252 305952
rect 234304 305940 234310 305992
rect 158714 305056 158720 305108
rect 158772 305096 158778 305108
rect 231210 305096 231216 305108
rect 158772 305068 231216 305096
rect 158772 305056 158778 305068
rect 231210 305056 231216 305068
rect 231268 305056 231274 305108
rect 234246 305056 234252 305108
rect 234304 305096 234310 305108
rect 274634 305096 274640 305108
rect 234304 305068 274640 305096
rect 234304 305056 234310 305068
rect 274634 305056 274640 305068
rect 274692 305056 274698 305108
rect 165062 304988 165068 305040
rect 165120 305028 165126 305040
rect 165522 305028 165528 305040
rect 165120 305000 165528 305028
rect 165120 304988 165126 305000
rect 165522 304988 165528 305000
rect 165580 305028 165586 305040
rect 262306 305028 262312 305040
rect 165580 305000 262312 305028
rect 165580 304988 165586 305000
rect 262306 304988 262312 305000
rect 262364 304988 262370 305040
rect 63218 304920 63224 304972
rect 63276 304960 63282 304972
rect 66806 304960 66812 304972
rect 63276 304932 66812 304960
rect 63276 304920 63282 304932
rect 66806 304920 66812 304932
rect 66864 304920 66870 304972
rect 158806 304920 158812 304972
rect 158864 304960 158870 304972
rect 168190 304960 168196 304972
rect 158864 304932 168196 304960
rect 158864 304920 158870 304932
rect 168190 304920 168196 304932
rect 168248 304920 168254 304972
rect 168190 304240 168196 304292
rect 168248 304280 168254 304292
rect 175918 304280 175924 304292
rect 168248 304252 175924 304280
rect 168248 304240 168254 304252
rect 175918 304240 175924 304252
rect 175976 304240 175982 304292
rect 182082 304240 182088 304292
rect 182140 304280 182146 304292
rect 206370 304280 206376 304292
rect 182140 304252 206376 304280
rect 182140 304240 182146 304252
rect 206370 304240 206376 304252
rect 206428 304240 206434 304292
rect 206646 303696 206652 303748
rect 206704 303736 206710 303748
rect 282270 303736 282276 303748
rect 206704 303708 282276 303736
rect 206704 303696 206710 303708
rect 282270 303696 282276 303708
rect 282328 303696 282334 303748
rect 211798 303628 211804 303680
rect 211856 303668 211862 303680
rect 304994 303668 305000 303680
rect 211856 303640 305000 303668
rect 211856 303628 211862 303640
rect 304994 303628 305000 303640
rect 305052 303628 305058 303680
rect 165614 302880 165620 302932
rect 165672 302920 165678 302932
rect 180150 302920 180156 302932
rect 165672 302892 180156 302920
rect 165672 302880 165678 302892
rect 180150 302880 180156 302892
rect 180208 302880 180214 302932
rect 329098 302880 329104 302932
rect 329156 302920 329162 302932
rect 357434 302920 357440 302932
rect 329156 302892 357440 302920
rect 329156 302880 329162 302892
rect 357434 302880 357440 302892
rect 357492 302880 357498 302932
rect 184382 302268 184388 302320
rect 184440 302308 184446 302320
rect 209958 302308 209964 302320
rect 184440 302280 209964 302308
rect 184440 302268 184446 302280
rect 209958 302268 209964 302280
rect 210016 302308 210022 302320
rect 210510 302308 210516 302320
rect 210016 302280 210516 302308
rect 210016 302268 210022 302280
rect 210510 302268 210516 302280
rect 210568 302268 210574 302320
rect 229830 302268 229836 302320
rect 229888 302308 229894 302320
rect 270586 302308 270592 302320
rect 229888 302280 270592 302308
rect 229888 302268 229894 302280
rect 270586 302268 270592 302280
rect 270644 302268 270650 302320
rect 208486 302200 208492 302252
rect 208544 302240 208550 302252
rect 209314 302240 209320 302252
rect 208544 302212 209320 302240
rect 208544 302200 208550 302212
rect 209314 302200 209320 302212
rect 209372 302240 209378 302252
rect 269850 302240 269856 302252
rect 209372 302212 269856 302240
rect 209372 302200 209378 302212
rect 269850 302200 269856 302212
rect 269908 302200 269914 302252
rect 59262 302132 59268 302184
rect 59320 302172 59326 302184
rect 66898 302172 66904 302184
rect 59320 302144 66904 302172
rect 59320 302132 59326 302144
rect 66898 302132 66904 302144
rect 66956 302132 66962 302184
rect 194134 301520 194140 301572
rect 194192 301560 194198 301572
rect 203518 301560 203524 301572
rect 194192 301532 203524 301560
rect 194192 301520 194198 301532
rect 203518 301520 203524 301532
rect 203576 301520 203582 301572
rect 207658 301520 207664 301572
rect 207716 301560 207722 301572
rect 221642 301560 221648 301572
rect 207716 301532 221648 301560
rect 207716 301520 207722 301532
rect 221642 301520 221648 301532
rect 221700 301520 221706 301572
rect 158714 301452 158720 301504
rect 158772 301492 158778 301504
rect 244550 301492 244556 301504
rect 158772 301464 244556 301492
rect 158772 301452 158778 301464
rect 244550 301452 244556 301464
rect 244608 301452 244614 301504
rect 274634 301452 274640 301504
rect 274692 301492 274698 301504
rect 302418 301492 302424 301504
rect 274692 301464 302424 301492
rect 274692 301452 274698 301464
rect 302418 301452 302424 301464
rect 302476 301492 302482 301504
rect 340230 301492 340236 301504
rect 302476 301464 340236 301492
rect 302476 301452 302482 301464
rect 340230 301452 340236 301464
rect 340288 301452 340294 301504
rect 57606 300840 57612 300892
rect 57664 300880 57670 300892
rect 66806 300880 66812 300892
rect 57664 300852 66812 300880
rect 57664 300840 57670 300852
rect 66806 300840 66812 300852
rect 66864 300840 66870 300892
rect 233142 300772 233148 300824
rect 233200 300812 233206 300824
rect 233694 300812 233700 300824
rect 233200 300784 233700 300812
rect 233200 300772 233206 300784
rect 233694 300772 233700 300784
rect 233752 300772 233758 300824
rect 159634 300092 159640 300144
rect 159692 300132 159698 300144
rect 180242 300132 180248 300144
rect 159692 300104 180248 300132
rect 159692 300092 159698 300104
rect 180242 300092 180248 300104
rect 180300 300092 180306 300144
rect 215294 299616 215300 299668
rect 215352 299656 215358 299668
rect 216030 299656 216036 299668
rect 215352 299628 216036 299656
rect 215352 299616 215358 299628
rect 216030 299616 216036 299628
rect 216088 299656 216094 299668
rect 216088 299628 219434 299656
rect 216088 299616 216094 299628
rect 219406 299588 219434 299628
rect 256786 299588 256792 299600
rect 219406 299560 256792 299588
rect 256786 299548 256792 299560
rect 256844 299548 256850 299600
rect 197170 299480 197176 299532
rect 197228 299520 197234 299532
rect 231302 299520 231308 299532
rect 197228 299492 231308 299520
rect 197228 299480 197234 299492
rect 231302 299480 231308 299492
rect 231360 299480 231366 299532
rect 233694 299480 233700 299532
rect 233752 299520 233758 299532
rect 582466 299520 582472 299532
rect 233752 299492 582472 299520
rect 233752 299480 233758 299492
rect 582466 299480 582472 299492
rect 582524 299480 582530 299532
rect 195790 298800 195796 298852
rect 195848 298840 195854 298852
rect 204346 298840 204352 298852
rect 195848 298812 204352 298840
rect 195848 298800 195854 298812
rect 204346 298800 204352 298812
rect 204404 298800 204410 298852
rect 159634 298732 159640 298784
rect 159692 298772 159698 298784
rect 174538 298772 174544 298784
rect 159692 298744 174544 298772
rect 159692 298732 159698 298744
rect 174538 298732 174544 298744
rect 174596 298732 174602 298784
rect 180610 298732 180616 298784
rect 180668 298772 180674 298784
rect 201494 298772 201500 298784
rect 180668 298744 201500 298772
rect 180668 298732 180674 298744
rect 201494 298732 201500 298744
rect 201552 298732 201558 298784
rect 221550 298732 221556 298784
rect 221608 298772 221614 298784
rect 241422 298772 241428 298784
rect 221608 298744 241428 298772
rect 221608 298732 221614 298744
rect 241422 298732 241428 298744
rect 241480 298732 241486 298784
rect 243722 298732 243728 298784
rect 243780 298772 243786 298784
rect 251174 298772 251180 298784
rect 243780 298744 251180 298772
rect 243780 298732 243786 298744
rect 251174 298732 251180 298744
rect 251232 298732 251238 298784
rect 292574 298732 292580 298784
rect 292632 298772 292638 298784
rect 361574 298772 361580 298784
rect 292632 298744 361580 298772
rect 292632 298732 292638 298744
rect 361574 298732 361580 298744
rect 361632 298732 361638 298784
rect 59262 298120 59268 298172
rect 59320 298160 59326 298172
rect 66622 298160 66628 298172
rect 59320 298132 66628 298160
rect 59320 298120 59326 298132
rect 66622 298120 66628 298132
rect 66680 298120 66686 298172
rect 243630 298120 243636 298172
rect 243688 298160 243694 298172
rect 292574 298160 292580 298172
rect 243688 298132 292580 298160
rect 243688 298120 243694 298132
rect 292574 298120 292580 298132
rect 292632 298120 292638 298172
rect 50890 298052 50896 298104
rect 50948 298092 50954 298104
rect 66806 298092 66812 298104
rect 50948 298064 66812 298092
rect 50948 298052 50954 298064
rect 66806 298052 66812 298064
rect 66864 298052 66870 298104
rect 158714 298052 158720 298104
rect 158772 298092 158778 298104
rect 175274 298092 175280 298104
rect 158772 298064 175280 298092
rect 158772 298052 158778 298064
rect 175274 298052 175280 298064
rect 175332 298092 175338 298104
rect 175734 298092 175740 298104
rect 175332 298064 175740 298092
rect 175332 298052 175338 298064
rect 175734 298052 175740 298064
rect 175792 298052 175798 298104
rect 201402 298052 201408 298104
rect 201460 298092 201466 298104
rect 202782 298092 202788 298104
rect 201460 298064 202788 298092
rect 201460 298052 201466 298064
rect 202782 298052 202788 298064
rect 202840 298052 202846 298104
rect 158622 297372 158628 297424
rect 158680 297412 158686 297424
rect 171134 297412 171140 297424
rect 158680 297384 171140 297412
rect 158680 297372 158686 297384
rect 171134 297372 171140 297384
rect 171192 297372 171198 297424
rect 188982 297372 188988 297424
rect 189040 297412 189046 297424
rect 194042 297412 194048 297424
rect 189040 297384 194048 297412
rect 189040 297372 189046 297384
rect 194042 297372 194048 297384
rect 194100 297372 194106 297424
rect 253198 297372 253204 297424
rect 253256 297412 253262 297424
rect 259454 297412 259460 297424
rect 253256 297384 259460 297412
rect 253256 297372 253262 297384
rect 259454 297372 259460 297384
rect 259512 297372 259518 297424
rect 206278 296760 206284 296812
rect 206336 296800 206342 296812
rect 211430 296800 211436 296812
rect 206336 296772 211436 296800
rect 206336 296760 206342 296772
rect 211430 296760 211436 296772
rect 211488 296760 211494 296812
rect 198366 296692 198372 296744
rect 198424 296732 198430 296744
rect 282914 296732 282920 296744
rect 198424 296704 282920 296732
rect 198424 296692 198430 296704
rect 282914 296692 282920 296704
rect 282972 296692 282978 296744
rect 164878 295944 164884 295996
rect 164936 295984 164942 295996
rect 184382 295984 184388 295996
rect 164936 295956 184388 295984
rect 164936 295944 164942 295956
rect 184382 295944 184388 295956
rect 184440 295944 184446 295996
rect 208026 295944 208032 295996
rect 208084 295984 208090 295996
rect 226334 295984 226340 295996
rect 208084 295956 226340 295984
rect 208084 295944 208090 295956
rect 226334 295944 226340 295956
rect 226392 295944 226398 295996
rect 231302 295944 231308 295996
rect 231360 295984 231366 295996
rect 272518 295984 272524 295996
rect 231360 295956 272524 295984
rect 231360 295944 231366 295956
rect 272518 295944 272524 295956
rect 272576 295944 272582 295996
rect 40678 295332 40684 295384
rect 40736 295372 40742 295384
rect 67726 295372 67732 295384
rect 40736 295344 67732 295372
rect 40736 295332 40742 295344
rect 67726 295332 67732 295344
rect 67784 295332 67790 295384
rect 158714 295332 158720 295384
rect 158772 295372 158778 295384
rect 169846 295372 169852 295384
rect 158772 295344 169852 295372
rect 158772 295332 158778 295344
rect 169846 295332 169852 295344
rect 169904 295332 169910 295384
rect 191282 295332 191288 295384
rect 191340 295372 191346 295384
rect 211062 295372 211068 295384
rect 191340 295344 211068 295372
rect 191340 295332 191346 295344
rect 211062 295332 211068 295344
rect 211120 295332 211126 295384
rect 211430 295332 211436 295384
rect 211488 295372 211494 295384
rect 278130 295372 278136 295384
rect 211488 295344 278136 295372
rect 211488 295332 211494 295344
rect 278130 295332 278136 295344
rect 278188 295332 278194 295384
rect 57790 295264 57796 295316
rect 57848 295304 57854 295316
rect 66806 295304 66812 295316
rect 57848 295276 66812 295304
rect 57848 295264 57854 295276
rect 66806 295264 66812 295276
rect 66864 295264 66870 295316
rect 162210 294652 162216 294704
rect 162268 294692 162274 294704
rect 213822 294692 213828 294704
rect 162268 294664 213828 294692
rect 162268 294652 162274 294664
rect 213822 294652 213828 294664
rect 213880 294652 213886 294704
rect 224218 294652 224224 294704
rect 224276 294692 224282 294704
rect 227438 294692 227444 294704
rect 224276 294664 227444 294692
rect 224276 294652 224282 294664
rect 227438 294652 227444 294664
rect 227496 294652 227502 294704
rect 160830 294584 160836 294636
rect 160888 294624 160894 294636
rect 164234 294624 164240 294636
rect 160888 294596 164240 294624
rect 160888 294584 160894 294596
rect 164234 294584 164240 294596
rect 164292 294624 164298 294636
rect 253198 294624 253204 294636
rect 164292 294596 253204 294624
rect 164292 294584 164298 294596
rect 253198 294584 253204 294596
rect 253256 294584 253262 294636
rect 221458 293972 221464 294024
rect 221516 294012 221522 294024
rect 223942 294012 223948 294024
rect 221516 293984 223948 294012
rect 221516 293972 221522 293984
rect 223942 293972 223948 293984
rect 224000 293972 224006 294024
rect 241974 293972 241980 294024
rect 242032 294012 242038 294024
rect 242250 294012 242256 294024
rect 242032 293984 242256 294012
rect 242032 293972 242038 293984
rect 242250 293972 242256 293984
rect 242308 294012 242314 294024
rect 283006 294012 283012 294024
rect 242308 293984 283012 294012
rect 242308 293972 242314 293984
rect 283006 293972 283012 293984
rect 283064 293972 283070 294024
rect 14458 293904 14464 293956
rect 14516 293944 14522 293956
rect 52362 293944 52368 293956
rect 14516 293916 52368 293944
rect 14516 293904 14522 293916
rect 52362 293904 52368 293916
rect 52420 293944 52426 293956
rect 66806 293944 66812 293956
rect 52420 293916 66812 293944
rect 52420 293904 52426 293916
rect 66806 293904 66812 293916
rect 66864 293904 66870 293956
rect 219710 292680 219716 292732
rect 219768 292720 219774 292732
rect 280798 292720 280804 292732
rect 219768 292692 280804 292720
rect 219768 292680 219774 292692
rect 280798 292680 280804 292692
rect 280856 292680 280862 292732
rect 158714 292612 158720 292664
rect 158772 292652 158778 292664
rect 220170 292652 220176 292664
rect 158772 292624 220176 292652
rect 158772 292612 158778 292624
rect 220170 292612 220176 292624
rect 220228 292612 220234 292664
rect 3510 292544 3516 292596
rect 3568 292584 3574 292596
rect 14550 292584 14556 292596
rect 3568 292556 14556 292584
rect 3568 292544 3574 292556
rect 14550 292544 14556 292556
rect 14608 292544 14614 292596
rect 183094 292544 183100 292596
rect 183152 292584 183158 292596
rect 254578 292584 254584 292596
rect 183152 292556 254584 292584
rect 183152 292544 183158 292556
rect 254578 292544 254584 292556
rect 254636 292544 254642 292596
rect 54938 292476 54944 292528
rect 54996 292516 55002 292528
rect 66806 292516 66812 292528
rect 54996 292488 66812 292516
rect 54996 292476 55002 292488
rect 66806 292476 66812 292488
rect 66864 292476 66870 292528
rect 158070 291796 158076 291848
rect 158128 291836 158134 291848
rect 194042 291836 194048 291848
rect 158128 291808 194048 291836
rect 158128 291796 158134 291808
rect 194042 291796 194048 291808
rect 194100 291796 194106 291848
rect 200022 291796 200028 291848
rect 200080 291836 200086 291848
rect 358078 291836 358084 291848
rect 200080 291808 358084 291836
rect 200080 291796 200086 291808
rect 358078 291796 358084 291808
rect 358136 291796 358142 291848
rect 158714 291184 158720 291236
rect 158772 291224 158778 291236
rect 247310 291224 247316 291236
rect 158772 291196 247316 291224
rect 158772 291184 158778 291196
rect 247310 291184 247316 291196
rect 247368 291184 247374 291236
rect 41322 290436 41328 290488
rect 41380 290476 41386 290488
rect 63494 290476 63500 290488
rect 41380 290448 63500 290476
rect 41380 290436 41386 290448
rect 63494 290436 63500 290448
rect 63552 290436 63558 290488
rect 166442 290436 166448 290488
rect 166500 290476 166506 290488
rect 177482 290476 177488 290488
rect 166500 290448 177488 290476
rect 166500 290436 166506 290448
rect 177482 290436 177488 290448
rect 177540 290436 177546 290488
rect 240502 290436 240508 290488
rect 240560 290476 240566 290488
rect 259546 290476 259552 290488
rect 240560 290448 259552 290476
rect 240560 290436 240566 290448
rect 259546 290436 259552 290448
rect 259604 290436 259610 290488
rect 313366 290436 313372 290488
rect 313424 290476 313430 290488
rect 358906 290476 358912 290488
rect 313424 290448 358912 290476
rect 313424 290436 313430 290448
rect 358906 290436 358912 290448
rect 358964 290436 358970 290488
rect 63494 289892 63500 289944
rect 63552 289932 63558 289944
rect 64690 289932 64696 289944
rect 63552 289904 64696 289932
rect 63552 289892 63558 289904
rect 64690 289892 64696 289904
rect 64748 289932 64754 289944
rect 66806 289932 66812 289944
rect 64748 289904 66812 289932
rect 64748 289892 64754 289904
rect 66806 289892 66812 289904
rect 66864 289892 66870 289944
rect 184014 289892 184020 289944
rect 184072 289932 184078 289944
rect 244642 289932 244648 289944
rect 184072 289904 244648 289932
rect 184072 289892 184078 289904
rect 244642 289892 244648 289904
rect 244700 289892 244706 289944
rect 158714 289824 158720 289876
rect 158772 289864 158778 289876
rect 223574 289864 223580 289876
rect 158772 289836 223580 289864
rect 158772 289824 158778 289836
rect 223574 289824 223580 289836
rect 223632 289824 223638 289876
rect 245010 289824 245016 289876
rect 245068 289864 245074 289876
rect 245930 289864 245936 289876
rect 245068 289836 245936 289864
rect 245068 289824 245074 289836
rect 245930 289824 245936 289836
rect 245988 289864 245994 289876
rect 313366 289864 313372 289876
rect 245988 289836 313372 289864
rect 245988 289824 245994 289836
rect 313366 289824 313372 289836
rect 313424 289824 313430 289876
rect 169846 289756 169852 289808
rect 169904 289796 169910 289808
rect 209038 289796 209044 289808
rect 169904 289768 209044 289796
rect 169904 289756 169910 289768
rect 209038 289756 209044 289768
rect 209096 289756 209102 289808
rect 50798 289076 50804 289128
rect 50856 289116 50862 289128
rect 66714 289116 66720 289128
rect 50856 289088 66720 289116
rect 50856 289076 50862 289088
rect 66714 289076 66720 289088
rect 66772 289076 66778 289128
rect 217318 288464 217324 288516
rect 217376 288504 217382 288516
rect 248506 288504 248512 288516
rect 217376 288476 248512 288504
rect 217376 288464 217382 288476
rect 248506 288464 248512 288476
rect 248564 288464 248570 288516
rect 50890 288396 50896 288448
rect 50948 288436 50954 288448
rect 66806 288436 66812 288448
rect 50948 288408 66812 288436
rect 50948 288396 50954 288408
rect 66806 288396 66812 288408
rect 66864 288396 66870 288448
rect 158806 288396 158812 288448
rect 158864 288436 158870 288448
rect 231302 288436 231308 288448
rect 158864 288408 231308 288436
rect 158864 288396 158870 288408
rect 231302 288396 231308 288408
rect 231360 288396 231366 288448
rect 239398 288396 239404 288448
rect 239456 288436 239462 288448
rect 582558 288436 582564 288448
rect 239456 288408 582564 288436
rect 239456 288396 239462 288408
rect 582558 288396 582564 288408
rect 582616 288396 582622 288448
rect 231210 288328 231216 288380
rect 231268 288368 231274 288380
rect 237006 288368 237012 288380
rect 231268 288340 237012 288368
rect 231268 288328 231274 288340
rect 237006 288328 237012 288340
rect 237064 288328 237070 288380
rect 238110 287648 238116 287700
rect 238168 287688 238174 287700
rect 242894 287688 242900 287700
rect 238168 287660 242900 287688
rect 238168 287648 238174 287660
rect 242894 287648 242900 287660
rect 242952 287648 242958 287700
rect 158714 287104 158720 287156
rect 158772 287144 158778 287156
rect 171962 287144 171968 287156
rect 158772 287116 171968 287144
rect 158772 287104 158778 287116
rect 171962 287104 171968 287116
rect 172020 287104 172026 287156
rect 184198 287104 184204 287156
rect 184256 287144 184262 287156
rect 216766 287144 216772 287156
rect 184256 287116 216772 287144
rect 184256 287104 184262 287116
rect 216766 287104 216772 287116
rect 216824 287104 216830 287156
rect 218054 287104 218060 287156
rect 218112 287144 218118 287156
rect 255406 287144 255412 287156
rect 218112 287116 255412 287144
rect 218112 287104 218118 287116
rect 255406 287104 255412 287116
rect 255464 287104 255470 287156
rect 63402 287036 63408 287088
rect 63460 287076 63466 287088
rect 64782 287076 64788 287088
rect 63460 287048 64788 287076
rect 63460 287036 63466 287048
rect 64782 287036 64788 287048
rect 64840 287076 64846 287088
rect 66622 287076 66628 287088
rect 64840 287048 66628 287076
rect 64840 287036 64846 287048
rect 66622 287036 66628 287048
rect 66680 287036 66686 287088
rect 170490 287036 170496 287088
rect 170548 287076 170554 287088
rect 223666 287076 223672 287088
rect 170548 287048 223672 287076
rect 170548 287036 170554 287048
rect 223666 287036 223672 287048
rect 223724 287036 223730 287088
rect 45462 286968 45468 287020
rect 45520 287008 45526 287020
rect 52454 287008 52460 287020
rect 45520 286980 52460 287008
rect 45520 286968 45526 286980
rect 52454 286968 52460 286980
rect 52512 286968 52518 287020
rect 57698 286968 57704 287020
rect 57756 287008 57762 287020
rect 66806 287008 66812 287020
rect 57756 286980 66812 287008
rect 57756 286968 57762 286980
rect 66806 286968 66812 286980
rect 66864 286968 66870 287020
rect 158714 286968 158720 287020
rect 158772 287008 158778 287020
rect 169110 287008 169116 287020
rect 158772 286980 169116 287008
rect 158772 286968 158778 286980
rect 169110 286968 169116 286980
rect 169168 286968 169174 287020
rect 210418 286968 210424 287020
rect 210476 287008 210482 287020
rect 218054 287008 218060 287020
rect 210476 286980 218060 287008
rect 210476 286968 210482 286980
rect 218054 286968 218060 286980
rect 218112 286968 218118 287020
rect 52454 286288 52460 286340
rect 52512 286328 52518 286340
rect 53558 286328 53564 286340
rect 52512 286300 53564 286328
rect 52512 286288 52518 286300
rect 53558 286288 53564 286300
rect 53616 286328 53622 286340
rect 66346 286328 66352 286340
rect 53616 286300 66352 286328
rect 53616 286288 53622 286300
rect 66346 286288 66352 286300
rect 66404 286288 66410 286340
rect 158714 286288 158720 286340
rect 158772 286328 158778 286340
rect 165062 286328 165068 286340
rect 158772 286300 165068 286328
rect 158772 286288 158778 286300
rect 165062 286288 165068 286300
rect 165120 286288 165126 286340
rect 166350 286288 166356 286340
rect 166408 286328 166414 286340
rect 188522 286328 188528 286340
rect 166408 286300 188528 286328
rect 166408 286288 166414 286300
rect 188522 286288 188528 286300
rect 188580 286288 188586 286340
rect 282270 286288 282276 286340
rect 282328 286328 282334 286340
rect 582834 286328 582840 286340
rect 282328 286300 582840 286328
rect 282328 286288 282334 286300
rect 582834 286288 582840 286300
rect 582892 286288 582898 286340
rect 223574 286084 223580 286136
rect 223632 286124 223638 286136
rect 224494 286124 224500 286136
rect 223632 286096 224500 286124
rect 223632 286084 223638 286096
rect 224494 286084 224500 286096
rect 224552 286084 224558 286136
rect 231118 285812 231124 285864
rect 231176 285852 231182 285864
rect 231670 285852 231676 285864
rect 231176 285824 231676 285852
rect 231176 285812 231182 285824
rect 231670 285812 231676 285824
rect 231728 285852 231734 285864
rect 231728 285824 238754 285852
rect 231728 285812 231734 285824
rect 190362 285744 190368 285796
rect 190420 285784 190426 285796
rect 210878 285784 210884 285796
rect 190420 285756 210884 285784
rect 190420 285744 190426 285756
rect 210878 285744 210884 285756
rect 210936 285744 210942 285796
rect 222102 285744 222108 285796
rect 222160 285784 222166 285796
rect 222838 285784 222844 285796
rect 222160 285756 222844 285784
rect 222160 285744 222166 285756
rect 222838 285744 222844 285756
rect 222896 285744 222902 285796
rect 225414 285744 225420 285796
rect 225472 285784 225478 285796
rect 226426 285784 226432 285796
rect 225472 285756 226432 285784
rect 225472 285744 225478 285756
rect 226426 285744 226432 285756
rect 226484 285744 226490 285796
rect 236086 285744 236092 285796
rect 236144 285784 236150 285796
rect 237282 285784 237288 285796
rect 236144 285756 237288 285784
rect 236144 285744 236150 285756
rect 237282 285744 237288 285756
rect 237340 285744 237346 285796
rect 238726 285784 238754 285824
rect 258718 285784 258724 285796
rect 238726 285756 258724 285784
rect 258718 285744 258724 285756
rect 258776 285744 258782 285796
rect 269022 285744 269028 285796
rect 269080 285784 269086 285796
rect 275278 285784 275284 285796
rect 269080 285756 275284 285784
rect 269080 285744 269086 285756
rect 275278 285744 275284 285756
rect 275336 285744 275342 285796
rect 198826 285676 198832 285728
rect 198884 285716 198890 285728
rect 204622 285716 204628 285728
rect 198884 285688 204628 285716
rect 198884 285676 198890 285688
rect 204622 285676 204628 285688
rect 204680 285676 204686 285728
rect 207566 285676 207572 285728
rect 207624 285716 207630 285728
rect 300946 285716 300952 285728
rect 207624 285688 300952 285716
rect 207624 285676 207630 285688
rect 300946 285676 300952 285688
rect 301004 285676 301010 285728
rect 56502 285608 56508 285660
rect 56560 285648 56566 285660
rect 66714 285648 66720 285660
rect 56560 285620 66720 285648
rect 56560 285608 56566 285620
rect 66714 285608 66720 285620
rect 66772 285608 66778 285660
rect 200114 285268 200120 285320
rect 200172 285308 200178 285320
rect 200942 285308 200948 285320
rect 200172 285280 200948 285308
rect 200172 285268 200178 285280
rect 200942 285268 200948 285280
rect 201000 285268 201006 285320
rect 240134 285268 240140 285320
rect 240192 285308 240198 285320
rect 241054 285308 241060 285320
rect 240192 285280 241060 285308
rect 240192 285268 240198 285280
rect 241054 285268 241060 285280
rect 241112 285268 241118 285320
rect 243170 285268 243176 285320
rect 243228 285308 243234 285320
rect 244090 285308 244096 285320
rect 243228 285280 244096 285308
rect 243228 285268 243234 285280
rect 244090 285268 244096 285280
rect 244148 285268 244154 285320
rect 240778 285132 240784 285184
rect 240836 285172 240842 285184
rect 243814 285172 243820 285184
rect 240836 285144 243820 285172
rect 240836 285132 240842 285144
rect 243814 285132 243820 285144
rect 243872 285132 243878 285184
rect 48222 284928 48228 284980
rect 48280 284968 48286 284980
rect 56502 284968 56508 284980
rect 48280 284940 56508 284968
rect 48280 284928 48286 284940
rect 56502 284928 56508 284940
rect 56560 284928 56566 284980
rect 169110 284928 169116 284980
rect 169168 284968 169174 284980
rect 198826 284968 198832 284980
rect 169168 284940 198832 284968
rect 169168 284928 169174 284940
rect 198826 284928 198832 284940
rect 198884 284928 198890 284980
rect 187602 284384 187608 284436
rect 187660 284424 187666 284436
rect 217686 284424 217692 284436
rect 187660 284396 217692 284424
rect 187660 284384 187666 284396
rect 217686 284384 217692 284396
rect 217744 284384 217750 284436
rect 244458 284356 244464 284368
rect 200086 284328 244464 284356
rect 158806 284248 158812 284300
rect 158864 284288 158870 284300
rect 200086 284288 200114 284328
rect 244458 284316 244464 284328
rect 244516 284316 244522 284368
rect 158864 284260 200114 284288
rect 158864 284248 158870 284260
rect 245654 283908 245660 283960
rect 245712 283948 245718 283960
rect 245930 283948 245936 283960
rect 245712 283920 245936 283948
rect 245712 283908 245718 283920
rect 245930 283908 245936 283920
rect 245988 283908 245994 283960
rect 245930 283772 245936 283824
rect 245988 283812 245994 283824
rect 248414 283812 248420 283824
rect 245988 283784 248420 283812
rect 245988 283772 245994 283784
rect 248414 283772 248420 283784
rect 248472 283772 248478 283824
rect 56502 283568 56508 283620
rect 56560 283608 56566 283620
rect 66990 283608 66996 283620
rect 56560 283580 66996 283608
rect 56560 283568 56566 283580
rect 66990 283568 66996 283580
rect 67048 283568 67054 283620
rect 158714 283568 158720 283620
rect 158772 283608 158778 283620
rect 178126 283608 178132 283620
rect 158772 283580 178132 283608
rect 158772 283568 158778 283580
rect 178126 283568 178132 283580
rect 178184 283568 178190 283620
rect 64598 282888 64604 282940
rect 64656 282928 64662 282940
rect 66806 282928 66812 282940
rect 64656 282900 66812 282928
rect 64656 282888 64662 282900
rect 66806 282888 66812 282900
rect 66864 282888 66870 282940
rect 178126 282888 178132 282940
rect 178184 282928 178190 282940
rect 179322 282928 179328 282940
rect 178184 282900 179328 282928
rect 178184 282888 178190 282900
rect 179322 282888 179328 282900
rect 179380 282928 179386 282940
rect 179380 282900 180794 282928
rect 179380 282888 179386 282900
rect 158714 282820 158720 282872
rect 158772 282860 158778 282872
rect 158772 282832 161474 282860
rect 158772 282820 158778 282832
rect 161446 282724 161474 282832
rect 180766 282792 180794 282900
rect 197262 282888 197268 282940
rect 197320 282928 197326 282940
rect 199470 282928 199476 282940
rect 197320 282900 199476 282928
rect 197320 282888 197326 282900
rect 199470 282888 199476 282900
rect 199528 282888 199534 282940
rect 195882 282820 195888 282872
rect 195940 282860 195946 282872
rect 197998 282860 198004 282872
rect 195940 282832 198004 282860
rect 195940 282820 195946 282832
rect 197998 282820 198004 282832
rect 198056 282820 198062 282872
rect 254578 282820 254584 282872
rect 254636 282860 254642 282872
rect 255130 282860 255136 282872
rect 254636 282832 255136 282860
rect 254636 282820 254642 282832
rect 255130 282820 255136 282832
rect 255188 282860 255194 282872
rect 383654 282860 383660 282872
rect 255188 282832 383660 282860
rect 255188 282820 255194 282832
rect 383654 282820 383660 282832
rect 383712 282820 383718 282872
rect 197354 282792 197360 282804
rect 180766 282764 197360 282792
rect 197354 282752 197360 282764
rect 197412 282752 197418 282804
rect 245746 282752 245752 282804
rect 245804 282792 245810 282804
rect 260926 282792 260932 282804
rect 245804 282764 260932 282792
rect 245804 282752 245810 282764
rect 260926 282752 260932 282764
rect 260984 282752 260990 282804
rect 183094 282724 183100 282736
rect 161446 282696 183100 282724
rect 183094 282684 183100 282696
rect 183152 282684 183158 282736
rect 182910 282140 182916 282192
rect 182968 282180 182974 282192
rect 192570 282180 192576 282192
rect 182968 282152 192576 282180
rect 182968 282140 182974 282152
rect 192570 282140 192576 282152
rect 192628 282140 192634 282192
rect 272610 282140 272616 282192
rect 272668 282180 272674 282192
rect 282178 282180 282184 282192
rect 272668 282152 282184 282180
rect 272668 282140 272674 282152
rect 282178 282140 282184 282152
rect 282236 282140 282242 282192
rect 282270 282140 282276 282192
rect 282328 282180 282334 282192
rect 302326 282180 302332 282192
rect 282328 282152 302332 282180
rect 282328 282140 282334 282152
rect 302326 282140 302332 282152
rect 302384 282140 302390 282192
rect 302878 282140 302884 282192
rect 302936 282180 302942 282192
rect 327718 282180 327724 282192
rect 302936 282152 327724 282180
rect 302936 282140 302942 282152
rect 327718 282140 327724 282152
rect 327776 282140 327782 282192
rect 192754 282072 192760 282124
rect 192812 282112 192818 282124
rect 194134 282112 194140 282124
rect 192812 282084 194140 282112
rect 192812 282072 192818 282084
rect 194134 282072 194140 282084
rect 194192 282072 194198 282124
rect 245930 281528 245936 281580
rect 245988 281568 245994 281580
rect 249886 281568 249892 281580
rect 245988 281540 249892 281568
rect 245988 281528 245994 281540
rect 249886 281528 249892 281540
rect 249944 281528 249950 281580
rect 180150 281460 180156 281512
rect 180208 281500 180214 281512
rect 197354 281500 197360 281512
rect 180208 281472 197360 281500
rect 180208 281460 180214 281472
rect 197354 281460 197360 281472
rect 197412 281460 197418 281512
rect 173250 280780 173256 280832
rect 173308 280820 173314 280832
rect 176010 280820 176016 280832
rect 173308 280792 176016 280820
rect 173308 280780 173314 280792
rect 176010 280780 176016 280792
rect 176068 280780 176074 280832
rect 245654 280780 245660 280832
rect 245712 280820 245718 280832
rect 250070 280820 250076 280832
rect 245712 280792 250076 280820
rect 245712 280780 245718 280792
rect 250070 280780 250076 280792
rect 250128 280820 250134 280832
rect 298278 280820 298284 280832
rect 250128 280792 298284 280820
rect 250128 280780 250134 280792
rect 298278 280780 298284 280792
rect 298336 280820 298342 280832
rect 378226 280820 378232 280832
rect 298336 280792 378232 280820
rect 298336 280780 298342 280792
rect 378226 280780 378232 280792
rect 378284 280780 378290 280832
rect 196710 280440 196716 280492
rect 196768 280480 196774 280492
rect 197262 280480 197268 280492
rect 196768 280452 197268 280480
rect 196768 280440 196774 280452
rect 197262 280440 197268 280452
rect 197320 280480 197326 280492
rect 198274 280480 198280 280492
rect 197320 280452 198280 280480
rect 197320 280440 197326 280452
rect 198274 280440 198280 280452
rect 198332 280440 198338 280492
rect 21358 280168 21364 280220
rect 21416 280208 21422 280220
rect 61838 280208 61844 280220
rect 21416 280180 61844 280208
rect 21416 280168 21422 280180
rect 61838 280168 61844 280180
rect 61896 280208 61902 280220
rect 67174 280208 67180 280220
rect 61896 280180 67180 280208
rect 61896 280168 61902 280180
rect 67174 280168 67180 280180
rect 67232 280168 67238 280220
rect 158714 280100 158720 280152
rect 158772 280140 158778 280152
rect 169294 280140 169300 280152
rect 158772 280112 169300 280140
rect 158772 280100 158778 280112
rect 169294 280100 169300 280112
rect 169352 280100 169358 280152
rect 196618 280100 196624 280152
rect 196676 280140 196682 280152
rect 199378 280140 199384 280152
rect 196676 280112 199384 280140
rect 196676 280100 196682 280112
rect 199378 280100 199384 280112
rect 199436 280100 199442 280152
rect 245746 279488 245752 279540
rect 245804 279528 245810 279540
rect 249978 279528 249984 279540
rect 245804 279500 249984 279528
rect 245804 279488 245810 279500
rect 249978 279488 249984 279500
rect 250036 279488 250042 279540
rect 54938 279420 54944 279472
rect 54996 279460 55002 279472
rect 67082 279460 67088 279472
rect 54996 279432 67088 279460
rect 54996 279420 55002 279432
rect 67082 279420 67088 279432
rect 67140 279420 67146 279472
rect 167638 279420 167644 279472
rect 167696 279460 167702 279472
rect 193214 279460 193220 279472
rect 167696 279432 193220 279460
rect 167696 279420 167702 279432
rect 193214 279420 193220 279432
rect 193272 279420 193278 279472
rect 245930 279420 245936 279472
rect 245988 279460 245994 279472
rect 255590 279460 255596 279472
rect 245988 279432 255596 279460
rect 245988 279420 245994 279432
rect 255590 279420 255596 279432
rect 255648 279420 255654 279472
rect 158714 278740 158720 278792
rect 158772 278780 158778 278792
rect 165062 278780 165068 278792
rect 158772 278752 165068 278780
rect 158772 278740 158778 278752
rect 165062 278740 165068 278752
rect 165120 278740 165126 278792
rect 193214 278740 193220 278792
rect 193272 278780 193278 278792
rect 197354 278780 197360 278792
rect 193272 278752 197360 278780
rect 193272 278740 193278 278752
rect 197354 278740 197360 278752
rect 197412 278740 197418 278792
rect 255590 278740 255596 278792
rect 255648 278780 255654 278792
rect 583110 278780 583116 278792
rect 255648 278752 583116 278780
rect 255648 278740 255654 278752
rect 583110 278740 583116 278752
rect 583168 278740 583174 278792
rect 196802 278672 196808 278724
rect 196860 278712 196866 278724
rect 197262 278712 197268 278724
rect 196860 278684 197268 278712
rect 196860 278672 196866 278684
rect 197262 278672 197268 278684
rect 197320 278672 197326 278724
rect 245746 278672 245752 278724
rect 245804 278712 245810 278724
rect 249978 278712 249984 278724
rect 245804 278684 249984 278712
rect 245804 278672 245810 278684
rect 249978 278672 249984 278684
rect 250036 278712 250042 278724
rect 389174 278712 389180 278724
rect 250036 278684 389180 278712
rect 250036 278672 250042 278684
rect 389174 278672 389180 278684
rect 389232 278672 389238 278724
rect 266262 278604 266268 278656
rect 266320 278644 266326 278656
rect 289078 278644 289084 278656
rect 266320 278616 289084 278644
rect 266320 278604 266326 278616
rect 289078 278604 289084 278616
rect 289136 278604 289142 278656
rect 180150 278060 180156 278112
rect 180208 278100 180214 278112
rect 198826 278100 198832 278112
rect 180208 278072 198832 278100
rect 180208 278060 180214 278072
rect 198826 278060 198832 278072
rect 198884 278060 198890 278112
rect 158806 277992 158812 278044
rect 158864 278032 158870 278044
rect 189074 278032 189080 278044
rect 158864 278004 189080 278032
rect 158864 277992 158870 278004
rect 189074 277992 189080 278004
rect 189132 277992 189138 278044
rect 389174 277992 389180 278044
rect 389232 278032 389238 278044
rect 583386 278032 583392 278044
rect 389232 278004 583392 278032
rect 389232 277992 389238 278004
rect 583386 277992 583392 278004
rect 583444 277992 583450 278044
rect 63218 277380 63224 277432
rect 63276 277420 63282 277432
rect 66806 277420 66812 277432
rect 63276 277392 66812 277420
rect 63276 277380 63282 277392
rect 66806 277380 66812 277392
rect 66864 277380 66870 277432
rect 158714 277312 158720 277364
rect 158772 277352 158778 277364
rect 165154 277352 165160 277364
rect 158772 277324 165160 277352
rect 158772 277312 158778 277324
rect 165154 277312 165160 277324
rect 165212 277312 165218 277364
rect 186038 277312 186044 277364
rect 186096 277352 186102 277364
rect 197354 277352 197360 277364
rect 186096 277324 197360 277352
rect 186096 277312 186102 277324
rect 197354 277312 197360 277324
rect 197412 277312 197418 277364
rect 49602 276632 49608 276684
rect 49660 276672 49666 276684
rect 60458 276672 60464 276684
rect 49660 276644 60464 276672
rect 49660 276632 49666 276644
rect 60458 276632 60464 276644
rect 60516 276672 60522 276684
rect 66806 276672 66812 276684
rect 60516 276644 66812 276672
rect 60516 276632 60522 276644
rect 66806 276632 66812 276644
rect 66864 276632 66870 276684
rect 189074 276632 189080 276684
rect 189132 276672 189138 276684
rect 190270 276672 190276 276684
rect 189132 276644 190276 276672
rect 189132 276632 189138 276644
rect 190270 276632 190276 276644
rect 190328 276672 190334 276684
rect 197354 276672 197360 276684
rect 190328 276644 197360 276672
rect 190328 276632 190334 276644
rect 197354 276632 197360 276644
rect 197412 276632 197418 276684
rect 246114 276632 246120 276684
rect 246172 276672 246178 276684
rect 318794 276672 318800 276684
rect 246172 276644 318800 276672
rect 246172 276632 246178 276644
rect 318794 276632 318800 276644
rect 318852 276672 318858 276684
rect 367186 276672 367192 276684
rect 318852 276644 367192 276672
rect 318852 276632 318858 276644
rect 367186 276632 367192 276644
rect 367244 276632 367250 276684
rect 244090 276020 244096 276072
rect 244148 276060 244154 276072
rect 245746 276060 245752 276072
rect 244148 276032 245752 276060
rect 244148 276020 244154 276032
rect 245746 276020 245752 276032
rect 245804 276020 245810 276072
rect 159358 275272 159364 275324
rect 159416 275312 159422 275324
rect 172054 275312 172060 275324
rect 159416 275284 172060 275312
rect 159416 275272 159422 275284
rect 172054 275272 172060 275284
rect 172112 275272 172118 275324
rect 262950 275272 262956 275324
rect 263008 275312 263014 275324
rect 278038 275312 278044 275324
rect 263008 275284 278044 275312
rect 263008 275272 263014 275284
rect 278038 275272 278044 275284
rect 278096 275272 278102 275324
rect 280982 275272 280988 275324
rect 281040 275312 281046 275324
rect 583294 275312 583300 275324
rect 281040 275284 583300 275312
rect 281040 275272 281046 275284
rect 583294 275272 583300 275284
rect 583352 275272 583358 275324
rect 175274 274728 175280 274780
rect 175332 274768 175338 274780
rect 178034 274768 178040 274780
rect 175332 274740 178040 274768
rect 175332 274728 175338 274740
rect 178034 274728 178040 274740
rect 178092 274728 178098 274780
rect 185670 274728 185676 274780
rect 185728 274768 185734 274780
rect 197446 274768 197452 274780
rect 185728 274740 197452 274768
rect 185728 274728 185734 274740
rect 197446 274728 197452 274740
rect 197504 274728 197510 274780
rect 66622 274700 66628 274712
rect 57900 274672 66628 274700
rect 35802 274592 35808 274644
rect 35860 274632 35866 274644
rect 57238 274632 57244 274644
rect 35860 274604 57244 274632
rect 35860 274592 35866 274604
rect 57238 274592 57244 274604
rect 57296 274632 57302 274644
rect 57900 274632 57928 274672
rect 66622 274660 66628 274672
rect 66680 274660 66686 274712
rect 158806 274660 158812 274712
rect 158864 274700 158870 274712
rect 167638 274700 167644 274712
rect 158864 274672 167644 274700
rect 158864 274660 158870 274672
rect 167638 274660 167644 274672
rect 167696 274660 167702 274712
rect 169294 274660 169300 274712
rect 169352 274700 169358 274712
rect 197354 274700 197360 274712
rect 169352 274672 197360 274700
rect 169352 274660 169358 274672
rect 197354 274660 197360 274672
rect 197412 274660 197418 274712
rect 57296 274604 57928 274632
rect 57296 274592 57302 274604
rect 158714 274592 158720 274644
rect 158772 274632 158778 274644
rect 191190 274632 191196 274644
rect 158772 274604 191196 274632
rect 158772 274592 158778 274604
rect 191190 274592 191196 274604
rect 191248 274592 191254 274644
rect 194042 274524 194048 274576
rect 194100 274564 194106 274576
rect 197078 274564 197084 274576
rect 194100 274536 197084 274564
rect 194100 274524 194106 274536
rect 197078 274524 197084 274536
rect 197136 274564 197142 274576
rect 197354 274564 197360 274576
rect 197136 274536 197360 274564
rect 197136 274524 197142 274536
rect 197354 274524 197360 274536
rect 197412 274524 197418 274576
rect 245930 273912 245936 273964
rect 245988 273952 245994 273964
rect 289814 273952 289820 273964
rect 245988 273924 289820 273952
rect 245988 273912 245994 273924
rect 289814 273912 289820 273924
rect 289872 273952 289878 273964
rect 369946 273952 369952 273964
rect 289872 273924 369952 273952
rect 289872 273912 289878 273924
rect 369946 273912 369952 273924
rect 370004 273912 370010 273964
rect 264330 273572 264336 273624
rect 264388 273612 264394 273624
rect 269114 273612 269120 273624
rect 264388 273584 269120 273612
rect 264388 273572 264394 273584
rect 269114 273572 269120 273584
rect 269172 273572 269178 273624
rect 180058 273300 180064 273352
rect 180116 273340 180122 273352
rect 197354 273340 197360 273352
rect 180116 273312 197360 273340
rect 180116 273300 180122 273312
rect 197354 273300 197360 273312
rect 197412 273300 197418 273352
rect 184842 273164 184848 273216
rect 184900 273204 184906 273216
rect 197354 273204 197360 273216
rect 184900 273176 197360 273204
rect 184900 273164 184906 273176
rect 197354 273164 197360 273176
rect 197412 273164 197418 273216
rect 245838 273164 245844 273216
rect 245896 273204 245902 273216
rect 251174 273204 251180 273216
rect 245896 273176 251180 273204
rect 245896 273164 245902 273176
rect 251174 273164 251180 273176
rect 251232 273204 251238 273216
rect 252462 273204 252468 273216
rect 251232 273176 252468 273204
rect 251232 273164 251238 273176
rect 252462 273164 252468 273176
rect 252520 273164 252526 273216
rect 192662 273096 192668 273148
rect 192720 273136 192726 273148
rect 197446 273136 197452 273148
rect 192720 273108 197452 273136
rect 192720 273096 192726 273108
rect 197446 273096 197452 273108
rect 197504 273096 197510 273148
rect 168282 272484 168288 272536
rect 168340 272524 168346 272536
rect 183554 272524 183560 272536
rect 168340 272496 183560 272524
rect 168340 272484 168346 272496
rect 183554 272484 183560 272496
rect 183612 272484 183618 272536
rect 252462 272484 252468 272536
rect 252520 272524 252526 272536
rect 288434 272524 288440 272536
rect 252520 272496 288440 272524
rect 252520 272484 252526 272496
rect 288434 272484 288440 272496
rect 288492 272524 288498 272536
rect 365714 272524 365720 272536
rect 288492 272496 365720 272524
rect 288492 272484 288498 272496
rect 365714 272484 365720 272496
rect 365772 272484 365778 272536
rect 52086 271872 52092 271924
rect 52144 271912 52150 271924
rect 66254 271912 66260 271924
rect 52144 271884 66260 271912
rect 52144 271872 52150 271884
rect 66254 271872 66260 271884
rect 66312 271872 66318 271924
rect 574738 271872 574744 271924
rect 574796 271912 574802 271924
rect 579798 271912 579804 271924
rect 574796 271884 579804 271912
rect 574796 271872 574802 271884
rect 579798 271872 579804 271884
rect 579856 271872 579862 271924
rect 191098 271804 191104 271856
rect 191156 271844 191162 271856
rect 191834 271844 191840 271856
rect 191156 271816 191840 271844
rect 191156 271804 191162 271816
rect 191834 271804 191840 271816
rect 191892 271804 191898 271856
rect 191190 271192 191196 271244
rect 191248 271232 191254 271244
rect 198734 271232 198740 271244
rect 191248 271204 198740 271232
rect 191248 271192 191254 271204
rect 198734 271192 198740 271204
rect 198792 271192 198798 271244
rect 158714 271124 158720 271176
rect 158772 271164 158778 271176
rect 181530 271164 181536 271176
rect 158772 271136 181536 271164
rect 158772 271124 158778 271136
rect 181530 271124 181536 271136
rect 181588 271124 181594 271176
rect 245930 271124 245936 271176
rect 245988 271164 245994 271176
rect 256970 271164 256976 271176
rect 245988 271136 256976 271164
rect 245988 271124 245994 271136
rect 256970 271124 256976 271136
rect 257028 271124 257034 271176
rect 286042 271124 286048 271176
rect 286100 271164 286106 271176
rect 372614 271164 372620 271176
rect 286100 271136 372620 271164
rect 286100 271124 286106 271136
rect 372614 271124 372620 271136
rect 372672 271124 372678 271176
rect 195146 270512 195152 270564
rect 195204 270552 195210 270564
rect 197354 270552 197360 270564
rect 195204 270524 197360 270552
rect 195204 270512 195210 270524
rect 197354 270512 197360 270524
rect 197412 270512 197418 270564
rect 245746 270444 245752 270496
rect 245804 270484 245810 270496
rect 254026 270484 254032 270496
rect 245804 270456 254032 270484
rect 245804 270444 245810 270456
rect 254026 270444 254032 270456
rect 254084 270444 254090 270496
rect 166902 269832 166908 269884
rect 166960 269872 166966 269884
rect 180242 269872 180248 269884
rect 166960 269844 180248 269872
rect 166960 269832 166966 269844
rect 180242 269832 180248 269844
rect 180300 269832 180306 269884
rect 180334 269832 180340 269884
rect 180392 269872 180398 269884
rect 196710 269872 196716 269884
rect 180392 269844 196716 269872
rect 180392 269832 180398 269844
rect 196710 269832 196716 269844
rect 196768 269832 196774 269884
rect 260098 269832 260104 269884
rect 260156 269872 260162 269884
rect 295334 269872 295340 269884
rect 260156 269844 295340 269872
rect 260156 269832 260162 269844
rect 295334 269832 295340 269844
rect 295392 269832 295398 269884
rect 4062 269764 4068 269816
rect 4120 269804 4126 269816
rect 11698 269804 11704 269816
rect 4120 269776 11704 269804
rect 4120 269764 4126 269776
rect 11698 269764 11704 269776
rect 11756 269764 11762 269816
rect 158530 269764 158536 269816
rect 158588 269804 158594 269816
rect 195146 269804 195152 269816
rect 158588 269776 195152 269804
rect 158588 269764 158594 269776
rect 195146 269764 195152 269776
rect 195204 269764 195210 269816
rect 245838 269764 245844 269816
rect 245896 269804 245902 269816
rect 287146 269804 287152 269816
rect 245896 269776 287152 269804
rect 245896 269764 245902 269776
rect 287146 269764 287152 269776
rect 287204 269764 287210 269816
rect 256878 269084 256884 269136
rect 256936 269084 256942 269136
rect 169202 269016 169208 269068
rect 169260 269056 169266 269068
rect 197354 269056 197360 269068
rect 169260 269028 197360 269056
rect 169260 269016 169266 269028
rect 197354 269016 197360 269028
rect 197412 269016 197418 269068
rect 249058 269016 249064 269068
rect 249116 269056 249122 269068
rect 250070 269056 250076 269068
rect 249116 269028 250076 269056
rect 249116 269016 249122 269028
rect 250070 269016 250076 269028
rect 250128 269016 250134 269068
rect 254394 269016 254400 269068
rect 254452 269056 254458 269068
rect 256896 269056 256924 269084
rect 583018 269056 583024 269068
rect 254452 269028 583024 269056
rect 254452 269016 254458 269028
rect 583018 269016 583024 269028
rect 583076 269016 583082 269068
rect 158714 268948 158720 269000
rect 158772 268988 158778 269000
rect 170490 268988 170496 269000
rect 158772 268960 170496 268988
rect 158772 268948 158778 268960
rect 170490 268948 170496 268960
rect 170548 268948 170554 269000
rect 189074 268948 189080 269000
rect 189132 268988 189138 269000
rect 189810 268988 189816 269000
rect 189132 268960 189816 268988
rect 189132 268948 189138 268960
rect 189810 268948 189816 268960
rect 189868 268988 189874 269000
rect 197446 268988 197452 269000
rect 189868 268960 197452 268988
rect 189868 268948 189874 268960
rect 197446 268948 197452 268960
rect 197504 268948 197510 269000
rect 178770 268336 178776 268388
rect 178828 268376 178834 268388
rect 189074 268376 189080 268388
rect 178828 268348 189080 268376
rect 178828 268336 178834 268348
rect 189074 268336 189080 268348
rect 189132 268336 189138 268388
rect 246758 268336 246764 268388
rect 246816 268376 246822 268388
rect 254394 268376 254400 268388
rect 246816 268348 254400 268376
rect 246816 268336 246822 268348
rect 254394 268336 254400 268348
rect 254452 268336 254458 268388
rect 158714 267928 158720 267980
rect 158772 267968 158778 267980
rect 162118 267968 162124 267980
rect 158772 267940 162124 267968
rect 158772 267928 158778 267940
rect 162118 267928 162124 267940
rect 162176 267928 162182 267980
rect 63310 267792 63316 267844
rect 63368 267832 63374 267844
rect 66806 267832 66812 267844
rect 63368 267804 66812 267832
rect 63368 267792 63374 267804
rect 66806 267792 66812 267804
rect 66864 267792 66870 267844
rect 3326 267724 3332 267776
rect 3384 267764 3390 267776
rect 22738 267764 22744 267776
rect 3384 267736 22744 267764
rect 3384 267724 3390 267736
rect 22738 267724 22744 267736
rect 22796 267724 22802 267776
rect 61930 267724 61936 267776
rect 61988 267764 61994 267776
rect 67174 267764 67180 267776
rect 61988 267736 67180 267764
rect 61988 267724 61994 267736
rect 67174 267724 67180 267736
rect 67232 267724 67238 267776
rect 170490 267656 170496 267708
rect 170548 267696 170554 267708
rect 182818 267696 182824 267708
rect 170548 267668 182824 267696
rect 170548 267656 170554 267668
rect 182818 267656 182824 267668
rect 182876 267656 182882 267708
rect 188338 267656 188344 267708
rect 188396 267696 188402 267708
rect 197354 267696 197360 267708
rect 188396 267668 197360 267696
rect 188396 267656 188402 267668
rect 197354 267656 197360 267668
rect 197412 267656 197418 267708
rect 246942 267520 246948 267572
rect 247000 267560 247006 267572
rect 248414 267560 248420 267572
rect 247000 267532 248420 267560
rect 247000 267520 247006 267532
rect 248414 267520 248420 267532
rect 248472 267520 248478 267572
rect 270402 266976 270408 267028
rect 270460 267016 270466 267028
rect 362954 267016 362960 267028
rect 270460 266988 362960 267016
rect 270460 266976 270466 266988
rect 362954 266976 362960 266988
rect 363012 266976 363018 267028
rect 189074 266364 189080 266416
rect 189132 266404 189138 266416
rect 195330 266404 195336 266416
rect 189132 266376 195336 266404
rect 189132 266364 189138 266376
rect 195330 266364 195336 266376
rect 195388 266364 195394 266416
rect 162210 265616 162216 265668
rect 162268 265656 162274 265668
rect 178862 265656 178868 265668
rect 162268 265628 178868 265656
rect 162268 265616 162274 265628
rect 178862 265616 178868 265628
rect 178920 265616 178926 265668
rect 245930 265616 245936 265668
rect 245988 265656 245994 265668
rect 248598 265656 248604 265668
rect 245988 265628 248604 265656
rect 245988 265616 245994 265628
rect 248598 265616 248604 265628
rect 248656 265656 248662 265668
rect 251266 265656 251272 265668
rect 248656 265628 251272 265656
rect 248656 265616 248662 265628
rect 251266 265616 251272 265628
rect 251324 265616 251330 265668
rect 53558 264936 53564 264988
rect 53616 264976 53622 264988
rect 66806 264976 66812 264988
rect 53616 264948 66812 264976
rect 53616 264936 53622 264948
rect 66806 264936 66812 264948
rect 66864 264936 66870 264988
rect 195330 264936 195336 264988
rect 195388 264976 195394 264988
rect 197446 264976 197452 264988
rect 195388 264948 197452 264976
rect 195388 264936 195394 264948
rect 197446 264936 197452 264948
rect 197504 264936 197510 264988
rect 187050 264868 187056 264920
rect 187108 264908 187114 264920
rect 197354 264908 197360 264920
rect 187108 264880 197360 264908
rect 187108 264868 187114 264880
rect 197354 264868 197360 264880
rect 197412 264868 197418 264920
rect 245838 264868 245844 264920
rect 245896 264908 245902 264920
rect 273254 264908 273260 264920
rect 245896 264880 273260 264908
rect 245896 264868 245902 264880
rect 273254 264868 273260 264880
rect 273312 264868 273318 264920
rect 167822 264188 167828 264240
rect 167880 264228 167886 264240
rect 183002 264228 183008 264240
rect 167880 264200 183008 264228
rect 167880 264188 167886 264200
rect 183002 264188 183008 264200
rect 183060 264188 183066 264240
rect 162762 263644 162768 263696
rect 162820 263684 162826 263696
rect 164234 263684 164240 263696
rect 162820 263656 164240 263684
rect 162820 263644 162826 263656
rect 164234 263644 164240 263656
rect 164292 263644 164298 263696
rect 182818 263644 182824 263696
rect 182876 263684 182882 263696
rect 197354 263684 197360 263696
rect 182876 263656 197360 263684
rect 182876 263644 182882 263656
rect 197354 263644 197360 263656
rect 197412 263644 197418 263696
rect 53742 263576 53748 263628
rect 53800 263616 53806 263628
rect 57698 263616 57704 263628
rect 53800 263588 57704 263616
rect 53800 263576 53806 263588
rect 57698 263576 57704 263588
rect 57756 263616 57762 263628
rect 66806 263616 66812 263628
rect 57756 263588 66812 263616
rect 57756 263576 57762 263588
rect 66806 263576 66812 263588
rect 66864 263576 66870 263628
rect 158714 263576 158720 263628
rect 158772 263616 158778 263628
rect 186958 263616 186964 263628
rect 158772 263588 186964 263616
rect 158772 263576 158778 263588
rect 186958 263576 186964 263588
rect 187016 263576 187022 263628
rect 253198 263508 253204 263560
rect 253256 263548 253262 263560
rect 385126 263548 385132 263560
rect 253256 263520 385132 263548
rect 253256 263508 253262 263520
rect 385126 263508 385132 263520
rect 385184 263508 385190 263560
rect 158070 262896 158076 262948
rect 158128 262936 158134 262948
rect 166442 262936 166448 262948
rect 158128 262908 166448 262936
rect 158128 262896 158134 262908
rect 166442 262896 166448 262908
rect 166500 262896 166506 262948
rect 169202 262896 169208 262948
rect 169260 262936 169266 262948
rect 191282 262936 191288 262948
rect 169260 262908 191288 262936
rect 169260 262896 169266 262908
rect 191282 262896 191288 262908
rect 191340 262896 191346 262948
rect 39850 262828 39856 262880
rect 39908 262868 39914 262880
rect 49602 262868 49608 262880
rect 39908 262840 49608 262868
rect 39908 262828 39914 262840
rect 49602 262828 49608 262840
rect 49660 262828 49666 262880
rect 159358 262828 159364 262880
rect 159416 262868 159422 262880
rect 196618 262868 196624 262880
rect 159416 262840 196624 262868
rect 159416 262828 159422 262840
rect 196618 262828 196624 262840
rect 196676 262828 196682 262880
rect 166534 262488 166540 262540
rect 166592 262528 166598 262540
rect 168650 262528 168656 262540
rect 166592 262500 168656 262528
rect 166592 262488 166598 262500
rect 168650 262488 168656 262500
rect 168708 262488 168714 262540
rect 49602 262216 49608 262268
rect 49660 262256 49666 262268
rect 66806 262256 66812 262268
rect 49660 262228 66812 262256
rect 49660 262216 49666 262228
rect 66806 262216 66812 262228
rect 66864 262216 66870 262268
rect 245930 262216 245936 262268
rect 245988 262256 245994 262268
rect 252646 262256 252652 262268
rect 245988 262228 252652 262256
rect 245988 262216 245994 262228
rect 252646 262216 252652 262228
rect 252704 262216 252710 262268
rect 11698 262148 11704 262200
rect 11756 262188 11762 262200
rect 66438 262188 66444 262200
rect 11756 262160 66444 262188
rect 11756 262148 11762 262160
rect 66438 262148 66444 262160
rect 66496 262148 66502 262200
rect 191374 262148 191380 262200
rect 191432 262188 191438 262200
rect 193214 262188 193220 262200
rect 191432 262160 193220 262188
rect 191432 262148 191438 262160
rect 193214 262148 193220 262160
rect 193272 262148 193278 262200
rect 175090 261536 175096 261588
rect 175148 261576 175154 261588
rect 184474 261576 184480 261588
rect 175148 261548 184480 261576
rect 175148 261536 175154 261548
rect 184474 261536 184480 261548
rect 184532 261536 184538 261588
rect 157978 261468 157984 261520
rect 158036 261508 158042 261520
rect 191834 261508 191840 261520
rect 158036 261480 191840 261508
rect 158036 261468 158042 261480
rect 191834 261468 191840 261480
rect 191892 261508 191898 261520
rect 197354 261508 197360 261520
rect 191892 261480 197360 261508
rect 191892 261468 191898 261480
rect 197354 261468 197360 261480
rect 197412 261468 197418 261520
rect 246390 261468 246396 261520
rect 246448 261508 246454 261520
rect 247310 261508 247316 261520
rect 246448 261480 247316 261508
rect 246448 261468 246454 261480
rect 247310 261468 247316 261480
rect 247368 261508 247374 261520
rect 251174 261508 251180 261520
rect 247368 261480 251180 261508
rect 247368 261468 247374 261480
rect 251174 261468 251180 261480
rect 251232 261468 251238 261520
rect 264238 261468 264244 261520
rect 264296 261508 264302 261520
rect 323578 261508 323584 261520
rect 264296 261480 323584 261508
rect 264296 261468 264302 261480
rect 323578 261468 323584 261480
rect 323636 261468 323642 261520
rect 245838 260788 245844 260840
rect 245896 260828 245902 260840
rect 253198 260828 253204 260840
rect 245896 260800 253204 260828
rect 245896 260788 245902 260800
rect 253198 260788 253204 260800
rect 253256 260788 253262 260840
rect 163498 260108 163504 260160
rect 163556 260148 163562 260160
rect 188338 260148 188344 260160
rect 163556 260120 188344 260148
rect 163556 260108 163562 260120
rect 188338 260108 188344 260120
rect 188396 260108 188402 260160
rect 260098 260108 260104 260160
rect 260156 260148 260162 260160
rect 282270 260148 282276 260160
rect 260156 260120 282276 260148
rect 260156 260108 260162 260120
rect 282270 260108 282276 260120
rect 282328 260108 282334 260160
rect 314654 260108 314660 260160
rect 314712 260148 314718 260160
rect 364334 260148 364340 260160
rect 314712 260120 364340 260148
rect 314712 260108 314718 260120
rect 364334 260108 364340 260120
rect 364392 260108 364398 260160
rect 64782 259428 64788 259480
rect 64840 259468 64846 259480
rect 66806 259468 66812 259480
rect 64840 259440 66812 259468
rect 64840 259428 64846 259440
rect 66806 259428 66812 259440
rect 66864 259428 66870 259480
rect 193122 259428 193128 259480
rect 193180 259468 193186 259480
rect 197354 259468 197360 259480
rect 193180 259440 197360 259468
rect 193180 259428 193186 259440
rect 197354 259428 197360 259440
rect 197412 259428 197418 259480
rect 245930 259428 245936 259480
rect 245988 259468 245994 259480
rect 314654 259468 314660 259480
rect 245988 259440 314660 259468
rect 245988 259428 245994 259440
rect 314654 259428 314660 259440
rect 314712 259428 314718 259480
rect 175182 259360 175188 259412
rect 175240 259400 175246 259412
rect 177390 259400 177396 259412
rect 175240 259372 177396 259400
rect 175240 259360 175246 259372
rect 177390 259360 177396 259372
rect 177448 259360 177454 259412
rect 191742 259360 191748 259412
rect 191800 259400 191806 259412
rect 197446 259400 197452 259412
rect 191800 259372 197452 259400
rect 191800 259360 191806 259372
rect 197446 259360 197452 259372
rect 197504 259360 197510 259412
rect 245838 259360 245844 259412
rect 245896 259400 245902 259412
rect 254118 259400 254124 259412
rect 245896 259372 254124 259400
rect 245896 259360 245902 259372
rect 254118 259360 254124 259372
rect 254176 259360 254182 259412
rect 381538 259360 381544 259412
rect 381596 259400 381602 259412
rect 580166 259400 580172 259412
rect 381596 259372 580172 259400
rect 381596 259360 381602 259372
rect 580166 259360 580172 259372
rect 580224 259360 580230 259412
rect 245930 259292 245936 259344
rect 245988 259332 245994 259344
rect 252738 259332 252744 259344
rect 245988 259304 252744 259332
rect 245988 259292 245994 259304
rect 252738 259292 252744 259304
rect 252796 259332 252802 259344
rect 253014 259332 253020 259344
rect 252796 259304 253020 259332
rect 252796 259292 252802 259304
rect 253014 259292 253020 259304
rect 253072 259292 253078 259344
rect 254118 258748 254124 258800
rect 254176 258788 254182 258800
rect 255130 258788 255136 258800
rect 254176 258760 255136 258788
rect 254176 258748 254182 258760
rect 255130 258748 255136 258760
rect 255188 258788 255194 258800
rect 278038 258788 278044 258800
rect 255188 258760 278044 258788
rect 255188 258748 255194 258760
rect 278038 258748 278044 258760
rect 278096 258748 278102 258800
rect 158714 258680 158720 258732
rect 158772 258720 158778 258732
rect 184198 258720 184204 258732
rect 158772 258692 184204 258720
rect 158772 258680 158778 258692
rect 184198 258680 184204 258692
rect 184256 258680 184262 258732
rect 187234 258680 187240 258732
rect 187292 258720 187298 258732
rect 194410 258720 194416 258732
rect 187292 258692 194416 258720
rect 187292 258680 187298 258692
rect 194410 258680 194416 258692
rect 194468 258720 194474 258732
rect 197354 258720 197360 258732
rect 194468 258692 197360 258720
rect 194468 258680 194474 258692
rect 197354 258680 197360 258692
rect 197412 258680 197418 258732
rect 253014 258680 253020 258732
rect 253072 258720 253078 258732
rect 294046 258720 294052 258732
rect 253072 258692 294052 258720
rect 253072 258680 253078 258692
rect 294046 258680 294052 258692
rect 294104 258720 294110 258732
rect 356698 258720 356704 258732
rect 294104 258692 356704 258720
rect 294104 258680 294110 258692
rect 356698 258680 356704 258692
rect 356756 258680 356762 258732
rect 159450 257320 159456 257372
rect 159508 257360 159514 257372
rect 177390 257360 177396 257372
rect 159508 257332 177396 257360
rect 159508 257320 159514 257332
rect 177390 257320 177396 257332
rect 177448 257320 177454 257372
rect 307662 257320 307668 257372
rect 307720 257360 307726 257372
rect 376846 257360 376852 257372
rect 307720 257332 376852 257360
rect 307720 257320 307726 257332
rect 376846 257320 376852 257332
rect 376904 257320 376910 257372
rect 187602 257048 187608 257100
rect 187660 257088 187666 257100
rect 188430 257088 188436 257100
rect 187660 257060 188436 257088
rect 187660 257048 187666 257060
rect 188430 257048 188436 257060
rect 188488 257048 188494 257100
rect 177942 256776 177948 256828
rect 178000 256816 178006 256828
rect 180794 256816 180800 256828
rect 178000 256788 180800 256816
rect 178000 256776 178006 256788
rect 180794 256776 180800 256788
rect 180852 256776 180858 256828
rect 196618 256776 196624 256828
rect 196676 256816 196682 256828
rect 197170 256816 197176 256828
rect 196676 256788 197176 256816
rect 196676 256776 196682 256788
rect 197170 256776 197176 256788
rect 197228 256816 197234 256828
rect 198090 256816 198096 256828
rect 197228 256788 198096 256816
rect 197228 256776 197234 256788
rect 198090 256776 198096 256788
rect 198148 256776 198154 256828
rect 160094 256708 160100 256760
rect 160152 256748 160158 256760
rect 186130 256748 186136 256760
rect 160152 256720 186136 256748
rect 160152 256708 160158 256720
rect 186130 256708 186136 256720
rect 186188 256748 186194 256760
rect 197446 256748 197452 256760
rect 186188 256720 197452 256748
rect 186188 256708 186194 256720
rect 197446 256708 197452 256720
rect 197504 256708 197510 256760
rect 246022 256708 246028 256760
rect 246080 256748 246086 256760
rect 262122 256748 262128 256760
rect 246080 256720 262128 256748
rect 246080 256708 246086 256720
rect 262122 256708 262128 256720
rect 262180 256708 262186 256760
rect 269022 256708 269028 256760
rect 269080 256748 269086 256760
rect 306558 256748 306564 256760
rect 269080 256720 306564 256748
rect 269080 256708 269086 256720
rect 306558 256708 306564 256720
rect 306616 256748 306622 256760
rect 307662 256748 307668 256760
rect 306616 256720 307668 256748
rect 306616 256708 306622 256720
rect 307662 256708 307668 256720
rect 307720 256708 307726 256760
rect 173158 256640 173164 256692
rect 173216 256680 173222 256692
rect 197354 256680 197360 256692
rect 173216 256652 197360 256680
rect 173216 256640 173222 256652
rect 197354 256640 197360 256652
rect 197412 256640 197418 256692
rect 245930 256640 245936 256692
rect 245988 256680 245994 256692
rect 259546 256680 259552 256692
rect 245988 256652 259552 256680
rect 245988 256640 245994 256652
rect 259546 256640 259552 256652
rect 259604 256680 259610 256692
rect 260742 256680 260748 256692
rect 259604 256652 260748 256680
rect 259604 256640 259610 256652
rect 260742 256640 260748 256652
rect 260800 256640 260806 256692
rect 61746 255960 61752 256012
rect 61804 256000 61810 256012
rect 66990 256000 66996 256012
rect 61804 255972 66996 256000
rect 61804 255960 61810 255972
rect 66990 255960 66996 255972
rect 67048 255960 67054 256012
rect 260742 255960 260748 256012
rect 260800 256000 260806 256012
rect 310606 256000 310612 256012
rect 260800 255972 310612 256000
rect 260800 255960 260806 255972
rect 310606 255960 310612 255972
rect 310664 256000 310670 256012
rect 379514 256000 379520 256012
rect 310664 255972 379520 256000
rect 310664 255960 310670 255972
rect 379514 255960 379520 255972
rect 379572 255960 379578 256012
rect 173710 255348 173716 255400
rect 173768 255388 173774 255400
rect 176654 255388 176660 255400
rect 173768 255360 176660 255388
rect 173768 255348 173774 255360
rect 176654 255348 176660 255360
rect 176712 255348 176718 255400
rect 58986 255280 58992 255332
rect 59044 255320 59050 255332
rect 66806 255320 66812 255332
rect 59044 255292 66812 255320
rect 59044 255280 59050 255292
rect 66806 255280 66812 255292
rect 66864 255280 66870 255332
rect 158806 255280 158812 255332
rect 158864 255320 158870 255332
rect 173802 255320 173808 255332
rect 158864 255292 173808 255320
rect 158864 255280 158870 255292
rect 173802 255280 173808 255292
rect 173860 255280 173866 255332
rect 3142 255212 3148 255264
rect 3200 255252 3206 255264
rect 18598 255252 18604 255264
rect 3200 255224 18604 255252
rect 3200 255212 3206 255224
rect 18598 255212 18604 255224
rect 18656 255212 18662 255264
rect 158714 255212 158720 255264
rect 158772 255252 158778 255264
rect 166994 255252 167000 255264
rect 158772 255224 167000 255252
rect 158772 255212 158778 255224
rect 166994 255212 167000 255224
rect 167052 255212 167058 255264
rect 176672 255252 176700 255348
rect 186222 255280 186228 255332
rect 186280 255320 186286 255332
rect 187786 255320 187792 255332
rect 186280 255292 187792 255320
rect 186280 255280 186286 255292
rect 187786 255280 187792 255292
rect 187844 255320 187850 255332
rect 197446 255320 197452 255332
rect 187844 255292 197452 255320
rect 187844 255280 187850 255292
rect 197446 255280 197452 255292
rect 197504 255280 197510 255332
rect 197354 255252 197360 255264
rect 176672 255224 197360 255252
rect 197354 255212 197360 255224
rect 197412 255212 197418 255264
rect 245930 255212 245936 255264
rect 245988 255252 245994 255264
rect 258166 255252 258172 255264
rect 245988 255224 258172 255252
rect 245988 255212 245994 255224
rect 258166 255212 258172 255224
rect 258224 255212 258230 255264
rect 166994 254532 167000 254584
rect 167052 254572 167058 254584
rect 191282 254572 191288 254584
rect 167052 254544 191288 254572
rect 167052 254532 167058 254544
rect 191282 254532 191288 254544
rect 191340 254532 191346 254584
rect 246942 254532 246948 254584
rect 247000 254572 247006 254584
rect 582926 254572 582932 254584
rect 247000 254544 582932 254572
rect 247000 254532 247006 254544
rect 582926 254532 582932 254544
rect 582984 254532 582990 254584
rect 245470 253852 245476 253904
rect 245528 253892 245534 253904
rect 269022 253892 269028 253904
rect 245528 253864 269028 253892
rect 245528 253852 245534 253864
rect 269022 253852 269028 253864
rect 269080 253852 269086 253904
rect 60366 253240 60372 253292
rect 60424 253280 60430 253292
rect 66898 253280 66904 253292
rect 60424 253252 66904 253280
rect 60424 253240 60430 253252
rect 66898 253240 66904 253252
rect 66956 253240 66962 253292
rect 160830 253172 160836 253224
rect 160888 253212 160894 253224
rect 164878 253212 164884 253224
rect 160888 253184 164884 253212
rect 160888 253172 160894 253184
rect 164878 253172 164884 253184
rect 164936 253172 164942 253224
rect 300762 253172 300768 253224
rect 300820 253212 300826 253224
rect 341518 253212 341524 253224
rect 300820 253184 341524 253212
rect 300820 253172 300826 253184
rect 341518 253172 341524 253184
rect 341576 253172 341582 253224
rect 60550 252968 60556 253020
rect 60608 253008 60614 253020
rect 66990 253008 66996 253020
rect 60608 252980 66996 253008
rect 60608 252968 60614 252980
rect 66990 252968 66996 252980
rect 67048 253008 67054 253020
rect 67358 253008 67364 253020
rect 67048 252980 67364 253008
rect 67048 252968 67054 252980
rect 67358 252968 67364 252980
rect 67416 252968 67422 253020
rect 158714 252560 158720 252612
rect 158772 252600 158778 252612
rect 176010 252600 176016 252612
rect 158772 252572 176016 252600
rect 158772 252560 158778 252572
rect 176010 252560 176016 252572
rect 176068 252560 176074 252612
rect 193030 252560 193036 252612
rect 193088 252600 193094 252612
rect 197354 252600 197360 252612
rect 193088 252572 197360 252600
rect 193088 252560 193094 252572
rect 197354 252560 197360 252572
rect 197412 252560 197418 252612
rect 245470 252560 245476 252612
rect 245528 252600 245534 252612
rect 299658 252600 299664 252612
rect 245528 252572 299664 252600
rect 245528 252560 245534 252572
rect 299658 252560 299664 252572
rect 299716 252600 299722 252612
rect 300762 252600 300768 252612
rect 299716 252572 300768 252600
rect 299716 252560 299722 252572
rect 300762 252560 300768 252572
rect 300820 252560 300826 252612
rect 165154 252492 165160 252544
rect 165212 252532 165218 252544
rect 166534 252532 166540 252544
rect 165212 252504 166540 252532
rect 165212 252492 165218 252504
rect 166534 252492 166540 252504
rect 166592 252492 166598 252544
rect 176562 252492 176568 252544
rect 176620 252532 176626 252544
rect 178034 252532 178040 252544
rect 176620 252504 178040 252532
rect 176620 252492 176626 252504
rect 178034 252492 178040 252504
rect 178092 252492 178098 252544
rect 245930 252492 245936 252544
rect 245988 252532 245994 252544
rect 251358 252532 251364 252544
rect 245988 252504 251364 252532
rect 245988 252492 245994 252504
rect 251358 252492 251364 252504
rect 251416 252532 251422 252544
rect 252462 252532 252468 252544
rect 251416 252504 252468 252532
rect 251416 252492 251422 252504
rect 252462 252492 252468 252504
rect 252520 252492 252526 252544
rect 187142 251880 187148 251932
rect 187200 251920 187206 251932
rect 194042 251920 194048 251932
rect 187200 251892 194048 251920
rect 187200 251880 187206 251892
rect 194042 251880 194048 251892
rect 194100 251880 194106 251932
rect 173802 251812 173808 251864
rect 173860 251852 173866 251864
rect 191650 251852 191656 251864
rect 173860 251824 191656 251852
rect 173860 251812 173866 251824
rect 191650 251812 191656 251824
rect 191708 251852 191714 251864
rect 195790 251852 195796 251864
rect 191708 251824 195796 251852
rect 191708 251812 191714 251824
rect 195790 251812 195796 251824
rect 195848 251852 195854 251864
rect 197354 251852 197360 251864
rect 195848 251824 197360 251852
rect 195848 251812 195854 251824
rect 197354 251812 197360 251824
rect 197412 251812 197418 251864
rect 252462 251812 252468 251864
rect 252520 251852 252526 251864
rect 566458 251852 566464 251864
rect 252520 251824 566464 251852
rect 252520 251812 252526 251824
rect 566458 251812 566464 251824
rect 566516 251812 566522 251864
rect 168282 251132 168288 251184
rect 168340 251172 168346 251184
rect 169294 251172 169300 251184
rect 168340 251144 169300 251172
rect 168340 251132 168346 251144
rect 169294 251132 169300 251144
rect 169352 251132 169358 251184
rect 179322 250520 179328 250572
rect 179380 250560 179386 250572
rect 187050 250560 187056 250572
rect 179380 250532 187056 250560
rect 179380 250520 179386 250532
rect 187050 250520 187056 250532
rect 187108 250520 187114 250572
rect 160738 250452 160744 250504
rect 160796 250492 160802 250504
rect 184842 250492 184848 250504
rect 160796 250464 184848 250492
rect 160796 250452 160802 250464
rect 184842 250452 184848 250464
rect 184900 250452 184906 250504
rect 309042 250452 309048 250504
rect 309100 250492 309106 250504
rect 340138 250492 340144 250504
rect 309100 250464 340144 250492
rect 309100 250452 309106 250464
rect 340138 250452 340144 250464
rect 340196 250452 340202 250504
rect 60550 249840 60556 249892
rect 60608 249880 60614 249892
rect 66898 249880 66904 249892
rect 60608 249852 66904 249880
rect 60608 249840 60614 249852
rect 66898 249840 66904 249852
rect 66956 249840 66962 249892
rect 195698 249840 195704 249892
rect 195756 249880 195762 249892
rect 197906 249880 197912 249892
rect 195756 249852 197912 249880
rect 195756 249840 195762 249852
rect 197906 249840 197912 249852
rect 197964 249840 197970 249892
rect 63126 249772 63132 249824
rect 63184 249812 63190 249824
rect 66806 249812 66812 249824
rect 63184 249784 66812 249812
rect 63184 249772 63190 249784
rect 66806 249772 66812 249784
rect 66864 249772 66870 249824
rect 187234 249772 187240 249824
rect 187292 249812 187298 249824
rect 197354 249812 197360 249824
rect 187292 249784 197360 249812
rect 187292 249772 187298 249784
rect 197354 249772 197360 249784
rect 197412 249772 197418 249824
rect 245746 249772 245752 249824
rect 245804 249812 245810 249824
rect 248598 249812 248604 249824
rect 245804 249784 248604 249812
rect 245804 249772 245810 249784
rect 248598 249772 248604 249784
rect 248656 249812 248662 249824
rect 307846 249812 307852 249824
rect 248656 249784 307852 249812
rect 248656 249772 248662 249784
rect 307846 249772 307852 249784
rect 307904 249812 307910 249824
rect 309042 249812 309048 249824
rect 307904 249784 309048 249812
rect 307904 249772 307910 249784
rect 309042 249772 309048 249784
rect 309100 249772 309106 249824
rect 181530 249704 181536 249756
rect 181588 249744 181594 249756
rect 183462 249744 183468 249756
rect 181588 249716 183468 249744
rect 181588 249704 181594 249716
rect 183462 249704 183468 249716
rect 183520 249704 183526 249756
rect 193858 249704 193864 249756
rect 193916 249744 193922 249756
rect 194502 249744 194508 249756
rect 193916 249716 194508 249744
rect 193916 249704 193922 249716
rect 194502 249704 194508 249716
rect 194560 249704 194566 249756
rect 245930 249500 245936 249552
rect 245988 249540 245994 249552
rect 249794 249540 249800 249552
rect 245988 249512 249800 249540
rect 245988 249500 245994 249512
rect 249794 249500 249800 249512
rect 249852 249500 249858 249552
rect 295978 249024 295984 249076
rect 296036 249064 296042 249076
rect 300854 249064 300860 249076
rect 296036 249036 300860 249064
rect 296036 249024 296042 249036
rect 300854 249024 300860 249036
rect 300912 249024 300918 249076
rect 194502 248684 194508 248736
rect 194560 248724 194566 248736
rect 197446 248724 197452 248736
rect 194560 248696 197452 248724
rect 194560 248684 194566 248696
rect 197446 248684 197452 248696
rect 197504 248684 197510 248736
rect 245930 248616 245936 248668
rect 245988 248656 245994 248668
rect 249978 248656 249984 248668
rect 245988 248628 249984 248656
rect 245988 248616 245994 248628
rect 249978 248616 249984 248628
rect 250036 248616 250042 248668
rect 158806 248480 158812 248532
rect 158864 248520 158870 248532
rect 176562 248520 176568 248532
rect 158864 248492 176568 248520
rect 158864 248480 158870 248492
rect 176562 248480 176568 248492
rect 176620 248480 176626 248532
rect 158714 248412 158720 248464
rect 158772 248452 158778 248464
rect 180702 248452 180708 248464
rect 158772 248424 180708 248452
rect 158772 248412 158778 248424
rect 180702 248412 180708 248424
rect 180760 248452 180766 248464
rect 182818 248452 182824 248464
rect 180760 248424 182824 248452
rect 180760 248412 180766 248424
rect 182818 248412 182824 248424
rect 182876 248412 182882 248464
rect 183462 248412 183468 248464
rect 183520 248452 183526 248464
rect 197354 248452 197360 248464
rect 183520 248424 197360 248452
rect 183520 248412 183526 248424
rect 197354 248412 197360 248424
rect 197412 248412 197418 248464
rect 169754 248344 169760 248396
rect 169812 248384 169818 248396
rect 185670 248384 185676 248396
rect 169812 248356 185676 248384
rect 169812 248344 169818 248356
rect 185670 248344 185676 248356
rect 185728 248344 185734 248396
rect 246942 247732 246948 247784
rect 247000 247772 247006 247784
rect 251358 247772 251364 247784
rect 247000 247744 251364 247772
rect 247000 247732 247006 247744
rect 251358 247732 251364 247744
rect 251416 247732 251422 247784
rect 329742 247732 329748 247784
rect 329800 247772 329806 247784
rect 354030 247772 354036 247784
rect 329800 247744 354036 247772
rect 329800 247732 329806 247744
rect 354030 247732 354036 247744
rect 354088 247732 354094 247784
rect 189718 247664 189724 247716
rect 189776 247704 189782 247716
rect 195698 247704 195704 247716
rect 189776 247676 195704 247704
rect 189776 247664 189782 247676
rect 195698 247664 195704 247676
rect 195756 247664 195762 247716
rect 244550 247664 244556 247716
rect 244608 247704 244614 247716
rect 264330 247704 264336 247716
rect 244608 247676 264336 247704
rect 244608 247664 244614 247676
rect 264330 247664 264336 247676
rect 264388 247664 264394 247716
rect 326338 247664 326344 247716
rect 326396 247704 326402 247716
rect 353294 247704 353300 247716
rect 326396 247676 353300 247704
rect 326396 247664 326402 247676
rect 353294 247664 353300 247676
rect 353352 247664 353358 247716
rect 162118 247460 162124 247512
rect 162176 247500 162182 247512
rect 168374 247500 168380 247512
rect 162176 247472 168380 247500
rect 162176 247460 162182 247472
rect 168374 247460 168380 247472
rect 168432 247460 168438 247512
rect 191742 247120 191748 247172
rect 191800 247160 191806 247172
rect 192754 247160 192760 247172
rect 191800 247132 192760 247160
rect 191800 247120 191806 247132
rect 192754 247120 192760 247132
rect 192812 247120 192818 247172
rect 52362 247052 52368 247104
rect 52420 247092 52426 247104
rect 66898 247092 66904 247104
rect 52420 247064 66904 247092
rect 52420 247052 52426 247064
rect 66898 247052 66904 247064
rect 66956 247052 66962 247104
rect 167730 247052 167736 247104
rect 167788 247092 167794 247104
rect 169754 247092 169760 247104
rect 167788 247064 169760 247092
rect 167788 247052 167794 247064
rect 169754 247052 169760 247064
rect 169812 247052 169818 247104
rect 192662 247052 192668 247104
rect 192720 247092 192726 247104
rect 197446 247092 197452 247104
rect 192720 247064 197452 247092
rect 192720 247052 192726 247064
rect 197446 247052 197452 247064
rect 197504 247052 197510 247104
rect 260190 247052 260196 247104
rect 260248 247092 260254 247104
rect 328454 247092 328460 247104
rect 260248 247064 328460 247092
rect 260248 247052 260254 247064
rect 328454 247052 328460 247064
rect 328512 247092 328518 247104
rect 329742 247092 329748 247104
rect 328512 247064 329748 247092
rect 328512 247052 328518 247064
rect 329742 247052 329748 247064
rect 329800 247052 329806 247104
rect 59170 246984 59176 247036
rect 59228 247024 59234 247036
rect 66806 247024 66812 247036
rect 59228 246996 66812 247024
rect 59228 246984 59234 246996
rect 66806 246984 66812 246996
rect 66864 246984 66870 247036
rect 184474 246984 184480 247036
rect 184532 247024 184538 247036
rect 197354 247024 197360 247036
rect 184532 246996 197360 247024
rect 184532 246984 184538 246996
rect 197354 246984 197360 246996
rect 197412 246984 197418 247036
rect 320634 246304 320640 246356
rect 320692 246344 320698 246356
rect 353938 246344 353944 246356
rect 320692 246316 353944 246344
rect 320692 246304 320698 246316
rect 353938 246304 353944 246316
rect 353996 246304 354002 246356
rect 197078 246100 197084 246152
rect 197136 246140 197142 246152
rect 199378 246140 199384 246152
rect 197136 246112 199384 246140
rect 197136 246100 197142 246112
rect 199378 246100 199384 246112
rect 199436 246100 199442 246152
rect 177850 245828 177856 245880
rect 177908 245868 177914 245880
rect 178678 245868 178684 245880
rect 177908 245840 178684 245868
rect 177908 245828 177914 245840
rect 178678 245828 178684 245840
rect 178736 245828 178742 245880
rect 162302 245692 162308 245744
rect 162360 245732 162366 245744
rect 166350 245732 166356 245744
rect 162360 245704 166356 245732
rect 162360 245692 162366 245704
rect 166350 245692 166356 245704
rect 166408 245692 166414 245744
rect 158806 245624 158812 245676
rect 158864 245664 158870 245676
rect 177850 245664 177856 245676
rect 158864 245636 177856 245664
rect 158864 245624 158870 245636
rect 177850 245624 177856 245636
rect 177908 245624 177914 245676
rect 245746 245624 245752 245676
rect 245804 245664 245810 245676
rect 266446 245664 266452 245676
rect 245804 245636 266452 245664
rect 245804 245624 245810 245636
rect 266446 245624 266452 245636
rect 266504 245664 266510 245676
rect 320266 245664 320272 245676
rect 266504 245636 320272 245664
rect 266504 245624 266510 245636
rect 320266 245624 320272 245636
rect 320324 245664 320330 245676
rect 320634 245664 320640 245676
rect 320324 245636 320640 245664
rect 320324 245624 320330 245636
rect 320634 245624 320640 245636
rect 320692 245624 320698 245676
rect 165062 244876 165068 244928
rect 165120 244916 165126 244928
rect 177482 244916 177488 244928
rect 165120 244888 177488 244916
rect 165120 244876 165126 244888
rect 177482 244876 177488 244888
rect 177540 244876 177546 244928
rect 184842 244876 184848 244928
rect 184900 244916 184906 244928
rect 197354 244916 197360 244928
rect 184900 244888 197360 244916
rect 184900 244876 184906 244888
rect 197354 244876 197360 244888
rect 197412 244876 197418 244928
rect 278130 244876 278136 244928
rect 278188 244916 278194 244928
rect 291838 244916 291844 244928
rect 278188 244888 291844 244916
rect 278188 244876 278194 244888
rect 291838 244876 291844 244888
rect 291896 244876 291902 244928
rect 303798 244876 303804 244928
rect 303856 244916 303862 244928
rect 342254 244916 342260 244928
rect 303856 244888 342260 244916
rect 303856 244876 303862 244888
rect 342254 244876 342260 244888
rect 342312 244876 342318 244928
rect 57882 244264 57888 244316
rect 57940 244304 57946 244316
rect 64506 244304 64512 244316
rect 57940 244276 64512 244304
rect 57940 244264 57946 244276
rect 64506 244264 64512 244276
rect 64564 244304 64570 244316
rect 66346 244304 66352 244316
rect 64564 244276 66352 244304
rect 64564 244264 64570 244276
rect 66346 244264 66352 244276
rect 66404 244264 66410 244316
rect 158714 244264 158720 244316
rect 158772 244304 158778 244316
rect 195606 244304 195612 244316
rect 158772 244276 195612 244304
rect 158772 244264 158778 244276
rect 195606 244264 195612 244276
rect 195664 244264 195670 244316
rect 250438 244264 250444 244316
rect 250496 244304 250502 244316
rect 303798 244304 303804 244316
rect 250496 244276 303804 244304
rect 250496 244264 250502 244276
rect 303798 244264 303804 244276
rect 303856 244264 303862 244316
rect 381538 244264 381544 244316
rect 381596 244304 381602 244316
rect 580166 244304 580172 244316
rect 381596 244276 580172 244304
rect 381596 244264 381602 244276
rect 580166 244264 580172 244276
rect 580224 244264 580230 244316
rect 182266 244196 182272 244248
rect 182324 244236 182330 244248
rect 197354 244236 197360 244248
rect 182324 244208 197360 244236
rect 182324 244196 182330 244208
rect 197354 244196 197360 244208
rect 197412 244196 197418 244248
rect 266354 244196 266360 244248
rect 266412 244236 266418 244248
rect 267642 244236 267648 244248
rect 266412 244208 267648 244236
rect 266412 244196 266418 244208
rect 267642 244196 267648 244208
rect 267700 244236 267706 244248
rect 267826 244236 267832 244248
rect 267700 244208 267832 244236
rect 267700 244196 267706 244208
rect 267826 244196 267832 244208
rect 267884 244196 267890 244248
rect 171962 243584 171968 243636
rect 172020 243624 172026 243636
rect 181622 243624 181628 243636
rect 172020 243596 181628 243624
rect 172020 243584 172026 243596
rect 181622 243584 181628 243596
rect 181680 243584 181686 243636
rect 156966 243516 156972 243568
rect 157024 243556 157030 243568
rect 168282 243556 168288 243568
rect 157024 243528 168288 243556
rect 157024 243516 157030 243528
rect 168282 243516 168288 243528
rect 168340 243556 168346 243568
rect 177390 243556 177396 243568
rect 168340 243528 177396 243556
rect 168340 243516 168346 243528
rect 177390 243516 177396 243528
rect 177448 243516 177454 243568
rect 181714 243516 181720 243568
rect 181772 243556 181778 243568
rect 197078 243556 197084 243568
rect 181772 243528 197084 243556
rect 181772 243516 181778 243528
rect 197078 243516 197084 243528
rect 197136 243516 197142 243568
rect 249058 243312 249064 243364
rect 249116 243352 249122 243364
rect 250070 243352 250076 243364
rect 249116 243324 250076 243352
rect 249116 243312 249122 243324
rect 250070 243312 250076 243324
rect 250128 243312 250134 243364
rect 158714 242904 158720 242956
rect 158772 242944 158778 242956
rect 164970 242944 164976 242956
rect 158772 242916 164976 242944
rect 158772 242904 158778 242916
rect 164970 242904 164976 242916
rect 165028 242904 165034 242956
rect 190270 242836 190276 242888
rect 190328 242876 190334 242888
rect 191098 242876 191104 242888
rect 190328 242848 191104 242876
rect 190328 242836 190334 242848
rect 191098 242836 191104 242848
rect 191156 242836 191162 242888
rect 300854 242156 300860 242208
rect 300912 242196 300918 242208
rect 352558 242196 352564 242208
rect 300912 242168 352564 242196
rect 300912 242156 300918 242168
rect 352558 242156 352564 242168
rect 352616 242156 352622 242208
rect 69750 241816 69756 241868
rect 69808 241856 69814 241868
rect 71038 241856 71044 241868
rect 69808 241828 71044 241856
rect 69808 241816 69814 241828
rect 71038 241816 71044 241828
rect 71096 241816 71102 241868
rect 156874 241544 156880 241596
rect 156932 241584 156938 241596
rect 184750 241584 184756 241596
rect 156932 241556 184756 241584
rect 156932 241544 156938 241556
rect 184750 241544 184756 241556
rect 184808 241544 184814 241596
rect 195974 241584 195980 241596
rect 190426 241556 195980 241584
rect 155310 241476 155316 241528
rect 155368 241516 155374 241528
rect 190426 241516 190454 241556
rect 195974 241544 195980 241556
rect 196032 241584 196038 241596
rect 196618 241584 196624 241596
rect 196032 241556 196624 241584
rect 196032 241544 196038 241556
rect 196618 241544 196624 241556
rect 196676 241544 196682 241596
rect 155368 241488 190454 241516
rect 155368 241476 155374 241488
rect 195514 241476 195520 241528
rect 195572 241516 195578 241528
rect 197814 241516 197820 241528
rect 195572 241488 197820 241516
rect 195572 241476 195578 241488
rect 197814 241476 197820 241488
rect 197872 241476 197878 241528
rect 246390 241476 246396 241528
rect 246448 241516 246454 241528
rect 247310 241516 247316 241528
rect 246448 241488 247316 241516
rect 246448 241476 246454 241488
rect 247310 241476 247316 241488
rect 247368 241516 247374 241528
rect 300854 241516 300860 241528
rect 247368 241488 300860 241516
rect 247368 241476 247374 241488
rect 300854 241476 300860 241488
rect 300912 241476 300918 241528
rect 3510 241408 3516 241460
rect 3568 241448 3574 241460
rect 25498 241448 25504 241460
rect 3568 241420 25504 241448
rect 3568 241408 3574 241420
rect 25498 241408 25504 241420
rect 25556 241408 25562 241460
rect 67818 241408 67824 241460
rect 67876 241448 67882 241460
rect 180058 241448 180064 241460
rect 67876 241420 180064 241448
rect 67876 241408 67882 241420
rect 180058 241408 180064 241420
rect 180116 241448 180122 241460
rect 180242 241448 180248 241460
rect 180116 241420 180248 241448
rect 180116 241408 180122 241420
rect 180242 241408 180248 241420
rect 180300 241408 180306 241460
rect 193950 241408 193956 241460
rect 194008 241448 194014 241460
rect 196986 241448 196992 241460
rect 194008 241420 196992 241448
rect 194008 241408 194014 241420
rect 196986 241408 196992 241420
rect 197044 241408 197050 241460
rect 288526 241408 288532 241460
rect 288584 241448 288590 241460
rect 291194 241448 291200 241460
rect 288584 241420 291200 241448
rect 288584 241408 288590 241420
rect 291194 241408 291200 241420
rect 291252 241408 291258 241460
rect 67450 240728 67456 240780
rect 67508 240768 67514 240780
rect 97902 240768 97908 240780
rect 67508 240740 97908 240768
rect 67508 240728 67514 240740
rect 97902 240728 97908 240740
rect 97960 240728 97966 240780
rect 111426 240728 111432 240780
rect 111484 240768 111490 240780
rect 136358 240768 136364 240780
rect 111484 240740 136364 240768
rect 111484 240728 111490 240740
rect 136358 240728 136364 240740
rect 136416 240728 136422 240780
rect 154482 240728 154488 240780
rect 154540 240768 154546 240780
rect 158530 240768 158536 240780
rect 154540 240740 158536 240768
rect 154540 240728 154546 240740
rect 158530 240728 158536 240740
rect 158588 240768 158594 240780
rect 164878 240768 164884 240780
rect 158588 240740 164884 240768
rect 158588 240728 158594 240740
rect 164878 240728 164884 240740
rect 164936 240728 164942 240780
rect 177850 240728 177856 240780
rect 177908 240768 177914 240780
rect 194318 240768 194324 240780
rect 177908 240740 194324 240768
rect 177908 240728 177914 240740
rect 194318 240728 194324 240740
rect 194376 240728 194382 240780
rect 200114 240320 200120 240372
rect 200172 240360 200178 240372
rect 200172 240332 204116 240360
rect 200172 240320 200178 240332
rect 192478 240252 192484 240304
rect 192536 240292 192542 240304
rect 192536 240264 201080 240292
rect 192536 240252 192542 240264
rect 201052 240168 201080 240264
rect 114554 240116 114560 240168
rect 114612 240156 114618 240168
rect 115198 240156 115204 240168
rect 114612 240128 115204 240156
rect 114612 240116 114618 240128
rect 115198 240116 115204 240128
rect 115256 240116 115262 240168
rect 126974 240116 126980 240168
rect 127032 240156 127038 240168
rect 127526 240156 127532 240168
rect 127032 240128 127532 240156
rect 127032 240116 127038 240128
rect 127526 240116 127532 240128
rect 127584 240116 127590 240168
rect 138014 240116 138020 240168
rect 138072 240156 138078 240168
rect 138566 240156 138572 240168
rect 138072 240128 138572 240156
rect 138072 240116 138078 240128
rect 138566 240116 138572 240128
rect 138624 240116 138630 240168
rect 195974 240116 195980 240168
rect 196032 240156 196038 240168
rect 200298 240156 200304 240168
rect 196032 240128 200304 240156
rect 196032 240116 196038 240128
rect 200298 240116 200304 240128
rect 200356 240116 200362 240168
rect 201034 240116 201040 240168
rect 201092 240116 201098 240168
rect 202138 240116 202144 240168
rect 202196 240156 202202 240168
rect 202782 240156 202788 240168
rect 202196 240128 202788 240156
rect 202196 240116 202202 240128
rect 202782 240116 202788 240128
rect 202840 240116 202846 240168
rect 204088 240156 204116 240332
rect 234586 240332 241514 240360
rect 207290 240156 207296 240168
rect 204088 240128 207296 240156
rect 207290 240116 207296 240128
rect 207348 240116 207354 240168
rect 213914 240116 213920 240168
rect 213972 240156 213978 240168
rect 221826 240156 221832 240168
rect 213972 240128 221832 240156
rect 213972 240116 213978 240128
rect 221826 240116 221832 240128
rect 221884 240116 221890 240168
rect 225322 240116 225328 240168
rect 225380 240156 225386 240168
rect 231946 240156 231952 240168
rect 225380 240128 231952 240156
rect 225380 240116 225386 240128
rect 231946 240116 231952 240128
rect 232004 240116 232010 240168
rect 233142 240116 233148 240168
rect 233200 240156 233206 240168
rect 234586 240156 234614 240332
rect 233200 240128 234614 240156
rect 241486 240156 241514 240332
rect 245654 240184 245660 240236
rect 245712 240224 245718 240236
rect 248598 240224 248604 240236
rect 245712 240196 248604 240224
rect 245712 240184 245718 240196
rect 248598 240184 248604 240196
rect 248656 240184 248662 240236
rect 288526 240156 288532 240168
rect 241486 240128 288532 240156
rect 233200 240116 233206 240128
rect 288526 240116 288532 240128
rect 288584 240116 288590 240168
rect 44082 240048 44088 240100
rect 44140 240088 44146 240100
rect 75914 240088 75920 240100
rect 44140 240060 75920 240088
rect 44140 240048 44146 240060
rect 75914 240048 75920 240060
rect 75972 240088 75978 240100
rect 76558 240088 76564 240100
rect 75972 240060 76564 240088
rect 75972 240048 75978 240060
rect 76558 240048 76564 240060
rect 76616 240048 76622 240100
rect 93210 240048 93216 240100
rect 93268 240088 93274 240100
rect 93762 240088 93768 240100
rect 93268 240060 93768 240088
rect 93268 240048 93274 240060
rect 93762 240048 93768 240060
rect 93820 240048 93826 240100
rect 96706 240048 96712 240100
rect 96764 240088 96770 240100
rect 97534 240088 97540 240100
rect 96764 240060 97540 240088
rect 96764 240048 96770 240060
rect 97534 240048 97540 240060
rect 97592 240048 97598 240100
rect 99650 240048 99656 240100
rect 99708 240088 99714 240100
rect 100662 240088 100668 240100
rect 99708 240060 100668 240088
rect 99708 240048 99714 240060
rect 100662 240048 100668 240060
rect 100720 240048 100726 240100
rect 102594 240048 102600 240100
rect 102652 240088 102658 240100
rect 103330 240088 103336 240100
rect 102652 240060 103336 240088
rect 102652 240048 102658 240060
rect 103330 240048 103336 240060
rect 103388 240048 103394 240100
rect 104066 240048 104072 240100
rect 104124 240088 104130 240100
rect 104802 240088 104808 240100
rect 104124 240060 104808 240088
rect 104124 240048 104130 240060
rect 104802 240048 104808 240060
rect 104860 240048 104866 240100
rect 110690 240048 110696 240100
rect 110748 240088 110754 240100
rect 218974 240088 218980 240100
rect 110748 240060 218980 240088
rect 110748 240048 110754 240060
rect 218974 240048 218980 240060
rect 219032 240048 219038 240100
rect 219894 240048 219900 240100
rect 219952 240088 219958 240100
rect 219952 240060 234614 240088
rect 219952 240048 219958 240060
rect 72602 239980 72608 240032
rect 72660 240020 72666 240032
rect 73062 240020 73068 240032
rect 72660 239992 73068 240020
rect 72660 239980 72666 239992
rect 73062 239980 73068 239992
rect 73120 239980 73126 240032
rect 119338 239980 119344 240032
rect 119396 240020 119402 240032
rect 119982 240020 119988 240032
rect 119396 239992 119988 240020
rect 119396 239980 119402 239992
rect 119982 239980 119988 239992
rect 120040 239980 120046 240032
rect 125962 239980 125968 240032
rect 126020 240020 126026 240032
rect 126790 240020 126796 240032
rect 126020 239992 126796 240020
rect 126020 239980 126026 239992
rect 126790 239980 126796 239992
rect 126848 239980 126854 240032
rect 131850 239980 131856 240032
rect 131908 240020 131914 240032
rect 132402 240020 132408 240032
rect 131908 239992 132408 240020
rect 131908 239980 131914 239992
rect 132402 239980 132408 239992
rect 132460 239980 132466 240032
rect 133322 239980 133328 240032
rect 133380 240020 133386 240032
rect 133782 240020 133788 240032
rect 133380 239992 133788 240020
rect 133380 239980 133386 239992
rect 133782 239980 133788 239992
rect 133840 239980 133846 240032
rect 149330 239980 149336 240032
rect 149388 240020 149394 240032
rect 150250 240020 150256 240032
rect 149388 239992 150256 240020
rect 149388 239980 149394 239992
rect 150250 239980 150256 239992
rect 150308 239980 150314 240032
rect 151998 239980 152004 240032
rect 152056 240020 152062 240032
rect 157334 240020 157340 240032
rect 152056 239992 157340 240020
rect 152056 239980 152062 239992
rect 157334 239980 157340 239992
rect 157392 239980 157398 240032
rect 197446 239980 197452 240032
rect 197504 240020 197510 240032
rect 201494 240020 201500 240032
rect 197504 239992 201500 240020
rect 197504 239980 197510 239992
rect 201494 239980 201500 239992
rect 201552 239980 201558 240032
rect 234586 240020 234614 240060
rect 244550 240020 244556 240032
rect 234586 239992 244556 240020
rect 244550 239980 244556 239992
rect 244608 239980 244614 240032
rect 79226 239912 79232 239964
rect 79284 239952 79290 239964
rect 79870 239952 79876 239964
rect 79284 239924 79876 239952
rect 79284 239912 79290 239924
rect 79870 239912 79876 239924
rect 79928 239912 79934 239964
rect 82170 239912 82176 239964
rect 82228 239952 82234 239964
rect 82722 239952 82728 239964
rect 82228 239924 82728 239952
rect 82228 239912 82234 239924
rect 82722 239912 82728 239924
rect 82780 239912 82786 239964
rect 117314 239912 117320 239964
rect 117372 239952 117378 239964
rect 117958 239952 117964 239964
rect 117372 239924 117964 239952
rect 117372 239912 117378 239924
rect 117958 239912 117964 239924
rect 118016 239912 118022 239964
rect 129826 239912 129832 239964
rect 129884 239952 129890 239964
rect 130470 239952 130476 239964
rect 129884 239924 130476 239952
rect 129884 239912 129890 239924
rect 130470 239912 130476 239924
rect 130528 239912 130534 239964
rect 132586 239912 132592 239964
rect 132644 239952 132650 239964
rect 133414 239952 133420 239964
rect 132644 239924 133420 239952
rect 132644 239912 132650 239924
rect 133414 239912 133420 239924
rect 133472 239912 133478 239964
rect 150802 239912 150808 239964
rect 150860 239952 150866 239964
rect 154482 239952 154488 239964
rect 150860 239924 154488 239952
rect 150860 239912 150866 239924
rect 154482 239912 154488 239924
rect 154540 239912 154546 239964
rect 85850 239844 85856 239896
rect 85908 239884 85914 239896
rect 86862 239884 86868 239896
rect 85908 239856 86868 239884
rect 85908 239844 85914 239856
rect 86862 239844 86868 239856
rect 86920 239844 86926 239896
rect 130378 239776 130384 239828
rect 130436 239816 130442 239828
rect 131022 239816 131028 239828
rect 130436 239788 131028 239816
rect 130436 239776 130442 239788
rect 131022 239776 131028 239788
rect 131080 239776 131086 239828
rect 112162 239640 112168 239692
rect 112220 239680 112226 239692
rect 112990 239680 112996 239692
rect 112220 239652 112996 239680
rect 112220 239640 112226 239652
rect 112990 239640 112996 239652
rect 113048 239640 113054 239692
rect 201494 239640 201500 239692
rect 201552 239680 201558 239692
rect 202414 239680 202420 239692
rect 201552 239652 202420 239680
rect 201552 239640 201558 239652
rect 202414 239640 202420 239652
rect 202472 239640 202478 239692
rect 116578 239504 116584 239556
rect 116636 239544 116642 239556
rect 117130 239544 117136 239556
rect 116636 239516 117136 239544
rect 116636 239504 116642 239516
rect 117130 239504 117136 239516
rect 117188 239504 117194 239556
rect 120810 239504 120816 239556
rect 120868 239544 120874 239556
rect 121362 239544 121368 239556
rect 120868 239516 121368 239544
rect 120868 239504 120874 239516
rect 121362 239504 121368 239516
rect 121420 239504 121426 239556
rect 108942 239436 108948 239488
rect 109000 239476 109006 239488
rect 129550 239476 129556 239488
rect 109000 239448 129556 239476
rect 109000 239436 109006 239448
rect 129550 239436 129556 239448
rect 129608 239436 129614 239488
rect 74074 239368 74080 239420
rect 74132 239408 74138 239420
rect 111058 239408 111064 239420
rect 74132 239380 111064 239408
rect 74132 239368 74138 239380
rect 111058 239368 111064 239380
rect 111116 239368 111122 239420
rect 141418 239368 141424 239420
rect 141476 239408 141482 239420
rect 141970 239408 141976 239420
rect 141476 239380 141976 239408
rect 141476 239368 141482 239380
rect 141970 239368 141976 239380
rect 142028 239368 142034 239420
rect 144178 239368 144184 239420
rect 144236 239408 144242 239420
rect 144822 239408 144828 239420
rect 144236 239380 144828 239408
rect 144236 239368 144242 239380
rect 144822 239368 144828 239380
rect 144880 239368 144886 239420
rect 145006 239368 145012 239420
rect 145064 239408 145070 239420
rect 145742 239408 145748 239420
rect 145064 239380 145748 239408
rect 145064 239368 145070 239380
rect 145742 239368 145748 239380
rect 145800 239368 145806 239420
rect 311986 239368 311992 239420
rect 312044 239408 312050 239420
rect 334066 239408 334072 239420
rect 312044 239380 334072 239408
rect 312044 239368 312050 239380
rect 334066 239368 334072 239380
rect 334124 239368 334130 239420
rect 95970 239232 95976 239284
rect 96028 239272 96034 239284
rect 96522 239272 96528 239284
rect 96028 239244 96528 239272
rect 96028 239232 96034 239244
rect 96522 239232 96528 239244
rect 96580 239232 96586 239284
rect 105538 239232 105544 239284
rect 105596 239272 105602 239284
rect 106182 239272 106188 239284
rect 105596 239244 106188 239272
rect 105596 239232 105602 239244
rect 106182 239232 106188 239244
rect 106240 239232 106246 239284
rect 128722 239232 128728 239284
rect 128780 239272 128786 239284
rect 129642 239272 129648 239284
rect 128780 239244 129648 239272
rect 128780 239232 128786 239244
rect 129642 239232 129648 239244
rect 129700 239232 129706 239284
rect 135530 239232 135536 239284
rect 135588 239272 135594 239284
rect 136450 239272 136456 239284
rect 135588 239244 136456 239272
rect 135588 239232 135594 239244
rect 136450 239232 136456 239244
rect 136508 239232 136514 239284
rect 143534 239232 143540 239284
rect 143592 239272 143598 239284
rect 144270 239272 144276 239284
rect 143592 239244 144276 239272
rect 143592 239232 143598 239244
rect 144270 239232 144276 239244
rect 144328 239232 144334 239284
rect 153746 239232 153752 239284
rect 153804 239272 153810 239284
rect 154482 239272 154488 239284
rect 153804 239244 154488 239272
rect 153804 239232 153810 239244
rect 154482 239232 154488 239244
rect 154540 239232 154546 239284
rect 82630 238756 82636 238808
rect 82688 238796 82694 238808
rect 84838 238796 84844 238808
rect 82688 238768 84844 238796
rect 82688 238756 82694 238768
rect 84838 238756 84844 238768
rect 84896 238756 84902 238808
rect 214558 238756 214564 238808
rect 214616 238796 214622 238808
rect 221458 238796 221464 238808
rect 214616 238768 221464 238796
rect 214616 238756 214622 238768
rect 221458 238756 221464 238768
rect 221516 238756 221522 238808
rect 224862 238756 224868 238808
rect 224920 238796 224926 238808
rect 224920 238768 231854 238796
rect 224920 238756 224926 238768
rect 67910 238688 67916 238740
rect 67968 238728 67974 238740
rect 190178 238728 190184 238740
rect 67968 238700 190184 238728
rect 67968 238688 67974 238700
rect 190178 238688 190184 238700
rect 190236 238728 190242 238740
rect 200206 238728 200212 238740
rect 190236 238700 200212 238728
rect 190236 238688 190242 238700
rect 200206 238688 200212 238700
rect 200264 238688 200270 238740
rect 205542 238688 205548 238740
rect 205600 238728 205606 238740
rect 222286 238728 222292 238740
rect 205600 238700 222292 238728
rect 205600 238688 205606 238700
rect 222286 238688 222292 238700
rect 222344 238728 222350 238740
rect 223298 238728 223304 238740
rect 222344 238700 223304 238728
rect 222344 238688 222350 238700
rect 223298 238688 223304 238700
rect 223356 238688 223362 238740
rect 231826 238728 231854 238768
rect 237374 238756 237380 238808
rect 237432 238796 237438 238808
rect 311986 238796 311992 238808
rect 237432 238768 311992 238796
rect 237432 238756 237438 238768
rect 311986 238756 311992 238768
rect 312044 238756 312050 238808
rect 258074 238728 258080 238740
rect 231826 238700 258080 238728
rect 258074 238688 258080 238700
rect 258132 238688 258138 238740
rect 259638 238688 259644 238740
rect 259696 238728 259702 238740
rect 361482 238728 361488 238740
rect 259696 238700 361488 238728
rect 259696 238688 259702 238700
rect 361482 238688 361488 238700
rect 361540 238728 361546 238740
rect 381538 238728 381544 238740
rect 361540 238700 381544 238728
rect 361540 238688 361546 238700
rect 381538 238688 381544 238700
rect 381596 238688 381602 238740
rect 129550 238620 129556 238672
rect 129608 238660 129614 238672
rect 219894 238660 219900 238672
rect 129608 238632 219900 238660
rect 129608 238620 129614 238632
rect 219894 238620 219900 238632
rect 219952 238620 219958 238672
rect 225782 238620 225788 238672
rect 225840 238660 225846 238672
rect 233142 238660 233148 238672
rect 225840 238632 233148 238660
rect 225840 238620 225846 238632
rect 233142 238620 233148 238632
rect 233200 238620 233206 238672
rect 240318 238620 240324 238672
rect 240376 238660 240382 238672
rect 240778 238660 240784 238672
rect 240376 238632 240784 238660
rect 240376 238620 240382 238632
rect 240778 238620 240784 238632
rect 240836 238660 240842 238672
rect 250438 238660 250444 238672
rect 240836 238632 250444 238660
rect 240836 238620 240842 238632
rect 250438 238620 250444 238632
rect 250496 238620 250502 238672
rect 151906 238552 151912 238604
rect 151964 238592 151970 238604
rect 157978 238592 157984 238604
rect 151964 238564 157984 238592
rect 151964 238552 151970 238564
rect 157978 238552 157984 238564
rect 158036 238552 158042 238604
rect 215662 238212 215668 238264
rect 215720 238252 215726 238264
rect 216490 238252 216496 238264
rect 215720 238224 216496 238252
rect 215720 238212 215726 238224
rect 216490 238212 216496 238224
rect 216548 238212 216554 238264
rect 63310 238008 63316 238060
rect 63368 238048 63374 238060
rect 69750 238048 69756 238060
rect 63368 238020 69756 238048
rect 63368 238008 63374 238020
rect 69750 238008 69756 238020
rect 69808 238008 69814 238060
rect 195238 238008 195244 238060
rect 195296 238048 195302 238060
rect 202322 238048 202328 238060
rect 195296 238020 202328 238048
rect 195296 238008 195302 238020
rect 202322 238008 202328 238020
rect 202380 238008 202386 238060
rect 202322 237668 202328 237720
rect 202380 237708 202386 237720
rect 204070 237708 204076 237720
rect 202380 237680 204076 237708
rect 202380 237668 202386 237680
rect 204070 237668 204076 237680
rect 204128 237668 204134 237720
rect 200206 237396 200212 237448
rect 200264 237436 200270 237448
rect 200758 237436 200764 237448
rect 200264 237408 200764 237436
rect 200264 237396 200270 237408
rect 200758 237396 200764 237408
rect 200816 237396 200822 237448
rect 201494 237396 201500 237448
rect 201552 237436 201558 237448
rect 202598 237436 202604 237448
rect 201552 237408 202604 237436
rect 201552 237396 201558 237408
rect 202598 237396 202604 237408
rect 202656 237396 202662 237448
rect 223390 237396 223396 237448
rect 223448 237436 223454 237448
rect 229646 237436 229652 237448
rect 223448 237408 229652 237436
rect 223448 237396 223454 237408
rect 229646 237396 229652 237408
rect 229704 237396 229710 237448
rect 14550 237328 14556 237380
rect 14608 237368 14614 237380
rect 55030 237368 55036 237380
rect 14608 237340 55036 237368
rect 14608 237328 14614 237340
rect 55030 237328 55036 237340
rect 55088 237368 55094 237380
rect 138014 237368 138020 237380
rect 55088 237340 138020 237368
rect 55088 237328 55094 237340
rect 138014 237328 138020 237340
rect 138072 237328 138078 237380
rect 138106 237328 138112 237380
rect 138164 237368 138170 237380
rect 156966 237368 156972 237380
rect 138164 237340 156972 237368
rect 138164 237328 138170 237340
rect 156966 237328 156972 237340
rect 157024 237328 157030 237380
rect 197078 237328 197084 237380
rect 197136 237368 197142 237380
rect 207658 237368 207664 237380
rect 197136 237340 207664 237368
rect 197136 237328 197142 237340
rect 207658 237328 207664 237340
rect 207716 237328 207722 237380
rect 241790 237328 241796 237380
rect 241848 237368 241854 237380
rect 242250 237368 242256 237380
rect 241848 237340 242256 237368
rect 241848 237328 241854 237340
rect 242250 237328 242256 237340
rect 242308 237368 242314 237380
rect 249058 237368 249064 237380
rect 242308 237340 249064 237368
rect 242308 237328 242314 237340
rect 249058 237328 249064 237340
rect 249116 237328 249122 237380
rect 242158 237260 242164 237312
rect 242216 237300 242222 237312
rect 252554 237300 252560 237312
rect 242216 237272 252560 237300
rect 242216 237260 242222 237272
rect 252554 237260 252560 237272
rect 252612 237260 252618 237312
rect 239398 237192 239404 237244
rect 239456 237232 239462 237244
rect 246298 237232 246304 237244
rect 239456 237204 246304 237232
rect 239456 237192 239462 237204
rect 246298 237192 246304 237204
rect 246356 237192 246362 237244
rect 157334 237124 157340 237176
rect 157392 237164 157398 237176
rect 162210 237164 162216 237176
rect 157392 237136 162216 237164
rect 157392 237124 157398 237136
rect 162210 237124 162216 237136
rect 162268 237124 162274 237176
rect 207014 236716 207020 236768
rect 207072 236756 207078 236768
rect 240686 236756 240692 236768
rect 207072 236728 240692 236756
rect 207072 236716 207078 236728
rect 240686 236716 240692 236728
rect 240744 236716 240750 236768
rect 64598 236648 64604 236700
rect 64656 236688 64662 236700
rect 73798 236688 73804 236700
rect 64656 236660 73804 236688
rect 64656 236648 64662 236660
rect 73798 236648 73804 236660
rect 73856 236648 73862 236700
rect 78490 236648 78496 236700
rect 78548 236688 78554 236700
rect 88334 236688 88340 236700
rect 78548 236660 88340 236688
rect 78548 236648 78554 236660
rect 88334 236648 88340 236660
rect 88392 236648 88398 236700
rect 97902 236648 97908 236700
rect 97960 236688 97966 236700
rect 239214 236688 239220 236700
rect 97960 236660 239220 236688
rect 97960 236648 97966 236660
rect 239214 236648 239220 236660
rect 239272 236648 239278 236700
rect 88334 235968 88340 236020
rect 88392 236008 88398 236020
rect 88978 236008 88984 236020
rect 88392 235980 88984 236008
rect 88392 235968 88398 235980
rect 88978 235968 88984 235980
rect 89036 235968 89042 236020
rect 162118 235968 162124 236020
rect 162176 236008 162182 236020
rect 164142 236008 164148 236020
rect 162176 235980 164148 236008
rect 162176 235968 162182 235980
rect 164142 235968 164148 235980
rect 164200 235968 164206 236020
rect 76098 235900 76104 235952
rect 76156 235940 76162 235952
rect 121638 235940 121644 235952
rect 76156 235912 121644 235940
rect 76156 235900 76162 235912
rect 121638 235900 121644 235912
rect 121696 235900 121702 235952
rect 147214 235900 147220 235952
rect 147272 235940 147278 235952
rect 147272 235912 180794 235940
rect 147272 235900 147278 235912
rect 136358 235832 136364 235884
rect 136416 235872 136422 235884
rect 155310 235872 155316 235884
rect 136416 235844 155316 235872
rect 136416 235832 136422 235844
rect 155310 235832 155316 235844
rect 155368 235832 155374 235884
rect 180766 235872 180794 235912
rect 195606 235900 195612 235952
rect 195664 235940 195670 235952
rect 241238 235940 241244 235952
rect 195664 235912 241244 235940
rect 195664 235900 195670 235912
rect 241238 235900 241244 235912
rect 241296 235900 241302 235952
rect 182082 235872 182088 235884
rect 180766 235844 182088 235872
rect 182082 235832 182088 235844
rect 182140 235872 182146 235884
rect 203610 235872 203616 235884
rect 182140 235844 203616 235872
rect 182140 235832 182146 235844
rect 203610 235832 203616 235844
rect 203668 235832 203674 235884
rect 240870 235560 240876 235612
rect 240928 235600 240934 235612
rect 243262 235600 243268 235612
rect 240928 235572 243268 235600
rect 240928 235560 240934 235572
rect 243262 235560 243268 235572
rect 243320 235560 243326 235612
rect 11698 235220 11704 235272
rect 11756 235260 11762 235272
rect 52178 235260 52184 235272
rect 11756 235232 52184 235260
rect 11756 235220 11762 235232
rect 52178 235220 52184 235232
rect 52236 235220 52242 235272
rect 60366 235220 60372 235272
rect 60424 235260 60430 235272
rect 146202 235260 146208 235272
rect 60424 235232 146208 235260
rect 60424 235220 60430 235232
rect 146202 235220 146208 235232
rect 146260 235220 146266 235272
rect 157426 235220 157432 235272
rect 157484 235260 157490 235272
rect 166902 235260 166908 235272
rect 157484 235232 166908 235260
rect 157484 235220 157490 235232
rect 166902 235220 166908 235232
rect 166960 235260 166966 235272
rect 171870 235260 171876 235272
rect 166960 235232 171876 235260
rect 166960 235220 166966 235232
rect 171870 235220 171876 235232
rect 171928 235220 171934 235272
rect 227714 235220 227720 235272
rect 227772 235260 227778 235272
rect 228726 235260 228732 235272
rect 227772 235232 228732 235260
rect 227772 235220 227778 235232
rect 228726 235220 228732 235232
rect 228784 235260 228790 235272
rect 295978 235260 295984 235272
rect 228784 235232 295984 235260
rect 228784 235220 228790 235232
rect 295978 235220 295984 235232
rect 296036 235220 296042 235272
rect 207382 235084 207388 235136
rect 207440 235124 207446 235136
rect 209038 235124 209044 235136
rect 207440 235096 209044 235124
rect 207440 235084 207446 235096
rect 209038 235084 209044 235096
rect 209096 235084 209102 235136
rect 211798 234608 211804 234660
rect 211856 234648 211862 234660
rect 212534 234648 212540 234660
rect 211856 234620 212540 234648
rect 211856 234608 211862 234620
rect 212534 234608 212540 234620
rect 212592 234608 212598 234660
rect 295518 234608 295524 234660
rect 295576 234648 295582 234660
rect 295978 234648 295984 234660
rect 295576 234620 295984 234648
rect 295576 234608 295582 234620
rect 295978 234608 295984 234620
rect 296036 234608 296042 234660
rect 22738 234540 22744 234592
rect 22796 234580 22802 234592
rect 92474 234580 92480 234592
rect 22796 234552 92480 234580
rect 22796 234540 22802 234552
rect 92474 234540 92480 234552
rect 92532 234540 92538 234592
rect 145006 234540 145012 234592
rect 145064 234580 145070 234592
rect 237374 234580 237380 234592
rect 145064 234552 237380 234580
rect 145064 234540 145070 234552
rect 237374 234540 237380 234552
rect 237432 234540 237438 234592
rect 96706 234472 96712 234524
rect 96764 234512 96770 234524
rect 150434 234512 150440 234524
rect 96764 234484 150440 234512
rect 96764 234472 96770 234484
rect 150434 234472 150440 234484
rect 150492 234472 150498 234524
rect 200298 234472 200304 234524
rect 200356 234512 200362 234524
rect 270494 234512 270500 234524
rect 200356 234484 270500 234512
rect 200356 234472 200362 234484
rect 270494 234472 270500 234484
rect 270552 234512 270558 234524
rect 271230 234512 271236 234524
rect 270552 234484 271236 234512
rect 270552 234472 270558 234484
rect 271230 234472 271236 234484
rect 271288 234472 271294 234524
rect 92474 234132 92480 234184
rect 92532 234172 92538 234184
rect 93118 234172 93124 234184
rect 92532 234144 93124 234172
rect 92532 234132 92538 234144
rect 93118 234132 93124 234144
rect 93176 234132 93182 234184
rect 163498 233860 163504 233912
rect 163556 233900 163562 233912
rect 187234 233900 187240 233912
rect 163556 233872 187240 233900
rect 163556 233860 163562 233872
rect 187234 233860 187240 233872
rect 187292 233860 187298 233912
rect 127066 233180 127072 233232
rect 127124 233220 127130 233232
rect 227714 233220 227720 233232
rect 127124 233192 227720 233220
rect 127124 233180 127130 233192
rect 227714 233180 227720 233192
rect 227772 233180 227778 233232
rect 235350 233180 235356 233232
rect 235408 233220 235414 233232
rect 253934 233220 253940 233232
rect 235408 233192 253940 233220
rect 235408 233180 235414 233192
rect 253934 233180 253940 233192
rect 253992 233180 253998 233232
rect 143350 233112 143356 233164
rect 143408 233152 143414 233164
rect 157334 233152 157340 233164
rect 143408 233124 157340 233152
rect 143408 233112 143414 233124
rect 157334 233112 157340 233124
rect 157392 233112 157398 233164
rect 65886 232568 65892 232620
rect 65944 232608 65950 232620
rect 128998 232608 129004 232620
rect 65944 232580 129004 232608
rect 65944 232568 65950 232580
rect 128998 232568 129004 232580
rect 129056 232568 129062 232620
rect 224310 232568 224316 232620
rect 224368 232608 224374 232620
rect 273898 232608 273904 232620
rect 224368 232580 273904 232608
rect 224368 232568 224374 232580
rect 273898 232568 273904 232580
rect 273956 232568 273962 232620
rect 61746 232500 61752 232552
rect 61804 232540 61810 232552
rect 126238 232540 126244 232552
rect 61804 232512 126244 232540
rect 61804 232500 61810 232512
rect 126238 232500 126244 232512
rect 126296 232500 126302 232552
rect 208394 232500 208400 232552
rect 208452 232540 208458 232552
rect 223390 232540 223396 232552
rect 208452 232512 223396 232540
rect 208452 232500 208458 232512
rect 223390 232500 223396 232512
rect 223448 232500 223454 232552
rect 253934 232500 253940 232552
rect 253992 232540 253998 232552
rect 582742 232540 582748 232552
rect 253992 232512 582748 232540
rect 253992 232500 253998 232512
rect 582742 232500 582748 232512
rect 582800 232500 582806 232552
rect 126790 231752 126796 231804
rect 126848 231792 126854 231804
rect 175182 231792 175188 231804
rect 126848 231764 175188 231792
rect 126848 231752 126854 231764
rect 175182 231752 175188 231764
rect 175240 231752 175246 231804
rect 176010 231752 176016 231804
rect 176068 231792 176074 231804
rect 247310 231792 247316 231804
rect 176068 231764 247316 231792
rect 176068 231752 176074 231764
rect 247310 231752 247316 231764
rect 247368 231752 247374 231804
rect 140682 231684 140688 231736
rect 140740 231724 140746 231736
rect 167730 231724 167736 231736
rect 140740 231696 167736 231724
rect 140740 231684 140746 231696
rect 167730 231684 167736 231696
rect 167788 231684 167794 231736
rect 200574 231684 200580 231736
rect 200632 231724 200638 231736
rect 202138 231724 202144 231736
rect 200632 231696 202144 231724
rect 200632 231684 200638 231696
rect 202138 231684 202144 231696
rect 202196 231684 202202 231736
rect 218974 231684 218980 231736
rect 219032 231724 219038 231736
rect 267734 231724 267740 231736
rect 219032 231696 267740 231724
rect 219032 231684 219038 231696
rect 267734 231684 267740 231696
rect 267792 231724 267798 231736
rect 269022 231724 269028 231736
rect 267792 231696 269028 231724
rect 267792 231684 267798 231696
rect 269022 231684 269028 231696
rect 269080 231684 269086 231736
rect 74534 231072 74540 231124
rect 74592 231112 74598 231124
rect 138382 231112 138388 231124
rect 74592 231084 138388 231112
rect 74592 231072 74598 231084
rect 138382 231072 138388 231084
rect 138440 231072 138446 231124
rect 269022 231072 269028 231124
rect 269080 231112 269086 231124
rect 288618 231112 288624 231124
rect 269080 231084 288624 231112
rect 269080 231072 269086 231084
rect 288618 231072 288624 231084
rect 288676 231072 288682 231124
rect 204162 230936 204168 230988
rect 204220 230976 204226 230988
rect 210418 230976 210424 230988
rect 204220 230948 210424 230976
rect 204220 230936 204226 230948
rect 210418 230936 210424 230948
rect 210476 230936 210482 230988
rect 142154 230392 142160 230444
rect 142212 230432 142218 230444
rect 234062 230432 234068 230444
rect 142212 230404 234068 230432
rect 142212 230392 142218 230404
rect 234062 230392 234068 230404
rect 234120 230392 234126 230444
rect 275922 230392 275928 230444
rect 275980 230432 275986 230444
rect 276658 230432 276664 230444
rect 275980 230404 276664 230432
rect 275980 230392 275986 230404
rect 276658 230392 276664 230404
rect 276716 230392 276722 230444
rect 293954 230392 293960 230444
rect 294012 230432 294018 230444
rect 294598 230432 294604 230444
rect 294012 230404 294604 230432
rect 294012 230392 294018 230404
rect 294598 230392 294604 230404
rect 294656 230392 294662 230444
rect 150250 230324 150256 230376
rect 150308 230364 150314 230376
rect 157426 230364 157432 230376
rect 150308 230336 157432 230364
rect 150308 230324 150314 230336
rect 157426 230324 157432 230336
rect 157484 230324 157490 230376
rect 188338 230324 188344 230376
rect 188396 230364 188402 230376
rect 206278 230364 206284 230376
rect 188396 230336 206284 230364
rect 188396 230324 188402 230336
rect 206278 230324 206284 230336
rect 206336 230364 206342 230376
rect 206830 230364 206836 230376
rect 206336 230336 206836 230364
rect 206336 230324 206342 230336
rect 206830 230324 206836 230336
rect 206888 230324 206894 230376
rect 66070 229712 66076 229764
rect 66128 229752 66134 229764
rect 147490 229752 147496 229764
rect 66128 229724 147496 229752
rect 66128 229712 66134 229724
rect 147490 229712 147496 229724
rect 147548 229712 147554 229764
rect 167638 229712 167644 229764
rect 167696 229752 167702 229764
rect 184198 229752 184204 229764
rect 167696 229724 184204 229752
rect 167696 229712 167702 229724
rect 184198 229712 184204 229724
rect 184256 229712 184262 229764
rect 208486 229712 208492 229764
rect 208544 229752 208550 229764
rect 275922 229752 275928 229764
rect 208544 229724 275928 229752
rect 208544 229712 208550 229724
rect 275922 229712 275928 229724
rect 275980 229712 275986 229764
rect 287698 229712 287704 229764
rect 287756 229752 287762 229764
rect 306466 229752 306472 229764
rect 287756 229724 306472 229752
rect 287756 229712 287762 229724
rect 306466 229712 306472 229724
rect 306524 229712 306530 229764
rect 262950 229100 262956 229152
rect 263008 229140 263014 229152
rect 293954 229140 293960 229152
rect 263008 229112 293960 229140
rect 263008 229100 263014 229112
rect 293954 229100 293960 229112
rect 294012 229100 294018 229152
rect 86218 229032 86224 229084
rect 86276 229072 86282 229084
rect 158162 229072 158168 229084
rect 86276 229044 158168 229072
rect 86276 229032 86282 229044
rect 158162 229032 158168 229044
rect 158220 229032 158226 229084
rect 181622 229032 181628 229084
rect 181680 229072 181686 229084
rect 223758 229072 223764 229084
rect 181680 229044 223764 229072
rect 181680 229032 181686 229044
rect 223758 229032 223764 229044
rect 223816 229032 223822 229084
rect 110322 228964 110328 229016
rect 110380 229004 110386 229016
rect 156782 229004 156788 229016
rect 110380 228976 156788 229004
rect 110380 228964 110386 228976
rect 156782 228964 156788 228976
rect 156840 228964 156846 229016
rect 156598 228352 156604 228404
rect 156656 228392 156662 228404
rect 166442 228392 166448 228404
rect 156656 228364 166448 228392
rect 156656 228352 156662 228364
rect 166442 228352 166448 228364
rect 166500 228352 166506 228404
rect 234062 228352 234068 228404
rect 234120 228392 234126 228404
rect 277578 228392 277584 228404
rect 234120 228364 277584 228392
rect 234120 228352 234126 228364
rect 277578 228352 277584 228364
rect 277636 228352 277642 228404
rect 223758 227740 223764 227792
rect 223816 227780 223822 227792
rect 226978 227780 226984 227792
rect 223816 227752 226984 227780
rect 223816 227740 223822 227752
rect 226978 227740 226984 227752
rect 227036 227740 227042 227792
rect 229094 227740 229100 227792
rect 229152 227780 229158 227792
rect 231946 227780 231952 227792
rect 229152 227752 231952 227780
rect 229152 227740 229158 227752
rect 231946 227740 231952 227752
rect 232004 227780 232010 227792
rect 259362 227780 259368 227792
rect 232004 227752 259368 227780
rect 232004 227740 232010 227752
rect 259362 227740 259368 227752
rect 259420 227780 259426 227792
rect 260098 227780 260104 227792
rect 259420 227752 260104 227780
rect 259420 227740 259426 227752
rect 260098 227740 260104 227752
rect 260156 227740 260162 227792
rect 60550 227672 60556 227724
rect 60608 227712 60614 227724
rect 156598 227712 156604 227724
rect 60608 227684 156604 227712
rect 60608 227672 60614 227684
rect 156598 227672 156604 227684
rect 156656 227672 156662 227724
rect 187142 227672 187148 227724
rect 187200 227712 187206 227724
rect 243538 227712 243544 227724
rect 187200 227684 243544 227712
rect 187200 227672 187206 227684
rect 243538 227672 243544 227684
rect 243596 227672 243602 227724
rect 126238 227604 126244 227656
rect 126296 227644 126302 227656
rect 187694 227644 187700 227656
rect 126296 227616 187700 227644
rect 126296 227604 126302 227616
rect 187694 227604 187700 227616
rect 187752 227604 187758 227656
rect 302142 227060 302148 227112
rect 302200 227100 302206 227112
rect 302878 227100 302884 227112
rect 302200 227072 302884 227100
rect 302200 227060 302206 227072
rect 302878 227060 302884 227072
rect 302936 227060 302942 227112
rect 196618 226992 196624 227044
rect 196676 227032 196682 227044
rect 245838 227032 245844 227044
rect 196676 227004 245844 227032
rect 196676 226992 196682 227004
rect 245838 226992 245844 227004
rect 245896 226992 245902 227044
rect 302326 226992 302332 227044
rect 302384 227032 302390 227044
rect 316034 227032 316040 227044
rect 302384 227004 316040 227032
rect 302384 226992 302390 227004
rect 316034 226992 316040 227004
rect 316092 226992 316098 227044
rect 156598 226584 156604 226636
rect 156656 226624 156662 226636
rect 162302 226624 162308 226636
rect 156656 226596 162308 226624
rect 156656 226584 156662 226596
rect 162302 226584 162308 226596
rect 162360 226584 162366 226636
rect 187694 226312 187700 226364
rect 187752 226352 187758 226364
rect 188522 226352 188528 226364
rect 187752 226324 188528 226352
rect 187752 226312 187758 226324
rect 188522 226312 188528 226324
rect 188580 226312 188586 226364
rect 279602 226312 279608 226364
rect 279660 226352 279666 226364
rect 302326 226352 302332 226364
rect 279660 226324 302332 226352
rect 279660 226312 279666 226324
rect 302326 226312 302332 226324
rect 302384 226312 302390 226364
rect 103330 226244 103336 226296
rect 103388 226284 103394 226296
rect 184750 226284 184756 226296
rect 103388 226256 184756 226284
rect 103388 226244 103394 226256
rect 184750 226244 184756 226256
rect 184808 226244 184814 226296
rect 220998 226244 221004 226296
rect 221056 226284 221062 226296
rect 276014 226284 276020 226296
rect 221056 226256 276020 226284
rect 221056 226244 221062 226256
rect 276014 226244 276020 226256
rect 276072 226244 276078 226296
rect 142798 226176 142804 226228
rect 142856 226216 142862 226228
rect 156874 226216 156880 226228
rect 142856 226188 156880 226216
rect 142856 226176 142862 226188
rect 156874 226176 156880 226188
rect 156932 226176 156938 226228
rect 194042 226176 194048 226228
rect 194100 226216 194106 226228
rect 222838 226216 222844 226228
rect 194100 226188 222844 226216
rect 194100 226176 194106 226188
rect 222838 226176 222844 226188
rect 222896 226176 222902 226228
rect 276014 225564 276020 225616
rect 276072 225604 276078 225616
rect 287238 225604 287244 225616
rect 276072 225576 287244 225604
rect 276072 225564 276078 225576
rect 287238 225564 287244 225576
rect 287296 225564 287302 225616
rect 184750 224952 184756 225004
rect 184808 224992 184814 225004
rect 195146 224992 195152 225004
rect 184808 224964 195152 224992
rect 184808 224952 184814 224964
rect 195146 224952 195152 224964
rect 195204 224952 195210 225004
rect 84838 224884 84844 224936
rect 84896 224924 84902 224936
rect 189718 224924 189724 224936
rect 84896 224896 189724 224924
rect 84896 224884 84902 224896
rect 189718 224884 189724 224896
rect 189776 224884 189782 224936
rect 195238 224884 195244 224936
rect 195296 224924 195302 224936
rect 249794 224924 249800 224936
rect 195296 224896 249800 224924
rect 195296 224884 195302 224896
rect 249794 224884 249800 224896
rect 249852 224884 249858 224936
rect 126974 224816 126980 224868
rect 127032 224856 127038 224868
rect 227254 224856 227260 224868
rect 127032 224828 227260 224856
rect 127032 224816 127038 224828
rect 227254 224816 227260 224828
rect 227312 224816 227318 224868
rect 277578 224204 277584 224256
rect 277636 224244 277642 224256
rect 309134 224244 309140 224256
rect 277636 224216 309140 224244
rect 277636 224204 277642 224216
rect 309134 224204 309140 224216
rect 309192 224244 309198 224256
rect 322934 224244 322940 224256
rect 309192 224216 322940 224244
rect 309192 224204 309198 224216
rect 322934 224204 322940 224216
rect 322992 224204 322998 224256
rect 269942 223632 269948 223644
rect 238726 223604 269948 223632
rect 69014 223524 69020 223576
rect 69072 223564 69078 223576
rect 231118 223564 231124 223576
rect 69072 223536 231124 223564
rect 69072 223524 69078 223536
rect 231118 223524 231124 223536
rect 231176 223564 231182 223576
rect 233234 223564 233240 223576
rect 231176 223536 233240 223564
rect 231176 223524 231182 223536
rect 233234 223524 233240 223536
rect 233292 223524 233298 223576
rect 138382 223456 138388 223508
rect 138440 223496 138446 223508
rect 155218 223496 155224 223508
rect 138440 223468 155224 223496
rect 138440 223456 138446 223468
rect 155218 223456 155224 223468
rect 155276 223456 155282 223508
rect 155770 223456 155776 223508
rect 155828 223496 155834 223508
rect 215110 223496 215116 223508
rect 155828 223468 215116 223496
rect 155828 223456 155834 223468
rect 215110 223456 215116 223468
rect 215168 223496 215174 223508
rect 238294 223496 238300 223508
rect 215168 223468 238300 223496
rect 215168 223456 215174 223468
rect 238294 223456 238300 223468
rect 238352 223496 238358 223508
rect 238726 223496 238754 223604
rect 269942 223592 269948 223604
rect 270000 223592 270006 223644
rect 238352 223468 238754 223496
rect 238352 223456 238358 223468
rect 279418 222844 279424 222896
rect 279476 222884 279482 222896
rect 295426 222884 295432 222896
rect 279476 222856 295432 222884
rect 279476 222844 279482 222856
rect 295426 222844 295432 222856
rect 295484 222844 295490 222896
rect 69658 222096 69664 222148
rect 69716 222136 69722 222148
rect 182910 222136 182916 222148
rect 69716 222108 182916 222136
rect 69716 222096 69722 222108
rect 182910 222096 182916 222108
rect 182968 222096 182974 222148
rect 184198 222096 184204 222148
rect 184256 222136 184262 222148
rect 244366 222136 244372 222148
rect 184256 222108 244372 222136
rect 184256 222096 184262 222108
rect 244366 222096 244372 222108
rect 244424 222096 244430 222148
rect 100754 221416 100760 221468
rect 100812 221456 100818 221468
rect 195882 221456 195888 221468
rect 100812 221428 195888 221456
rect 100812 221416 100818 221428
rect 195882 221416 195888 221428
rect 195940 221416 195946 221468
rect 202414 221416 202420 221468
rect 202472 221456 202478 221468
rect 276658 221456 276664 221468
rect 202472 221428 276664 221456
rect 202472 221416 202478 221428
rect 276658 221416 276664 221428
rect 276716 221416 276722 221468
rect 91186 220736 91192 220788
rect 91244 220776 91250 220788
rect 211338 220776 211344 220788
rect 91244 220748 211344 220776
rect 91244 220736 91250 220748
rect 211338 220736 211344 220748
rect 211396 220736 211402 220788
rect 227254 220736 227260 220788
rect 227312 220776 227318 220788
rect 262950 220776 262956 220788
rect 227312 220748 262956 220776
rect 227312 220736 227318 220748
rect 262950 220736 262956 220748
rect 263008 220736 263014 220788
rect 104894 220668 104900 220720
rect 104952 220708 104958 220720
rect 193122 220708 193128 220720
rect 104952 220680 193128 220708
rect 104952 220668 104958 220680
rect 193122 220668 193128 220680
rect 193180 220668 193186 220720
rect 193122 220056 193128 220108
rect 193180 220096 193186 220108
rect 227070 220096 227076 220108
rect 193180 220068 227076 220096
rect 193180 220056 193186 220068
rect 227070 220056 227076 220068
rect 227128 220056 227134 220108
rect 215202 219444 215208 219496
rect 215260 219484 215266 219496
rect 228358 219484 228364 219496
rect 215260 219456 228364 219484
rect 215260 219444 215266 219456
rect 228358 219444 228364 219456
rect 228416 219444 228422 219496
rect 124214 219376 124220 219428
rect 124272 219416 124278 219428
rect 227714 219416 227720 219428
rect 124272 219388 227720 219416
rect 124272 219376 124278 219388
rect 227714 219376 227720 219388
rect 227772 219376 227778 219428
rect 231854 219376 231860 219428
rect 231912 219416 231918 219428
rect 279602 219416 279608 219428
rect 231912 219388 279608 219416
rect 231912 219376 231918 219388
rect 279602 219376 279608 219388
rect 279660 219376 279666 219428
rect 73062 219308 73068 219360
rect 73120 219348 73126 219360
rect 156598 219348 156604 219360
rect 73120 219320 156604 219348
rect 73120 219308 73126 219320
rect 156598 219308 156604 219320
rect 156656 219308 156662 219360
rect 170398 219308 170404 219360
rect 170456 219348 170462 219360
rect 215202 219348 215208 219360
rect 170456 219320 215208 219348
rect 170456 219308 170462 219320
rect 215202 219308 215208 219320
rect 215260 219308 215266 219360
rect 95234 217948 95240 218000
rect 95292 217988 95298 218000
rect 244274 217988 244280 218000
rect 95292 217960 244280 217988
rect 95292 217948 95298 217960
rect 244274 217948 244280 217960
rect 244332 217948 244338 218000
rect 132310 217880 132316 217932
rect 132368 217920 132374 217932
rect 192662 217920 192668 217932
rect 132368 217892 192668 217920
rect 132368 217880 132374 217892
rect 192662 217880 192668 217892
rect 192720 217880 192726 217932
rect 195882 217880 195888 217932
rect 195940 217920 195946 217932
rect 212534 217920 212540 217932
rect 195940 217892 212540 217920
rect 195940 217880 195946 217892
rect 212534 217880 212540 217892
rect 212592 217880 212598 217932
rect 192478 216656 192484 216708
rect 192536 216696 192542 216708
rect 192662 216696 192668 216708
rect 192536 216668 192668 216696
rect 192536 216656 192542 216668
rect 192662 216656 192668 216668
rect 192720 216656 192726 216708
rect 212534 216656 212540 216708
rect 212592 216696 212598 216708
rect 213178 216696 213184 216708
rect 212592 216668 213184 216696
rect 212592 216656 212598 216668
rect 213178 216656 213184 216668
rect 213236 216656 213242 216708
rect 117314 216588 117320 216640
rect 117372 216628 117378 216640
rect 224218 216628 224224 216640
rect 117372 216600 224224 216628
rect 117372 216588 117378 216600
rect 224218 216588 224224 216600
rect 224276 216588 224282 216640
rect 177482 216520 177488 216572
rect 177540 216560 177546 216572
rect 220170 216560 220176 216572
rect 177540 216532 220176 216560
rect 177540 216520 177546 216532
rect 220170 216520 220176 216532
rect 220228 216560 220234 216572
rect 220446 216560 220452 216572
rect 220228 216532 220452 216560
rect 220228 216520 220234 216532
rect 220446 216520 220452 216532
rect 220504 216520 220510 216572
rect 91094 215908 91100 215960
rect 91152 215948 91158 215960
rect 92382 215948 92388 215960
rect 91152 215920 92388 215948
rect 91152 215908 91158 215920
rect 92382 215908 92388 215920
rect 92440 215948 92446 215960
rect 175274 215948 175280 215960
rect 92440 215920 175280 215948
rect 92440 215908 92446 215920
rect 175274 215908 175280 215920
rect 175332 215908 175338 215960
rect 164970 215228 164976 215280
rect 165028 215268 165034 215280
rect 249886 215268 249892 215280
rect 165028 215240 249892 215268
rect 165028 215228 165034 215240
rect 249886 215228 249892 215240
rect 249944 215228 249950 215280
rect 114462 214616 114468 214668
rect 114520 214656 114526 214668
rect 187142 214656 187148 214668
rect 114520 214628 187148 214656
rect 114520 214616 114526 214628
rect 187142 214616 187148 214628
rect 187200 214616 187206 214668
rect 35158 214548 35164 214600
rect 35216 214588 35222 214600
rect 159358 214588 159364 214600
rect 35216 214560 159364 214588
rect 35216 214548 35222 214560
rect 159358 214548 159364 214560
rect 159416 214548 159422 214600
rect 197170 214548 197176 214600
rect 197228 214588 197234 214600
rect 233326 214588 233332 214600
rect 197228 214560 233332 214588
rect 197228 214548 197234 214560
rect 233326 214548 233332 214560
rect 233384 214548 233390 214600
rect 260742 214548 260748 214600
rect 260800 214588 260806 214600
rect 291286 214588 291292 214600
rect 260800 214560 291292 214588
rect 260800 214548 260806 214560
rect 291286 214548 291292 214560
rect 291344 214548 291350 214600
rect 100570 213868 100576 213920
rect 100628 213908 100634 213920
rect 183278 213908 183284 213920
rect 100628 213880 183284 213908
rect 100628 213868 100634 213880
rect 183278 213868 183284 213880
rect 183336 213908 183342 213920
rect 184474 213908 184480 213920
rect 183336 213880 184480 213908
rect 183336 213868 183342 213880
rect 184474 213868 184480 213880
rect 184532 213868 184538 213920
rect 198642 213868 198648 213920
rect 198700 213908 198706 213920
rect 199470 213908 199476 213920
rect 198700 213880 199476 213908
rect 198700 213868 198706 213880
rect 199470 213868 199476 213880
rect 199528 213868 199534 213920
rect 124306 213188 124312 213240
rect 124364 213228 124370 213240
rect 198642 213228 198648 213240
rect 124364 213200 198648 213228
rect 124364 213188 124370 213200
rect 198642 213188 198648 213200
rect 198700 213188 198706 213240
rect 189074 212576 189080 212628
rect 189132 212616 189138 212628
rect 190362 212616 190368 212628
rect 189132 212588 190368 212616
rect 189132 212576 189138 212588
rect 190362 212576 190368 212588
rect 190420 212616 190426 212628
rect 232130 212616 232136 212628
rect 190420 212588 232136 212616
rect 190420 212576 190426 212588
rect 232130 212576 232136 212588
rect 232188 212576 232194 212628
rect 207750 212508 207756 212560
rect 207808 212548 207814 212560
rect 208210 212548 208216 212560
rect 207808 212520 208216 212548
rect 207808 212508 207814 212520
rect 208210 212508 208216 212520
rect 208268 212548 208274 212560
rect 278130 212548 278136 212560
rect 208268 212520 278136 212548
rect 208268 212508 208274 212520
rect 278130 212508 278136 212520
rect 278188 212508 278194 212560
rect 86954 212440 86960 212492
rect 87012 212480 87018 212492
rect 209682 212480 209688 212492
rect 87012 212452 209688 212480
rect 87012 212440 87018 212452
rect 209682 212440 209688 212452
rect 209740 212440 209746 212492
rect 144822 211760 144828 211812
rect 144880 211800 144886 211812
rect 237374 211800 237380 211812
rect 144880 211772 237380 211800
rect 144880 211760 144886 211772
rect 237374 211760 237380 211772
rect 237432 211760 237438 211812
rect 209682 211148 209688 211200
rect 209740 211188 209746 211200
rect 214650 211188 214656 211200
rect 209740 211160 214656 211188
rect 209740 211148 209746 211160
rect 214650 211148 214656 211160
rect 214708 211148 214714 211200
rect 184842 210468 184848 210520
rect 184900 210508 184906 210520
rect 244458 210508 244464 210520
rect 184900 210480 244464 210508
rect 184900 210468 184906 210480
rect 244458 210468 244464 210480
rect 244516 210468 244522 210520
rect 71038 210400 71044 210452
rect 71096 210440 71102 210452
rect 188338 210440 188344 210452
rect 71096 210412 188344 210440
rect 71096 210400 71102 210412
rect 188338 210400 188344 210412
rect 188396 210400 188402 210452
rect 216490 209788 216496 209840
rect 216548 209828 216554 209840
rect 245930 209828 245936 209840
rect 216548 209800 245936 209828
rect 216548 209788 216554 209800
rect 245930 209788 245936 209800
rect 245988 209788 245994 209840
rect 67726 209720 67732 209772
rect 67784 209760 67790 209772
rect 206370 209760 206376 209772
rect 67784 209732 206376 209760
rect 67784 209720 67790 209732
rect 206370 209720 206376 209732
rect 206428 209720 206434 209772
rect 132402 209652 132408 209704
rect 132460 209692 132466 209704
rect 248506 209692 248512 209704
rect 132460 209664 248512 209692
rect 132460 209652 132466 209664
rect 248506 209652 248512 209664
rect 248564 209652 248570 209704
rect 216674 208360 216680 208412
rect 216732 208400 216738 208412
rect 217962 208400 217968 208412
rect 216732 208372 217968 208400
rect 216732 208360 216738 208372
rect 217962 208360 217968 208372
rect 218020 208400 218026 208412
rect 307846 208400 307852 208412
rect 218020 208372 307852 208400
rect 218020 208360 218026 208372
rect 307846 208360 307852 208372
rect 307904 208360 307910 208412
rect 70394 208292 70400 208344
rect 70452 208332 70458 208344
rect 216490 208332 216496 208344
rect 70452 208304 216496 208332
rect 70452 208292 70458 208304
rect 216490 208292 216496 208304
rect 216548 208292 216554 208344
rect 187142 208224 187148 208276
rect 187200 208264 187206 208276
rect 245746 208264 245752 208276
rect 187200 208236 245752 208264
rect 187200 208224 187206 208236
rect 245746 208224 245752 208236
rect 245804 208224 245810 208276
rect 133782 206932 133788 206984
rect 133840 206972 133846 206984
rect 248690 206972 248696 206984
rect 133840 206944 248696 206972
rect 133840 206932 133846 206944
rect 248690 206932 248696 206944
rect 248748 206932 248754 206984
rect 122834 206864 122840 206916
rect 122892 206904 122898 206916
rect 225598 206904 225604 206916
rect 122892 206876 225604 206904
rect 122892 206864 122898 206876
rect 225598 206864 225604 206876
rect 225656 206864 225662 206916
rect 82722 205572 82728 205624
rect 82780 205612 82786 205624
rect 253934 205612 253940 205624
rect 82780 205584 253940 205612
rect 82780 205572 82786 205584
rect 253934 205572 253940 205584
rect 253992 205572 253998 205624
rect 106182 205504 106188 205556
rect 106240 205544 106246 205556
rect 216674 205544 216680 205556
rect 106240 205516 216680 205544
rect 106240 205504 106246 205516
rect 216674 205504 216680 205516
rect 216732 205504 216738 205556
rect 218054 204280 218060 204332
rect 218112 204320 218118 204332
rect 218238 204320 218244 204332
rect 218112 204292 218244 204320
rect 218112 204280 218118 204292
rect 218238 204280 218244 204292
rect 218296 204320 218302 204332
rect 229370 204320 229376 204332
rect 218296 204292 229376 204320
rect 218296 204280 218302 204292
rect 229370 204280 229376 204292
rect 229428 204280 229434 204332
rect 73798 204212 73804 204264
rect 73856 204252 73862 204264
rect 217134 204252 217140 204264
rect 73856 204224 217140 204252
rect 73856 204212 73862 204224
rect 217134 204212 217140 204224
rect 217192 204212 217198 204264
rect 188338 204144 188344 204196
rect 188396 204184 188402 204196
rect 234614 204184 234620 204196
rect 188396 204156 234620 204184
rect 188396 204144 188402 204156
rect 234614 204144 234620 204156
rect 234672 204144 234678 204196
rect 173158 203532 173164 203584
rect 173216 203572 173222 203584
rect 184198 203572 184204 203584
rect 173216 203544 184204 203572
rect 173216 203532 173222 203544
rect 184198 203532 184204 203544
rect 184256 203532 184262 203584
rect 225690 203532 225696 203584
rect 225748 203572 225754 203584
rect 284386 203572 284392 203584
rect 225748 203544 284392 203572
rect 225748 203532 225754 203544
rect 284386 203532 284392 203544
rect 284444 203532 284450 203584
rect 3418 202784 3424 202836
rect 3476 202824 3482 202836
rect 137278 202824 137284 202836
rect 3476 202796 137284 202824
rect 3476 202784 3482 202796
rect 137278 202784 137284 202796
rect 137336 202784 137342 202836
rect 147582 202784 147588 202836
rect 147640 202824 147646 202836
rect 247126 202824 247132 202836
rect 147640 202796 247132 202824
rect 147640 202784 147646 202796
rect 247126 202784 247132 202796
rect 247184 202784 247190 202836
rect 168282 202716 168288 202768
rect 168340 202756 168346 202768
rect 169110 202756 169116 202768
rect 168340 202728 169116 202756
rect 168340 202716 168346 202728
rect 169110 202716 169116 202728
rect 169168 202716 169174 202768
rect 141970 202104 141976 202156
rect 142028 202144 142034 202156
rect 168282 202144 168288 202156
rect 142028 202116 168288 202144
rect 142028 202104 142034 202116
rect 168282 202104 168288 202116
rect 168340 202104 168346 202156
rect 194410 202104 194416 202156
rect 194468 202144 194474 202156
rect 245654 202144 245660 202156
rect 194468 202116 245660 202144
rect 194468 202104 194474 202116
rect 245654 202104 245660 202116
rect 245712 202104 245718 202156
rect 117222 200812 117228 200864
rect 117280 200852 117286 200864
rect 190454 200852 190460 200864
rect 117280 200824 190460 200852
rect 117280 200812 117286 200824
rect 190454 200812 190460 200824
rect 190512 200812 190518 200864
rect 236822 200812 236828 200864
rect 236880 200852 236886 200864
rect 245746 200852 245752 200864
rect 236880 200824 245752 200852
rect 236880 200812 236886 200824
rect 245746 200812 245752 200824
rect 245804 200812 245810 200864
rect 272518 200812 272524 200864
rect 272576 200852 272582 200864
rect 289998 200852 290004 200864
rect 272576 200824 290004 200852
rect 272576 200812 272582 200824
rect 289998 200812 290004 200824
rect 290056 200812 290062 200864
rect 3418 200744 3424 200796
rect 3476 200784 3482 200796
rect 169018 200784 169024 200796
rect 3476 200756 169024 200784
rect 3476 200744 3482 200756
rect 169018 200744 169024 200756
rect 169076 200744 169082 200796
rect 209038 200744 209044 200796
rect 209096 200784 209102 200796
rect 238110 200784 238116 200796
rect 209096 200756 238116 200784
rect 209096 200744 209102 200756
rect 238110 200744 238116 200756
rect 238168 200744 238174 200796
rect 262858 200744 262864 200796
rect 262916 200784 262922 200796
rect 281534 200784 281540 200796
rect 262916 200756 281540 200784
rect 262916 200744 262922 200756
rect 281534 200744 281540 200756
rect 281592 200744 281598 200796
rect 49602 200064 49608 200116
rect 49660 200104 49666 200116
rect 177298 200104 177304 200116
rect 49660 200076 177304 200104
rect 49660 200064 49666 200076
rect 177298 200064 177304 200076
rect 177356 200064 177362 200116
rect 128998 199996 129004 200048
rect 129056 200036 129062 200048
rect 195514 200036 195520 200048
rect 129056 200008 195520 200036
rect 129056 199996 129062 200008
rect 195514 199996 195520 200008
rect 195572 199996 195578 200048
rect 215202 199452 215208 199504
rect 215260 199492 215266 199504
rect 242342 199492 242348 199504
rect 215260 199464 242348 199492
rect 215260 199452 215266 199464
rect 242342 199452 242348 199464
rect 242400 199452 242406 199504
rect 202322 199384 202328 199436
rect 202380 199424 202386 199436
rect 238754 199424 238760 199436
rect 202380 199396 238760 199424
rect 202380 199384 202386 199396
rect 238754 199384 238760 199396
rect 238812 199384 238818 199436
rect 284294 198704 284300 198756
rect 284352 198744 284358 198756
rect 294598 198744 294604 198756
rect 284352 198716 294604 198744
rect 284352 198704 284358 198716
rect 294598 198704 294604 198716
rect 294656 198704 294662 198756
rect 76558 198636 76564 198688
rect 76616 198676 76622 198688
rect 238938 198676 238944 198688
rect 76616 198648 238944 198676
rect 76616 198636 76622 198648
rect 238938 198636 238944 198648
rect 238996 198636 239002 198688
rect 126882 198568 126888 198620
rect 126940 198608 126946 198620
rect 252554 198608 252560 198620
rect 126940 198580 252560 198608
rect 126940 198568 126946 198580
rect 252554 198568 252560 198580
rect 252612 198568 252618 198620
rect 260190 198024 260196 198076
rect 260248 198064 260254 198076
rect 270586 198064 270592 198076
rect 260248 198036 270592 198064
rect 260248 198024 260254 198036
rect 270586 198024 270592 198036
rect 270644 198024 270650 198076
rect 241422 197956 241428 198008
rect 241480 197996 241486 198008
rect 306650 197996 306656 198008
rect 241480 197968 306656 197996
rect 241480 197956 241486 197968
rect 306650 197956 306656 197968
rect 306708 197956 306714 198008
rect 103422 197276 103428 197328
rect 103480 197316 103486 197328
rect 163498 197316 163504 197328
rect 103480 197288 163504 197316
rect 103480 197276 103486 197288
rect 163498 197276 163504 197288
rect 163556 197276 163562 197328
rect 201402 196664 201408 196716
rect 201460 196704 201466 196716
rect 232590 196704 232596 196716
rect 201460 196676 232596 196704
rect 201460 196664 201466 196676
rect 232590 196664 232596 196676
rect 232648 196664 232654 196716
rect 50890 196596 50896 196648
rect 50948 196636 50954 196648
rect 204254 196636 204260 196648
rect 50948 196608 204260 196636
rect 50948 196596 50954 196608
rect 204254 196596 204260 196608
rect 204312 196596 204318 196648
rect 206462 196596 206468 196648
rect 206520 196636 206526 196648
rect 284294 196636 284300 196648
rect 206520 196608 284300 196636
rect 206520 196596 206526 196608
rect 284294 196596 284300 196608
rect 284352 196596 284358 196648
rect 106274 195916 106280 195968
rect 106332 195956 106338 195968
rect 162762 195956 162768 195968
rect 106332 195928 162768 195956
rect 106332 195916 106338 195928
rect 162762 195916 162768 195928
rect 162820 195916 162826 195968
rect 162762 195304 162768 195356
rect 162820 195344 162826 195356
rect 192662 195344 192668 195356
rect 162820 195316 192668 195344
rect 162820 195304 162826 195316
rect 192662 195304 192668 195316
rect 192720 195304 192726 195356
rect 119982 195236 119988 195288
rect 120040 195276 120046 195288
rect 177298 195276 177304 195288
rect 120040 195248 177304 195276
rect 120040 195236 120046 195248
rect 177298 195236 177304 195248
rect 177356 195236 177362 195288
rect 191374 195236 191380 195288
rect 191432 195276 191438 195288
rect 200850 195276 200856 195288
rect 191432 195248 200856 195276
rect 191432 195236 191438 195248
rect 200850 195236 200856 195248
rect 200908 195236 200914 195288
rect 206278 195236 206284 195288
rect 206336 195276 206342 195288
rect 245838 195276 245844 195288
rect 206336 195248 245844 195276
rect 206336 195236 206342 195248
rect 245838 195236 245844 195248
rect 245896 195236 245902 195288
rect 207658 193944 207664 193996
rect 207716 193984 207722 193996
rect 227714 193984 227720 193996
rect 207716 193956 227720 193984
rect 207716 193944 207722 193956
rect 227714 193944 227720 193956
rect 227772 193944 227778 193996
rect 188522 193876 188528 193928
rect 188580 193916 188586 193928
rect 217410 193916 217416 193928
rect 188580 193888 217416 193916
rect 188580 193876 188586 193888
rect 217410 193876 217416 193888
rect 217468 193876 217474 193928
rect 113082 193808 113088 193860
rect 113140 193848 113146 193860
rect 191190 193848 191196 193860
rect 113140 193820 191196 193848
rect 113140 193808 113146 193820
rect 191190 193808 191196 193820
rect 191248 193808 191254 193860
rect 220262 193808 220268 193860
rect 220320 193848 220326 193860
rect 276842 193848 276848 193860
rect 220320 193820 276848 193848
rect 220320 193808 220326 193820
rect 276842 193808 276848 193820
rect 276900 193808 276906 193860
rect 291838 193808 291844 193860
rect 291896 193848 291902 193860
rect 301130 193848 301136 193860
rect 291896 193820 301136 193848
rect 291896 193808 291902 193820
rect 301130 193808 301136 193820
rect 301188 193808 301194 193860
rect 214650 192516 214656 192568
rect 214708 192556 214714 192568
rect 233878 192556 233884 192568
rect 214708 192528 233884 192556
rect 214708 192516 214714 192528
rect 233878 192516 233884 192528
rect 233936 192516 233942 192568
rect 177390 192448 177396 192500
rect 177448 192488 177454 192500
rect 247126 192488 247132 192500
rect 177448 192460 247132 192488
rect 177448 192448 177454 192460
rect 247126 192448 247132 192460
rect 247184 192448 247190 192500
rect 266998 192448 267004 192500
rect 267056 192488 267062 192500
rect 292666 192488 292672 192500
rect 267056 192460 292672 192488
rect 267056 192448 267062 192460
rect 292666 192448 292672 192460
rect 292724 192448 292730 192500
rect 115198 191836 115204 191888
rect 115256 191876 115262 191888
rect 196802 191876 196808 191888
rect 115256 191848 196808 191876
rect 115256 191836 115262 191848
rect 196802 191836 196808 191848
rect 196860 191836 196866 191888
rect 227714 191224 227720 191276
rect 227772 191264 227778 191276
rect 253198 191264 253204 191276
rect 227772 191236 253204 191264
rect 227772 191224 227778 191236
rect 253198 191224 253204 191236
rect 253256 191224 253262 191276
rect 90358 191156 90364 191208
rect 90416 191196 90422 191208
rect 192570 191196 192576 191208
rect 90416 191168 192576 191196
rect 90416 191156 90422 191168
rect 192570 191156 192576 191168
rect 192628 191156 192634 191208
rect 202138 191156 202144 191208
rect 202196 191196 202202 191208
rect 232498 191196 232504 191208
rect 202196 191168 232504 191196
rect 202196 191156 202202 191168
rect 232498 191156 232504 191168
rect 232556 191156 232562 191208
rect 259362 191156 259368 191208
rect 259420 191196 259426 191208
rect 305086 191196 305092 191208
rect 259420 191168 305092 191196
rect 259420 191156 259426 191168
rect 305086 191156 305092 191168
rect 305144 191156 305150 191208
rect 52086 191088 52092 191140
rect 52144 191128 52150 191140
rect 166994 191128 167000 191140
rect 52144 191100 167000 191128
rect 52144 191088 52150 191100
rect 166994 191088 167000 191100
rect 167052 191088 167058 191140
rect 192478 191088 192484 191140
rect 192536 191128 192542 191140
rect 228450 191128 228456 191140
rect 192536 191100 228456 191128
rect 192536 191088 192542 191100
rect 228450 191088 228456 191100
rect 228508 191088 228514 191140
rect 238110 191088 238116 191140
rect 238168 191128 238174 191140
rect 303890 191128 303896 191140
rect 238168 191100 303896 191128
rect 238168 191088 238174 191100
rect 303890 191088 303896 191100
rect 303948 191088 303954 191140
rect 136634 190408 136640 190460
rect 136692 190448 136698 190460
rect 243906 190448 243912 190460
rect 136692 190420 243912 190448
rect 136692 190408 136698 190420
rect 243906 190408 243912 190420
rect 243964 190408 243970 190460
rect 217318 189728 217324 189780
rect 217376 189768 217382 189780
rect 238846 189768 238852 189780
rect 217376 189740 238852 189768
rect 217376 189728 217382 189740
rect 238846 189728 238852 189740
rect 238904 189728 238910 189780
rect 125502 189048 125508 189100
rect 125560 189088 125566 189100
rect 174630 189088 174636 189100
rect 125560 189060 174636 189088
rect 125560 189048 125566 189060
rect 174630 189048 174636 189060
rect 174688 189048 174694 189100
rect 3510 188980 3516 189032
rect 3568 189020 3574 189032
rect 15838 189020 15844 189032
rect 3568 188992 15844 189020
rect 3568 188980 3574 188992
rect 15838 188980 15844 188992
rect 15896 188980 15902 189032
rect 164878 188368 164884 188420
rect 164936 188408 164942 188420
rect 241606 188408 241612 188420
rect 164936 188380 241612 188408
rect 164936 188368 164942 188380
rect 241606 188368 241612 188380
rect 241664 188368 241670 188420
rect 275922 188368 275928 188420
rect 275980 188408 275986 188420
rect 295610 188408 295616 188420
rect 275980 188380 295616 188408
rect 275980 188368 275986 188380
rect 295610 188368 295616 188380
rect 295668 188368 295674 188420
rect 89622 188300 89628 188352
rect 89680 188340 89686 188352
rect 220262 188340 220268 188352
rect 89680 188312 220268 188340
rect 89680 188300 89686 188312
rect 220262 188300 220268 188312
rect 220320 188300 220326 188352
rect 262122 188300 262128 188352
rect 262180 188340 262186 188352
rect 299474 188340 299480 188352
rect 262180 188312 299480 188340
rect 262180 188300 262186 188312
rect 299474 188300 299480 188312
rect 299532 188300 299538 188352
rect 302142 188300 302148 188352
rect 302200 188340 302206 188352
rect 314746 188340 314752 188352
rect 302200 188312 314752 188340
rect 302200 188300 302206 188312
rect 314746 188300 314752 188312
rect 314804 188300 314810 188352
rect 133138 187688 133144 187740
rect 133196 187728 133202 187740
rect 164970 187728 164976 187740
rect 133196 187700 164976 187728
rect 133196 187688 133202 187700
rect 164970 187688 164976 187700
rect 165028 187688 165034 187740
rect 255958 187620 255964 187672
rect 256016 187660 256022 187672
rect 258074 187660 258080 187672
rect 256016 187632 258080 187660
rect 256016 187620 256022 187632
rect 258074 187620 258080 187632
rect 258132 187620 258138 187672
rect 198642 186940 198648 186992
rect 198700 186980 198706 186992
rect 242986 186980 242992 186992
rect 198700 186952 242992 186980
rect 198700 186940 198706 186952
rect 242986 186940 242992 186952
rect 243044 186940 243050 186992
rect 223482 186668 223488 186720
rect 223540 186708 223546 186720
rect 227162 186708 227168 186720
rect 223540 186680 227168 186708
rect 223540 186668 223546 186680
rect 227162 186668 227168 186680
rect 227220 186668 227226 186720
rect 113082 186396 113088 186448
rect 113140 186436 113146 186448
rect 177390 186436 177396 186448
rect 113140 186408 177396 186436
rect 113140 186396 113146 186408
rect 177390 186396 177396 186408
rect 177448 186396 177454 186448
rect 133782 186328 133788 186380
rect 133840 186368 133846 186380
rect 210510 186368 210516 186380
rect 133840 186340 210516 186368
rect 133840 186328 133846 186340
rect 210510 186328 210516 186340
rect 210568 186328 210574 186380
rect 292850 186368 292856 186380
rect 229066 186340 292856 186368
rect 53466 186260 53472 186312
rect 53524 186300 53530 186312
rect 169386 186300 169392 186312
rect 53524 186272 169392 186300
rect 53524 186260 53530 186272
rect 169386 186260 169392 186272
rect 169444 186260 169450 186312
rect 202230 186260 202236 186312
rect 202288 186300 202294 186312
rect 229066 186300 229094 186340
rect 292850 186328 292856 186340
rect 292908 186328 292914 186380
rect 202288 186272 229094 186300
rect 202288 186260 202294 186272
rect 232590 185716 232596 185768
rect 232648 185756 232654 185768
rect 242894 185756 242900 185768
rect 232648 185728 242900 185756
rect 232648 185716 232654 185728
rect 242894 185716 242900 185728
rect 242952 185716 242958 185768
rect 230198 185648 230204 185700
rect 230256 185688 230262 185700
rect 233050 185688 233056 185700
rect 230256 185660 233056 185688
rect 230256 185648 230262 185660
rect 233050 185648 233056 185660
rect 233108 185648 233114 185700
rect 213178 185580 213184 185632
rect 213236 185620 213242 185632
rect 238938 185620 238944 185632
rect 213236 185592 238944 185620
rect 213236 185580 213242 185592
rect 238938 185580 238944 185592
rect 238996 185580 239002 185632
rect 269758 185580 269764 185632
rect 269816 185620 269822 185632
rect 285950 185620 285956 185632
rect 269816 185592 285956 185620
rect 269816 185580 269822 185592
rect 285950 185580 285956 185592
rect 286008 185580 286014 185632
rect 118602 184900 118608 184952
rect 118660 184940 118666 184952
rect 185578 184940 185584 184952
rect 118660 184912 185584 184940
rect 118660 184900 118666 184912
rect 185578 184900 185584 184912
rect 185636 184900 185642 184952
rect 227070 184220 227076 184272
rect 227128 184260 227134 184272
rect 244550 184260 244556 184272
rect 227128 184232 244556 184260
rect 227128 184220 227134 184232
rect 244550 184220 244556 184232
rect 244608 184220 244614 184272
rect 191098 184152 191104 184204
rect 191156 184192 191162 184204
rect 230566 184192 230572 184204
rect 191156 184164 230572 184192
rect 191156 184152 191162 184164
rect 230566 184152 230572 184164
rect 230624 184152 230630 184204
rect 244182 184152 244188 184204
rect 244240 184192 244246 184204
rect 283558 184192 283564 184204
rect 244240 184164 283564 184192
rect 244240 184152 244246 184164
rect 283558 184152 283564 184164
rect 283616 184152 283622 184204
rect 316770 184152 316776 184204
rect 316828 184192 316834 184204
rect 326338 184192 326344 184204
rect 316828 184164 326344 184192
rect 316828 184152 316834 184164
rect 326338 184152 326344 184164
rect 326396 184152 326402 184204
rect 128998 183608 129004 183660
rect 129056 183648 129062 183660
rect 167822 183648 167828 183660
rect 129056 183620 167828 183648
rect 129056 183608 129062 183620
rect 167822 183608 167828 183620
rect 167880 183608 167886 183660
rect 107562 183540 107568 183592
rect 107620 183580 107626 183592
rect 166350 183580 166356 183592
rect 107620 183552 166356 183580
rect 107620 183540 107626 183552
rect 166350 183540 166356 183552
rect 166408 183540 166414 183592
rect 180702 182860 180708 182912
rect 180760 182900 180766 182912
rect 229462 182900 229468 182912
rect 180760 182872 229468 182900
rect 180760 182860 180766 182872
rect 229462 182860 229468 182872
rect 229520 182860 229526 182912
rect 199378 182792 199384 182844
rect 199436 182832 199442 182844
rect 248598 182832 248604 182844
rect 199436 182804 248604 182832
rect 199436 182792 199442 182804
rect 248598 182792 248604 182804
rect 248656 182792 248662 182844
rect 280890 182792 280896 182844
rect 280948 182832 280954 182844
rect 291378 182832 291384 182844
rect 280948 182804 291384 182832
rect 280948 182792 280954 182804
rect 291378 182792 291384 182804
rect 291436 182792 291442 182844
rect 134794 182248 134800 182300
rect 134852 182288 134858 182300
rect 162854 182288 162860 182300
rect 134852 182260 162860 182288
rect 134852 182248 134858 182260
rect 162854 182248 162860 182260
rect 162912 182248 162918 182300
rect 121914 182180 121920 182232
rect 121972 182220 121978 182232
rect 173250 182220 173256 182232
rect 121972 182192 173256 182220
rect 121972 182180 121978 182192
rect 173250 182180 173256 182192
rect 173308 182180 173314 182232
rect 271230 181500 271236 181552
rect 271288 181540 271294 181552
rect 283190 181540 283196 181552
rect 271288 181512 283196 181540
rect 271288 181500 271294 181512
rect 283190 181500 283196 181512
rect 283248 181500 283254 181552
rect 184290 181432 184296 181484
rect 184348 181472 184354 181484
rect 237466 181472 237472 181484
rect 184348 181444 237472 181472
rect 184348 181432 184354 181444
rect 237466 181432 237472 181444
rect 237524 181432 237530 181484
rect 273898 181432 273904 181484
rect 273956 181472 273962 181484
rect 288710 181472 288716 181484
rect 273956 181444 288716 181472
rect 273956 181432 273962 181444
rect 288710 181432 288716 181444
rect 288768 181432 288774 181484
rect 105906 180888 105912 180940
rect 105964 180928 105970 180940
rect 170398 180928 170404 180940
rect 105964 180900 170404 180928
rect 105964 180888 105970 180900
rect 170398 180888 170404 180900
rect 170456 180888 170462 180940
rect 132402 180820 132408 180872
rect 132460 180860 132466 180872
rect 214926 180860 214932 180872
rect 132460 180832 214932 180860
rect 132460 180820 132466 180832
rect 214926 180820 214932 180832
rect 214984 180820 214990 180872
rect 226242 180820 226248 180872
rect 226300 180860 226306 180872
rect 251358 180860 251364 180872
rect 226300 180832 251364 180860
rect 226300 180820 226306 180832
rect 251358 180820 251364 180832
rect 251416 180820 251422 180872
rect 220262 180140 220268 180192
rect 220320 180180 220326 180192
rect 232222 180180 232228 180192
rect 220320 180152 232228 180180
rect 220320 180140 220326 180152
rect 232222 180140 232228 180152
rect 232280 180140 232286 180192
rect 278130 180140 278136 180192
rect 278188 180180 278194 180192
rect 280246 180180 280252 180192
rect 278188 180152 280252 180180
rect 278188 180140 278194 180152
rect 280246 180140 280252 180152
rect 280304 180140 280310 180192
rect 187050 180072 187056 180124
rect 187108 180112 187114 180124
rect 226426 180112 226432 180124
rect 187108 180084 226432 180112
rect 187108 180072 187114 180084
rect 226426 180072 226432 180084
rect 226484 180072 226490 180124
rect 233878 180072 233884 180124
rect 233936 180112 233942 180124
rect 241514 180112 241520 180124
rect 233936 180084 241520 180112
rect 233936 180072 233942 180084
rect 241514 180072 241520 180084
rect 241572 180072 241578 180124
rect 253198 180072 253204 180124
rect 253256 180112 253262 180124
rect 276014 180112 276020 180124
rect 253256 180084 276020 180112
rect 253256 180072 253262 180084
rect 276014 180072 276020 180084
rect 276072 180072 276078 180124
rect 284938 180072 284944 180124
rect 284996 180112 285002 180124
rect 298370 180112 298376 180124
rect 284996 180084 298376 180112
rect 284996 180072 285002 180084
rect 298370 180072 298376 180084
rect 298428 180072 298434 180124
rect 119890 179460 119896 179512
rect 119948 179500 119954 179512
rect 167730 179500 167736 179512
rect 119948 179472 167736 179500
rect 119948 179460 119954 179472
rect 167730 179460 167736 179472
rect 167788 179460 167794 179512
rect 126790 179392 126796 179444
rect 126848 179432 126854 179444
rect 206278 179432 206284 179444
rect 126848 179404 206284 179432
rect 126848 179392 126854 179404
rect 206278 179392 206284 179404
rect 206336 179392 206342 179444
rect 227162 179392 227168 179444
rect 227220 179432 227226 179444
rect 229278 179432 229284 179444
rect 227220 179404 229284 179432
rect 227220 179392 227226 179404
rect 229278 179392 229284 179404
rect 229336 179392 229342 179444
rect 276842 179392 276848 179444
rect 276900 179432 276906 179444
rect 279142 179432 279148 179444
rect 276900 179404 279148 179432
rect 276900 179392 276906 179404
rect 279142 179392 279148 179404
rect 279200 179392 279206 179444
rect 281442 179392 281448 179444
rect 281500 179432 281506 179444
rect 284478 179432 284484 179444
rect 281500 179404 284484 179432
rect 281500 179392 281506 179404
rect 284478 179392 284484 179404
rect 284536 179392 284542 179444
rect 220170 178712 220176 178764
rect 220228 178752 220234 178764
rect 233234 178752 233240 178764
rect 220228 178724 233240 178752
rect 220228 178712 220234 178724
rect 233234 178712 233240 178724
rect 233292 178712 233298 178764
rect 279418 178712 279424 178764
rect 279476 178752 279482 178764
rect 296990 178752 296996 178764
rect 279476 178724 296996 178752
rect 279476 178712 279482 178724
rect 296990 178712 296996 178724
rect 297048 178712 297054 178764
rect 200850 178644 200856 178696
rect 200908 178684 200914 178696
rect 231946 178684 231952 178696
rect 200908 178656 231952 178684
rect 200908 178644 200914 178656
rect 231946 178644 231952 178656
rect 232004 178644 232010 178696
rect 232498 178644 232504 178696
rect 232556 178684 232562 178696
rect 292758 178684 292764 178696
rect 232556 178656 292764 178684
rect 232556 178644 232562 178656
rect 292758 178644 292764 178656
rect 292816 178644 292822 178696
rect 123294 178100 123300 178152
rect 123352 178140 123358 178152
rect 169110 178140 169116 178152
rect 123352 178112 169116 178140
rect 123352 178100 123358 178112
rect 169110 178100 169116 178112
rect 169168 178100 169174 178152
rect 148226 178032 148232 178084
rect 148284 178072 148290 178084
rect 203610 178072 203616 178084
rect 148284 178044 203616 178072
rect 148284 178032 148290 178044
rect 203610 178032 203616 178044
rect 203668 178032 203674 178084
rect 129458 177964 129464 178016
rect 129516 178004 129522 178016
rect 133138 178004 133144 178016
rect 129516 177976 133144 178004
rect 129516 177964 129522 177976
rect 133138 177964 133144 177976
rect 133196 177964 133202 178016
rect 203518 177964 203524 178016
rect 203576 178004 203582 178016
rect 226334 178004 226340 178016
rect 203576 177976 226340 178004
rect 203576 177964 203582 177976
rect 226334 177964 226340 177976
rect 226392 177964 226398 178016
rect 114186 177556 114192 177608
rect 114244 177596 114250 177608
rect 115198 177596 115204 177608
rect 114244 177568 115204 177596
rect 114244 177556 114250 177568
rect 115198 177556 115204 177568
rect 115256 177556 115262 177608
rect 127986 177556 127992 177608
rect 128044 177596 128050 177608
rect 128998 177596 129004 177608
rect 128044 177568 129004 177596
rect 128044 177556 128050 177568
rect 128998 177556 129004 177568
rect 129056 177556 129062 177608
rect 278038 177352 278044 177404
rect 278096 177392 278102 177404
rect 287330 177392 287336 177404
rect 278096 177364 287336 177392
rect 278096 177352 278102 177364
rect 287330 177352 287336 177364
rect 287388 177352 287394 177404
rect 228358 177284 228364 177336
rect 228416 177324 228422 177336
rect 233418 177324 233424 177336
rect 228416 177296 233424 177324
rect 228416 177284 228422 177296
rect 233418 177284 233424 177296
rect 233476 177284 233482 177336
rect 268378 177284 268384 177336
rect 268436 177324 268442 177336
rect 281810 177324 281816 177336
rect 268436 177296 281816 177324
rect 268436 177284 268442 177296
rect 281810 177284 281816 177296
rect 281868 177284 281874 177336
rect 158990 176740 158996 176792
rect 159048 176780 159054 176792
rect 173158 176780 173164 176792
rect 159048 176752 173164 176780
rect 159048 176740 159054 176752
rect 173158 176740 173164 176752
rect 173216 176740 173222 176792
rect 128170 176672 128176 176724
rect 128228 176712 128234 176724
rect 207014 176712 207020 176724
rect 128228 176684 207020 176712
rect 128228 176672 128234 176684
rect 207014 176672 207020 176684
rect 207072 176672 207078 176724
rect 229094 176712 229100 176724
rect 224972 176684 229100 176712
rect 135714 176604 135720 176656
rect 135772 176644 135778 176656
rect 213914 176644 213920 176656
rect 135772 176616 213920 176644
rect 135772 176604 135778 176616
rect 213914 176604 213920 176616
rect 213972 176604 213978 176656
rect 197262 176536 197268 176588
rect 197320 176576 197326 176588
rect 224972 176576 225000 176684
rect 229094 176672 229100 176684
rect 229152 176672 229158 176724
rect 269942 176604 269948 176656
rect 270000 176644 270006 176656
rect 281718 176644 281724 176656
rect 270000 176616 281724 176644
rect 270000 176604 270006 176616
rect 281718 176604 281724 176616
rect 281776 176644 281782 176656
rect 334618 176644 334624 176656
rect 281776 176616 334624 176644
rect 281776 176604 281782 176616
rect 334618 176604 334624 176616
rect 334676 176604 334682 176656
rect 197320 176548 225000 176576
rect 197320 176536 197326 176548
rect 283558 175992 283564 176044
rect 283616 176032 283622 176044
rect 284570 176032 284576 176044
rect 283616 176004 284576 176032
rect 283616 175992 283622 176004
rect 284570 175992 284576 176004
rect 284628 175992 284634 176044
rect 130746 175924 130752 175976
rect 130804 175964 130810 175976
rect 165522 175964 165528 175976
rect 130804 175936 165528 175964
rect 130804 175924 130810 175936
rect 165522 175924 165528 175936
rect 165580 175924 165586 175976
rect 226426 175924 226432 175976
rect 226484 175964 226490 175976
rect 233510 175964 233516 175976
rect 226484 175936 233516 175964
rect 226484 175924 226490 175936
rect 233510 175924 233516 175936
rect 233568 175924 233574 175976
rect 276658 175924 276664 175976
rect 276716 175964 276722 175976
rect 276716 175936 277394 175964
rect 276716 175924 276722 175936
rect 226518 175788 226524 175840
rect 226576 175788 226582 175840
rect 228450 175788 228456 175840
rect 228508 175828 228514 175840
rect 231854 175828 231860 175840
rect 228508 175800 231860 175828
rect 228508 175788 228514 175800
rect 231854 175788 231860 175800
rect 231912 175788 231918 175840
rect 277366 175828 277394 175936
rect 283006 175924 283012 175976
rect 283064 175964 283070 175976
rect 283190 175964 283196 175976
rect 283064 175936 283196 175964
rect 283064 175924 283070 175936
rect 283190 175924 283196 175936
rect 283248 175924 283254 175976
rect 283190 175828 283196 175840
rect 277366 175800 283196 175828
rect 283190 175788 283196 175800
rect 283248 175788 283254 175840
rect 210510 175176 210516 175228
rect 210568 175216 210574 175228
rect 214006 175216 214012 175228
rect 210568 175188 214012 175216
rect 210568 175176 210574 175188
rect 214006 175176 214012 175188
rect 214064 175176 214070 175228
rect 214558 175176 214564 175228
rect 214616 175216 214622 175228
rect 226536 175216 226564 175788
rect 239582 175244 239588 175296
rect 239640 175284 239646 175296
rect 264974 175284 264980 175296
rect 239640 175256 264980 175284
rect 239640 175244 239646 175256
rect 264974 175244 264980 175256
rect 265032 175244 265038 175296
rect 230658 175216 230664 175228
rect 214616 175188 219434 175216
rect 226536 175188 230664 175216
rect 214616 175176 214622 175188
rect 219406 175148 219434 175188
rect 230658 175176 230664 175188
rect 230716 175176 230722 175228
rect 232222 175176 232228 175228
rect 232280 175216 232286 175228
rect 256970 175216 256976 175228
rect 232280 175188 256976 175216
rect 232280 175176 232286 175188
rect 256970 175176 256976 175188
rect 257028 175176 257034 175228
rect 280982 175176 280988 175228
rect 281040 175216 281046 175228
rect 281902 175216 281908 175228
rect 281040 175188 281908 175216
rect 281040 175176 281046 175188
rect 281902 175176 281908 175188
rect 281960 175176 281966 175228
rect 282178 175176 282184 175228
rect 282236 175216 282242 175228
rect 285766 175216 285772 175228
rect 282236 175188 285772 175216
rect 282236 175176 282242 175188
rect 285766 175176 285772 175188
rect 285824 175176 285830 175228
rect 229370 175148 229376 175160
rect 219406 175120 229376 175148
rect 229370 175108 229376 175120
rect 229428 175108 229434 175160
rect 162854 175040 162860 175092
rect 162912 175080 162918 175092
rect 213914 175080 213920 175092
rect 162912 175052 213920 175080
rect 162912 175040 162918 175052
rect 213914 175040 213920 175052
rect 213972 175040 213978 175092
rect 280798 175040 280804 175092
rect 280856 175080 280862 175092
rect 285766 175080 285772 175092
rect 280856 175052 285772 175080
rect 280856 175040 280862 175052
rect 285766 175040 285772 175052
rect 285824 175040 285830 175092
rect 229002 174972 229008 175024
rect 229060 175012 229066 175024
rect 231946 175012 231952 175024
rect 229060 174984 231952 175012
rect 229060 174972 229066 174984
rect 231946 174972 231952 174984
rect 232004 174972 232010 175024
rect 260282 173952 260288 174004
rect 260340 173992 260346 174004
rect 265066 173992 265072 174004
rect 260340 173964 265072 173992
rect 260340 173952 260346 173964
rect 265066 173952 265072 173964
rect 265124 173952 265130 174004
rect 236638 173884 236644 173936
rect 236696 173924 236702 173936
rect 264974 173924 264980 173936
rect 236696 173896 264980 173924
rect 236696 173884 236702 173896
rect 264974 173884 264980 173896
rect 265032 173884 265038 173936
rect 165522 173816 165528 173868
rect 165580 173856 165586 173868
rect 213914 173856 213920 173868
rect 165580 173828 213920 173856
rect 165580 173816 165586 173828
rect 213914 173816 213920 173828
rect 213972 173816 213978 173868
rect 282454 173816 282460 173868
rect 282512 173856 282518 173868
rect 302418 173856 302424 173868
rect 282512 173828 302424 173856
rect 282512 173816 282518 173828
rect 302418 173816 302424 173828
rect 302476 173816 302482 173868
rect 230750 173136 230756 173188
rect 230808 173176 230814 173188
rect 247218 173176 247224 173188
rect 230808 173148 247224 173176
rect 230808 173136 230814 173148
rect 247218 173136 247224 173148
rect 247276 173136 247282 173188
rect 230382 172524 230388 172576
rect 230440 172564 230446 172576
rect 233326 172564 233332 172576
rect 230440 172536 233332 172564
rect 230440 172524 230446 172536
rect 233326 172524 233332 172536
rect 233384 172524 233390 172576
rect 249242 172524 249248 172576
rect 249300 172564 249306 172576
rect 264974 172564 264980 172576
rect 249300 172536 264980 172564
rect 249300 172524 249306 172536
rect 264974 172524 264980 172536
rect 265032 172524 265038 172576
rect 164970 172456 164976 172508
rect 165028 172496 165034 172508
rect 213914 172496 213920 172508
rect 165028 172468 213920 172496
rect 165028 172456 165034 172468
rect 213914 172456 213920 172468
rect 213972 172456 213978 172508
rect 231394 172456 231400 172508
rect 231452 172496 231458 172508
rect 252554 172496 252560 172508
rect 231452 172468 252560 172496
rect 231452 172456 231458 172468
rect 252554 172456 252560 172468
rect 252612 172456 252618 172508
rect 207014 172388 207020 172440
rect 207072 172428 207078 172440
rect 214006 172428 214012 172440
rect 207072 172400 214012 172428
rect 207072 172388 207078 172400
rect 214006 172388 214012 172400
rect 214064 172388 214070 172440
rect 231302 172388 231308 172440
rect 231360 172428 231366 172440
rect 240134 172428 240140 172440
rect 231360 172400 240140 172428
rect 231360 172388 231366 172400
rect 240134 172388 240140 172400
rect 240192 172388 240198 172440
rect 254670 171164 254676 171216
rect 254728 171204 254734 171216
rect 264974 171204 264980 171216
rect 254728 171176 264980 171204
rect 254728 171164 254734 171176
rect 264974 171164 264980 171176
rect 265032 171164 265038 171216
rect 167914 171096 167920 171148
rect 167972 171136 167978 171148
rect 182910 171136 182916 171148
rect 167972 171108 182916 171136
rect 167972 171096 167978 171108
rect 182910 171096 182916 171108
rect 182968 171096 182974 171148
rect 247678 171096 247684 171148
rect 247736 171136 247742 171148
rect 265066 171136 265072 171148
rect 247736 171108 265072 171136
rect 247736 171096 247742 171108
rect 265066 171096 265072 171108
rect 265124 171096 265130 171148
rect 167822 171028 167828 171080
rect 167880 171068 167886 171080
rect 213914 171068 213920 171080
rect 167880 171040 213920 171068
rect 167880 171028 167886 171040
rect 213914 171028 213920 171040
rect 213972 171028 213978 171080
rect 206278 170960 206284 171012
rect 206336 171000 206342 171012
rect 214006 171000 214012 171012
rect 206336 170972 214012 171000
rect 206336 170960 206342 170972
rect 214006 170960 214012 170972
rect 214064 170960 214070 171012
rect 282270 170892 282276 170944
rect 282328 170932 282334 170944
rect 285766 170932 285772 170944
rect 282328 170904 285772 170932
rect 282328 170892 282334 170904
rect 285766 170892 285772 170904
rect 285824 170892 285830 170944
rect 246666 170348 246672 170400
rect 246724 170388 246730 170400
rect 256786 170388 256792 170400
rect 246724 170360 256792 170388
rect 246724 170348 246730 170360
rect 256786 170348 256792 170360
rect 256844 170348 256850 170400
rect 261478 169804 261484 169856
rect 261536 169844 261542 169856
rect 265066 169844 265072 169856
rect 261536 169816 265072 169844
rect 261536 169804 261542 169816
rect 265066 169804 265072 169816
rect 265124 169804 265130 169856
rect 231210 169736 231216 169788
rect 231268 169776 231274 169788
rect 234614 169776 234620 169788
rect 231268 169748 234620 169776
rect 231268 169736 231274 169748
rect 234614 169736 234620 169748
rect 234672 169736 234678 169788
rect 234890 169736 234896 169788
rect 234948 169776 234954 169788
rect 238018 169776 238024 169788
rect 234948 169748 238024 169776
rect 234948 169736 234954 169748
rect 238018 169736 238024 169748
rect 238076 169736 238082 169788
rect 238294 169736 238300 169788
rect 238352 169776 238358 169788
rect 264974 169776 264980 169788
rect 238352 169748 264980 169776
rect 238352 169736 238358 169748
rect 264974 169736 264980 169748
rect 265032 169736 265038 169788
rect 169110 169668 169116 169720
rect 169168 169708 169174 169720
rect 214006 169708 214012 169720
rect 169168 169680 214012 169708
rect 169168 169668 169174 169680
rect 214006 169668 214012 169680
rect 214064 169668 214070 169720
rect 282822 169668 282828 169720
rect 282880 169708 282886 169720
rect 292850 169708 292856 169720
rect 282880 169680 292856 169708
rect 282880 169668 282886 169680
rect 292850 169668 292856 169680
rect 292908 169668 292914 169720
rect 174630 169600 174636 169652
rect 174688 169640 174694 169652
rect 213914 169640 213920 169652
rect 174688 169612 213920 169640
rect 174688 169600 174694 169612
rect 213914 169600 213920 169612
rect 213972 169600 213978 169652
rect 230566 169464 230572 169516
rect 230624 169504 230630 169516
rect 233234 169504 233240 169516
rect 230624 169476 233240 169504
rect 230624 169464 230630 169476
rect 233234 169464 233240 169476
rect 233292 169464 233298 169516
rect 231118 169396 231124 169448
rect 231176 169436 231182 169448
rect 234798 169436 234804 169448
rect 231176 169408 234804 169436
rect 231176 169396 231182 169408
rect 234798 169396 234804 169408
rect 234856 169396 234862 169448
rect 233878 168512 233884 168564
rect 233936 168552 233942 168564
rect 238754 168552 238760 168564
rect 233936 168524 238760 168552
rect 233936 168512 233942 168524
rect 238754 168512 238760 168524
rect 238812 168512 238818 168564
rect 243538 168444 243544 168496
rect 243596 168484 243602 168496
rect 264974 168484 264980 168496
rect 243596 168456 264980 168484
rect 243596 168444 243602 168456
rect 264974 168444 264980 168456
rect 265032 168444 265038 168496
rect 238018 168376 238024 168428
rect 238076 168416 238082 168428
rect 265066 168416 265072 168428
rect 238076 168388 265072 168416
rect 238076 168376 238082 168388
rect 265066 168376 265072 168388
rect 265124 168376 265130 168428
rect 166534 168308 166540 168360
rect 166592 168348 166598 168360
rect 214006 168348 214012 168360
rect 166592 168320 214012 168348
rect 166592 168308 166598 168320
rect 214006 168308 214012 168320
rect 214064 168308 214070 168360
rect 282270 168308 282276 168360
rect 282328 168348 282334 168360
rect 290090 168348 290096 168360
rect 282328 168320 290096 168348
rect 282328 168308 282334 168320
rect 290090 168308 290096 168320
rect 290148 168308 290154 168360
rect 173250 168240 173256 168292
rect 173308 168280 173314 168292
rect 213914 168280 213920 168292
rect 173308 168252 213920 168280
rect 173308 168240 173314 168252
rect 213914 168240 213920 168252
rect 213972 168240 213978 168292
rect 231394 168036 231400 168088
rect 231452 168076 231458 168088
rect 237466 168076 237472 168088
rect 231452 168048 237472 168076
rect 231452 168036 231458 168048
rect 237466 168036 237472 168048
rect 237524 168036 237530 168088
rect 231394 167084 231400 167136
rect 231452 167124 231458 167136
rect 236822 167124 236828 167136
rect 231452 167096 236828 167124
rect 231452 167084 231458 167096
rect 236822 167084 236828 167096
rect 236880 167084 236886 167136
rect 239766 167084 239772 167136
rect 239824 167124 239830 167136
rect 264974 167124 264980 167136
rect 239824 167096 264980 167124
rect 239824 167084 239830 167096
rect 264974 167084 264980 167096
rect 265032 167084 265038 167136
rect 236730 167016 236736 167068
rect 236788 167056 236794 167068
rect 265066 167056 265072 167068
rect 236788 167028 265072 167056
rect 236788 167016 236794 167028
rect 265066 167016 265072 167028
rect 265124 167016 265130 167068
rect 167730 166948 167736 167000
rect 167788 166988 167794 167000
rect 213914 166988 213920 167000
rect 167788 166960 213920 166988
rect 167788 166948 167794 166960
rect 213914 166948 213920 166960
rect 213972 166948 213978 167000
rect 566458 166948 566464 167000
rect 566516 166988 566522 167000
rect 580166 166988 580172 167000
rect 566516 166960 580172 166988
rect 566516 166948 566522 166960
rect 580166 166948 580172 166960
rect 580224 166948 580230 167000
rect 171778 166880 171784 166932
rect 171836 166920 171842 166932
rect 214006 166920 214012 166932
rect 171836 166892 214012 166920
rect 171836 166880 171842 166892
rect 214006 166880 214012 166892
rect 214064 166880 214070 166932
rect 231762 166676 231768 166728
rect 231820 166716 231826 166728
rect 234890 166716 234896 166728
rect 231820 166688 234896 166716
rect 231820 166676 231826 166688
rect 234890 166676 234896 166688
rect 234948 166676 234954 166728
rect 234062 166064 234068 166116
rect 234120 166104 234126 166116
rect 238938 166104 238944 166116
rect 234120 166076 238944 166104
rect 234120 166064 234126 166076
rect 238938 166064 238944 166076
rect 238996 166064 239002 166116
rect 245102 165656 245108 165708
rect 245160 165696 245166 165708
rect 265066 165696 265072 165708
rect 245160 165668 265072 165696
rect 245160 165656 245166 165668
rect 265066 165656 265072 165668
rect 265124 165656 265130 165708
rect 235258 165588 235264 165640
rect 235316 165628 235322 165640
rect 264974 165628 264980 165640
rect 235316 165600 264980 165628
rect 235316 165588 235322 165600
rect 264974 165588 264980 165600
rect 265032 165588 265038 165640
rect 166442 165520 166448 165572
rect 166500 165560 166506 165572
rect 214006 165560 214012 165572
rect 166500 165532 214012 165560
rect 166500 165520 166506 165532
rect 214006 165520 214012 165532
rect 214064 165520 214070 165572
rect 180150 165452 180156 165504
rect 180208 165492 180214 165504
rect 213914 165492 213920 165504
rect 180208 165464 213920 165492
rect 180208 165452 180214 165464
rect 213914 165452 213920 165464
rect 213972 165452 213978 165504
rect 281902 165316 281908 165368
rect 281960 165356 281966 165368
rect 284570 165356 284576 165368
rect 281960 165328 284576 165356
rect 281960 165316 281966 165328
rect 284570 165316 284576 165328
rect 284628 165316 284634 165368
rect 231486 165180 231492 165232
rect 231544 165220 231550 165232
rect 235442 165220 235448 165232
rect 231544 165192 235448 165220
rect 231544 165180 231550 165192
rect 235442 165180 235448 165192
rect 235500 165180 235506 165232
rect 253382 164296 253388 164348
rect 253440 164336 253446 164348
rect 264974 164336 264980 164348
rect 253440 164308 264980 164336
rect 253440 164296 253446 164308
rect 264974 164296 264980 164308
rect 265032 164296 265038 164348
rect 240778 164228 240784 164280
rect 240836 164268 240842 164280
rect 265066 164268 265072 164280
rect 240836 164240 265072 164268
rect 240836 164228 240842 164240
rect 265066 164228 265072 164240
rect 265124 164228 265130 164280
rect 3234 164160 3240 164212
rect 3292 164200 3298 164212
rect 40678 164200 40684 164212
rect 3292 164172 40684 164200
rect 3292 164160 3298 164172
rect 40678 164160 40684 164172
rect 40736 164160 40742 164212
rect 177390 164160 177396 164212
rect 177448 164200 177454 164212
rect 214006 164200 214012 164212
rect 177448 164172 214012 164200
rect 177448 164160 177454 164172
rect 214006 164160 214012 164172
rect 214064 164160 214070 164212
rect 230014 164160 230020 164212
rect 230072 164200 230078 164212
rect 230658 164200 230664 164212
rect 230072 164172 230664 164200
rect 230072 164160 230078 164172
rect 230658 164160 230664 164172
rect 230716 164160 230722 164212
rect 231026 164160 231032 164212
rect 231084 164200 231090 164212
rect 255406 164200 255412 164212
rect 231084 164172 255412 164200
rect 231084 164160 231090 164172
rect 255406 164160 255412 164172
rect 255464 164160 255470 164212
rect 196802 164092 196808 164144
rect 196860 164132 196866 164144
rect 213914 164132 213920 164144
rect 196860 164104 213920 164132
rect 196860 164092 196866 164104
rect 213914 164092 213920 164104
rect 213972 164092 213978 164144
rect 231670 164092 231676 164144
rect 231728 164132 231734 164144
rect 244366 164132 244372 164144
rect 231728 164104 244372 164132
rect 231728 164092 231734 164104
rect 244366 164092 244372 164104
rect 244424 164092 244430 164144
rect 282822 163276 282828 163328
rect 282880 163316 282886 163328
rect 288710 163316 288716 163328
rect 282880 163288 288716 163316
rect 282880 163276 282886 163288
rect 288710 163276 288716 163288
rect 288768 163276 288774 163328
rect 258902 162936 258908 162988
rect 258960 162976 258966 162988
rect 265066 162976 265072 162988
rect 258960 162948 265072 162976
rect 258960 162936 258966 162948
rect 265066 162936 265072 162948
rect 265124 162936 265130 162988
rect 245010 162868 245016 162920
rect 245068 162908 245074 162920
rect 264974 162908 264980 162920
rect 245068 162880 264980 162908
rect 245068 162868 245074 162880
rect 264974 162868 264980 162880
rect 265032 162868 265038 162920
rect 164878 162800 164884 162852
rect 164936 162840 164942 162852
rect 213914 162840 213920 162852
rect 164936 162812 213920 162840
rect 164936 162800 164942 162812
rect 213914 162800 213920 162812
rect 213972 162800 213978 162852
rect 230382 162800 230388 162852
rect 230440 162840 230446 162852
rect 230842 162840 230848 162852
rect 230440 162812 230848 162840
rect 230440 162800 230446 162812
rect 230842 162800 230848 162812
rect 230900 162800 230906 162852
rect 230934 162800 230940 162852
rect 230992 162840 230998 162852
rect 233510 162840 233516 162852
rect 230992 162812 233516 162840
rect 230992 162800 230998 162812
rect 233510 162800 233516 162812
rect 233568 162800 233574 162852
rect 282822 162800 282828 162852
rect 282880 162840 282886 162852
rect 296898 162840 296904 162852
rect 282880 162812 296904 162840
rect 282880 162800 282886 162812
rect 296898 162800 296904 162812
rect 296956 162800 296962 162852
rect 207750 162732 207756 162784
rect 207808 162772 207814 162784
rect 214006 162772 214012 162784
rect 207808 162744 214012 162772
rect 207808 162732 207814 162744
rect 214006 162732 214012 162744
rect 214064 162732 214070 162784
rect 184474 162120 184480 162172
rect 184532 162160 184538 162172
rect 207658 162160 207664 162172
rect 184532 162132 207664 162160
rect 184532 162120 184538 162132
rect 207658 162120 207664 162132
rect 207716 162120 207722 162172
rect 231118 162120 231124 162172
rect 231176 162160 231182 162172
rect 260282 162160 260288 162172
rect 231176 162132 260288 162160
rect 231176 162120 231182 162132
rect 260282 162120 260288 162132
rect 260340 162120 260346 162172
rect 262858 161644 262864 161696
rect 262916 161684 262922 161696
rect 265066 161684 265072 161696
rect 262916 161656 265072 161684
rect 262916 161644 262922 161656
rect 265066 161644 265072 161656
rect 265124 161644 265130 161696
rect 243906 161440 243912 161492
rect 243964 161480 243970 161492
rect 264974 161480 264980 161492
rect 243964 161452 264980 161480
rect 243964 161440 243970 161452
rect 264974 161440 264980 161452
rect 265032 161440 265038 161492
rect 166350 161372 166356 161424
rect 166408 161412 166414 161424
rect 214006 161412 214012 161424
rect 166408 161384 214012 161412
rect 166408 161372 166414 161384
rect 214006 161372 214012 161384
rect 214064 161372 214070 161424
rect 282822 161372 282828 161424
rect 282880 161412 282886 161424
rect 303798 161412 303804 161424
rect 282880 161384 303804 161412
rect 282880 161372 282886 161384
rect 303798 161372 303804 161384
rect 303856 161372 303862 161424
rect 170490 161304 170496 161356
rect 170548 161344 170554 161356
rect 213914 161344 213920 161356
rect 170548 161316 213920 161344
rect 170548 161304 170554 161316
rect 213914 161304 213920 161316
rect 213972 161304 213978 161356
rect 231670 160692 231676 160744
rect 231728 160732 231734 160744
rect 242986 160732 242992 160744
rect 231728 160704 242992 160732
rect 231728 160692 231734 160704
rect 242986 160692 242992 160704
rect 243044 160692 243050 160744
rect 281718 160556 281724 160608
rect 281776 160596 281782 160608
rect 284478 160596 284484 160608
rect 281776 160568 284484 160596
rect 281776 160556 281782 160568
rect 284478 160556 284484 160568
rect 284536 160556 284542 160608
rect 257430 160148 257436 160200
rect 257488 160188 257494 160200
rect 264974 160188 264980 160200
rect 257488 160160 264980 160188
rect 257488 160148 257494 160160
rect 264974 160148 264980 160160
rect 265032 160148 265038 160200
rect 234154 160080 234160 160132
rect 234212 160120 234218 160132
rect 265066 160120 265072 160132
rect 234212 160092 265072 160120
rect 234212 160080 234218 160092
rect 265066 160080 265072 160092
rect 265124 160080 265130 160132
rect 170398 160012 170404 160064
rect 170456 160052 170462 160064
rect 213914 160052 213920 160064
rect 170456 160024 213920 160052
rect 170456 160012 170462 160024
rect 213914 160012 213920 160024
rect 213972 160012 213978 160064
rect 231762 160012 231768 160064
rect 231820 160052 231826 160064
rect 248414 160052 248420 160064
rect 231820 160024 248420 160052
rect 231820 160012 231826 160024
rect 248414 160012 248420 160024
rect 248472 160012 248478 160064
rect 281902 160012 281908 160064
rect 281960 160052 281966 160064
rect 318794 160052 318800 160064
rect 281960 160024 318800 160052
rect 281960 160012 281966 160024
rect 318794 160012 318800 160024
rect 318852 160012 318858 160064
rect 231394 159944 231400 159996
rect 231452 159984 231458 159996
rect 240962 159984 240968 159996
rect 231452 159956 240968 159984
rect 231452 159944 231458 159956
rect 240962 159944 240968 159956
rect 241020 159944 241026 159996
rect 282362 159944 282368 159996
rect 282420 159984 282426 159996
rect 292758 159984 292764 159996
rect 282420 159956 292764 159984
rect 282420 159944 282426 159956
rect 292758 159944 292764 159956
rect 292816 159944 292822 159996
rect 254578 158788 254584 158840
rect 254636 158828 254642 158840
rect 264974 158828 264980 158840
rect 254636 158800 264980 158828
rect 254636 158788 254642 158800
rect 264974 158788 264980 158800
rect 265032 158788 265038 158840
rect 240870 158720 240876 158772
rect 240928 158760 240934 158772
rect 265066 158760 265072 158772
rect 240928 158732 265072 158760
rect 240928 158720 240934 158732
rect 265066 158720 265072 158732
rect 265124 158720 265130 158772
rect 169018 158652 169024 158704
rect 169076 158692 169082 158704
rect 214006 158692 214012 158704
rect 169076 158664 214012 158692
rect 169076 158652 169082 158664
rect 214006 158652 214012 158664
rect 214064 158652 214070 158704
rect 192478 158584 192484 158636
rect 192536 158624 192542 158636
rect 213914 158624 213920 158636
rect 192536 158596 213920 158624
rect 192536 158584 192542 158596
rect 213914 158584 213920 158596
rect 213972 158584 213978 158636
rect 231210 158584 231216 158636
rect 231268 158624 231274 158636
rect 235994 158624 236000 158636
rect 231268 158596 236000 158624
rect 231268 158584 231274 158596
rect 235994 158584 236000 158596
rect 236052 158584 236058 158636
rect 282822 157564 282828 157616
rect 282880 157604 282886 157616
rect 287330 157604 287336 157616
rect 282880 157576 287336 157604
rect 282880 157564 282886 157576
rect 287330 157564 287336 157576
rect 287388 157564 287394 157616
rect 249334 157428 249340 157480
rect 249392 157468 249398 157480
rect 264974 157468 264980 157480
rect 249392 157440 264980 157468
rect 249392 157428 249398 157440
rect 264974 157428 264980 157440
rect 265032 157428 265038 157480
rect 240962 157360 240968 157412
rect 241020 157400 241026 157412
rect 265066 157400 265072 157412
rect 241020 157372 265072 157400
rect 241020 157360 241026 157372
rect 265066 157360 265072 157372
rect 265124 157360 265130 157412
rect 167638 157292 167644 157344
rect 167696 157332 167702 157344
rect 214006 157332 214012 157344
rect 167696 157304 214012 157332
rect 167696 157292 167702 157304
rect 214006 157292 214012 157304
rect 214064 157292 214070 157344
rect 188522 157224 188528 157276
rect 188580 157264 188586 157276
rect 213914 157264 213920 157276
rect 188580 157236 213920 157264
rect 188580 157224 188586 157236
rect 213914 157224 213920 157236
rect 213972 157224 213978 157276
rect 231762 157224 231768 157276
rect 231820 157264 231826 157276
rect 244274 157264 244280 157276
rect 231820 157236 244280 157264
rect 231820 157224 231826 157236
rect 244274 157224 244280 157236
rect 244332 157224 244338 157276
rect 280062 156612 280068 156664
rect 280120 156652 280126 156664
rect 285858 156652 285864 156664
rect 280120 156624 285864 156652
rect 280120 156612 280126 156624
rect 285858 156612 285864 156624
rect 285916 156612 285922 156664
rect 247862 156000 247868 156052
rect 247920 156040 247926 156052
rect 264974 156040 264980 156052
rect 247920 156012 264980 156040
rect 247920 156000 247926 156012
rect 264974 156000 264980 156012
rect 265032 156000 265038 156052
rect 235534 155932 235540 155984
rect 235592 155972 235598 155984
rect 265066 155972 265072 155984
rect 235592 155944 265072 155972
rect 235592 155932 235598 155944
rect 265066 155932 265072 155944
rect 265124 155932 265130 155984
rect 166258 155864 166264 155916
rect 166316 155904 166322 155916
rect 214006 155904 214012 155916
rect 166316 155876 214012 155904
rect 166316 155864 166322 155876
rect 214006 155864 214012 155876
rect 214064 155864 214070 155916
rect 281626 155864 281632 155916
rect 281684 155904 281690 155916
rect 321554 155904 321560 155916
rect 281684 155876 321560 155904
rect 281684 155864 281690 155876
rect 321554 155864 321560 155876
rect 321612 155864 321618 155916
rect 184566 155796 184572 155848
rect 184624 155836 184630 155848
rect 213914 155836 213920 155848
rect 184624 155808 213920 155836
rect 184624 155796 184630 155808
rect 213914 155796 213920 155808
rect 213972 155796 213978 155848
rect 231486 155796 231492 155848
rect 231544 155836 231550 155848
rect 234062 155836 234068 155848
rect 231544 155808 234068 155836
rect 231544 155796 231550 155808
rect 234062 155796 234068 155808
rect 234120 155796 234126 155848
rect 231670 155184 231676 155236
rect 231728 155224 231734 155236
rect 240410 155224 240416 155236
rect 231728 155196 240416 155224
rect 231728 155184 231734 155196
rect 240410 155184 240416 155196
rect 240468 155184 240474 155236
rect 250530 154640 250536 154692
rect 250588 154680 250594 154692
rect 264974 154680 264980 154692
rect 250588 154652 264980 154680
rect 250588 154640 250594 154652
rect 264974 154640 264980 154652
rect 265032 154640 265038 154692
rect 238110 154572 238116 154624
rect 238168 154612 238174 154624
rect 265158 154612 265164 154624
rect 238168 154584 265164 154612
rect 238168 154572 238174 154584
rect 265158 154572 265164 154584
rect 265216 154572 265222 154624
rect 231486 154504 231492 154556
rect 231544 154544 231550 154556
rect 242894 154544 242900 154556
rect 231544 154516 242900 154544
rect 231544 154504 231550 154516
rect 242894 154504 242900 154516
rect 242952 154504 242958 154556
rect 231762 154436 231768 154488
rect 231820 154476 231826 154488
rect 241606 154476 241612 154488
rect 231820 154448 241612 154476
rect 231820 154436 231826 154448
rect 241606 154436 241612 154448
rect 241664 154436 241670 154488
rect 281626 154436 281632 154488
rect 281684 154476 281690 154488
rect 295610 154476 295616 154488
rect 281684 154448 295616 154476
rect 281684 154436 281690 154448
rect 295610 154436 295616 154448
rect 295668 154436 295674 154488
rect 206370 153280 206376 153332
rect 206428 153320 206434 153332
rect 213914 153320 213920 153332
rect 206428 153292 213920 153320
rect 206428 153280 206434 153292
rect 213914 153280 213920 153292
rect 213972 153280 213978 153332
rect 249058 153280 249064 153332
rect 249116 153320 249122 153332
rect 264974 153320 264980 153332
rect 249116 153292 264980 153320
rect 249116 153280 249122 153292
rect 264974 153280 264980 153292
rect 265032 153280 265038 153332
rect 198182 153212 198188 153264
rect 198240 153252 198246 153264
rect 214006 153252 214012 153264
rect 198240 153224 214012 153252
rect 198240 153212 198246 153224
rect 214006 153212 214012 153224
rect 214064 153212 214070 153264
rect 243722 153212 243728 153264
rect 243780 153252 243786 153264
rect 265066 153252 265072 153264
rect 243780 153224 265072 153252
rect 243780 153212 243786 153224
rect 265066 153212 265072 153224
rect 265124 153212 265130 153264
rect 281626 153144 281632 153196
rect 281684 153184 281690 153196
rect 296990 153184 296996 153196
rect 281684 153156 296996 153184
rect 281684 153144 281690 153156
rect 296990 153144 296996 153156
rect 297048 153144 297054 153196
rect 231486 152940 231492 152992
rect 231544 152980 231550 152992
rect 237374 152980 237380 152992
rect 231544 152952 237380 152980
rect 231544 152940 231550 152952
rect 237374 152940 237380 152952
rect 237432 152940 237438 152992
rect 236914 152464 236920 152516
rect 236972 152504 236978 152516
rect 265342 152504 265348 152516
rect 236972 152476 265348 152504
rect 236972 152464 236978 152476
rect 265342 152464 265348 152476
rect 265400 152464 265406 152516
rect 281626 152464 281632 152516
rect 281684 152504 281690 152516
rect 295518 152504 295524 152516
rect 281684 152476 295524 152504
rect 281684 152464 281690 152476
rect 295518 152464 295524 152476
rect 295576 152464 295582 152516
rect 211798 152192 211804 152244
rect 211856 152232 211862 152244
rect 214006 152232 214012 152244
rect 211856 152204 214012 152232
rect 211856 152192 211862 152204
rect 214006 152192 214012 152204
rect 214064 152192 214070 152244
rect 252002 151784 252008 151836
rect 252060 151824 252066 151836
rect 264974 151824 264980 151836
rect 252060 151796 264980 151824
rect 252060 151784 252066 151796
rect 264974 151784 264980 151796
rect 265032 151784 265038 151836
rect 231486 151716 231492 151768
rect 231544 151756 231550 151768
rect 245930 151756 245936 151768
rect 231544 151728 245936 151756
rect 231544 151716 231550 151728
rect 245930 151716 245936 151728
rect 245988 151716 245994 151768
rect 281810 151036 281816 151088
rect 281868 151076 281874 151088
rect 300854 151076 300860 151088
rect 281868 151048 300860 151076
rect 281868 151036 281874 151048
rect 300854 151036 300860 151048
rect 300912 151036 300918 151088
rect 231670 150900 231676 150952
rect 231728 150940 231734 150952
rect 234706 150940 234712 150952
rect 231728 150912 234712 150940
rect 231728 150900 231734 150912
rect 234706 150900 234712 150912
rect 234764 150900 234770 150952
rect 187142 150492 187148 150544
rect 187200 150532 187206 150544
rect 213914 150532 213920 150544
rect 187200 150504 213920 150532
rect 187200 150492 187206 150504
rect 213914 150492 213920 150504
rect 213972 150492 213978 150544
rect 247770 150492 247776 150544
rect 247828 150532 247834 150544
rect 264974 150532 264980 150544
rect 247828 150504 264980 150532
rect 247828 150492 247834 150504
rect 264974 150492 264980 150504
rect 265032 150492 265038 150544
rect 169110 150424 169116 150476
rect 169168 150464 169174 150476
rect 214006 150464 214012 150476
rect 169168 150436 214012 150464
rect 169168 150424 169174 150436
rect 214006 150424 214012 150436
rect 214064 150424 214070 150476
rect 235442 150424 235448 150476
rect 235500 150464 235506 150476
rect 265066 150464 265072 150476
rect 235500 150436 265072 150464
rect 235500 150424 235506 150436
rect 265066 150424 265072 150436
rect 265124 150424 265130 150476
rect 3510 150356 3516 150408
rect 3568 150396 3574 150408
rect 11698 150396 11704 150408
rect 3568 150368 11704 150396
rect 3568 150356 3574 150368
rect 11698 150356 11704 150368
rect 11756 150356 11762 150408
rect 182910 150356 182916 150408
rect 182968 150396 182974 150408
rect 214098 150396 214104 150408
rect 182968 150368 214104 150396
rect 182968 150356 182974 150368
rect 214098 150356 214104 150368
rect 214156 150356 214162 150408
rect 281626 150356 281632 150408
rect 281684 150396 281690 150408
rect 294138 150396 294144 150408
rect 281684 150368 294144 150396
rect 281684 150356 281690 150368
rect 294138 150356 294144 150368
rect 294196 150356 294202 150408
rect 281718 150288 281724 150340
rect 281776 150328 281782 150340
rect 292666 150328 292672 150340
rect 281776 150300 292672 150328
rect 281776 150288 281782 150300
rect 292666 150288 292672 150300
rect 292724 150288 292730 150340
rect 173158 149676 173164 149728
rect 173216 149716 173222 149728
rect 213914 149716 213920 149728
rect 173216 149688 213920 149716
rect 173216 149676 173222 149688
rect 213914 149676 213920 149688
rect 213972 149676 213978 149728
rect 232682 149676 232688 149728
rect 232740 149716 232746 149728
rect 265618 149716 265624 149728
rect 232740 149688 265624 149716
rect 232740 149676 232746 149688
rect 265618 149676 265624 149688
rect 265676 149676 265682 149728
rect 244918 149064 244924 149116
rect 244976 149104 244982 149116
rect 264974 149104 264980 149116
rect 244976 149076 264980 149104
rect 244976 149064 244982 149076
rect 264974 149064 264980 149076
rect 265032 149064 265038 149116
rect 281626 148996 281632 149048
rect 281684 149036 281690 149048
rect 294046 149036 294052 149048
rect 281684 149008 294052 149036
rect 281684 148996 281690 149008
rect 294046 148996 294052 149008
rect 294104 148996 294110 149048
rect 231486 148792 231492 148844
rect 231544 148832 231550 148844
rect 233878 148832 233884 148844
rect 231544 148804 233884 148832
rect 231544 148792 231550 148804
rect 233878 148792 233884 148804
rect 233936 148792 233942 148844
rect 232866 148316 232872 148368
rect 232924 148356 232930 148368
rect 265158 148356 265164 148368
rect 232924 148328 265164 148356
rect 232924 148316 232930 148328
rect 265158 148316 265164 148328
rect 265216 148316 265222 148368
rect 173250 147636 173256 147688
rect 173308 147676 173314 147688
rect 213914 147676 213920 147688
rect 173308 147648 213920 147676
rect 173308 147636 173314 147648
rect 213914 147636 213920 147648
rect 213972 147636 213978 147688
rect 229922 147636 229928 147688
rect 229980 147676 229986 147688
rect 232130 147676 232136 147688
rect 229980 147648 232136 147676
rect 229980 147636 229986 147648
rect 232130 147636 232136 147648
rect 232188 147636 232194 147688
rect 238202 147636 238208 147688
rect 238260 147676 238266 147688
rect 264974 147676 264980 147688
rect 238260 147648 264980 147676
rect 238260 147636 238266 147648
rect 264974 147636 264980 147648
rect 265032 147636 265038 147688
rect 282822 147568 282828 147620
rect 282880 147608 282886 147620
rect 306650 147608 306656 147620
rect 282880 147580 306656 147608
rect 282880 147568 282886 147580
rect 306650 147568 306656 147580
rect 306708 147568 306714 147620
rect 181438 146888 181444 146940
rect 181496 146928 181502 146940
rect 192478 146928 192484 146940
rect 181496 146900 192484 146928
rect 181496 146888 181502 146900
rect 192478 146888 192484 146900
rect 192536 146888 192542 146940
rect 192570 146888 192576 146940
rect 192628 146928 192634 146940
rect 204990 146928 204996 146940
rect 192628 146900 204996 146928
rect 192628 146888 192634 146900
rect 204990 146888 204996 146900
rect 205048 146888 205054 146940
rect 206278 146888 206284 146940
rect 206336 146928 206342 146940
rect 214558 146928 214564 146940
rect 206336 146900 214564 146928
rect 206336 146888 206342 146900
rect 214558 146888 214564 146900
rect 214616 146888 214622 146940
rect 262766 146344 262772 146396
rect 262824 146384 262830 146396
rect 265066 146384 265072 146396
rect 262824 146356 265072 146384
rect 262824 146344 262830 146356
rect 265066 146344 265072 146356
rect 265124 146344 265130 146396
rect 166258 146276 166264 146328
rect 166316 146316 166322 146328
rect 213914 146316 213920 146328
rect 166316 146288 213920 146316
rect 166316 146276 166322 146288
rect 213914 146276 213920 146288
rect 213972 146276 213978 146328
rect 256050 146276 256056 146328
rect 256108 146316 256114 146328
rect 264974 146316 264980 146328
rect 256108 146288 264980 146316
rect 256108 146276 256114 146288
rect 264974 146276 264980 146288
rect 265032 146276 265038 146328
rect 231670 146208 231676 146260
rect 231728 146248 231734 146260
rect 245838 146248 245844 146260
rect 231728 146220 245844 146248
rect 231728 146208 231734 146220
rect 245838 146208 245844 146220
rect 245896 146208 245902 146260
rect 282362 146208 282368 146260
rect 282420 146248 282426 146260
rect 291470 146248 291476 146260
rect 282420 146220 291476 146248
rect 282420 146208 282426 146220
rect 291470 146208 291476 146220
rect 291528 146208 291534 146260
rect 184290 145528 184296 145580
rect 184348 145568 184354 145580
rect 214006 145568 214012 145580
rect 184348 145540 214012 145568
rect 184348 145528 184354 145540
rect 214006 145528 214012 145540
rect 214064 145528 214070 145580
rect 262582 144984 262588 145036
rect 262640 145024 262646 145036
rect 265066 145024 265072 145036
rect 262640 144996 265072 145024
rect 262640 144984 262646 144996
rect 265066 144984 265072 144996
rect 265124 144984 265130 145036
rect 201402 144916 201408 144968
rect 201460 144956 201466 144968
rect 213914 144956 213920 144968
rect 201460 144928 213920 144956
rect 201460 144916 201466 144928
rect 213914 144916 213920 144928
rect 213972 144916 213978 144968
rect 246574 144916 246580 144968
rect 246632 144956 246638 144968
rect 264974 144956 264980 144968
rect 246632 144928 264980 144956
rect 246632 144916 246638 144928
rect 264974 144916 264980 144928
rect 265032 144916 265038 144968
rect 231210 144848 231216 144900
rect 231268 144888 231274 144900
rect 238294 144888 238300 144900
rect 231268 144860 238300 144888
rect 231268 144848 231274 144860
rect 238294 144848 238300 144860
rect 238352 144848 238358 144900
rect 167638 144168 167644 144220
rect 167696 144208 167702 144220
rect 201402 144208 201408 144220
rect 167696 144180 201408 144208
rect 167696 144168 167702 144180
rect 201402 144168 201408 144180
rect 201460 144168 201466 144220
rect 236822 144168 236828 144220
rect 236880 144208 236886 144220
rect 262766 144208 262772 144220
rect 236880 144180 262772 144208
rect 236880 144168 236886 144180
rect 262766 144168 262772 144180
rect 262824 144168 262830 144220
rect 209038 143624 209044 143676
rect 209096 143664 209102 143676
rect 213914 143664 213920 143676
rect 209096 143636 213920 143664
rect 209096 143624 209102 143636
rect 213914 143624 213920 143636
rect 213972 143624 213978 143676
rect 184382 143556 184388 143608
rect 184440 143596 184446 143608
rect 214006 143596 214012 143608
rect 184440 143568 214012 143596
rect 184440 143556 184446 143568
rect 214006 143556 214012 143568
rect 214064 143556 214070 143608
rect 252094 143556 252100 143608
rect 252152 143596 252158 143608
rect 264974 143596 264980 143608
rect 252152 143568 264980 143596
rect 252152 143556 252158 143568
rect 264974 143556 264980 143568
rect 265032 143556 265038 143608
rect 282822 143488 282828 143540
rect 282880 143528 282886 143540
rect 289998 143528 290004 143540
rect 282880 143500 290004 143528
rect 282880 143488 282886 143500
rect 289998 143488 290004 143500
rect 290056 143488 290062 143540
rect 231670 143420 231676 143472
rect 231728 143460 231734 143472
rect 234246 143460 234252 143472
rect 231728 143432 234252 143460
rect 231728 143420 231734 143432
rect 234246 143420 234252 143432
rect 234304 143420 234310 143472
rect 231302 142876 231308 142928
rect 231360 142916 231366 142928
rect 254670 142916 254676 142928
rect 231360 142888 254676 142916
rect 231360 142876 231366 142888
rect 254670 142876 254676 142888
rect 254728 142876 254734 142928
rect 238386 142808 238392 142860
rect 238444 142848 238450 142860
rect 262582 142848 262588 142860
rect 238444 142820 262588 142848
rect 238444 142808 238450 142820
rect 262582 142808 262588 142820
rect 262640 142808 262646 142860
rect 258810 142740 258816 142792
rect 258868 142780 258874 142792
rect 264974 142780 264980 142792
rect 258868 142752 264980 142780
rect 258868 142740 258874 142752
rect 264974 142740 264980 142752
rect 265032 142740 265038 142792
rect 177482 142128 177488 142180
rect 177540 142168 177546 142180
rect 213914 142168 213920 142180
rect 177540 142140 213920 142168
rect 177540 142128 177546 142140
rect 213914 142128 213920 142140
rect 213972 142128 213978 142180
rect 282086 142060 282092 142112
rect 282144 142100 282150 142112
rect 299474 142100 299480 142112
rect 282144 142072 299480 142100
rect 282144 142060 282150 142072
rect 299474 142060 299480 142072
rect 299532 142060 299538 142112
rect 282822 141992 282828 142044
rect 282880 142032 282886 142044
rect 298278 142032 298284 142044
rect 282880 142004 298284 142032
rect 282880 141992 282886 142004
rect 298278 141992 298284 142004
rect 298336 141992 298342 142044
rect 180058 141380 180064 141432
rect 180116 141420 180122 141432
rect 200758 141420 200764 141432
rect 180116 141392 200764 141420
rect 180116 141380 180122 141392
rect 200758 141380 200764 141392
rect 200816 141380 200822 141432
rect 250806 141380 250812 141432
rect 250864 141420 250870 141432
rect 265710 141420 265716 141432
rect 250864 141392 265716 141420
rect 250864 141380 250870 141392
rect 265710 141380 265716 141392
rect 265768 141380 265774 141432
rect 231118 141312 231124 141364
rect 231176 141352 231182 141364
rect 233878 141352 233884 141364
rect 231176 141324 233884 141352
rect 231176 141312 231182 141324
rect 233878 141312 233884 141324
rect 233936 141312 233942 141364
rect 203518 140768 203524 140820
rect 203576 140808 203582 140820
rect 213914 140808 213920 140820
rect 203576 140780 213920 140808
rect 203576 140768 203582 140780
rect 213914 140768 213920 140780
rect 213972 140768 213978 140820
rect 231762 140700 231768 140752
rect 231820 140740 231826 140752
rect 247126 140740 247132 140752
rect 231820 140712 247132 140740
rect 231820 140700 231826 140712
rect 247126 140700 247132 140712
rect 247184 140700 247190 140752
rect 282822 140700 282828 140752
rect 282880 140740 282886 140752
rect 313366 140740 313372 140752
rect 282880 140712 313372 140740
rect 282880 140700 282886 140712
rect 313366 140700 313372 140712
rect 313424 140700 313430 140752
rect 231670 140020 231676 140072
rect 231728 140060 231734 140072
rect 247678 140060 247684 140072
rect 231728 140032 247684 140060
rect 231728 140020 231734 140032
rect 247678 140020 247684 140032
rect 247736 140020 247742 140072
rect 189718 139408 189724 139460
rect 189776 139448 189782 139460
rect 213914 139448 213920 139460
rect 189776 139420 213920 139448
rect 189776 139408 189782 139420
rect 213914 139408 213920 139420
rect 213972 139408 213978 139460
rect 263042 139408 263048 139460
rect 263100 139448 263106 139460
rect 265342 139448 265348 139460
rect 263100 139420 265348 139448
rect 263100 139408 263106 139420
rect 265342 139408 265348 139420
rect 265400 139408 265406 139460
rect 282822 139340 282828 139392
rect 282880 139380 282886 139392
rect 302510 139380 302516 139392
rect 282880 139352 302516 139380
rect 282880 139340 282886 139352
rect 302510 139340 302516 139352
rect 302568 139340 302574 139392
rect 231486 138864 231492 138916
rect 231544 138904 231550 138916
rect 235350 138904 235356 138916
rect 231544 138876 235356 138904
rect 231544 138864 231550 138876
rect 235350 138864 235356 138876
rect 235408 138864 235414 138916
rect 176010 138660 176016 138712
rect 176068 138700 176074 138712
rect 214006 138700 214012 138712
rect 176068 138672 214012 138700
rect 176068 138660 176074 138672
rect 214006 138660 214012 138672
rect 214064 138660 214070 138712
rect 202138 137980 202144 138032
rect 202196 138020 202202 138032
rect 213914 138020 213920 138032
rect 202196 137992 213920 138020
rect 202196 137980 202202 137992
rect 213914 137980 213920 137992
rect 213972 137980 213978 138032
rect 233878 137980 233884 138032
rect 233936 138020 233942 138032
rect 264974 138020 264980 138032
rect 233936 137992 264980 138020
rect 233936 137980 233942 137992
rect 264974 137980 264980 137992
rect 265032 137980 265038 138032
rect 265710 137980 265716 138032
rect 265768 138020 265774 138032
rect 267090 138020 267096 138032
rect 265768 137992 267096 138020
rect 265768 137980 265774 137992
rect 267090 137980 267096 137992
rect 267148 137980 267154 138032
rect 3510 137912 3516 137964
rect 3568 137952 3574 137964
rect 17218 137952 17224 137964
rect 3568 137924 17224 137952
rect 3568 137912 3574 137924
rect 17218 137912 17224 137924
rect 17276 137912 17282 137964
rect 231578 137912 231584 137964
rect 231636 137952 231642 137964
rect 251358 137952 251364 137964
rect 231636 137924 251364 137952
rect 231636 137912 231642 137924
rect 251358 137912 251364 137924
rect 251416 137912 251422 137964
rect 282822 137912 282828 137964
rect 282880 137952 282886 137964
rect 299658 137952 299664 137964
rect 282880 137924 299664 137952
rect 282880 137912 282886 137924
rect 299658 137912 299664 137924
rect 299716 137912 299722 137964
rect 198090 136688 198096 136740
rect 198148 136728 198154 136740
rect 213914 136728 213920 136740
rect 198148 136700 213920 136728
rect 198148 136688 198154 136700
rect 213914 136688 213920 136700
rect 213972 136688 213978 136740
rect 171778 136620 171784 136672
rect 171836 136660 171842 136672
rect 214006 136660 214012 136672
rect 171836 136632 214012 136660
rect 171836 136620 171842 136632
rect 214006 136620 214012 136632
rect 214064 136620 214070 136672
rect 247678 136620 247684 136672
rect 247736 136660 247742 136672
rect 264974 136660 264980 136672
rect 247736 136632 264980 136660
rect 247736 136620 247742 136632
rect 264974 136620 264980 136632
rect 265032 136620 265038 136672
rect 230566 136552 230572 136604
rect 230624 136592 230630 136604
rect 232682 136592 232688 136604
rect 230624 136564 232688 136592
rect 230624 136552 230630 136564
rect 232682 136552 232688 136564
rect 232740 136552 232746 136604
rect 282822 136552 282828 136604
rect 282880 136592 282886 136604
rect 303890 136592 303896 136604
rect 282880 136564 303896 136592
rect 282880 136552 282886 136564
rect 303890 136552 303896 136564
rect 303948 136552 303954 136604
rect 167822 135872 167828 135924
rect 167880 135912 167886 135924
rect 213178 135912 213184 135924
rect 167880 135884 213184 135912
rect 167880 135872 167886 135884
rect 213178 135872 213184 135884
rect 213236 135872 213242 135924
rect 231486 135872 231492 135924
rect 231544 135912 231550 135924
rect 236638 135912 236644 135924
rect 231544 135884 236644 135912
rect 231544 135872 231550 135884
rect 236638 135872 236644 135884
rect 236696 135872 236702 135924
rect 243630 135328 243636 135380
rect 243688 135368 243694 135380
rect 264974 135368 264980 135380
rect 243688 135340 264980 135368
rect 243688 135328 243694 135340
rect 264974 135328 264980 135340
rect 265032 135328 265038 135380
rect 180058 135260 180064 135312
rect 180116 135300 180122 135312
rect 213914 135300 213920 135312
rect 180116 135272 213920 135300
rect 180116 135260 180122 135272
rect 213914 135260 213920 135272
rect 213972 135260 213978 135312
rect 235350 135260 235356 135312
rect 235408 135300 235414 135312
rect 265066 135300 265072 135312
rect 235408 135272 265072 135300
rect 235408 135260 235414 135272
rect 265066 135260 265072 135272
rect 265124 135260 265130 135312
rect 231578 135192 231584 135244
rect 231636 135232 231642 135244
rect 264238 135232 264244 135244
rect 231636 135204 264244 135232
rect 231636 135192 231642 135204
rect 264238 135192 264244 135204
rect 264296 135192 264302 135244
rect 282454 135124 282460 135176
rect 282512 135164 282518 135176
rect 285950 135164 285956 135176
rect 282512 135136 285956 135164
rect 282512 135124 282518 135136
rect 285950 135124 285956 135136
rect 286008 135124 286014 135176
rect 192570 134512 192576 134564
rect 192628 134552 192634 134564
rect 214098 134552 214104 134564
rect 192628 134524 214104 134552
rect 192628 134512 192634 134524
rect 214098 134512 214104 134524
rect 214156 134512 214162 134564
rect 230750 134512 230756 134564
rect 230808 134552 230814 134564
rect 239766 134552 239772 134564
rect 230808 134524 239772 134552
rect 230808 134512 230814 134524
rect 239766 134512 239772 134524
rect 239824 134512 239830 134564
rect 173158 133900 173164 133952
rect 173216 133940 173222 133952
rect 213914 133940 213920 133952
rect 173216 133912 213920 133940
rect 173216 133900 173222 133912
rect 213914 133900 213920 133912
rect 213972 133900 213978 133952
rect 239490 133900 239496 133952
rect 239548 133940 239554 133952
rect 264974 133940 264980 133952
rect 239548 133912 264980 133940
rect 239548 133900 239554 133912
rect 264974 133900 264980 133912
rect 265032 133900 265038 133952
rect 230842 133832 230848 133884
rect 230900 133872 230906 133884
rect 257614 133872 257620 133884
rect 230900 133844 257620 133872
rect 230900 133832 230906 133844
rect 257614 133832 257620 133844
rect 257672 133832 257678 133884
rect 282730 133832 282736 133884
rect 282788 133872 282794 133884
rect 311986 133872 311992 133884
rect 282788 133844 311992 133872
rect 282788 133832 282794 133844
rect 311986 133832 311992 133844
rect 312044 133832 312050 133884
rect 231762 133764 231768 133816
rect 231820 133804 231826 133816
rect 249242 133804 249248 133816
rect 231820 133776 249248 133804
rect 231820 133764 231826 133776
rect 249242 133764 249248 133776
rect 249300 133764 249306 133816
rect 282822 133764 282828 133816
rect 282880 133804 282886 133816
rect 300946 133804 300952 133816
rect 282880 133776 300952 133804
rect 282880 133764 282886 133776
rect 300946 133764 300952 133776
rect 301004 133764 301010 133816
rect 174630 133152 174636 133204
rect 174688 133192 174694 133204
rect 206370 133192 206376 133204
rect 174688 133164 206376 133192
rect 174688 133152 174694 133164
rect 206370 133152 206376 133164
rect 206428 133152 206434 133204
rect 249426 133152 249432 133204
rect 249484 133192 249490 133204
rect 265802 133192 265808 133204
rect 249484 133164 265808 133192
rect 249484 133152 249490 133164
rect 265802 133152 265808 133164
rect 265860 133152 265866 133204
rect 209130 132540 209136 132592
rect 209188 132580 209194 132592
rect 213914 132580 213920 132592
rect 209188 132552 213920 132580
rect 209188 132540 209194 132552
rect 213914 132540 213920 132552
rect 213972 132540 213978 132592
rect 181438 132472 181444 132524
rect 181496 132512 181502 132524
rect 214006 132512 214012 132524
rect 181496 132484 214012 132512
rect 181496 132472 181502 132484
rect 214006 132472 214012 132484
rect 214064 132472 214070 132524
rect 257338 132472 257344 132524
rect 257396 132512 257402 132524
rect 264974 132512 264980 132524
rect 257396 132484 264980 132512
rect 257396 132472 257402 132484
rect 264974 132472 264980 132484
rect 265032 132472 265038 132524
rect 231670 132404 231676 132456
rect 231728 132444 231734 132456
rect 261478 132444 261484 132456
rect 231728 132416 261484 132444
rect 231728 132404 231734 132416
rect 261478 132404 261484 132416
rect 261536 132404 261542 132456
rect 282822 132404 282828 132456
rect 282880 132444 282886 132456
rect 316126 132444 316132 132456
rect 282880 132416 316132 132444
rect 282880 132404 282886 132416
rect 316126 132404 316132 132416
rect 316184 132404 316190 132456
rect 231118 131724 231124 131776
rect 231176 131764 231182 131776
rect 253474 131764 253480 131776
rect 231176 131736 253480 131764
rect 231176 131724 231182 131736
rect 253474 131724 253480 131736
rect 253532 131724 253538 131776
rect 210510 131180 210516 131232
rect 210568 131220 210574 131232
rect 214006 131220 214012 131232
rect 210568 131192 214012 131220
rect 210568 131180 210574 131192
rect 214006 131180 214012 131192
rect 214064 131180 214070 131232
rect 195514 131112 195520 131164
rect 195572 131152 195578 131164
rect 213914 131152 213920 131164
rect 195572 131124 213920 131152
rect 195572 131112 195578 131124
rect 213914 131112 213920 131124
rect 213972 131112 213978 131164
rect 260466 131112 260472 131164
rect 260524 131152 260530 131164
rect 264974 131152 264980 131164
rect 260524 131124 264980 131152
rect 260524 131112 260530 131124
rect 264974 131112 264980 131124
rect 265032 131112 265038 131164
rect 230566 131044 230572 131096
rect 230624 131084 230630 131096
rect 243538 131084 243544 131096
rect 230624 131056 243544 131084
rect 230624 131044 230630 131056
rect 243538 131044 243544 131056
rect 243596 131044 243602 131096
rect 282822 131044 282828 131096
rect 282880 131084 282886 131096
rect 307754 131084 307760 131096
rect 282880 131056 307760 131084
rect 282880 131044 282886 131056
rect 307754 131044 307760 131056
rect 307812 131044 307818 131096
rect 282730 130976 282736 131028
rect 282788 131016 282794 131028
rect 307846 131016 307852 131028
rect 282788 130988 307852 131016
rect 282788 130976 282794 130988
rect 307846 130976 307852 130988
rect 307904 130976 307910 131028
rect 231670 129888 231676 129940
rect 231728 129928 231734 129940
rect 238018 129928 238024 129940
rect 231728 129900 238024 129928
rect 231728 129888 231734 129900
rect 238018 129888 238024 129900
rect 238076 129888 238082 129940
rect 180150 129752 180156 129804
rect 180208 129792 180214 129804
rect 213914 129792 213920 129804
rect 180208 129764 213920 129792
rect 180208 129752 180214 129764
rect 213914 129752 213920 129764
rect 213972 129752 213978 129804
rect 254670 129752 254676 129804
rect 254728 129792 254734 129804
rect 264974 129792 264980 129804
rect 254728 129764 264980 129792
rect 254728 129752 254734 129764
rect 264974 129752 264980 129764
rect 265032 129752 265038 129804
rect 231762 129684 231768 129736
rect 231820 129724 231826 129736
rect 239674 129724 239680 129736
rect 231820 129696 239680 129724
rect 231820 129684 231826 129696
rect 239674 129684 239680 129696
rect 239732 129684 239738 129736
rect 281810 129684 281816 129736
rect 281868 129724 281874 129736
rect 284294 129724 284300 129736
rect 281868 129696 284300 129724
rect 281868 129684 281874 129696
rect 284294 129684 284300 129696
rect 284352 129684 284358 129736
rect 178770 129004 178776 129056
rect 178828 129044 178834 129056
rect 214834 129044 214840 129056
rect 178828 129016 214840 129044
rect 178828 129004 178834 129016
rect 214834 129004 214840 129016
rect 214892 129004 214898 129056
rect 230934 129004 230940 129056
rect 230992 129044 230998 129056
rect 258902 129044 258908 129056
rect 230992 129016 258908 129044
rect 230992 129004 230998 129016
rect 258902 129004 258908 129016
rect 258960 129004 258966 129056
rect 283558 129004 283564 129056
rect 283616 129044 283622 129056
rect 301130 129044 301136 129056
rect 283616 129016 301136 129044
rect 283616 129004 283622 129016
rect 301130 129004 301136 129016
rect 301188 129004 301194 129056
rect 207750 128324 207756 128376
rect 207808 128364 207814 128376
rect 213914 128364 213920 128376
rect 207808 128336 213920 128364
rect 207808 128324 207814 128336
rect 213914 128324 213920 128336
rect 213972 128324 213978 128376
rect 243814 128324 243820 128376
rect 243872 128364 243878 128376
rect 247678 128364 247684 128376
rect 243872 128336 247684 128364
rect 243872 128324 243878 128336
rect 247678 128324 247684 128336
rect 247736 128324 247742 128376
rect 261478 128324 261484 128376
rect 261536 128364 261542 128376
rect 265158 128364 265164 128376
rect 261536 128336 265164 128364
rect 261536 128324 261542 128336
rect 265158 128324 265164 128336
rect 265216 128324 265222 128376
rect 282822 128256 282828 128308
rect 282880 128296 282886 128308
rect 314746 128296 314752 128308
rect 282880 128268 314752 128296
rect 282880 128256 282886 128268
rect 314746 128256 314752 128268
rect 314804 128256 314810 128308
rect 282730 128188 282736 128240
rect 282788 128228 282794 128240
rect 305086 128228 305092 128240
rect 282788 128200 305092 128228
rect 282788 128188 282794 128200
rect 305086 128188 305092 128200
rect 305144 128188 305150 128240
rect 231762 127916 231768 127968
rect 231820 127956 231826 127968
rect 236730 127956 236736 127968
rect 231820 127928 236736 127956
rect 231820 127916 231826 127928
rect 236730 127916 236736 127928
rect 236788 127916 236794 127968
rect 230566 127644 230572 127696
rect 230624 127684 230630 127696
rect 245102 127684 245108 127696
rect 230624 127656 245108 127684
rect 230624 127644 230630 127656
rect 245102 127644 245108 127656
rect 245160 127644 245166 127696
rect 241054 127576 241060 127628
rect 241112 127616 241118 127628
rect 264974 127616 264980 127628
rect 241112 127588 264980 127616
rect 241112 127576 241118 127588
rect 264974 127576 264980 127588
rect 265032 127576 265038 127628
rect 203610 127032 203616 127084
rect 203668 127072 203674 127084
rect 213914 127072 213920 127084
rect 203668 127044 213920 127072
rect 203668 127032 203674 127044
rect 213914 127032 213920 127044
rect 213972 127032 213978 127084
rect 170398 126964 170404 127016
rect 170456 127004 170462 127016
rect 214006 127004 214012 127016
rect 170456 126976 214012 127004
rect 170456 126964 170462 126976
rect 214006 126964 214012 126976
rect 214064 126964 214070 127016
rect 247678 126964 247684 127016
rect 247736 127004 247742 127016
rect 264974 127004 264980 127016
rect 247736 126976 264980 127004
rect 247736 126964 247742 126976
rect 264974 126964 264980 126976
rect 265032 126964 265038 127016
rect 231762 126896 231768 126948
rect 231820 126936 231826 126948
rect 260098 126936 260104 126948
rect 231820 126908 260104 126936
rect 231820 126896 231826 126908
rect 260098 126896 260104 126908
rect 260156 126896 260162 126948
rect 282362 126896 282368 126948
rect 282420 126936 282426 126948
rect 287146 126936 287152 126948
rect 282420 126908 287152 126936
rect 282420 126896 282426 126908
rect 287146 126896 287152 126908
rect 287204 126896 287210 126948
rect 230842 126828 230848 126880
rect 230900 126868 230906 126880
rect 235258 126868 235264 126880
rect 230900 126840 235264 126868
rect 230900 126828 230906 126840
rect 235258 126828 235264 126840
rect 235316 126828 235322 126880
rect 282086 126216 282092 126268
rect 282144 126256 282150 126268
rect 306558 126256 306564 126268
rect 282144 126228 306564 126256
rect 282144 126216 282150 126228
rect 306558 126216 306564 126228
rect 306616 126216 306622 126268
rect 193858 125672 193864 125724
rect 193916 125712 193922 125724
rect 213914 125712 213920 125724
rect 193916 125684 213920 125712
rect 193916 125672 193922 125684
rect 213914 125672 213920 125684
rect 213972 125672 213978 125724
rect 182910 125604 182916 125656
rect 182968 125644 182974 125656
rect 214006 125644 214012 125656
rect 182968 125616 214012 125644
rect 182968 125604 182974 125616
rect 214006 125604 214012 125616
rect 214064 125604 214070 125656
rect 261570 125604 261576 125656
rect 261628 125644 261634 125656
rect 264974 125644 264980 125656
rect 261628 125616 264980 125644
rect 261628 125604 261634 125616
rect 264974 125604 264980 125616
rect 265032 125604 265038 125656
rect 231486 125536 231492 125588
rect 231544 125576 231550 125588
rect 253382 125576 253388 125588
rect 231544 125548 253388 125576
rect 231544 125536 231550 125548
rect 253382 125536 253388 125548
rect 253440 125536 253446 125588
rect 282822 125536 282828 125588
rect 282880 125576 282886 125588
rect 320266 125576 320272 125588
rect 282880 125548 320272 125576
rect 282880 125536 282886 125548
rect 320266 125536 320272 125548
rect 320324 125536 320330 125588
rect 231762 125468 231768 125520
rect 231820 125508 231826 125520
rect 240778 125508 240784 125520
rect 231820 125480 240784 125508
rect 231820 125468 231826 125480
rect 240778 125468 240784 125480
rect 240836 125468 240842 125520
rect 282730 125468 282736 125520
rect 282788 125508 282794 125520
rect 292574 125508 292580 125520
rect 282788 125480 292580 125508
rect 282788 125468 282794 125480
rect 292574 125468 292580 125480
rect 292632 125468 292638 125520
rect 177574 124856 177580 124908
rect 177632 124896 177638 124908
rect 214742 124896 214748 124908
rect 177632 124868 214748 124896
rect 177632 124856 177638 124868
rect 214742 124856 214748 124868
rect 214800 124856 214806 124908
rect 253474 124856 253480 124908
rect 253532 124896 253538 124908
rect 265618 124896 265624 124908
rect 253532 124868 265624 124896
rect 253532 124856 253538 124868
rect 265618 124856 265624 124868
rect 265676 124856 265682 124908
rect 167730 124176 167736 124228
rect 167788 124216 167794 124228
rect 213914 124216 213920 124228
rect 167788 124188 213920 124216
rect 167788 124176 167794 124188
rect 213914 124176 213920 124188
rect 213972 124176 213978 124228
rect 260190 124176 260196 124228
rect 260248 124216 260254 124228
rect 264974 124216 264980 124228
rect 260248 124188 264980 124216
rect 260248 124176 260254 124188
rect 264974 124176 264980 124188
rect 265032 124176 265038 124228
rect 231762 124108 231768 124160
rect 231820 124148 231826 124160
rect 260374 124148 260380 124160
rect 231820 124120 260380 124148
rect 231820 124108 231826 124120
rect 260374 124108 260380 124120
rect 260432 124108 260438 124160
rect 231670 124040 231676 124092
rect 231728 124080 231734 124092
rect 245010 124080 245016 124092
rect 231728 124052 245016 124080
rect 231728 124040 231734 124052
rect 245010 124040 245016 124052
rect 245068 124040 245074 124092
rect 282822 123632 282828 123684
rect 282880 123672 282886 123684
rect 288434 123672 288440 123684
rect 282880 123644 288440 123672
rect 282880 123632 282886 123644
rect 288434 123632 288440 123644
rect 288492 123632 288498 123684
rect 188522 123428 188528 123480
rect 188580 123468 188586 123480
rect 214006 123468 214012 123480
rect 188580 123440 214012 123468
rect 188580 123428 188586 123440
rect 214006 123428 214012 123440
rect 214064 123428 214070 123480
rect 282178 123428 282184 123480
rect 282236 123468 282242 123480
rect 314654 123468 314660 123480
rect 282236 123440 314660 123468
rect 282236 123428 282242 123440
rect 314654 123428 314660 123440
rect 314712 123428 314718 123480
rect 170490 122816 170496 122868
rect 170548 122856 170554 122868
rect 213914 122856 213920 122868
rect 170548 122828 213920 122856
rect 170548 122816 170554 122828
rect 213914 122816 213920 122828
rect 213972 122816 213978 122868
rect 250714 122816 250720 122868
rect 250772 122856 250778 122868
rect 264974 122856 264980 122868
rect 250772 122828 264980 122856
rect 250772 122816 250778 122828
rect 264974 122816 264980 122828
rect 265032 122816 265038 122868
rect 231762 122748 231768 122800
rect 231820 122788 231826 122800
rect 242250 122788 242256 122800
rect 231820 122760 242256 122788
rect 231820 122748 231826 122760
rect 242250 122748 242256 122760
rect 242308 122748 242314 122800
rect 282822 122748 282828 122800
rect 282880 122788 282886 122800
rect 298186 122788 298192 122800
rect 282880 122760 298192 122788
rect 282880 122748 282886 122760
rect 298186 122748 298192 122760
rect 298244 122748 298250 122800
rect 230750 122068 230756 122120
rect 230808 122108 230814 122120
rect 253198 122108 253204 122120
rect 230808 122080 253204 122108
rect 230808 122068 230814 122080
rect 253198 122068 253204 122080
rect 253256 122068 253262 122120
rect 282638 122068 282644 122120
rect 282696 122108 282702 122120
rect 303706 122108 303712 122120
rect 282696 122080 303712 122108
rect 282696 122068 282702 122080
rect 303706 122068 303712 122080
rect 303764 122068 303770 122120
rect 199470 121524 199476 121576
rect 199528 121564 199534 121576
rect 214006 121564 214012 121576
rect 199528 121536 214012 121564
rect 199528 121524 199534 121536
rect 214006 121524 214012 121536
rect 214064 121524 214070 121576
rect 260098 121524 260104 121576
rect 260156 121564 260162 121576
rect 265066 121564 265072 121576
rect 260156 121536 265072 121564
rect 260156 121524 260162 121536
rect 265066 121524 265072 121536
rect 265124 121524 265130 121576
rect 178678 121456 178684 121508
rect 178736 121496 178742 121508
rect 213914 121496 213920 121508
rect 178736 121468 213920 121496
rect 178736 121456 178742 121468
rect 213914 121456 213920 121468
rect 213972 121456 213978 121508
rect 255958 121456 255964 121508
rect 256016 121496 256022 121508
rect 264974 121496 264980 121508
rect 256016 121468 264980 121496
rect 256016 121456 256022 121468
rect 264974 121456 264980 121468
rect 265032 121456 265038 121508
rect 282822 121388 282828 121440
rect 282880 121428 282886 121440
rect 289906 121428 289912 121440
rect 282880 121400 289912 121428
rect 282880 121388 282886 121400
rect 289906 121388 289912 121400
rect 289964 121388 289970 121440
rect 230566 121184 230572 121236
rect 230624 121224 230630 121236
rect 234154 121224 234160 121236
rect 230624 121196 234160 121224
rect 230624 121184 230630 121196
rect 234154 121184 234160 121196
rect 234212 121184 234218 121236
rect 282086 120912 282092 120964
rect 282144 120952 282150 120964
rect 285674 120952 285680 120964
rect 282144 120924 285680 120952
rect 282144 120912 282150 120924
rect 285674 120912 285680 120924
rect 285732 120912 285738 120964
rect 231578 120708 231584 120760
rect 231636 120748 231642 120760
rect 252002 120748 252008 120760
rect 231636 120720 252008 120748
rect 231636 120708 231642 120720
rect 252002 120708 252008 120720
rect 252060 120708 252066 120760
rect 174722 120164 174728 120216
rect 174780 120204 174786 120216
rect 213914 120204 213920 120216
rect 174780 120176 213920 120204
rect 174780 120164 174786 120176
rect 213914 120164 213920 120176
rect 213972 120164 213978 120216
rect 261662 120164 261668 120216
rect 261720 120204 261726 120216
rect 265066 120204 265072 120216
rect 261720 120176 265072 120204
rect 261720 120164 261726 120176
rect 265066 120164 265072 120176
rect 265124 120164 265130 120216
rect 169202 120096 169208 120148
rect 169260 120136 169266 120148
rect 214006 120136 214012 120148
rect 169260 120108 214012 120136
rect 169260 120096 169266 120108
rect 214006 120096 214012 120108
rect 214064 120096 214070 120148
rect 238294 120096 238300 120148
rect 238352 120136 238358 120148
rect 264974 120136 264980 120148
rect 238352 120108 264980 120136
rect 238352 120096 238358 120108
rect 264974 120096 264980 120108
rect 265032 120096 265038 120148
rect 231486 120028 231492 120080
rect 231544 120068 231550 120080
rect 240870 120068 240876 120080
rect 231544 120040 240876 120068
rect 231544 120028 231550 120040
rect 240870 120028 240876 120040
rect 240928 120028 240934 120080
rect 282822 120028 282828 120080
rect 282880 120068 282886 120080
rect 298370 120068 298376 120080
rect 282880 120040 298376 120068
rect 282880 120028 282886 120040
rect 298370 120028 298376 120040
rect 298428 120028 298434 120080
rect 241146 119348 241152 119400
rect 241204 119388 241210 119400
rect 264606 119388 264612 119400
rect 241204 119360 264612 119388
rect 241204 119348 241210 119360
rect 264606 119348 264612 119360
rect 264664 119348 264670 119400
rect 284938 119348 284944 119400
rect 284996 119388 285002 119400
rect 304994 119388 305000 119400
rect 284996 119360 305000 119388
rect 284996 119348 285002 119360
rect 304994 119348 305000 119360
rect 305052 119348 305058 119400
rect 210418 118736 210424 118788
rect 210476 118776 210482 118788
rect 214006 118776 214012 118788
rect 210476 118748 214012 118776
rect 210476 118736 210482 118748
rect 214006 118736 214012 118748
rect 214064 118736 214070 118788
rect 205174 118668 205180 118720
rect 205232 118708 205238 118720
rect 213914 118708 213920 118720
rect 205232 118680 213920 118708
rect 205232 118668 205238 118680
rect 213914 118668 213920 118680
rect 213972 118668 213978 118720
rect 231486 118668 231492 118720
rect 231544 118708 231550 118720
rect 238386 118708 238392 118720
rect 231544 118680 238392 118708
rect 231544 118668 231550 118680
rect 238386 118668 238392 118680
rect 238444 118668 238450 118720
rect 247954 118668 247960 118720
rect 248012 118708 248018 118720
rect 264974 118708 264980 118720
rect 248012 118680 264980 118708
rect 248012 118668 248018 118680
rect 264974 118668 264980 118680
rect 265032 118668 265038 118720
rect 231394 118600 231400 118652
rect 231452 118640 231458 118652
rect 254578 118640 254584 118652
rect 231452 118612 254584 118640
rect 231452 118600 231458 118612
rect 254578 118600 254584 118612
rect 254636 118600 254642 118652
rect 282822 118600 282828 118652
rect 282880 118640 282886 118652
rect 293954 118640 293960 118652
rect 282880 118612 293960 118640
rect 282880 118600 282886 118612
rect 293954 118600 293960 118612
rect 294012 118600 294018 118652
rect 231762 118532 231768 118584
rect 231820 118572 231826 118584
rect 240962 118572 240968 118584
rect 231820 118544 240968 118572
rect 231820 118532 231826 118544
rect 240962 118532 240968 118544
rect 241020 118532 241026 118584
rect 282822 117920 282828 117972
rect 282880 117960 282886 117972
rect 288618 117960 288624 117972
rect 282880 117932 288624 117960
rect 282880 117920 282886 117932
rect 288618 117920 288624 117932
rect 288676 117920 288682 117972
rect 184474 117376 184480 117428
rect 184532 117416 184538 117428
rect 214006 117416 214012 117428
rect 184532 117388 214012 117416
rect 184532 117376 184538 117388
rect 214006 117376 214012 117388
rect 214064 117376 214070 117428
rect 170582 117308 170588 117360
rect 170640 117348 170646 117360
rect 213914 117348 213920 117360
rect 170640 117320 213920 117348
rect 170640 117308 170646 117320
rect 213914 117308 213920 117320
rect 213972 117308 213978 117360
rect 252002 117308 252008 117360
rect 252060 117348 252066 117360
rect 264974 117348 264980 117360
rect 252060 117320 264980 117348
rect 252060 117308 252066 117320
rect 264974 117308 264980 117320
rect 265032 117308 265038 117360
rect 230934 117240 230940 117292
rect 230992 117280 230998 117292
rect 236914 117280 236920 117292
rect 230992 117252 236920 117280
rect 230992 117240 230998 117252
rect 236914 117240 236920 117252
rect 236972 117240 236978 117292
rect 290642 117240 290648 117292
rect 290700 117280 290706 117292
rect 360194 117280 360200 117292
rect 290700 117252 360200 117280
rect 290700 117240 290706 117252
rect 360194 117240 360200 117252
rect 360252 117240 360258 117292
rect 230750 116696 230756 116748
rect 230808 116736 230814 116748
rect 235534 116736 235540 116748
rect 230808 116708 235540 116736
rect 230808 116696 230814 116708
rect 235534 116696 235540 116708
rect 235592 116696 235598 116748
rect 177390 116560 177396 116612
rect 177448 116600 177454 116612
rect 195514 116600 195520 116612
rect 177448 116572 195520 116600
rect 177448 116560 177454 116572
rect 195514 116560 195520 116572
rect 195572 116560 195578 116612
rect 282822 116560 282828 116612
rect 282880 116600 282886 116612
rect 290642 116600 290648 116612
rect 282880 116572 290648 116600
rect 282880 116560 282886 116572
rect 290642 116560 290648 116572
rect 290700 116560 290706 116612
rect 195422 116016 195428 116068
rect 195480 116056 195486 116068
rect 213914 116056 213920 116068
rect 195480 116028 213920 116056
rect 195480 116016 195486 116028
rect 213914 116016 213920 116028
rect 213972 116016 213978 116068
rect 254578 116016 254584 116068
rect 254636 116056 254642 116068
rect 265066 116056 265072 116068
rect 254636 116028 265072 116056
rect 254636 116016 254642 116028
rect 265066 116016 265072 116028
rect 265124 116016 265130 116068
rect 187050 115948 187056 116000
rect 187108 115988 187114 116000
rect 214006 115988 214012 116000
rect 187108 115960 214012 115988
rect 187108 115948 187114 115960
rect 214006 115948 214012 115960
rect 214064 115948 214070 116000
rect 236730 115948 236736 116000
rect 236788 115988 236794 116000
rect 264974 115988 264980 116000
rect 236788 115960 264980 115988
rect 236788 115948 236794 115960
rect 264974 115948 264980 115960
rect 265032 115948 265038 116000
rect 231762 115880 231768 115932
rect 231820 115920 231826 115932
rect 251910 115920 251916 115932
rect 231820 115892 251916 115920
rect 231820 115880 231826 115892
rect 251910 115880 251916 115892
rect 251968 115880 251974 115932
rect 282822 115880 282828 115932
rect 282880 115920 282886 115932
rect 301038 115920 301044 115932
rect 282880 115892 301044 115920
rect 282880 115880 282886 115892
rect 301038 115880 301044 115892
rect 301096 115920 301102 115932
rect 382274 115920 382280 115932
rect 301096 115892 382280 115920
rect 301096 115880 301102 115892
rect 382274 115880 382280 115892
rect 382332 115880 382338 115932
rect 231026 115812 231032 115864
rect 231084 115852 231090 115864
rect 238110 115852 238116 115864
rect 231084 115824 238116 115852
rect 231084 115812 231090 115824
rect 238110 115812 238116 115824
rect 238168 115812 238174 115864
rect 187234 114588 187240 114640
rect 187292 114628 187298 114640
rect 213914 114628 213920 114640
rect 187292 114600 213920 114628
rect 187292 114588 187298 114600
rect 213914 114588 213920 114600
rect 213972 114588 213978 114640
rect 257430 114588 257436 114640
rect 257488 114628 257494 114640
rect 265066 114628 265072 114640
rect 257488 114600 265072 114628
rect 257488 114588 257494 114600
rect 265066 114588 265072 114600
rect 265124 114588 265130 114640
rect 171870 114520 171876 114572
rect 171928 114560 171934 114572
rect 214006 114560 214012 114572
rect 171928 114532 214012 114560
rect 171928 114520 171934 114532
rect 214006 114520 214012 114532
rect 214064 114520 214070 114572
rect 242250 114520 242256 114572
rect 242308 114560 242314 114572
rect 264974 114560 264980 114572
rect 242308 114532 264980 114560
rect 242308 114520 242314 114532
rect 264974 114520 264980 114532
rect 265032 114520 265038 114572
rect 230566 114452 230572 114504
rect 230624 114492 230630 114504
rect 250530 114492 250536 114504
rect 230624 114464 250536 114492
rect 230624 114452 230630 114464
rect 250530 114452 250536 114464
rect 250588 114452 250594 114504
rect 231578 114316 231584 114368
rect 231636 114356 231642 114368
rect 233970 114356 233976 114368
rect 231636 114328 233976 114356
rect 231636 114316 231642 114328
rect 233970 114316 233976 114328
rect 234028 114316 234034 114368
rect 282822 114112 282828 114164
rect 282880 114152 282886 114164
rect 287238 114152 287244 114164
rect 282880 114124 287244 114152
rect 282880 114112 282886 114124
rect 287238 114112 287244 114124
rect 287296 114112 287302 114164
rect 173434 113772 173440 113824
rect 173492 113812 173498 113824
rect 214098 113812 214104 113824
rect 173492 113784 214104 113812
rect 173492 113772 173498 113784
rect 214098 113772 214104 113784
rect 214156 113772 214162 113824
rect 281718 113772 281724 113824
rect 281776 113812 281782 113824
rect 299566 113812 299572 113824
rect 281776 113784 299572 113812
rect 281776 113772 281782 113784
rect 299566 113772 299572 113784
rect 299624 113772 299630 113824
rect 257614 113228 257620 113280
rect 257672 113268 257678 113280
rect 265066 113268 265072 113280
rect 257672 113240 265072 113268
rect 257672 113228 257678 113240
rect 265066 113228 265072 113240
rect 265124 113228 265130 113280
rect 193950 113160 193956 113212
rect 194008 113200 194014 113212
rect 213914 113200 213920 113212
rect 194008 113172 213920 113200
rect 194008 113160 194014 113172
rect 213914 113160 213920 113172
rect 213972 113160 213978 113212
rect 250438 113160 250444 113212
rect 250496 113200 250502 113212
rect 264974 113200 264980 113212
rect 250496 113172 264980 113200
rect 250496 113160 250502 113172
rect 264974 113160 264980 113172
rect 265032 113160 265038 113212
rect 231762 113092 231768 113144
rect 231820 113132 231826 113144
rect 250806 113132 250812 113144
rect 231820 113104 250812 113132
rect 231820 113092 231826 113104
rect 250806 113092 250812 113104
rect 250864 113092 250870 113144
rect 282822 113092 282828 113144
rect 282880 113132 282886 113144
rect 317506 113132 317512 113144
rect 282880 113104 317512 113132
rect 282880 113092 282886 113104
rect 317506 113092 317512 113104
rect 317564 113132 317570 113144
rect 368474 113132 368480 113144
rect 317564 113104 368480 113132
rect 317564 113092 317570 113104
rect 368474 113092 368480 113104
rect 368532 113092 368538 113144
rect 231670 113024 231676 113076
rect 231728 113064 231734 113076
rect 243722 113064 243728 113076
rect 231728 113036 243728 113064
rect 231728 113024 231734 113036
rect 243722 113024 243728 113036
rect 243780 113024 243786 113076
rect 169018 112412 169024 112464
rect 169076 112452 169082 112464
rect 211798 112452 211804 112464
rect 169076 112424 211804 112452
rect 169076 112412 169082 112424
rect 211798 112412 211804 112424
rect 211856 112412 211862 112464
rect 211890 111868 211896 111920
rect 211948 111908 211954 111920
rect 214006 111908 214012 111920
rect 211948 111880 214012 111908
rect 211948 111868 211954 111880
rect 214006 111868 214012 111880
rect 214064 111868 214070 111920
rect 260374 111868 260380 111920
rect 260432 111908 260438 111920
rect 265894 111908 265900 111920
rect 260432 111880 265900 111908
rect 260432 111868 260438 111880
rect 265894 111868 265900 111880
rect 265952 111868 265958 111920
rect 172146 111800 172152 111852
rect 172204 111840 172210 111852
rect 213914 111840 213920 111852
rect 172204 111812 213920 111840
rect 172204 111800 172210 111812
rect 213914 111800 213920 111812
rect 213972 111800 213978 111852
rect 247862 111800 247868 111852
rect 247920 111840 247926 111852
rect 264974 111840 264980 111852
rect 247920 111812 264980 111840
rect 247920 111800 247926 111812
rect 264974 111800 264980 111812
rect 265032 111800 265038 111852
rect 3142 111732 3148 111784
rect 3200 111772 3206 111784
rect 35158 111772 35164 111784
rect 3200 111744 35164 111772
rect 3200 111732 3206 111744
rect 35158 111732 35164 111744
rect 35216 111732 35222 111784
rect 167822 111732 167828 111784
rect 167880 111772 167886 111784
rect 187142 111772 187148 111784
rect 167880 111744 187148 111772
rect 167880 111732 167886 111744
rect 187142 111732 187148 111744
rect 187200 111732 187206 111784
rect 282822 111732 282828 111784
rect 282880 111772 282886 111784
rect 295426 111772 295432 111784
rect 282880 111744 295432 111772
rect 282880 111732 282886 111744
rect 295426 111732 295432 111744
rect 295484 111732 295490 111784
rect 282086 111596 282092 111648
rect 282144 111636 282150 111648
rect 284938 111636 284944 111648
rect 282144 111608 284944 111636
rect 282144 111596 282150 111608
rect 284938 111596 284944 111608
rect 284996 111596 285002 111648
rect 230934 111052 230940 111104
rect 230992 111092 230998 111104
rect 256050 111092 256056 111104
rect 230992 111064 256056 111092
rect 230992 111052 230998 111064
rect 256050 111052 256056 111064
rect 256108 111052 256114 111104
rect 230566 110848 230572 110900
rect 230624 110888 230630 110900
rect 232866 110888 232872 110900
rect 230624 110860 232872 110888
rect 230624 110848 230630 110860
rect 232866 110848 232872 110860
rect 232924 110848 232930 110900
rect 196802 110508 196808 110560
rect 196860 110548 196866 110560
rect 213914 110548 213920 110560
rect 196860 110520 213920 110548
rect 196860 110508 196866 110520
rect 213914 110508 213920 110520
rect 213972 110508 213978 110560
rect 176194 110440 176200 110492
rect 176252 110480 176258 110492
rect 214006 110480 214012 110492
rect 176252 110452 214012 110480
rect 176252 110440 176258 110452
rect 214006 110440 214012 110452
rect 214064 110440 214070 110492
rect 245010 110440 245016 110492
rect 245068 110480 245074 110492
rect 264974 110480 264980 110492
rect 245068 110452 264980 110480
rect 245068 110440 245074 110452
rect 264974 110440 264980 110452
rect 265032 110440 265038 110492
rect 168190 110372 168196 110424
rect 168248 110412 168254 110424
rect 169110 110412 169116 110424
rect 168248 110384 169116 110412
rect 168248 110372 168254 110384
rect 169110 110372 169116 110384
rect 169168 110372 169174 110424
rect 231762 110372 231768 110424
rect 231820 110412 231826 110424
rect 247770 110412 247776 110424
rect 231820 110384 247776 110412
rect 231820 110372 231826 110384
rect 247770 110372 247776 110384
rect 247828 110372 247834 110424
rect 282638 110372 282644 110424
rect 282696 110412 282702 110424
rect 295334 110412 295340 110424
rect 282696 110384 295340 110412
rect 282696 110372 282702 110384
rect 295334 110372 295340 110384
rect 295392 110372 295398 110424
rect 230750 109964 230756 110016
rect 230808 110004 230814 110016
rect 235442 110004 235448 110016
rect 230808 109976 235448 110004
rect 230808 109964 230814 109976
rect 235442 109964 235448 109976
rect 235500 109964 235506 110016
rect 199378 109080 199384 109132
rect 199436 109120 199442 109132
rect 214006 109120 214012 109132
rect 199436 109092 214012 109120
rect 199436 109080 199442 109092
rect 214006 109080 214012 109092
rect 214064 109080 214070 109132
rect 170674 109012 170680 109064
rect 170732 109052 170738 109064
rect 213914 109052 213920 109064
rect 170732 109024 213920 109052
rect 170732 109012 170738 109024
rect 213914 109012 213920 109024
rect 213972 109012 213978 109064
rect 235534 109012 235540 109064
rect 235592 109052 235598 109064
rect 265066 109052 265072 109064
rect 235592 109024 265072 109052
rect 235592 109012 235598 109024
rect 265066 109012 265072 109024
rect 265124 109012 265130 109064
rect 231762 108944 231768 108996
rect 231820 108984 231826 108996
rect 257522 108984 257528 108996
rect 231820 108956 257528 108984
rect 231820 108944 231826 108956
rect 257522 108944 257528 108956
rect 257580 108944 257586 108996
rect 281718 108944 281724 108996
rect 281776 108984 281782 108996
rect 328454 108984 328460 108996
rect 281776 108956 328460 108984
rect 281776 108944 281782 108956
rect 328454 108944 328460 108956
rect 328512 108944 328518 108996
rect 231486 108876 231492 108928
rect 231544 108916 231550 108928
rect 244918 108916 244924 108928
rect 231544 108888 244924 108916
rect 231544 108876 231550 108888
rect 244918 108876 244924 108888
rect 244976 108876 244982 108928
rect 282822 108876 282828 108928
rect 282880 108916 282886 108928
rect 309134 108916 309140 108928
rect 282880 108888 309140 108916
rect 282880 108876 282886 108888
rect 309134 108876 309140 108888
rect 309192 108876 309198 108928
rect 167914 107720 167920 107772
rect 167972 107760 167978 107772
rect 213914 107760 213920 107772
rect 167972 107732 213920 107760
rect 167972 107720 167978 107732
rect 213914 107720 213920 107732
rect 213972 107720 213978 107772
rect 262950 107720 262956 107772
rect 263008 107760 263014 107772
rect 265342 107760 265348 107772
rect 263008 107732 265348 107760
rect 263008 107720 263014 107732
rect 265342 107720 265348 107732
rect 265400 107720 265406 107772
rect 166350 107652 166356 107704
rect 166408 107692 166414 107704
rect 214006 107692 214012 107704
rect 166408 107664 214012 107692
rect 166408 107652 166414 107664
rect 214006 107652 214012 107664
rect 214064 107652 214070 107704
rect 256142 107652 256148 107704
rect 256200 107692 256206 107704
rect 264974 107692 264980 107704
rect 256200 107664 264980 107692
rect 256200 107652 256206 107664
rect 264974 107652 264980 107664
rect 265032 107652 265038 107704
rect 231762 107584 231768 107636
rect 231820 107624 231826 107636
rect 265710 107624 265716 107636
rect 231820 107596 265716 107624
rect 231820 107584 231826 107596
rect 265710 107584 265716 107596
rect 265768 107584 265774 107636
rect 231486 107516 231492 107568
rect 231544 107556 231550 107568
rect 249426 107556 249432 107568
rect 231544 107528 249432 107556
rect 231544 107516 231550 107528
rect 249426 107516 249432 107528
rect 249484 107516 249490 107568
rect 282822 106904 282828 106956
rect 282880 106944 282886 106956
rect 287054 106944 287060 106956
rect 282880 106916 287060 106944
rect 282880 106904 282886 106916
rect 287054 106904 287060 106916
rect 287112 106904 287118 106956
rect 202322 106360 202328 106412
rect 202380 106400 202386 106412
rect 214006 106400 214012 106412
rect 202380 106372 214012 106400
rect 202380 106360 202386 106372
rect 214006 106360 214012 106372
rect 214064 106360 214070 106412
rect 167822 106292 167828 106344
rect 167880 106332 167886 106344
rect 213914 106332 213920 106344
rect 167880 106304 213920 106332
rect 167880 106292 167886 106304
rect 213914 106292 213920 106304
rect 213972 106292 213978 106344
rect 249242 106292 249248 106344
rect 249300 106332 249306 106344
rect 264974 106332 264980 106344
rect 249300 106304 264980 106332
rect 249300 106292 249306 106304
rect 264974 106292 264980 106304
rect 265032 106292 265038 106344
rect 282822 106224 282828 106276
rect 282880 106264 282886 106276
rect 291194 106264 291200 106276
rect 282880 106236 291200 106264
rect 282880 106224 282886 106236
rect 291194 106224 291200 106236
rect 291252 106224 291258 106276
rect 231762 106020 231768 106072
rect 231820 106060 231826 106072
rect 238202 106060 238208 106072
rect 231820 106032 238208 106060
rect 231820 106020 231826 106032
rect 238202 106020 238208 106032
rect 238260 106020 238266 106072
rect 245194 105612 245200 105664
rect 245252 105652 245258 105664
rect 262122 105652 262128 105664
rect 245252 105624 262128 105652
rect 245252 105612 245258 105624
rect 262122 105612 262128 105624
rect 262180 105612 262186 105664
rect 230750 105544 230756 105596
rect 230808 105584 230814 105596
rect 264422 105584 264428 105596
rect 230808 105556 264428 105584
rect 230808 105544 230814 105556
rect 264422 105544 264428 105556
rect 264480 105544 264486 105596
rect 282822 105272 282828 105324
rect 282880 105312 282886 105324
rect 288526 105312 288532 105324
rect 282880 105284 288532 105312
rect 282880 105272 282886 105284
rect 288526 105272 288532 105284
rect 288584 105272 288590 105324
rect 191282 104932 191288 104984
rect 191340 104972 191346 104984
rect 214006 104972 214012 104984
rect 191340 104944 214012 104972
rect 191340 104932 191346 104944
rect 214006 104932 214012 104944
rect 214064 104932 214070 104984
rect 169110 104864 169116 104916
rect 169168 104904 169174 104916
rect 213914 104904 213920 104916
rect 169168 104876 213920 104904
rect 169168 104864 169174 104876
rect 213914 104864 213920 104876
rect 213972 104864 213978 104916
rect 263134 104864 263140 104916
rect 263192 104904 263198 104916
rect 264974 104904 264980 104916
rect 263192 104876 264980 104904
rect 263192 104864 263198 104876
rect 264974 104864 264980 104876
rect 265032 104864 265038 104916
rect 230934 104796 230940 104848
rect 230992 104836 230998 104848
rect 236822 104836 236828 104848
rect 230992 104808 236828 104836
rect 230992 104796 230998 104808
rect 236822 104796 236828 104808
rect 236880 104796 236886 104848
rect 282822 104796 282828 104848
rect 282880 104836 282886 104848
rect 291378 104836 291384 104848
rect 282880 104808 291384 104836
rect 282880 104796 282886 104808
rect 291378 104796 291384 104808
rect 291436 104796 291442 104848
rect 281534 104728 281540 104780
rect 281592 104768 281598 104780
rect 284386 104768 284392 104780
rect 281592 104740 284392 104768
rect 281592 104728 281598 104740
rect 284386 104728 284392 104740
rect 284444 104728 284450 104780
rect 250622 104184 250628 104236
rect 250680 104224 250686 104236
rect 263042 104224 263048 104236
rect 250680 104196 263048 104224
rect 250680 104184 250686 104196
rect 263042 104184 263048 104196
rect 263100 104184 263106 104236
rect 164878 104116 164884 104168
rect 164936 104156 164942 104168
rect 177482 104156 177488 104168
rect 164936 104128 177488 104156
rect 164936 104116 164942 104128
rect 177482 104116 177488 104128
rect 177540 104116 177546 104168
rect 230566 104116 230572 104168
rect 230624 104156 230630 104168
rect 252094 104156 252100 104168
rect 230624 104128 252100 104156
rect 230624 104116 230630 104128
rect 252094 104116 252100 104128
rect 252152 104116 252158 104168
rect 261754 103912 261760 103964
rect 261812 103952 261818 103964
rect 264974 103952 264980 103964
rect 261812 103924 264980 103952
rect 261812 103912 261818 103924
rect 264974 103912 264980 103924
rect 265032 103912 265038 103964
rect 178862 103504 178868 103556
rect 178920 103544 178926 103556
rect 213914 103544 213920 103556
rect 178920 103516 213920 103544
rect 178920 103504 178926 103516
rect 213914 103504 213920 103516
rect 213972 103504 213978 103556
rect 231762 103436 231768 103488
rect 231820 103476 231826 103488
rect 246574 103476 246580 103488
rect 231820 103448 246580 103476
rect 231820 103436 231826 103448
rect 246574 103436 246580 103448
rect 246632 103436 246638 103488
rect 282086 103436 282092 103488
rect 282144 103476 282150 103488
rect 291286 103476 291292 103488
rect 282144 103448 291292 103476
rect 282144 103436 282150 103448
rect 291286 103436 291292 103448
rect 291344 103436 291350 103488
rect 231486 103368 231492 103420
rect 231544 103408 231550 103420
rect 241146 103408 241152 103420
rect 231544 103380 241152 103408
rect 231544 103368 231550 103380
rect 241146 103368 241152 103380
rect 241204 103368 241210 103420
rect 181622 102756 181628 102808
rect 181680 102796 181686 102808
rect 209038 102796 209044 102808
rect 181680 102768 209044 102796
rect 181680 102756 181686 102768
rect 209038 102756 209044 102768
rect 209096 102756 209102 102808
rect 212442 102212 212448 102264
rect 212500 102252 212506 102264
rect 214006 102252 214012 102264
rect 212500 102224 214012 102252
rect 212500 102212 212506 102224
rect 214006 102212 214012 102224
rect 214064 102212 214070 102264
rect 258902 102212 258908 102264
rect 258960 102252 258966 102264
rect 265066 102252 265072 102264
rect 258960 102224 265072 102252
rect 258960 102212 258966 102224
rect 265066 102212 265072 102224
rect 265124 102212 265130 102264
rect 185578 102144 185584 102196
rect 185636 102184 185642 102196
rect 213914 102184 213920 102196
rect 185636 102156 213920 102184
rect 185636 102144 185642 102156
rect 213914 102144 213920 102156
rect 213972 102144 213978 102196
rect 240870 102144 240876 102196
rect 240928 102184 240934 102196
rect 264974 102184 264980 102196
rect 240928 102156 264980 102184
rect 240928 102144 240934 102156
rect 264974 102144 264980 102156
rect 265032 102144 265038 102196
rect 231670 102076 231676 102128
rect 231728 102116 231734 102128
rect 258810 102116 258816 102128
rect 231728 102088 258816 102116
rect 231728 102076 231734 102088
rect 258810 102076 258816 102088
rect 258868 102076 258874 102128
rect 282270 102076 282276 102128
rect 282328 102116 282334 102128
rect 296806 102116 296812 102128
rect 282328 102088 296812 102116
rect 282328 102076 282334 102088
rect 296806 102076 296812 102088
rect 296864 102076 296870 102128
rect 230658 102008 230664 102060
rect 230716 102048 230722 102060
rect 242342 102048 242348 102060
rect 230716 102020 242348 102048
rect 230716 102008 230722 102020
rect 242342 102008 242348 102020
rect 242400 102008 242406 102060
rect 196710 101396 196716 101448
rect 196768 101436 196774 101448
rect 217226 101436 217232 101448
rect 196768 101408 217232 101436
rect 196768 101396 196774 101408
rect 217226 101396 217232 101408
rect 217284 101396 217290 101448
rect 258718 100784 258724 100836
rect 258776 100824 258782 100836
rect 264974 100824 264980 100836
rect 258776 100796 264980 100824
rect 258776 100784 258782 100796
rect 264974 100784 264980 100796
rect 265032 100784 265038 100836
rect 177482 100716 177488 100768
rect 177540 100756 177546 100768
rect 213914 100756 213920 100768
rect 177540 100728 213920 100756
rect 177540 100716 177546 100728
rect 213914 100716 213920 100728
rect 213972 100716 213978 100768
rect 263042 100716 263048 100768
rect 263100 100756 263106 100768
rect 265066 100756 265072 100768
rect 263100 100728 265072 100756
rect 263100 100716 263106 100728
rect 265066 100716 265072 100728
rect 265124 100716 265130 100768
rect 230658 100648 230664 100700
rect 230716 100688 230722 100700
rect 254762 100688 254768 100700
rect 230716 100660 254768 100688
rect 230716 100648 230722 100660
rect 254762 100648 254768 100660
rect 254820 100648 254826 100700
rect 231762 100580 231768 100632
rect 231820 100620 231826 100632
rect 253474 100620 253480 100632
rect 231820 100592 253480 100620
rect 231820 100580 231826 100592
rect 253474 100580 253480 100592
rect 253532 100580 253538 100632
rect 169294 99968 169300 100020
rect 169352 100008 169358 100020
rect 202138 100008 202144 100020
rect 169352 99980 202144 100008
rect 169352 99968 169358 99980
rect 202138 99968 202144 99980
rect 202196 99968 202202 100020
rect 205082 99968 205088 100020
rect 205140 100008 205146 100020
rect 214834 100008 214840 100020
rect 205140 99980 214840 100008
rect 205140 99968 205146 99980
rect 214834 99968 214840 99980
rect 214892 99968 214898 100020
rect 281994 99968 282000 100020
rect 282052 100008 282058 100020
rect 310606 100008 310612 100020
rect 282052 99980 310612 100008
rect 282052 99968 282058 99980
rect 310606 99968 310612 99980
rect 310664 99968 310670 100020
rect 166442 99356 166448 99408
rect 166500 99396 166506 99408
rect 213914 99396 213920 99408
rect 166500 99368 213920 99396
rect 166500 99356 166506 99368
rect 213914 99356 213920 99368
rect 213972 99356 213978 99408
rect 264422 99356 264428 99408
rect 264480 99396 264486 99408
rect 265986 99396 265992 99408
rect 264480 99368 265992 99396
rect 264480 99356 264486 99368
rect 265986 99356 265992 99368
rect 266044 99356 266050 99408
rect 281626 99288 281632 99340
rect 281684 99328 281690 99340
rect 283558 99328 283564 99340
rect 281684 99300 283564 99328
rect 281684 99288 281690 99300
rect 283558 99288 283564 99300
rect 283616 99288 283622 99340
rect 173342 98608 173348 98660
rect 173400 98648 173406 98660
rect 214098 98648 214104 98660
rect 173400 98620 214104 98648
rect 173400 98608 173406 98620
rect 214098 98608 214104 98620
rect 214156 98608 214162 98660
rect 242342 98064 242348 98116
rect 242400 98104 242406 98116
rect 265066 98104 265072 98116
rect 242400 98076 265072 98104
rect 242400 98064 242406 98076
rect 265066 98064 265072 98076
rect 265124 98064 265130 98116
rect 166534 97996 166540 98048
rect 166592 98036 166598 98048
rect 213914 98036 213920 98048
rect 166592 98008 213920 98036
rect 166592 97996 166598 98008
rect 213914 97996 213920 98008
rect 213972 97996 213978 98048
rect 231210 97996 231216 98048
rect 231268 98036 231274 98048
rect 264974 98036 264980 98048
rect 231268 98008 264980 98036
rect 231268 97996 231274 98008
rect 264974 97996 264980 98008
rect 265032 97996 265038 98048
rect 3510 97928 3516 97980
rect 3568 97968 3574 97980
rect 33778 97968 33784 97980
rect 3568 97940 33784 97968
rect 3568 97928 3574 97940
rect 33778 97928 33784 97940
rect 33836 97928 33842 97980
rect 204898 97928 204904 97980
rect 204956 97968 204962 97980
rect 229094 97968 229100 97980
rect 204956 97940 229100 97968
rect 204956 97928 204962 97940
rect 229094 97928 229100 97940
rect 229152 97928 229158 97980
rect 229186 97316 229192 97368
rect 229244 97356 229250 97368
rect 264974 97356 264980 97368
rect 229244 97328 264980 97356
rect 229244 97316 229250 97328
rect 264974 97316 264980 97328
rect 265032 97316 265038 97368
rect 265066 97288 265072 97300
rect 219406 97260 265072 97288
rect 165522 96636 165528 96688
rect 165580 96676 165586 96688
rect 213914 96676 213920 96688
rect 165580 96648 213920 96676
rect 165580 96636 165586 96648
rect 213914 96636 213920 96648
rect 213972 96636 213978 96688
rect 219406 96076 219434 97260
rect 265066 97248 265072 97260
rect 265124 97248 265130 97300
rect 282178 97248 282184 97300
rect 282236 97288 282242 97300
rect 310514 97288 310520 97300
rect 282236 97260 310520 97288
rect 282236 97248 282242 97260
rect 310514 97248 310520 97260
rect 310572 97248 310578 97300
rect 219342 96024 219348 96076
rect 219400 96036 219434 96076
rect 219400 96024 219406 96036
rect 165430 95888 165436 95940
rect 165488 95928 165494 95940
rect 216030 95928 216036 95940
rect 165488 95900 216036 95928
rect 165488 95888 165494 95900
rect 216030 95888 216036 95900
rect 216088 95888 216094 95940
rect 255866 95888 255872 95940
rect 255924 95928 255930 95940
rect 267826 95928 267832 95940
rect 255924 95900 267832 95928
rect 255924 95888 255930 95900
rect 267826 95888 267832 95900
rect 267884 95888 267890 95940
rect 230474 95276 230480 95328
rect 230532 95316 230538 95328
rect 232590 95316 232596 95328
rect 230532 95288 232596 95316
rect 230532 95276 230538 95288
rect 232590 95276 232596 95288
rect 232648 95276 232654 95328
rect 206370 95208 206376 95260
rect 206428 95248 206434 95260
rect 213914 95248 213920 95260
rect 206428 95220 213920 95248
rect 206428 95208 206434 95220
rect 213914 95208 213920 95220
rect 213972 95208 213978 95260
rect 225690 95208 225696 95260
rect 225748 95248 225754 95260
rect 264974 95248 264980 95260
rect 225748 95220 264980 95248
rect 225748 95208 225754 95220
rect 264974 95208 264980 95220
rect 265032 95208 265038 95260
rect 267642 95208 267648 95260
rect 267700 95248 267706 95260
rect 269206 95248 269212 95260
rect 267700 95220 269212 95248
rect 267700 95208 267706 95220
rect 269206 95208 269212 95220
rect 269264 95208 269270 95260
rect 259362 95140 259368 95192
rect 259420 95180 259426 95192
rect 279326 95180 279332 95192
rect 259420 95152 279332 95180
rect 259420 95140 259426 95152
rect 279326 95140 279332 95152
rect 279384 95140 279390 95192
rect 176102 94528 176108 94580
rect 176160 94568 176166 94580
rect 214558 94568 214564 94580
rect 176160 94540 214564 94568
rect 176160 94528 176166 94540
rect 214558 94528 214564 94540
rect 214616 94528 214622 94580
rect 209038 94460 209044 94512
rect 209096 94500 209102 94512
rect 260374 94500 260380 94512
rect 209096 94472 260380 94500
rect 209096 94460 209102 94472
rect 260374 94460 260380 94472
rect 260432 94460 260438 94512
rect 117130 93916 117136 93968
rect 117188 93956 117194 93968
rect 169202 93956 169208 93968
rect 117188 93928 169208 93956
rect 117188 93916 117194 93928
rect 169202 93916 169208 93928
rect 169260 93916 169266 93968
rect 107746 93848 107752 93900
rect 107804 93888 107810 93900
rect 195422 93888 195428 93900
rect 107804 93860 195428 93888
rect 107804 93848 107810 93860
rect 195422 93848 195428 93860
rect 195480 93848 195486 93900
rect 224218 93848 224224 93900
rect 224276 93888 224282 93900
rect 230014 93888 230020 93900
rect 224276 93860 230020 93888
rect 224276 93848 224282 93860
rect 230014 93848 230020 93860
rect 230072 93848 230078 93900
rect 264882 93848 264888 93900
rect 264940 93888 264946 93900
rect 267918 93888 267924 93900
rect 264940 93860 267924 93888
rect 264940 93848 264946 93860
rect 267918 93848 267924 93860
rect 267976 93848 267982 93900
rect 267826 93780 267832 93832
rect 267884 93820 267890 93832
rect 273990 93820 273996 93832
rect 267884 93792 273996 93820
rect 267884 93780 267890 93792
rect 273990 93780 273996 93792
rect 274048 93780 274054 93832
rect 115842 93168 115848 93220
rect 115900 93208 115906 93220
rect 174722 93208 174728 93220
rect 115900 93180 174728 93208
rect 115900 93168 115906 93180
rect 174722 93168 174728 93180
rect 174780 93168 174786 93220
rect 216030 93168 216036 93220
rect 216088 93208 216094 93220
rect 234154 93208 234160 93220
rect 216088 93180 234160 93208
rect 216088 93168 216094 93180
rect 234154 93168 234160 93180
rect 234212 93168 234218 93220
rect 60642 93100 60648 93152
rect 60700 93140 60706 93152
rect 90358 93140 90364 93152
rect 60700 93112 90364 93140
rect 60700 93100 60706 93112
rect 90358 93100 90364 93112
rect 90416 93100 90422 93152
rect 95050 93100 95056 93152
rect 95108 93140 95114 93152
rect 166350 93140 166356 93152
rect 95108 93112 166356 93140
rect 95108 93100 95114 93112
rect 166350 93100 166356 93112
rect 166408 93100 166414 93152
rect 211798 93100 211804 93152
rect 211856 93140 211862 93152
rect 243814 93140 243820 93152
rect 211856 93112 243820 93140
rect 211856 93100 211862 93112
rect 243814 93100 243820 93112
rect 243872 93100 243878 93152
rect 276750 93100 276756 93152
rect 276808 93140 276814 93152
rect 305638 93140 305644 93152
rect 276808 93112 305644 93140
rect 276808 93100 276814 93112
rect 305638 93100 305644 93112
rect 305696 93100 305702 93152
rect 86770 92488 86776 92540
rect 86828 92528 86834 92540
rect 115290 92528 115296 92540
rect 86828 92500 115296 92528
rect 86828 92488 86834 92500
rect 115290 92488 115296 92500
rect 115348 92488 115354 92540
rect 136082 92420 136088 92472
rect 136140 92460 136146 92472
rect 173250 92460 173256 92472
rect 136140 92432 173256 92460
rect 136140 92420 136146 92432
rect 173250 92420 173256 92432
rect 173308 92420 173314 92472
rect 217318 91808 217324 91860
rect 217376 91848 217382 91860
rect 245194 91848 245200 91860
rect 217376 91820 245200 91848
rect 217376 91808 217382 91820
rect 245194 91808 245200 91820
rect 245252 91808 245258 91860
rect 62022 91740 62028 91792
rect 62080 91780 62086 91792
rect 88978 91780 88984 91792
rect 62080 91752 88984 91780
rect 62080 91740 62086 91752
rect 88978 91740 88984 91752
rect 89036 91740 89042 91792
rect 160738 91740 160744 91792
rect 160796 91780 160802 91792
rect 171778 91780 171784 91792
rect 160796 91752 171784 91780
rect 160796 91740 160802 91752
rect 171778 91740 171784 91752
rect 171836 91740 171842 91792
rect 202138 91740 202144 91792
rect 202196 91780 202202 91792
rect 231302 91780 231308 91792
rect 202196 91752 231308 91780
rect 202196 91740 202202 91752
rect 231302 91740 231308 91752
rect 231360 91740 231366 91792
rect 102042 91128 102048 91180
rect 102100 91168 102106 91180
rect 115198 91168 115204 91180
rect 102100 91140 115204 91168
rect 102100 91128 102106 91140
rect 115198 91128 115204 91140
rect 115256 91128 115262 91180
rect 152090 91128 152096 91180
rect 152148 91168 152154 91180
rect 158714 91168 158720 91180
rect 152148 91140 158720 91168
rect 152148 91128 152154 91140
rect 158714 91128 158720 91140
rect 158772 91128 158778 91180
rect 89070 91060 89076 91112
rect 89128 91100 89134 91112
rect 122098 91100 122104 91112
rect 89128 91072 122104 91100
rect 89128 91060 89134 91072
rect 122098 91060 122104 91072
rect 122156 91060 122162 91112
rect 132402 91060 132408 91112
rect 132460 91100 132466 91112
rect 134518 91100 134524 91112
rect 132460 91072 134524 91100
rect 132460 91060 132466 91072
rect 134518 91060 134524 91072
rect 134576 91060 134582 91112
rect 134702 91060 134708 91112
rect 134760 91100 134766 91112
rect 153102 91100 153108 91112
rect 134760 91072 153108 91100
rect 134760 91060 134766 91072
rect 153102 91060 153108 91072
rect 153160 91060 153166 91112
rect 112346 90992 112352 91044
rect 112404 91032 112410 91044
rect 210418 91032 210424 91044
rect 112404 91004 210424 91032
rect 112404 90992 112410 91004
rect 210418 90992 210424 91004
rect 210476 90992 210482 91044
rect 110322 90924 110328 90976
rect 110380 90964 110386 90976
rect 170582 90964 170588 90976
rect 110380 90936 170588 90964
rect 110380 90924 110386 90936
rect 170582 90924 170588 90936
rect 170640 90924 170646 90976
rect 222838 90380 222844 90432
rect 222896 90420 222902 90432
rect 235350 90420 235356 90432
rect 222896 90392 235356 90420
rect 222896 90380 222902 90392
rect 235350 90380 235356 90392
rect 235408 90380 235414 90432
rect 65978 90312 65984 90364
rect 66036 90352 66042 90364
rect 111058 90352 111064 90364
rect 66036 90324 111064 90352
rect 66036 90312 66042 90324
rect 111058 90312 111064 90324
rect 111116 90312 111122 90364
rect 220078 90312 220084 90364
rect 220136 90352 220142 90364
rect 263134 90352 263140 90364
rect 220136 90324 263140 90352
rect 220136 90312 220142 90324
rect 263134 90312 263140 90324
rect 263192 90312 263198 90364
rect 119706 89632 119712 89684
rect 119764 89672 119770 89684
rect 199470 89672 199476 89684
rect 119764 89644 199476 89672
rect 119764 89632 119770 89644
rect 199470 89632 199476 89644
rect 199528 89632 199534 89684
rect 121730 89564 121736 89616
rect 121788 89604 121794 89616
rect 170490 89604 170496 89616
rect 121788 89576 170496 89604
rect 121788 89564 121794 89576
rect 170490 89564 170496 89576
rect 170548 89564 170554 89616
rect 218698 89020 218704 89072
rect 218756 89060 218762 89072
rect 239674 89060 239680 89072
rect 218756 89032 239680 89060
rect 218756 89020 218762 89032
rect 239674 89020 239680 89032
rect 239732 89020 239738 89072
rect 103330 88952 103336 89004
rect 103388 88992 103394 89004
rect 120074 88992 120080 89004
rect 103388 88964 120080 88992
rect 103388 88952 103394 88964
rect 120074 88952 120080 88964
rect 120132 88952 120138 89004
rect 171778 88952 171784 89004
rect 171836 88992 171842 89004
rect 209222 88992 209228 89004
rect 171836 88964 209228 88992
rect 171836 88952 171842 88964
rect 209222 88952 209228 88964
rect 209280 88952 209286 89004
rect 214558 88952 214564 89004
rect 214616 88992 214622 89004
rect 261754 88992 261760 89004
rect 214616 88964 261760 88992
rect 214616 88952 214622 88964
rect 261754 88952 261760 88964
rect 261812 88952 261818 89004
rect 120810 88272 120816 88324
rect 120868 88312 120874 88324
rect 216122 88312 216128 88324
rect 120868 88284 216128 88312
rect 120868 88272 120874 88284
rect 216122 88272 216128 88284
rect 216180 88272 216186 88324
rect 114370 88204 114376 88256
rect 114428 88244 114434 88256
rect 205174 88244 205180 88256
rect 114428 88216 205180 88244
rect 114428 88204 114434 88216
rect 205174 88204 205180 88216
rect 205232 88204 205238 88256
rect 209130 87660 209136 87712
rect 209188 87700 209194 87712
rect 232774 87700 232780 87712
rect 209188 87672 232780 87700
rect 209188 87660 209194 87672
rect 232774 87660 232780 87672
rect 232832 87660 232838 87712
rect 67726 87592 67732 87644
rect 67784 87632 67790 87644
rect 105538 87632 105544 87644
rect 67784 87604 105544 87632
rect 67784 87592 67790 87604
rect 105538 87592 105544 87604
rect 105596 87592 105602 87644
rect 227070 87592 227076 87644
rect 227128 87632 227134 87644
rect 253382 87632 253388 87644
rect 227128 87604 253388 87632
rect 227128 87592 227134 87604
rect 253382 87592 253388 87604
rect 253440 87592 253446 87644
rect 111242 86912 111248 86964
rect 111300 86952 111306 86964
rect 184474 86952 184480 86964
rect 111300 86924 184480 86952
rect 111300 86912 111306 86924
rect 184474 86912 184480 86924
rect 184532 86912 184538 86964
rect 158714 86844 158720 86896
rect 158772 86884 158778 86896
rect 206278 86884 206284 86896
rect 158772 86856 206284 86884
rect 158772 86844 158778 86856
rect 206278 86844 206284 86856
rect 206336 86844 206342 86896
rect 3234 86232 3240 86284
rect 3292 86272 3298 86284
rect 21358 86272 21364 86284
rect 3292 86244 21364 86272
rect 3292 86232 3298 86244
rect 21358 86232 21364 86244
rect 21416 86232 21422 86284
rect 66070 86232 66076 86284
rect 66128 86272 66134 86284
rect 111150 86272 111156 86284
rect 66128 86244 111156 86272
rect 66128 86232 66134 86244
rect 111150 86232 111156 86244
rect 111208 86232 111214 86284
rect 184290 86232 184296 86284
rect 184348 86272 184354 86284
rect 261662 86272 261668 86284
rect 184348 86244 261668 86272
rect 184348 86232 184354 86244
rect 261662 86232 261668 86244
rect 261720 86232 261726 86284
rect 104250 85484 104256 85536
rect 104308 85524 104314 85536
rect 193950 85524 193956 85536
rect 104308 85496 193956 85524
rect 104308 85484 104314 85496
rect 193950 85484 193956 85496
rect 194008 85484 194014 85536
rect 151538 85416 151544 85468
rect 151596 85456 151602 85468
rect 174630 85456 174636 85468
rect 151596 85428 174636 85456
rect 151596 85416 151602 85428
rect 174630 85416 174636 85428
rect 174688 85416 174694 85468
rect 206278 84872 206284 84924
rect 206336 84912 206342 84924
rect 231210 84912 231216 84924
rect 206336 84884 231216 84912
rect 206336 84872 206342 84884
rect 231210 84872 231216 84884
rect 231268 84872 231274 84924
rect 67358 84804 67364 84856
rect 67416 84844 67422 84856
rect 120718 84844 120724 84856
rect 67416 84816 120724 84844
rect 67416 84804 67422 84816
rect 120718 84804 120724 84816
rect 120776 84804 120782 84856
rect 204990 84804 204996 84856
rect 205048 84844 205054 84856
rect 264422 84844 264428 84856
rect 205048 84816 264428 84844
rect 205048 84804 205054 84816
rect 264422 84804 264428 84816
rect 264480 84804 264486 84856
rect 93762 84124 93768 84176
rect 93820 84164 93826 84176
rect 202322 84164 202328 84176
rect 93820 84136 202328 84164
rect 93820 84124 93826 84136
rect 202322 84124 202328 84136
rect 202380 84124 202386 84176
rect 126698 84056 126704 84108
rect 126756 84096 126762 84108
rect 182910 84096 182916 84108
rect 126756 84068 182916 84096
rect 126756 84056 126762 84068
rect 182910 84056 182916 84068
rect 182968 84056 182974 84108
rect 207658 83444 207664 83496
rect 207716 83484 207722 83496
rect 284938 83484 284944 83496
rect 207716 83456 284944 83484
rect 207716 83444 207722 83456
rect 284938 83444 284944 83456
rect 284996 83444 285002 83496
rect 85482 82764 85488 82816
rect 85540 82804 85546 82816
rect 177482 82804 177488 82816
rect 85540 82776 177488 82804
rect 85540 82764 85546 82776
rect 177482 82764 177488 82776
rect 177540 82764 177546 82816
rect 126790 82696 126796 82748
rect 126848 82736 126854 82748
rect 162210 82736 162216 82748
rect 126848 82708 162216 82736
rect 126848 82696 126854 82708
rect 162210 82696 162216 82708
rect 162268 82696 162274 82748
rect 204898 82084 204904 82136
rect 204956 82124 204962 82136
rect 238294 82124 238300 82136
rect 204956 82096 238300 82124
rect 204956 82084 204962 82096
rect 238294 82084 238300 82096
rect 238352 82084 238358 82136
rect 99190 81336 99196 81388
rect 99248 81376 99254 81388
rect 196802 81376 196808 81388
rect 99248 81348 196808 81376
rect 99248 81336 99254 81348
rect 196802 81336 196808 81348
rect 196860 81336 196866 81388
rect 126882 81268 126888 81320
rect 126940 81308 126946 81320
rect 164878 81308 164884 81320
rect 126940 81280 164884 81308
rect 126940 81268 126946 81280
rect 164878 81268 164884 81280
rect 164936 81268 164942 81320
rect 115842 79976 115848 80028
rect 115900 80016 115906 80028
rect 173434 80016 173440 80028
rect 115900 79988 173440 80016
rect 115900 79976 115906 79988
rect 173434 79976 173440 79988
rect 173492 79976 173498 80028
rect 133782 79908 133788 79960
rect 133840 79948 133846 79960
rect 166258 79948 166264 79960
rect 133840 79920 166264 79948
rect 133840 79908 133846 79920
rect 166258 79908 166264 79920
rect 166316 79908 166322 79960
rect 151630 78616 151636 78668
rect 151688 78656 151694 78668
rect 198182 78656 198188 78668
rect 151688 78628 198188 78656
rect 151688 78616 151694 78628
rect 198182 78616 198188 78628
rect 198240 78616 198246 78668
rect 128998 78548 129004 78600
rect 129056 78588 129062 78600
rect 157978 78588 157984 78600
rect 129056 78560 157984 78588
rect 129056 78548 129062 78560
rect 157978 78548 157984 78560
rect 158036 78548 158042 78600
rect 159358 77936 159364 77988
rect 159416 77976 159422 77988
rect 254762 77976 254768 77988
rect 159416 77948 254768 77976
rect 159416 77936 159422 77948
rect 254762 77936 254768 77948
rect 254820 77936 254826 77988
rect 64782 77188 64788 77240
rect 64840 77228 64846 77240
rect 171962 77228 171968 77240
rect 64840 77200 171968 77228
rect 64840 77188 64846 77200
rect 171962 77188 171968 77200
rect 172020 77188 172026 77240
rect 117222 77120 117228 77172
rect 117280 77160 117286 77172
rect 160738 77160 160744 77172
rect 117280 77132 160744 77160
rect 117280 77120 117286 77132
rect 160738 77120 160744 77132
rect 160796 77120 160802 77172
rect 115290 75828 115296 75880
rect 115348 75868 115354 75880
rect 200850 75868 200856 75880
rect 115348 75840 200856 75868
rect 115348 75828 115354 75840
rect 200850 75828 200856 75840
rect 200908 75828 200914 75880
rect 111150 75760 111156 75812
rect 111208 75800 111214 75812
rect 185578 75800 185584 75812
rect 111208 75772 185584 75800
rect 111208 75760 111214 75772
rect 185578 75760 185584 75772
rect 185636 75760 185642 75812
rect 106090 74468 106096 74520
rect 106148 74508 106154 74520
rect 177390 74508 177396 74520
rect 106148 74480 177396 74508
rect 106148 74468 106154 74480
rect 177390 74468 177396 74480
rect 177448 74468 177454 74520
rect 124030 74400 124036 74452
rect 124088 74440 124094 74452
rect 167730 74440 167736 74452
rect 124088 74412 167736 74440
rect 124088 74400 124094 74412
rect 167730 74400 167736 74412
rect 167788 74400 167794 74452
rect 111702 73108 111708 73160
rect 111760 73148 111766 73160
rect 173158 73148 173164 73160
rect 111760 73120 173164 73148
rect 111760 73108 111766 73120
rect 173158 73108 173164 73120
rect 173216 73108 173222 73160
rect 123478 73040 123484 73092
rect 123536 73080 123542 73092
rect 178862 73080 178868 73092
rect 123536 73052 178868 73080
rect 123536 73040 123542 73052
rect 178862 73040 178868 73052
rect 178920 73040 178926 73092
rect 3510 71680 3516 71732
rect 3568 71720 3574 71732
rect 36538 71720 36544 71732
rect 3568 71692 36544 71720
rect 3568 71680 3574 71692
rect 36538 71680 36544 71692
rect 36596 71680 36602 71732
rect 101950 71680 101956 71732
rect 102008 71720 102014 71732
rect 164970 71720 164976 71732
rect 102008 71692 164976 71720
rect 102008 71680 102014 71692
rect 164970 71680 164976 71692
rect 165028 71680 165034 71732
rect 128262 71612 128268 71664
rect 128320 71652 128326 71664
rect 181622 71652 181628 71664
rect 128320 71624 181628 71652
rect 128320 71612 128326 71624
rect 181622 71612 181628 71624
rect 181680 71612 181686 71664
rect 120718 70320 120724 70372
rect 120776 70360 120782 70372
rect 196710 70360 196716 70372
rect 120776 70332 196716 70360
rect 120776 70320 120782 70332
rect 196710 70320 196716 70332
rect 196768 70320 196774 70372
rect 112990 70252 112996 70304
rect 113048 70292 113054 70304
rect 180058 70292 180064 70304
rect 113048 70264 180064 70292
rect 113048 70252 113054 70264
rect 180058 70252 180064 70264
rect 180116 70252 180122 70304
rect 115198 68960 115204 69012
rect 115256 69000 115262 69012
rect 205082 69000 205088 69012
rect 115256 68972 205088 69000
rect 115256 68960 115262 68972
rect 205082 68960 205088 68972
rect 205140 68960 205146 69012
rect 110230 68892 110236 68944
rect 110288 68932 110294 68944
rect 187050 68932 187056 68944
rect 110288 68904 187056 68932
rect 110288 68892 110294 68904
rect 187050 68892 187056 68904
rect 187108 68892 187114 68944
rect 105538 67532 105544 67584
rect 105596 67572 105602 67584
rect 214650 67572 214656 67584
rect 105596 67544 214656 67572
rect 105596 67532 105602 67544
rect 214650 67532 214656 67544
rect 214708 67532 214714 67584
rect 151722 67464 151728 67516
rect 151780 67504 151786 67516
rect 169018 67504 169024 67516
rect 151780 67476 169024 67504
rect 151780 67464 151786 67476
rect 169018 67464 169024 67476
rect 169076 67464 169082 67516
rect 101858 66172 101864 66224
rect 101916 66212 101922 66224
rect 176102 66212 176108 66224
rect 101916 66184 176108 66212
rect 101916 66172 101922 66184
rect 176102 66172 176108 66184
rect 176160 66172 176166 66224
rect 307754 66172 307760 66224
rect 307812 66212 307818 66224
rect 338758 66212 338764 66224
rect 307812 66184 338764 66212
rect 307812 66172 307818 66184
rect 338758 66172 338764 66184
rect 338816 66172 338822 66224
rect 125410 66104 125416 66156
rect 125468 66144 125474 66156
rect 193858 66144 193864 66156
rect 125468 66116 193864 66144
rect 125468 66104 125474 66116
rect 193858 66104 193864 66116
rect 193916 66104 193922 66156
rect 110138 64812 110144 64864
rect 110196 64852 110202 64864
rect 213270 64852 213276 64864
rect 110196 64824 213276 64852
rect 110196 64812 110202 64824
rect 213270 64812 213276 64824
rect 213328 64812 213334 64864
rect 86862 64132 86868 64184
rect 86920 64172 86926 64184
rect 249150 64172 249156 64184
rect 86920 64144 249156 64172
rect 86920 64132 86926 64144
rect 249150 64132 249156 64144
rect 249208 64132 249214 64184
rect 97902 63452 97908 63504
rect 97960 63492 97966 63504
rect 199378 63492 199384 63504
rect 97960 63464 199384 63492
rect 97960 63452 97966 63464
rect 199378 63452 199384 63464
rect 199436 63452 199442 63504
rect 122098 63384 122104 63436
rect 122156 63424 122162 63436
rect 173342 63424 173348 63436
rect 122156 63396 173348 63424
rect 122156 63384 122162 63396
rect 173342 63384 173348 63396
rect 173400 63384 173406 63436
rect 134518 62024 134524 62076
rect 134576 62064 134582 62076
rect 215938 62064 215944 62076
rect 134576 62036 215944 62064
rect 134576 62024 134582 62036
rect 215938 62024 215944 62036
rect 215996 62024 216002 62076
rect 119890 61956 119896 62008
rect 119948 61996 119954 62008
rect 178770 61996 178776 62008
rect 119948 61968 178776 61996
rect 119948 61956 119954 61968
rect 178770 61956 178776 61968
rect 178828 61956 178834 62008
rect 125502 60664 125508 60716
rect 125560 60704 125566 60716
rect 203518 60704 203524 60716
rect 125560 60676 203524 60704
rect 125560 60664 125566 60676
rect 203518 60664 203524 60676
rect 203576 60664 203582 60716
rect 244274 60052 244280 60104
rect 244332 60092 244338 60104
rect 302234 60092 302240 60104
rect 244332 60064 302240 60092
rect 244332 60052 244338 60064
rect 302234 60052 302240 60064
rect 302292 60052 302298 60104
rect 97902 59984 97908 60036
rect 97960 60024 97966 60036
rect 245102 60024 245108 60036
rect 97960 59996 245108 60024
rect 97960 59984 97966 59996
rect 245102 59984 245108 59996
rect 245160 59984 245166 60036
rect 99282 59304 99288 59356
rect 99340 59344 99346 59356
rect 170398 59344 170404 59356
rect 99340 59316 170404 59344
rect 99340 59304 99346 59316
rect 170398 59304 170404 59316
rect 170456 59304 170462 59356
rect 3326 58828 3332 58880
rect 3384 58868 3390 58880
rect 7558 58868 7564 58880
rect 3384 58840 7564 58868
rect 3384 58828 3390 58840
rect 7558 58828 7564 58840
rect 7616 58828 7622 58880
rect 102042 58624 102048 58676
rect 102100 58664 102106 58676
rect 264330 58664 264336 58676
rect 102100 58636 264336 58664
rect 102100 58624 102106 58636
rect 264330 58624 264336 58636
rect 264388 58624 264394 58676
rect 106918 57876 106924 57928
rect 106976 57916 106982 57928
rect 207750 57916 207756 57928
rect 106976 57888 207756 57916
rect 106976 57876 106982 57888
rect 207750 57876 207756 57888
rect 207808 57876 207814 57928
rect 111702 57196 111708 57248
rect 111760 57236 111766 57248
rect 267734 57236 267740 57248
rect 111760 57208 267740 57236
rect 111760 57196 111766 57208
rect 267734 57196 267740 57208
rect 267792 57196 267798 57248
rect 91002 56516 91008 56568
rect 91060 56556 91066 56568
rect 191282 56556 191288 56568
rect 91060 56528 191288 56556
rect 91060 56516 91066 56528
rect 191282 56516 191288 56528
rect 191340 56516 191346 56568
rect 115842 55836 115848 55888
rect 115900 55876 115906 55888
rect 245010 55876 245016 55888
rect 115900 55848 245016 55876
rect 115900 55836 115906 55848
rect 245010 55836 245016 55848
rect 245068 55836 245074 55888
rect 75730 55156 75736 55208
rect 75788 55196 75794 55208
rect 206370 55196 206376 55208
rect 75788 55168 206376 55196
rect 75788 55156 75794 55168
rect 206370 55156 206376 55168
rect 206428 55156 206434 55208
rect 123478 54476 123484 54528
rect 123536 54516 123542 54528
rect 209130 54516 209136 54528
rect 123536 54488 209136 54516
rect 123536 54476 123542 54488
rect 209130 54476 209136 54488
rect 209188 54476 209194 54528
rect 118602 53728 118608 53780
rect 118660 53768 118666 53780
rect 178678 53768 178684 53780
rect 118660 53740 178684 53768
rect 118660 53728 118666 53740
rect 178678 53728 178684 53740
rect 178736 53728 178742 53780
rect 88978 53116 88984 53168
rect 89036 53156 89042 53168
rect 112438 53156 112444 53168
rect 89036 53128 112444 53156
rect 89036 53116 89042 53128
rect 112438 53116 112444 53128
rect 112496 53116 112502 53168
rect 84102 53048 84108 53100
rect 84160 53088 84166 53100
rect 217318 53088 217324 53100
rect 84160 53060 217324 53088
rect 84160 53048 84166 53060
rect 217318 53048 217324 53060
rect 217376 53048 217382 53100
rect 103422 52368 103428 52420
rect 103480 52408 103486 52420
rect 202230 52408 202236 52420
rect 103480 52380 202236 52408
rect 103480 52368 103486 52380
rect 202230 52368 202236 52380
rect 202288 52368 202294 52420
rect 121362 51688 121368 51740
rect 121420 51728 121426 51740
rect 246390 51728 246396 51740
rect 121420 51700 246396 51728
rect 121420 51688 121426 51700
rect 246390 51688 246396 51700
rect 246448 51688 246454 51740
rect 114462 51008 114468 51060
rect 114520 51048 114526 51060
rect 198090 51048 198096 51060
rect 114520 51020 198096 51048
rect 114520 51008 114526 51020
rect 198090 51008 198096 51020
rect 198148 51008 198154 51060
rect 34422 50328 34428 50380
rect 34480 50368 34486 50380
rect 258718 50368 258724 50380
rect 34480 50340 258724 50368
rect 34480 50328 34486 50340
rect 258718 50328 258724 50340
rect 258776 50328 258782 50380
rect 123938 49648 123944 49700
rect 123996 49688 124002 49700
rect 188522 49688 188528 49700
rect 123996 49660 188528 49688
rect 123996 49648 124002 49660
rect 188522 49648 188528 49660
rect 188580 49648 188586 49700
rect 37182 48968 37188 49020
rect 37240 49008 37246 49020
rect 246482 49008 246488 49020
rect 37240 48980 246488 49008
rect 37240 48968 37246 48980
rect 246482 48968 246488 48980
rect 246540 48968 246546 49020
rect 90358 47608 90364 47660
rect 90416 47648 90422 47660
rect 274634 47648 274640 47660
rect 90416 47620 274640 47648
rect 90416 47608 90422 47620
rect 274634 47608 274640 47620
rect 274692 47608 274698 47660
rect 12342 47540 12348 47592
rect 12400 47580 12406 47592
rect 251910 47580 251916 47592
rect 12400 47552 251916 47580
rect 12400 47540 12406 47552
rect 251910 47540 251916 47552
rect 251968 47540 251974 47592
rect 98638 46248 98644 46300
rect 98696 46288 98702 46300
rect 270586 46288 270592 46300
rect 98696 46260 270592 46288
rect 98696 46248 98702 46260
rect 270586 46248 270592 46260
rect 270644 46248 270650 46300
rect 49602 46180 49608 46232
rect 49660 46220 49666 46232
rect 254578 46220 254584 46232
rect 49660 46192 254584 46220
rect 49660 46180 49666 46192
rect 254578 46180 254584 46192
rect 254636 46180 254642 46232
rect 3510 45500 3516 45552
rect 3568 45540 3574 45552
rect 43438 45540 43444 45552
rect 3568 45512 43444 45540
rect 3568 45500 3574 45512
rect 43438 45500 43444 45512
rect 43496 45500 43502 45552
rect 86770 44820 86776 44872
rect 86828 44860 86834 44872
rect 250530 44860 250536 44872
rect 86828 44832 250536 44860
rect 86828 44820 86834 44832
rect 250530 44820 250536 44832
rect 250588 44820 250594 44872
rect 87598 43460 87604 43512
rect 87656 43500 87662 43512
rect 210418 43500 210424 43512
rect 87656 43472 210424 43500
rect 87656 43460 87662 43472
rect 210418 43460 210424 43472
rect 210476 43460 210482 43512
rect 9582 43392 9588 43444
rect 9640 43432 9646 43444
rect 253198 43432 253204 43444
rect 9640 43404 253204 43432
rect 9640 43392 9646 43404
rect 253198 43392 253204 43404
rect 253256 43392 253262 43444
rect 91002 42032 91008 42084
rect 91060 42072 91066 42084
rect 262950 42072 262956 42084
rect 91060 42044 262956 42072
rect 91060 42032 91066 42044
rect 262950 42032 262956 42044
rect 263008 42032 263014 42084
rect 77202 40740 77208 40792
rect 77260 40780 77266 40792
rect 256050 40780 256056 40792
rect 77260 40752 256056 40780
rect 77260 40740 77266 40752
rect 256050 40740 256056 40752
rect 256108 40740 256114 40792
rect 28902 40672 28908 40724
rect 28960 40712 28966 40724
rect 270494 40712 270500 40724
rect 28960 40684 270500 40712
rect 28960 40672 28966 40684
rect 270494 40672 270500 40684
rect 270552 40672 270558 40724
rect 103422 39380 103428 39432
rect 103480 39420 103486 39432
rect 239398 39420 239404 39432
rect 103480 39392 239404 39420
rect 103480 39380 103486 39392
rect 239398 39380 239404 39392
rect 239456 39380 239462 39432
rect 59262 39312 59268 39364
rect 59320 39352 59326 39364
rect 238202 39352 238208 39364
rect 59320 39324 238208 39352
rect 59320 39312 59326 39324
rect 238202 39312 238208 39324
rect 238260 39312 238266 39364
rect 71038 37884 71044 37936
rect 71096 37924 71102 37936
rect 228358 37924 228364 37936
rect 71096 37896 228364 37924
rect 71096 37884 71102 37896
rect 228358 37884 228364 37896
rect 228416 37884 228422 37936
rect 125502 36592 125508 36644
rect 125560 36632 125566 36644
rect 151078 36632 151084 36644
rect 125560 36604 151084 36632
rect 125560 36592 125566 36604
rect 151078 36592 151084 36604
rect 151136 36592 151142 36644
rect 26142 36524 26148 36576
rect 26200 36564 26206 36576
rect 206278 36564 206284 36576
rect 26200 36536 206284 36564
rect 26200 36524 26206 36536
rect 206278 36524 206284 36536
rect 206336 36524 206342 36576
rect 206370 36524 206376 36576
rect 206428 36564 206434 36576
rect 224218 36564 224224 36576
rect 206428 36536 224224 36564
rect 206428 36524 206434 36536
rect 224218 36524 224224 36536
rect 224276 36524 224282 36576
rect 116578 35232 116584 35284
rect 116636 35272 116642 35284
rect 184290 35272 184296 35284
rect 116636 35244 184296 35272
rect 116636 35232 116642 35244
rect 184290 35232 184296 35244
rect 184348 35232 184354 35284
rect 192478 35232 192484 35284
rect 192536 35272 192542 35284
rect 220170 35272 220176 35284
rect 192536 35244 220176 35272
rect 192536 35232 192542 35244
rect 220170 35232 220176 35244
rect 220228 35232 220234 35284
rect 182910 35164 182916 35216
rect 182968 35204 182974 35216
rect 269114 35204 269120 35216
rect 182968 35176 269120 35204
rect 182968 35164 182974 35176
rect 269114 35164 269120 35176
rect 269172 35164 269178 35216
rect 2866 33056 2872 33108
rect 2924 33096 2930 33108
rect 32398 33096 32404 33108
rect 2924 33068 32404 33096
rect 2924 33056 2930 33068
rect 32398 33056 32404 33068
rect 32456 33056 32462 33108
rect 583386 33056 583392 33108
rect 583444 33096 583450 33108
rect 583662 33096 583668 33108
rect 583444 33068 583668 33096
rect 583444 33056 583450 33068
rect 583662 33056 583668 33068
rect 583720 33056 583726 33108
rect 110322 32444 110328 32496
rect 110380 32484 110386 32496
rect 260190 32484 260196 32496
rect 110380 32456 260196 32484
rect 110380 32444 110386 32456
rect 260190 32444 260196 32456
rect 260248 32444 260254 32496
rect 52362 32376 52368 32428
rect 52420 32416 52426 32428
rect 250530 32416 250536 32428
rect 52420 32388 250536 32416
rect 52420 32376 52426 32388
rect 250530 32376 250536 32388
rect 250588 32376 250594 32428
rect 61930 31084 61936 31136
rect 61988 31124 61994 31136
rect 220078 31124 220084 31136
rect 61988 31096 220084 31124
rect 61988 31084 61994 31096
rect 220078 31084 220084 31096
rect 220136 31084 220142 31136
rect 74442 31016 74448 31068
rect 74500 31056 74506 31068
rect 251818 31056 251824 31068
rect 74500 31028 251824 31056
rect 74500 31016 74506 31028
rect 251818 31016 251824 31028
rect 251876 31016 251882 31068
rect 13722 29656 13728 29708
rect 13780 29696 13786 29708
rect 250438 29696 250444 29708
rect 13780 29668 250444 29696
rect 13780 29656 13786 29668
rect 250438 29656 250444 29668
rect 250496 29656 250502 29708
rect 63402 29588 63408 29640
rect 63460 29628 63466 29640
rect 310514 29628 310520 29640
rect 63460 29600 310520 29628
rect 63460 29588 63466 29600
rect 310514 29588 310520 29600
rect 310572 29588 310578 29640
rect 85482 28296 85488 28348
rect 85540 28336 85546 28348
rect 260098 28336 260104 28348
rect 85540 28308 260104 28336
rect 85540 28296 85546 28308
rect 260098 28296 260104 28308
rect 260156 28296 260162 28348
rect 1394 28228 1400 28280
rect 1452 28268 1458 28280
rect 231118 28268 231124 28280
rect 1452 28240 231124 28268
rect 1452 28228 1458 28240
rect 231118 28228 231124 28240
rect 231176 28228 231182 28280
rect 48222 26868 48228 26920
rect 48280 26908 48286 26920
rect 251174 26908 251180 26920
rect 48280 26880 251180 26908
rect 48280 26868 48286 26880
rect 251174 26868 251180 26880
rect 251232 26868 251238 26920
rect 92382 25576 92388 25628
rect 92440 25616 92446 25628
rect 240778 25616 240784 25628
rect 92440 25588 240784 25616
rect 92440 25576 92446 25588
rect 240778 25576 240784 25588
rect 240836 25576 240842 25628
rect 73062 25508 73068 25560
rect 73120 25548 73126 25560
rect 267826 25548 267832 25560
rect 73120 25520 267832 25548
rect 73120 25508 73126 25520
rect 267826 25508 267832 25520
rect 267884 25508 267890 25560
rect 322198 25508 322204 25560
rect 322256 25548 322262 25560
rect 328454 25548 328460 25560
rect 322256 25520 328460 25548
rect 322256 25508 322262 25520
rect 328454 25508 328460 25520
rect 328512 25508 328518 25560
rect 20622 24148 20628 24200
rect 20680 24188 20686 24200
rect 247678 24188 247684 24200
rect 20680 24160 247684 24188
rect 20680 24148 20686 24160
rect 247678 24148 247684 24160
rect 247736 24148 247742 24200
rect 57238 24080 57244 24132
rect 57296 24120 57302 24132
rect 324406 24120 324412 24132
rect 57296 24092 324412 24120
rect 57296 24080 57302 24092
rect 324406 24080 324412 24092
rect 324464 24080 324470 24132
rect 56502 22788 56508 22840
rect 56560 22828 56566 22840
rect 216030 22828 216036 22840
rect 56560 22800 216036 22828
rect 56560 22788 56566 22800
rect 216030 22788 216036 22800
rect 216088 22788 216094 22840
rect 88242 22720 88248 22772
rect 88300 22760 88306 22772
rect 255958 22760 255964 22772
rect 88300 22732 255964 22760
rect 88300 22720 88306 22732
rect 255958 22720 255964 22732
rect 256016 22720 256022 22772
rect 37090 21428 37096 21480
rect 37148 21468 37154 21480
rect 225598 21468 225604 21480
rect 37148 21440 225604 21468
rect 37148 21428 37154 21440
rect 225598 21428 225604 21440
rect 225656 21428 225662 21480
rect 46842 21360 46848 21412
rect 46900 21400 46906 21412
rect 238110 21400 238116 21412
rect 46900 21372 238116 21400
rect 46900 21360 46906 21372
rect 238110 21360 238116 21372
rect 238168 21360 238174 21412
rect 114462 20000 114468 20052
rect 114520 20040 114526 20052
rect 182910 20040 182916 20052
rect 114520 20012 182916 20040
rect 114520 20000 114526 20012
rect 182910 20000 182916 20012
rect 182968 20000 182974 20052
rect 187050 20000 187056 20052
rect 187108 20040 187114 20052
rect 209038 20040 209044 20052
rect 187108 20012 209044 20040
rect 187108 20000 187114 20012
rect 209038 20000 209044 20012
rect 209096 20000 209102 20052
rect 24762 19932 24768 19984
rect 24820 19972 24826 19984
rect 159358 19972 159364 19984
rect 24820 19944 159364 19972
rect 24820 19932 24826 19944
rect 159358 19932 159364 19944
rect 159416 19932 159422 19984
rect 184198 19932 184204 19984
rect 184256 19972 184262 19984
rect 291838 19972 291844 19984
rect 184256 19944 291844 19972
rect 184256 19932 184262 19944
rect 291838 19932 291844 19944
rect 291896 19932 291902 19984
rect 319438 19932 319444 19984
rect 319496 19972 319502 19984
rect 378134 19972 378140 19984
rect 319496 19944 378140 19972
rect 319496 19932 319502 19944
rect 378134 19932 378140 19944
rect 378192 19932 378198 19984
rect 6822 18640 6828 18692
rect 6880 18680 6886 18692
rect 98638 18680 98644 18692
rect 6880 18652 98644 18680
rect 6880 18640 6886 18652
rect 98638 18640 98644 18652
rect 98696 18640 98702 18692
rect 99282 18640 99288 18692
rect 99340 18680 99346 18692
rect 206370 18680 206376 18692
rect 99340 18652 206376 18680
rect 99340 18640 99346 18652
rect 206370 18640 206376 18652
rect 206428 18640 206434 18692
rect 65518 18572 65524 18624
rect 65576 18612 65582 18624
rect 262858 18612 262864 18624
rect 65576 18584 262864 18612
rect 65576 18572 65582 18584
rect 262858 18572 262864 18584
rect 262916 18572 262922 18624
rect 119890 17212 119896 17264
rect 119948 17252 119954 17264
rect 204990 17252 204996 17264
rect 119948 17224 204996 17252
rect 119948 17212 119954 17224
rect 204990 17212 204996 17224
rect 205048 17212 205054 17264
rect 259546 17212 259552 17264
rect 259604 17252 259610 17264
rect 276014 17252 276020 17264
rect 259604 17224 276020 17252
rect 259604 17212 259610 17224
rect 276014 17212 276020 17224
rect 276072 17212 276078 17264
rect 96246 15920 96252 15972
rect 96304 15960 96310 15972
rect 222838 15960 222844 15972
rect 96304 15932 222844 15960
rect 96304 15920 96310 15932
rect 222838 15920 222844 15932
rect 222896 15920 222902 15972
rect 309778 15920 309784 15972
rect 309836 15960 309842 15972
rect 322106 15960 322112 15972
rect 309836 15932 322112 15960
rect 309836 15920 309842 15932
rect 322106 15920 322112 15932
rect 322164 15920 322170 15972
rect 50982 15852 50988 15904
rect 51040 15892 51046 15904
rect 297266 15892 297272 15904
rect 51040 15864 297272 15892
rect 51040 15852 51046 15864
rect 297266 15852 297272 15864
rect 297324 15852 297330 15904
rect 313918 15852 313924 15904
rect 313976 15892 313982 15904
rect 345290 15892 345296 15904
rect 313976 15864 345296 15892
rect 313976 15852 313982 15864
rect 345290 15852 345296 15864
rect 345348 15852 345354 15904
rect 118602 14492 118608 14544
rect 118660 14532 118666 14544
rect 233878 14532 233884 14544
rect 118660 14504 233884 14532
rect 118660 14492 118666 14504
rect 233878 14492 233884 14504
rect 233936 14492 233942 14544
rect 27522 14424 27528 14476
rect 27580 14464 27586 14476
rect 227070 14464 227076 14476
rect 27580 14436 227076 14464
rect 27580 14424 27586 14436
rect 227070 14424 227076 14436
rect 227128 14424 227134 14476
rect 331214 14424 331220 14476
rect 331272 14464 331278 14476
rect 373994 14464 374000 14476
rect 331272 14436 374000 14464
rect 331272 14424 331278 14436
rect 373994 14424 374000 14436
rect 374052 14424 374058 14476
rect 300118 13744 300124 13796
rect 300176 13784 300182 13796
rect 349154 13784 349160 13796
rect 300176 13756 349160 13784
rect 300176 13744 300182 13756
rect 349154 13744 349160 13756
rect 349212 13744 349218 13796
rect 100662 13132 100668 13184
rect 100720 13172 100726 13184
rect 242158 13172 242164 13184
rect 100720 13144 242164 13172
rect 100720 13132 100726 13144
rect 242158 13132 242164 13144
rect 242216 13132 242222 13184
rect 28810 13064 28816 13116
rect 28868 13104 28874 13116
rect 242250 13104 242256 13116
rect 28868 13076 242256 13104
rect 28868 13064 28874 13076
rect 242250 13064 242256 13076
rect 242308 13064 242314 13116
rect 299658 12452 299664 12504
rect 299716 12492 299722 12504
rect 300118 12492 300124 12504
rect 299716 12464 300124 12492
rect 299716 12452 299722 12464
rect 300118 12452 300124 12464
rect 300176 12452 300182 12504
rect 81342 11772 81348 11824
rect 81400 11812 81406 11824
rect 204898 11812 204904 11824
rect 81400 11784 204904 11812
rect 81400 11772 81406 11784
rect 204898 11772 204904 11784
rect 204956 11772 204962 11824
rect 340966 11772 340972 11824
rect 341024 11812 341030 11824
rect 342162 11812 342168 11824
rect 341024 11784 342168 11812
rect 341024 11772 341030 11784
rect 342162 11772 342168 11784
rect 342220 11772 342226 11824
rect 53650 11704 53656 11756
rect 53708 11744 53714 11756
rect 238018 11744 238024 11756
rect 53708 11716 238024 11744
rect 53708 11704 53714 11716
rect 238018 11704 238024 11716
rect 238076 11704 238082 11756
rect 257062 11704 257068 11756
rect 257120 11744 257126 11756
rect 358814 11744 358820 11756
rect 257120 11716 358820 11744
rect 257120 11704 257126 11716
rect 358814 11704 358820 11716
rect 358872 11704 358878 11756
rect 67542 10344 67548 10396
rect 67600 10384 67606 10396
rect 264238 10384 264244 10396
rect 67600 10356 264244 10384
rect 67600 10344 67606 10356
rect 264238 10344 264244 10356
rect 264296 10344 264302 10396
rect 42702 10276 42708 10328
rect 42760 10316 42766 10328
rect 243538 10316 243544 10328
rect 42760 10288 243544 10316
rect 42760 10276 42766 10288
rect 243538 10276 243544 10288
rect 243596 10276 243602 10328
rect 249978 9596 249984 9648
rect 250036 9636 250042 9648
rect 250530 9636 250536 9648
rect 250036 9608 250536 9636
rect 250036 9596 250042 9608
rect 250530 9596 250536 9608
rect 250588 9636 250594 9648
rect 376754 9636 376760 9648
rect 250588 9608 376760 9636
rect 250588 9596 250594 9608
rect 376754 9596 376760 9608
rect 376812 9596 376818 9648
rect 106918 8916 106924 8968
rect 106976 8956 106982 8968
rect 211798 8956 211804 8968
rect 106976 8928 211804 8956
rect 106976 8916 106982 8928
rect 211798 8916 211804 8928
rect 211856 8916 211862 8968
rect 71498 7624 71504 7676
rect 71556 7664 71562 7676
rect 226978 7664 226984 7676
rect 71556 7636 226984 7664
rect 71556 7624 71562 7636
rect 226978 7624 226984 7636
rect 227036 7624 227042 7676
rect 55122 7556 55128 7608
rect 55180 7596 55186 7608
rect 262950 7596 262956 7608
rect 55180 7568 262956 7596
rect 55180 7556 55186 7568
rect 262950 7556 262956 7568
rect 263008 7596 263014 7608
rect 375374 7596 375380 7608
rect 263008 7568 375380 7596
rect 263008 7556 263014 7568
rect 375374 7556 375380 7568
rect 375432 7556 375438 7608
rect 302878 6808 302884 6860
rect 302936 6848 302942 6860
rect 369854 6848 369860 6860
rect 302936 6820 369860 6848
rect 302936 6808 302942 6820
rect 369854 6808 369860 6820
rect 369912 6808 369918 6860
rect 574738 6808 574744 6860
rect 574796 6848 574802 6860
rect 580166 6848 580172 6860
rect 574796 6820 580172 6848
rect 574796 6808 574802 6820
rect 580166 6808 580172 6820
rect 580224 6808 580230 6860
rect 102226 6196 102232 6248
rect 102284 6236 102290 6248
rect 202138 6236 202144 6248
rect 102284 6208 202144 6236
rect 102284 6196 102290 6208
rect 202138 6196 202144 6208
rect 202196 6196 202202 6248
rect 17034 6128 17040 6180
rect 17092 6168 17098 6180
rect 249058 6168 249064 6180
rect 17092 6140 249064 6168
rect 17092 6128 17098 6140
rect 249058 6128 249064 6140
rect 249116 6128 249122 6180
rect 284938 6128 284944 6180
rect 284996 6168 285002 6180
rect 301958 6168 301964 6180
rect 284996 6140 301964 6168
rect 284996 6128 285002 6140
rect 301958 6128 301964 6140
rect 302016 6128 302022 6180
rect 325602 6128 325608 6180
rect 325660 6168 325666 6180
rect 332686 6168 332692 6180
rect 325660 6140 332692 6168
rect 325660 6128 325666 6140
rect 332686 6128 332692 6140
rect 332744 6128 332750 6180
rect 241698 5516 241704 5568
rect 241756 5556 241762 5568
rect 246298 5556 246304 5568
rect 241756 5528 246304 5556
rect 241756 5516 241762 5528
rect 246298 5516 246304 5528
rect 246356 5516 246362 5568
rect 305730 5516 305736 5568
rect 305788 5556 305794 5568
rect 307938 5556 307944 5568
rect 305788 5528 307944 5556
rect 305788 5516 305794 5528
rect 307938 5516 307944 5528
rect 307996 5516 308002 5568
rect 338666 5448 338672 5500
rect 338724 5488 338730 5500
rect 367094 5488 367100 5500
rect 338724 5460 367100 5488
rect 338724 5448 338730 5460
rect 367094 5448 367100 5460
rect 367152 5448 367158 5500
rect 54938 4836 54944 4888
rect 54996 4876 55002 4888
rect 214558 4876 214564 4888
rect 54996 4848 214564 4876
rect 54996 4836 55002 4848
rect 214558 4836 214564 4848
rect 214616 4836 214622 4888
rect 60826 4768 60832 4820
rect 60884 4808 60890 4820
rect 232498 4808 232504 4820
rect 60884 4780 232504 4808
rect 60884 4768 60890 4780
rect 232498 4768 232504 4780
rect 232556 4768 232562 4820
rect 232590 4156 232596 4208
rect 232648 4196 232654 4208
rect 235810 4196 235816 4208
rect 232648 4168 235816 4196
rect 232648 4156 232654 4168
rect 235810 4156 235816 4168
rect 235868 4156 235874 4208
rect 177298 4088 177304 4140
rect 177356 4128 177362 4140
rect 257062 4128 257068 4140
rect 177356 4100 257068 4128
rect 177356 4088 177362 4100
rect 257062 4088 257068 4100
rect 257120 4088 257126 4140
rect 296070 4088 296076 4140
rect 296128 4128 296134 4140
rect 298094 4128 298100 4140
rect 296128 4100 298100 4128
rect 296128 4088 296134 4100
rect 298094 4088 298100 4100
rect 298152 4088 298158 4140
rect 316678 4088 316684 4140
rect 316736 4128 316742 4140
rect 319714 4128 319720 4140
rect 316736 4100 319720 4128
rect 316736 4088 316742 4100
rect 319714 4088 319720 4100
rect 319772 4088 319778 4140
rect 116394 4020 116400 4072
rect 116452 4060 116458 4072
rect 123478 4060 123484 4072
rect 116452 4032 123484 4060
rect 116452 4020 116458 4032
rect 123478 4020 123484 4032
rect 123536 4020 123542 4072
rect 255866 4020 255872 4072
rect 255924 4060 255930 4072
rect 282178 4060 282184 4072
rect 255924 4032 282184 4060
rect 255924 4020 255930 4032
rect 282178 4020 282184 4032
rect 282236 4020 282242 4072
rect 310238 4020 310244 4072
rect 310296 4060 310302 4072
rect 317414 4060 317420 4072
rect 310296 4032 317420 4060
rect 310296 4020 310302 4032
rect 317414 4020 317420 4032
rect 317472 4020 317478 4072
rect 63218 3816 63224 3868
rect 63276 3856 63282 3868
rect 65518 3856 65524 3868
rect 63276 3828 65524 3856
rect 63276 3816 63282 3828
rect 65518 3816 65524 3828
rect 65576 3816 65582 3868
rect 305546 3748 305552 3800
rect 305604 3788 305610 3800
rect 306466 3788 306472 3800
rect 305604 3760 306472 3788
rect 305604 3748 305610 3760
rect 306466 3748 306472 3760
rect 306524 3748 306530 3800
rect 71038 3652 71044 3664
rect 64846 3624 71044 3652
rect 2866 3544 2872 3596
rect 2924 3584 2930 3596
rect 3970 3584 3976 3596
rect 2924 3556 3976 3584
rect 2924 3544 2930 3556
rect 3970 3544 3976 3556
rect 4028 3544 4034 3596
rect 8754 3476 8760 3528
rect 8812 3516 8818 3528
rect 9582 3516 9588 3528
rect 8812 3488 9588 3516
rect 8812 3476 8818 3488
rect 9582 3476 9588 3488
rect 9640 3476 9646 3528
rect 9950 3476 9956 3528
rect 10008 3516 10014 3528
rect 10962 3516 10968 3528
rect 10008 3488 10968 3516
rect 10008 3476 10014 3488
rect 10962 3476 10968 3488
rect 11020 3476 11026 3528
rect 15930 3476 15936 3528
rect 15988 3516 15994 3528
rect 16482 3516 16488 3528
rect 15988 3488 16488 3516
rect 15988 3476 15994 3488
rect 16482 3476 16488 3488
rect 16540 3476 16546 3528
rect 18230 3476 18236 3528
rect 18288 3516 18294 3528
rect 19242 3516 19248 3528
rect 18288 3488 19248 3516
rect 18288 3476 18294 3488
rect 19242 3476 19248 3488
rect 19300 3476 19306 3528
rect 24210 3476 24216 3528
rect 24268 3516 24274 3528
rect 24762 3516 24768 3528
rect 24268 3488 24768 3516
rect 24268 3476 24274 3488
rect 24762 3476 24768 3488
rect 24820 3476 24826 3528
rect 25314 3476 25320 3528
rect 25372 3516 25378 3528
rect 26142 3516 26148 3528
rect 25372 3488 26148 3516
rect 25372 3476 25378 3488
rect 26142 3476 26148 3488
rect 26200 3476 26206 3528
rect 26510 3476 26516 3528
rect 26568 3516 26574 3528
rect 27522 3516 27528 3528
rect 26568 3488 27528 3516
rect 26568 3476 26574 3488
rect 27522 3476 27528 3488
rect 27580 3476 27586 3528
rect 27706 3476 27712 3528
rect 27764 3516 27770 3528
rect 28810 3516 28816 3528
rect 27764 3488 28816 3516
rect 27764 3476 27770 3488
rect 28810 3476 28816 3488
rect 28868 3476 28874 3528
rect 32398 3476 32404 3528
rect 32456 3516 32462 3528
rect 33042 3516 33048 3528
rect 32456 3488 33048 3516
rect 32456 3476 32462 3488
rect 33042 3476 33048 3488
rect 33100 3476 33106 3528
rect 33594 3476 33600 3528
rect 33652 3516 33658 3528
rect 34422 3516 34428 3528
rect 33652 3488 34428 3516
rect 33652 3476 33658 3488
rect 34422 3476 34428 3488
rect 34480 3476 34486 3528
rect 34790 3476 34796 3528
rect 34848 3516 34854 3528
rect 35802 3516 35808 3528
rect 34848 3488 35808 3516
rect 34848 3476 34854 3488
rect 35802 3476 35808 3488
rect 35860 3476 35866 3528
rect 35986 3476 35992 3528
rect 36044 3516 36050 3528
rect 37090 3516 37096 3528
rect 36044 3488 37096 3516
rect 36044 3476 36050 3488
rect 37090 3476 37096 3488
rect 37148 3476 37154 3528
rect 40678 3476 40684 3528
rect 40736 3516 40742 3528
rect 41322 3516 41328 3528
rect 40736 3488 41328 3516
rect 40736 3476 40742 3488
rect 41322 3476 41328 3488
rect 41380 3476 41386 3528
rect 41874 3476 41880 3528
rect 41932 3516 41938 3528
rect 42702 3516 42708 3528
rect 41932 3488 42708 3516
rect 41932 3476 41938 3488
rect 42702 3476 42708 3488
rect 42760 3476 42766 3528
rect 43070 3476 43076 3528
rect 43128 3516 43134 3528
rect 44082 3516 44088 3528
rect 43128 3488 44088 3516
rect 43128 3476 43134 3488
rect 44082 3476 44088 3488
rect 44140 3476 44146 3528
rect 44266 3476 44272 3528
rect 44324 3516 44330 3528
rect 64846 3516 64874 3624
rect 71038 3612 71044 3624
rect 71096 3612 71102 3664
rect 87598 3652 87604 3664
rect 84166 3624 87604 3652
rect 70210 3544 70216 3596
rect 70268 3584 70274 3596
rect 84166 3584 84194 3624
rect 87598 3612 87604 3624
rect 87656 3612 87662 3664
rect 70268 3556 84194 3584
rect 70268 3544 70274 3556
rect 85666 3544 85672 3596
rect 85724 3584 85730 3596
rect 86770 3584 86776 3596
rect 85724 3556 86776 3584
rect 85724 3544 85730 3556
rect 86770 3544 86776 3556
rect 86828 3544 86834 3596
rect 95050 3544 95056 3596
rect 95108 3584 95114 3596
rect 126238 3584 126244 3596
rect 95108 3556 103514 3584
rect 95108 3544 95114 3556
rect 44324 3488 64874 3516
rect 44324 3476 44330 3488
rect 66714 3476 66720 3528
rect 66772 3516 66778 3528
rect 67542 3516 67548 3528
rect 66772 3488 67548 3516
rect 66772 3476 66778 3488
rect 67542 3476 67548 3488
rect 67600 3476 67606 3528
rect 67910 3476 67916 3528
rect 67968 3516 67974 3528
rect 68922 3516 68928 3528
rect 67968 3488 68928 3516
rect 67968 3476 67974 3488
rect 68922 3476 68928 3488
rect 68980 3476 68986 3528
rect 69106 3476 69112 3528
rect 69164 3516 69170 3528
rect 70302 3516 70308 3528
rect 69164 3488 70308 3516
rect 69164 3476 69170 3488
rect 70302 3476 70308 3488
rect 70360 3476 70366 3528
rect 72602 3476 72608 3528
rect 72660 3516 72666 3528
rect 73062 3516 73068 3528
rect 72660 3488 73068 3516
rect 72660 3476 72666 3488
rect 73062 3476 73068 3488
rect 73120 3476 73126 3528
rect 73798 3476 73804 3528
rect 73856 3516 73862 3528
rect 74442 3516 74448 3528
rect 73856 3488 74448 3516
rect 73856 3476 73862 3488
rect 74442 3476 74448 3488
rect 74500 3476 74506 3528
rect 76190 3476 76196 3528
rect 76248 3516 76254 3528
rect 77202 3516 77208 3528
rect 76248 3488 77208 3516
rect 76248 3476 76254 3488
rect 77202 3476 77208 3488
rect 77260 3476 77266 3528
rect 80882 3476 80888 3528
rect 80940 3516 80946 3528
rect 81342 3516 81348 3528
rect 80940 3488 81348 3516
rect 80940 3476 80946 3488
rect 81342 3476 81348 3488
rect 81400 3476 81406 3528
rect 84470 3476 84476 3528
rect 84528 3516 84534 3528
rect 85482 3516 85488 3528
rect 84528 3488 85488 3516
rect 84528 3476 84534 3488
rect 85482 3476 85488 3488
rect 85540 3476 85546 3528
rect 89162 3476 89168 3528
rect 89220 3516 89226 3528
rect 89622 3516 89628 3528
rect 89220 3488 89628 3516
rect 89220 3476 89226 3488
rect 89622 3476 89628 3488
rect 89680 3476 89686 3528
rect 90358 3476 90364 3528
rect 90416 3516 90422 3528
rect 91002 3516 91008 3528
rect 90416 3488 91008 3516
rect 90416 3476 90422 3488
rect 91002 3476 91008 3488
rect 91060 3476 91066 3528
rect 91554 3476 91560 3528
rect 91612 3516 91618 3528
rect 92382 3516 92388 3528
rect 91612 3488 92388 3516
rect 91612 3476 91618 3488
rect 92382 3476 92388 3488
rect 92440 3476 92446 3528
rect 92750 3476 92756 3528
rect 92808 3516 92814 3528
rect 93762 3516 93768 3528
rect 92808 3488 93768 3516
rect 92808 3476 92814 3488
rect 93762 3476 93768 3488
rect 93820 3476 93826 3528
rect 93946 3476 93952 3528
rect 94004 3516 94010 3528
rect 95142 3516 95148 3528
rect 94004 3488 95148 3516
rect 94004 3476 94010 3488
rect 95142 3476 95148 3488
rect 95200 3476 95206 3528
rect 97442 3476 97448 3528
rect 97500 3516 97506 3528
rect 97902 3516 97908 3528
rect 97500 3488 97908 3516
rect 97500 3476 97506 3488
rect 97902 3476 97908 3488
rect 97960 3476 97966 3528
rect 98638 3476 98644 3528
rect 98696 3516 98702 3528
rect 99282 3516 99288 3528
rect 98696 3488 99288 3516
rect 98696 3476 98702 3488
rect 99282 3476 99288 3488
rect 99340 3476 99346 3528
rect 99834 3476 99840 3528
rect 99892 3516 99898 3528
rect 100662 3516 100668 3528
rect 99892 3488 100668 3516
rect 99892 3476 99898 3488
rect 100662 3476 100668 3488
rect 100720 3476 100726 3528
rect 101030 3476 101036 3528
rect 101088 3516 101094 3528
rect 102042 3516 102048 3528
rect 101088 3488 102048 3516
rect 101088 3476 101094 3488
rect 102042 3476 102048 3488
rect 102100 3476 102106 3528
rect 103486 3516 103514 3556
rect 122806 3556 126244 3584
rect 122806 3516 122834 3556
rect 126238 3544 126244 3556
rect 126296 3544 126302 3596
rect 103486 3488 122834 3516
rect 124674 3476 124680 3528
rect 124732 3516 124738 3528
rect 125502 3516 125508 3528
rect 124732 3488 125508 3516
rect 124732 3476 124738 3488
rect 125502 3476 125508 3488
rect 125560 3476 125566 3528
rect 129366 3476 129372 3528
rect 129424 3516 129430 3528
rect 130378 3516 130384 3528
rect 129424 3488 130384 3516
rect 129424 3476 129430 3488
rect 130378 3476 130384 3488
rect 130436 3476 130442 3528
rect 291838 3476 291844 3528
rect 291896 3516 291902 3528
rect 292574 3516 292580 3528
rect 291896 3488 292580 3516
rect 291896 3476 291902 3488
rect 292574 3476 292580 3488
rect 292632 3476 292638 3528
rect 307754 3476 307760 3528
rect 307812 3516 307818 3528
rect 309042 3516 309048 3528
rect 307812 3488 309048 3516
rect 307812 3476 307818 3488
rect 309042 3476 309048 3488
rect 309100 3476 309106 3528
rect 324314 3476 324320 3528
rect 324372 3516 324378 3528
rect 325602 3516 325608 3528
rect 324372 3488 325608 3516
rect 324372 3476 324378 3488
rect 325602 3476 325608 3488
rect 325660 3476 325666 3528
rect 335998 3476 336004 3528
rect 336056 3516 336062 3528
rect 337470 3516 337476 3528
rect 336056 3488 337476 3516
rect 336056 3476 336062 3488
rect 337470 3476 337476 3488
rect 337528 3476 337534 3528
rect 349246 3476 349252 3528
rect 349304 3516 349310 3528
rect 357434 3516 357440 3528
rect 349304 3488 357440 3516
rect 349304 3476 349310 3488
rect 357434 3476 357440 3488
rect 357492 3476 357498 3528
rect 580994 3476 581000 3528
rect 581052 3516 581058 3528
rect 583478 3516 583484 3528
rect 581052 3488 583484 3516
rect 581052 3476 581058 3488
rect 583478 3476 583484 3488
rect 583536 3476 583542 3528
rect 20530 3408 20536 3460
rect 20588 3448 20594 3460
rect 20588 3420 45554 3448
rect 20588 3408 20594 3420
rect 45526 3380 45554 3420
rect 48958 3408 48964 3460
rect 49016 3448 49022 3460
rect 49602 3448 49608 3460
rect 49016 3420 49608 3448
rect 49016 3408 49022 3420
rect 49602 3408 49608 3420
rect 49660 3408 49666 3460
rect 52546 3408 52552 3460
rect 52604 3448 52610 3460
rect 53650 3448 53656 3460
rect 52604 3420 53656 3448
rect 52604 3408 52610 3420
rect 53650 3408 53656 3420
rect 53708 3408 53714 3460
rect 56042 3408 56048 3460
rect 56100 3448 56106 3460
rect 56502 3448 56508 3460
rect 56100 3420 56508 3448
rect 56100 3408 56106 3420
rect 56502 3408 56508 3420
rect 56560 3408 56566 3460
rect 57238 3408 57244 3460
rect 57296 3448 57302 3460
rect 57882 3448 57888 3460
rect 57296 3420 57888 3448
rect 57296 3408 57302 3420
rect 57882 3408 57888 3420
rect 57940 3408 57946 3460
rect 58434 3408 58440 3460
rect 58492 3448 58498 3460
rect 59262 3448 59268 3460
rect 58492 3420 59268 3448
rect 58492 3408 58498 3420
rect 59262 3408 59268 3420
rect 59320 3408 59326 3460
rect 59630 3408 59636 3460
rect 59688 3448 59694 3460
rect 60642 3448 60648 3460
rect 59688 3420 60648 3448
rect 59688 3408 59694 3420
rect 60642 3408 60648 3420
rect 60700 3408 60706 3460
rect 64322 3408 64328 3460
rect 64380 3448 64386 3460
rect 64782 3448 64788 3460
rect 64380 3420 64788 3448
rect 64380 3408 64386 3420
rect 64782 3408 64788 3420
rect 64840 3408 64846 3460
rect 83274 3408 83280 3460
rect 83332 3448 83338 3460
rect 84102 3448 84108 3460
rect 83332 3420 84108 3448
rect 83332 3408 83338 3420
rect 84102 3408 84108 3420
rect 84160 3408 84166 3460
rect 93826 3420 103514 3448
rect 61378 3380 61384 3392
rect 45526 3352 61384 3380
rect 61378 3340 61384 3352
rect 61436 3340 61442 3392
rect 77386 3340 77392 3392
rect 77444 3380 77450 3392
rect 93826 3380 93854 3420
rect 77444 3352 93854 3380
rect 103486 3380 103514 3420
rect 105722 3408 105728 3460
rect 105780 3448 105786 3460
rect 106182 3448 106188 3460
rect 105780 3420 106188 3448
rect 105780 3408 105786 3420
rect 106182 3408 106188 3420
rect 106240 3408 106246 3460
rect 108114 3408 108120 3460
rect 108172 3448 108178 3460
rect 108942 3448 108948 3460
rect 108172 3420 108948 3448
rect 108172 3408 108178 3420
rect 108942 3408 108948 3420
rect 109000 3408 109006 3460
rect 109310 3408 109316 3460
rect 109368 3448 109374 3460
rect 110322 3448 110328 3460
rect 109368 3420 110328 3448
rect 109368 3408 109374 3420
rect 110322 3408 110328 3420
rect 110380 3408 110386 3460
rect 114002 3408 114008 3460
rect 114060 3448 114066 3460
rect 114462 3448 114468 3460
rect 114060 3420 114468 3448
rect 114060 3408 114066 3420
rect 114462 3408 114468 3420
rect 114520 3408 114526 3460
rect 115198 3408 115204 3460
rect 115256 3448 115262 3460
rect 115842 3448 115848 3460
rect 115256 3420 115848 3448
rect 115256 3408 115262 3420
rect 115842 3408 115848 3420
rect 115900 3408 115906 3460
rect 117590 3408 117596 3460
rect 117648 3448 117654 3460
rect 118602 3448 118608 3460
rect 117648 3420 118608 3448
rect 117648 3408 117654 3420
rect 118602 3408 118608 3420
rect 118660 3408 118666 3460
rect 118786 3408 118792 3460
rect 118844 3448 118850 3460
rect 119798 3448 119804 3460
rect 118844 3420 119804 3448
rect 118844 3408 118850 3420
rect 119798 3408 119804 3420
rect 119856 3408 119862 3460
rect 122282 3408 122288 3460
rect 122340 3448 122346 3460
rect 122742 3448 122748 3460
rect 122340 3420 122748 3448
rect 122340 3408 122346 3420
rect 122742 3408 122748 3420
rect 122800 3408 122806 3460
rect 123478 3408 123484 3460
rect 123536 3448 123542 3460
rect 187050 3448 187056 3460
rect 123536 3420 187056 3448
rect 123536 3408 123542 3420
rect 187050 3408 187056 3420
rect 187108 3408 187114 3460
rect 195238 3408 195244 3460
rect 195296 3448 195302 3460
rect 246390 3448 246396 3460
rect 195296 3420 246396 3448
rect 195296 3408 195302 3420
rect 246390 3408 246396 3420
rect 246448 3408 246454 3460
rect 288986 3408 288992 3460
rect 289044 3448 289050 3460
rect 296714 3448 296720 3460
rect 289044 3420 296720 3448
rect 289044 3408 289050 3420
rect 296714 3408 296720 3420
rect 296772 3408 296778 3460
rect 323578 3408 323584 3460
rect 323636 3448 323642 3460
rect 348050 3448 348056 3460
rect 323636 3420 348056 3448
rect 323636 3408 323642 3420
rect 348050 3408 348056 3420
rect 348108 3408 348114 3460
rect 350442 3408 350448 3460
rect 350500 3448 350506 3460
rect 360286 3448 360292 3460
rect 350500 3420 360292 3448
rect 350500 3408 350506 3420
rect 360286 3408 360292 3420
rect 360344 3408 360350 3460
rect 116578 3380 116584 3392
rect 103486 3352 116584 3380
rect 77444 3340 77450 3352
rect 116578 3340 116584 3352
rect 116636 3340 116642 3392
rect 582190 3272 582196 3324
rect 582248 3312 582254 3324
rect 583570 3312 583576 3324
rect 582248 3284 583576 3312
rect 582248 3272 582254 3284
rect 583570 3272 583576 3284
rect 583628 3272 583634 3324
rect 74994 3204 75000 3256
rect 75052 3244 75058 3256
rect 75822 3244 75828 3256
rect 75052 3216 75828 3244
rect 75052 3204 75058 3216
rect 75822 3204 75828 3216
rect 75880 3204 75886 3256
rect 268378 3136 268384 3188
rect 268436 3176 268442 3188
rect 276014 3176 276020 3188
rect 268436 3148 276020 3176
rect 268436 3136 268442 3148
rect 276014 3136 276020 3148
rect 276072 3136 276078 3188
rect 280798 3136 280804 3188
rect 280856 3176 280862 3188
rect 283098 3176 283104 3188
rect 280856 3148 283104 3176
rect 280856 3136 280862 3148
rect 283098 3136 283104 3148
rect 283156 3136 283162 3188
rect 337378 3136 337384 3188
rect 337436 3176 337442 3188
rect 339862 3176 339868 3188
rect 337436 3148 339868 3176
rect 337436 3136 337442 3148
rect 339862 3136 339868 3148
rect 339920 3136 339926 3188
rect 11146 3000 11152 3052
rect 11204 3040 11210 3052
rect 15838 3040 15844 3052
rect 11204 3012 15844 3040
rect 11204 3000 11210 3012
rect 15838 3000 15844 3012
rect 15896 3000 15902 3052
rect 50154 3000 50160 3052
rect 50212 3040 50218 3052
rect 50890 3040 50896 3052
rect 50212 3012 50896 3040
rect 50212 3000 50218 3012
rect 50890 3000 50896 3012
rect 50948 3000 50954 3052
rect 82078 3000 82084 3052
rect 82136 3040 82142 3052
rect 82722 3040 82728 3052
rect 82136 3012 82728 3040
rect 82136 3000 82142 3012
rect 82722 3000 82728 3012
rect 82780 3000 82786 3052
rect 110506 3000 110512 3052
rect 110564 3040 110570 3052
rect 111518 3040 111524 3052
rect 110564 3012 111524 3040
rect 110564 3000 110570 3012
rect 111518 3000 111524 3012
rect 111576 3000 111582 3052
rect 19426 2932 19432 2984
rect 19484 2972 19490 2984
rect 20622 2972 20628 2984
rect 19484 2944 20628 2972
rect 19484 2932 19490 2944
rect 20622 2932 20628 2944
rect 20680 2932 20686 2984
rect 309870 2932 309876 2984
rect 309928 2972 309934 2984
rect 315022 2972 315028 2984
rect 309928 2944 315028 2972
rect 309928 2932 309934 2944
rect 315022 2932 315028 2944
rect 315080 2932 315086 2984
rect 112806 2116 112812 2168
rect 112864 2156 112870 2168
rect 218698 2156 218704 2168
rect 112864 2128 218704 2156
rect 112864 2116 112870 2128
rect 218698 2116 218704 2128
rect 218756 2116 218762 2168
rect 220170 2116 220176 2168
rect 220228 2156 220234 2168
rect 240502 2156 240508 2168
rect 220228 2128 240508 2156
rect 220228 2116 220234 2128
rect 240502 2116 240508 2128
rect 240560 2116 240566 2168
rect 51350 2048 51356 2100
rect 51408 2088 51414 2100
rect 58618 2088 58624 2100
rect 51408 2060 58624 2088
rect 51408 2048 51414 2060
rect 58618 2048 58624 2060
rect 58676 2048 58682 2100
rect 65518 2048 65524 2100
rect 65576 2088 65582 2100
rect 233970 2088 233976 2100
rect 65576 2060 233976 2088
rect 65576 2048 65582 2060
rect 233970 2048 233976 2060
rect 234028 2048 234034 2100
rect 253198 2048 253204 2100
rect 253256 2088 253262 2100
rect 272426 2088 272432 2100
rect 253256 2060 272432 2088
rect 253256 2048 253262 2060
rect 272426 2048 272432 2060
rect 272484 2048 272490 2100
rect 331858 2048 331864 2100
rect 331916 2088 331922 2100
rect 340966 2088 340972 2100
rect 331916 2060 340972 2088
rect 331916 2048 331922 2060
rect 340966 2048 340972 2060
rect 341024 2048 341030 2100
rect 332594 552 332600 604
rect 332652 592 332658 604
rect 333882 592 333888 604
rect 332652 564 333888 592
rect 332652 552 332658 564
rect 333882 552 333888 564
rect 333940 552 333946 604
<< via1 >>
rect 331220 702992 331272 703044
rect 332508 702992 332560 703044
rect 170312 702924 170364 702976
rect 281540 702924 281592 702976
rect 62028 702856 62080 702908
rect 267648 702856 267700 702908
rect 276020 702856 276072 702908
rect 478512 702856 478564 702908
rect 202788 702788 202840 702840
rect 273260 702788 273312 702840
rect 349804 702788 349856 702840
rect 494796 702788 494848 702840
rect 233884 702720 233936 702772
rect 397368 702720 397420 702772
rect 197268 702652 197320 702704
rect 364984 702652 365036 702704
rect 382924 702652 382976 702704
rect 462320 702652 462372 702704
rect 95148 702584 95200 702636
rect 300124 702584 300176 702636
rect 300768 702584 300820 702636
rect 363604 702584 363656 702636
rect 543464 702584 543516 702636
rect 86868 702516 86920 702568
rect 235172 702516 235224 702568
rect 264244 702516 264296 702568
rect 559656 702516 559708 702568
rect 8116 702448 8168 702500
rect 88800 702448 88852 702500
rect 99288 702448 99340 702500
rect 527180 702448 527232 702500
rect 129648 700340 129700 700392
rect 137836 700340 137888 700392
rect 68284 700272 68336 700324
rect 105452 700272 105504 700324
rect 130384 700272 130436 700324
rect 218980 700272 219032 700324
rect 283840 700272 283892 700324
rect 295340 700272 295392 700324
rect 300768 700272 300820 700324
rect 360200 700272 360252 700324
rect 374644 700272 374696 700324
rect 429844 700272 429896 700324
rect 24308 699660 24360 699712
rect 25504 699660 25556 699712
rect 65800 699660 65852 699712
rect 72976 699660 73028 699712
rect 87604 699660 87656 699712
rect 89168 699660 89220 699712
rect 327724 698912 327776 698964
rect 348792 698912 348844 698964
rect 3424 683136 3476 683188
rect 11704 683136 11756 683188
rect 3516 670692 3568 670744
rect 14464 670692 14516 670744
rect 3424 658112 3476 658164
rect 7564 658112 7616 658164
rect 3424 632068 3476 632120
rect 17224 632068 17276 632120
rect 3148 618264 3200 618316
rect 15844 618264 15896 618316
rect 3240 605820 3292 605872
rect 90364 605820 90416 605872
rect 74632 598952 74684 599004
rect 98644 598952 98696 599004
rect 349160 598884 349212 598936
rect 349804 598884 349856 598936
rect 70308 597524 70360 597576
rect 349160 597524 349212 597576
rect 67456 596776 67508 596828
rect 170404 596776 170456 596828
rect 86868 594872 86920 594924
rect 113180 594872 113232 594924
rect 65984 594804 66036 594856
rect 295340 594804 295392 594856
rect 295984 594804 296036 594856
rect 90364 594396 90416 594448
rect 91100 594396 91152 594448
rect 40040 594056 40092 594108
rect 89812 594056 89864 594108
rect 73988 593376 74040 593428
rect 116584 593376 116636 593428
rect 25504 592628 25556 592680
rect 80336 592628 80388 592680
rect 75644 592084 75696 592136
rect 96620 592084 96672 592136
rect 84108 592016 84160 592068
rect 112536 592016 112588 592068
rect 7564 591268 7616 591320
rect 69112 591268 69164 591320
rect 70124 590724 70176 590776
rect 73160 590724 73212 590776
rect 86776 590724 86828 590776
rect 115296 590724 115348 590776
rect 69112 590656 69164 590708
rect 70400 590656 70452 590708
rect 73068 590656 73120 590708
rect 81716 590656 81768 590708
rect 85028 590656 85080 590708
rect 86868 590656 86920 590708
rect 86224 590588 86276 590640
rect 204260 590656 204312 590708
rect 70400 589908 70452 589960
rect 89076 589908 89128 589960
rect 100760 589908 100812 589960
rect 111064 589908 111116 589960
rect 3424 589296 3476 589348
rect 74908 589296 74960 589348
rect 75644 589296 75696 589348
rect 76748 589296 76800 589348
rect 100760 589296 100812 589348
rect 187608 589296 187660 589348
rect 255964 589296 256016 589348
rect 79784 588480 79836 588532
rect 72424 588412 72476 588464
rect 72884 588412 72936 588464
rect 80704 588412 80756 588464
rect 89168 588412 89220 588464
rect 55036 587868 55088 587920
rect 66812 587868 66864 587920
rect 105544 587868 105596 587920
rect 93124 587664 93176 587716
rect 88892 587392 88944 587444
rect 88892 587120 88944 587172
rect 89168 586576 89220 586628
rect 106924 586576 106976 586628
rect 59084 586508 59136 586560
rect 66260 586508 66312 586560
rect 91744 586508 91796 586560
rect 95240 586508 95292 586560
rect 57888 585148 57940 585200
rect 66812 585148 66864 585200
rect 67548 585148 67600 585200
rect 68284 585148 68336 585200
rect 91376 584400 91428 584452
rect 95148 584400 95200 584452
rect 132500 584400 132552 584452
rect 91192 583652 91244 583704
rect 99288 583652 99340 583704
rect 104164 583652 104216 583704
rect 48136 582360 48188 582412
rect 66812 582360 66864 582412
rect 64696 581000 64748 581052
rect 66444 581000 66496 581052
rect 91744 581000 91796 581052
rect 142804 581000 142856 581052
rect 52276 579640 52328 579692
rect 66812 579640 66864 579692
rect 91744 579640 91796 579692
rect 108304 579640 108356 579692
rect 91744 578212 91796 578264
rect 120724 578212 120776 578264
rect 17224 576104 17276 576156
rect 67364 576104 67416 576156
rect 91100 576104 91152 576156
rect 123024 576104 123076 576156
rect 61844 574064 61896 574116
rect 67088 574064 67140 574116
rect 91100 574064 91152 574116
rect 97264 574064 97316 574116
rect 60648 571344 60700 571396
rect 66812 571344 66864 571396
rect 91100 571344 91152 571396
rect 115204 571344 115256 571396
rect 149704 571344 149756 571396
rect 266360 571344 266412 571396
rect 91100 569984 91152 570036
rect 94504 569984 94556 570036
rect 93124 569916 93176 569968
rect 353300 569916 353352 569968
rect 67364 569848 67416 569900
rect 68284 569848 68336 569900
rect 91192 569168 91244 569220
rect 126980 569168 127032 569220
rect 63316 568556 63368 568608
rect 66812 568556 66864 568608
rect 91100 568556 91152 568608
rect 100024 568556 100076 568608
rect 126980 568556 127032 568608
rect 213920 568556 213972 568608
rect 273260 567672 273312 567724
rect 273904 567672 273956 567724
rect 64788 567196 64840 567248
rect 66720 567196 66772 567248
rect 89812 567196 89864 567248
rect 133880 567264 133932 567316
rect 209044 567264 209096 567316
rect 197176 567196 197228 567248
rect 273260 567196 273312 567248
rect 53104 566448 53156 566500
rect 67456 566448 67508 566500
rect 94504 566448 94556 566500
rect 137100 566448 137152 566500
rect 3424 565836 3476 565888
rect 43444 565836 43496 565888
rect 91376 565836 91428 565888
rect 102784 565836 102836 565888
rect 136640 565836 136692 565888
rect 137100 565836 137152 565888
rect 291200 565836 291252 565888
rect 177304 564476 177356 564528
rect 259460 564476 259512 564528
rect 50896 564408 50948 564460
rect 66812 564408 66864 564460
rect 91376 564408 91428 564460
rect 107016 564408 107068 564460
rect 115296 564408 115348 564460
rect 117964 564408 118016 564460
rect 166816 564408 166868 564460
rect 298100 564408 298152 564460
rect 195888 563116 195940 563168
rect 271880 563116 271932 563168
rect 50988 563048 51040 563100
rect 66812 563048 66864 563100
rect 91376 563048 91428 563100
rect 134708 563048 134760 563100
rect 206284 563048 206336 563100
rect 582840 563048 582892 563100
rect 52368 561688 52420 561740
rect 66812 561688 66864 561740
rect 111064 561688 111116 561740
rect 111708 561688 111760 561740
rect 358912 561688 358964 561740
rect 263600 561620 263652 561672
rect 264244 561620 264296 561672
rect 197084 560328 197136 560380
rect 288440 560328 288492 560380
rect 41328 560260 41380 560312
rect 66812 560260 66864 560312
rect 146944 560260 146996 560312
rect 263600 560260 263652 560312
rect 192484 558968 192536 559020
rect 287060 558968 287112 559020
rect 63408 558900 63460 558952
rect 66812 558900 66864 558952
rect 89628 558900 89680 558952
rect 122104 558900 122156 558952
rect 160008 558900 160060 558952
rect 309140 558900 309192 558952
rect 59176 558424 59228 558476
rect 62028 558424 62080 558476
rect 97264 558152 97316 558204
rect 122932 558152 122984 558204
rect 198832 558152 198884 558204
rect 331220 558152 331272 558204
rect 62028 557540 62080 557592
rect 66812 557540 66864 557592
rect 195428 557540 195480 557592
rect 357440 557540 357492 557592
rect 92388 556792 92440 556844
rect 152464 556792 152516 556844
rect 204260 556792 204312 556844
rect 582380 556792 582432 556844
rect 91192 556180 91244 556232
rect 121460 556180 121512 556232
rect 181536 556180 181588 556232
rect 251824 556180 251876 556232
rect 324320 555228 324372 555280
rect 324872 555228 324924 555280
rect 327724 555228 327776 555280
rect 187056 554820 187108 554872
rect 324320 554820 324372 554872
rect 53656 554752 53708 554804
rect 66812 554752 66864 554804
rect 91744 554752 91796 554804
rect 106188 554752 106240 554804
rect 244924 554752 244976 554804
rect 49608 554004 49660 554056
rect 65984 554004 66036 554056
rect 66536 554004 66588 554056
rect 198556 554004 198608 554056
rect 583024 554004 583076 554056
rect 91744 553392 91796 553444
rect 112444 553392 112496 553444
rect 188344 553392 188396 553444
rect 270500 553392 270552 553444
rect 91744 552100 91796 552152
rect 97356 552100 97408 552152
rect 193864 552100 193916 552152
rect 296720 552100 296772 552152
rect 91192 552032 91244 552084
rect 100116 552032 100168 552084
rect 112536 552032 112588 552084
rect 226984 552032 227036 552084
rect 198648 551284 198700 551336
rect 582748 551284 582800 551336
rect 91192 550604 91244 550656
rect 108948 550604 109000 550656
rect 124864 550604 124916 550656
rect 180156 550604 180208 550656
rect 229100 550604 229152 550656
rect 295984 549856 296036 549908
rect 351920 549856 351972 549908
rect 161388 549312 161440 549364
rect 215392 549312 215444 549364
rect 56508 549244 56560 549296
rect 66444 549244 66496 549296
rect 189816 549244 189868 549296
rect 305000 549244 305052 549296
rect 180064 547952 180116 548004
rect 285128 547952 285180 548004
rect 59268 547884 59320 547936
rect 66444 547884 66496 547936
rect 91468 547884 91520 547936
rect 95332 547884 95384 547936
rect 184204 547884 184256 547936
rect 343640 547884 343692 547936
rect 95332 547136 95384 547188
rect 245660 547136 245712 547188
rect 91192 546456 91244 546508
rect 97264 546456 97316 546508
rect 126888 546456 126940 546508
rect 339960 546456 340012 546508
rect 185584 545164 185636 545216
rect 220820 545164 220872 545216
rect 48228 545096 48280 545148
rect 66812 545096 66864 545148
rect 91192 545096 91244 545148
rect 94504 545096 94556 545148
rect 188436 545096 188488 545148
rect 290096 545096 290148 545148
rect 328460 545096 328512 545148
rect 375472 545096 375524 545148
rect 194140 543804 194192 543856
rect 223672 543804 223724 543856
rect 330024 543804 330076 543856
rect 364432 543804 364484 543856
rect 55128 543736 55180 543788
rect 66812 543736 66864 543788
rect 91836 543736 91888 543788
rect 93676 543736 93728 543788
rect 284300 543736 284352 543788
rect 311900 543736 311952 543788
rect 356244 543736 356296 543788
rect 11704 542988 11756 543040
rect 36544 542988 36596 543040
rect 166908 542444 166960 542496
rect 306656 542444 306708 542496
rect 338304 542444 338356 542496
rect 363052 542444 363104 542496
rect 36544 542376 36596 542428
rect 37188 542376 37240 542428
rect 66812 542376 66864 542428
rect 91192 542376 91244 542428
rect 98736 542376 98788 542428
rect 195244 542376 195296 542428
rect 356152 542376 356204 542428
rect 209044 542308 209096 542360
rect 210424 542308 210476 542360
rect 244924 542308 244976 542360
rect 247040 542308 247092 542360
rect 14464 541628 14516 541680
rect 67088 541628 67140 541680
rect 67364 541628 67416 541680
rect 91192 541628 91244 541680
rect 128360 541628 128412 541680
rect 199476 541628 199528 541680
rect 204260 541628 204312 541680
rect 207020 541628 207072 541680
rect 331680 541016 331732 541068
rect 360292 541016 360344 541068
rect 128360 540948 128412 541000
rect 129648 540948 129700 541000
rect 258448 540948 258500 541000
rect 316592 540948 316644 541000
rect 364524 540948 364576 541000
rect 3424 540200 3476 540252
rect 67272 539724 67324 539776
rect 61936 539588 61988 539640
rect 67548 539588 67600 539640
rect 70400 539588 70452 539640
rect 71872 539588 71924 539640
rect 88156 539588 88208 539640
rect 92388 539588 92440 539640
rect 93216 539588 93268 539640
rect 129648 539656 129700 539708
rect 357532 539656 357584 539708
rect 250628 539588 250680 539640
rect 347688 539588 347740 539640
rect 580264 539588 580316 539640
rect 67456 539520 67508 539572
rect 273904 539520 273956 539572
rect 275652 539520 275704 539572
rect 278044 539520 278096 539572
rect 278964 539520 279016 539572
rect 270868 539452 270920 539504
rect 273996 539452 274048 539504
rect 67456 539316 67508 539368
rect 57796 538908 57848 538960
rect 65800 538908 65852 538960
rect 65984 538908 66036 538960
rect 175924 538908 175976 538960
rect 194140 538908 194192 538960
rect 3424 538840 3476 538892
rect 89720 538840 89772 538892
rect 157984 538840 158036 538892
rect 195244 538840 195296 538892
rect 199384 538296 199436 538348
rect 255596 538296 255648 538348
rect 347044 538296 347096 538348
rect 359096 538296 359148 538348
rect 65984 538228 66036 538280
rect 76748 538228 76800 538280
rect 195244 538228 195296 538280
rect 216680 538228 216732 538280
rect 220912 538228 220964 538280
rect 356336 538228 356388 538280
rect 88616 538160 88668 538212
rect 89628 538160 89680 538212
rect 86868 538092 86920 538144
rect 130384 538160 130436 538212
rect 8208 537480 8260 537532
rect 91284 537480 91336 537532
rect 198096 537480 198148 537532
rect 220912 537480 220964 537532
rect 323676 537480 323728 537532
rect 580172 537480 580224 537532
rect 178776 536800 178828 536852
rect 233884 536800 233936 536852
rect 234068 536800 234120 536852
rect 337108 536800 337160 536852
rect 371332 536800 371384 536852
rect 43444 536732 43496 536784
rect 69572 536732 69624 536784
rect 75184 536732 75236 536784
rect 129648 536732 129700 536784
rect 84292 536460 84344 536512
rect 89076 536460 89128 536512
rect 15844 536052 15896 536104
rect 43996 536052 44048 536104
rect 73160 536052 73212 536104
rect 81532 535576 81584 535628
rect 83464 535576 83516 535628
rect 198740 535576 198792 535628
rect 200396 535576 200448 535628
rect 130476 535508 130528 535560
rect 308404 535508 308456 535560
rect 327448 535508 327500 535560
rect 361672 535508 361724 535560
rect 89628 535440 89680 535492
rect 90456 535440 90508 535492
rect 201408 535440 201460 535492
rect 208676 535440 208728 535492
rect 247592 535440 247644 535492
rect 582380 535440 582432 535492
rect 175188 534760 175240 534812
rect 202052 535236 202104 535288
rect 11704 534692 11756 534744
rect 91192 534692 91244 534744
rect 67732 534012 67784 534064
rect 76564 534012 76616 534064
rect 164148 533332 164200 533384
rect 191196 533332 191248 533384
rect 77852 532788 77904 532840
rect 100944 532788 100996 532840
rect 48136 532720 48188 532772
rect 162860 532720 162912 532772
rect 164148 532720 164200 532772
rect 100944 532652 100996 532704
rect 197360 532652 197412 532704
rect 17868 531972 17920 532024
rect 91100 531972 91152 532024
rect 358728 531972 358780 532024
rect 358912 531972 358964 532024
rect 582748 531972 582800 532024
rect 41328 531224 41380 531276
rect 195428 531224 195480 531276
rect 64696 530544 64748 530596
rect 79324 530544 79376 530596
rect 177396 529864 177448 529916
rect 197360 529864 197412 529916
rect 59084 529252 59136 529304
rect 85580 529252 85632 529304
rect 80060 529184 80112 529236
rect 129740 529184 129792 529236
rect 129740 528572 129792 528624
rect 177304 528572 177356 528624
rect 124864 528504 124916 528556
rect 197360 528504 197412 528556
rect 70492 527484 70544 527536
rect 71044 527484 71096 527536
rect 71044 527144 71096 527196
rect 124956 527144 125008 527196
rect 358728 527144 358780 527196
rect 367100 527144 367152 527196
rect 34428 525036 34480 525088
rect 198004 525036 198056 525088
rect 358728 524424 358780 524476
rect 378232 524424 378284 524476
rect 66904 523676 66956 523728
rect 188436 523676 188488 523728
rect 189724 522248 189776 522300
rect 197452 522248 197504 522300
rect 358728 522248 358780 522300
rect 582380 522248 582432 522300
rect 147588 521636 147640 521688
rect 197360 521636 197412 521688
rect 46848 520888 46900 520940
rect 195336 520888 195388 520940
rect 56508 520208 56560 520260
rect 189816 520208 189868 520260
rect 357900 520004 357952 520056
rect 360200 520004 360252 520056
rect 162124 518916 162176 518968
rect 197360 518916 197412 518968
rect 39948 518168 40000 518220
rect 184388 518168 184440 518220
rect 66168 517420 66220 517472
rect 187056 517420 187108 517472
rect 176016 516128 176068 516180
rect 197360 516128 197412 516180
rect 358728 516128 358780 516180
rect 375380 516128 375432 516180
rect 2780 514768 2832 514820
rect 4804 514768 4856 514820
rect 358636 514768 358688 514820
rect 360200 514768 360252 514820
rect 45468 514020 45520 514072
rect 191104 514020 191156 514072
rect 156604 512592 156656 512644
rect 199476 512592 199528 512644
rect 124956 510552 125008 510604
rect 197360 510552 197412 510604
rect 169024 506472 169076 506524
rect 197360 506472 197412 506524
rect 357624 505724 357676 505776
rect 367192 505724 367244 505776
rect 358728 505112 358780 505164
rect 385040 505112 385092 505164
rect 358728 502324 358780 502376
rect 369952 502324 370004 502376
rect 3516 502256 3568 502308
rect 11704 502256 11756 502308
rect 177304 500896 177356 500948
rect 197360 500896 197412 500948
rect 358728 499536 358780 499588
rect 371424 499536 371476 499588
rect 356336 496748 356388 496800
rect 357164 496748 357216 496800
rect 582932 496748 582984 496800
rect 188436 495456 188488 495508
rect 197360 495456 197412 495508
rect 358636 493960 358688 494012
rect 412640 493960 412692 494012
rect 130384 492668 130436 492720
rect 197360 492668 197412 492720
rect 152556 489880 152608 489932
rect 197360 489880 197412 489932
rect 152464 487772 152516 487824
rect 180800 487772 180852 487824
rect 182088 487772 182140 487824
rect 182088 487160 182140 487212
rect 197360 487160 197412 487212
rect 358728 487160 358780 487212
rect 372620 487160 372672 487212
rect 358728 484372 358780 484424
rect 369860 484372 369912 484424
rect 191104 480428 191156 480480
rect 197360 480428 197412 480480
rect 116584 478116 116636 478168
rect 128452 478116 128504 478168
rect 128452 477504 128504 477556
rect 176660 477504 176712 477556
rect 197360 477504 197412 477556
rect 358728 477504 358780 477556
rect 362960 477504 363012 477556
rect 147128 476756 147180 476808
rect 198096 476756 198148 476808
rect 68284 476076 68336 476128
rect 68928 476076 68980 476128
rect 147128 476076 147180 476128
rect 147496 476076 147548 476128
rect 3332 475328 3384 475380
rect 8208 475328 8260 475380
rect 25504 475328 25556 475380
rect 144184 474716 144236 474768
rect 197360 474716 197412 474768
rect 358728 474716 358780 474768
rect 375564 474716 375616 474768
rect 140044 473356 140096 473408
rect 197360 473356 197412 473408
rect 358728 471996 358780 472048
rect 368572 471996 368624 472048
rect 195796 470704 195848 470756
rect 197636 470704 197688 470756
rect 358728 470568 358780 470620
rect 380900 470568 380952 470620
rect 165528 467848 165580 467900
rect 197360 467848 197412 467900
rect 358728 467848 358780 467900
rect 363144 467848 363196 467900
rect 105544 467780 105596 467832
rect 187516 467780 187568 467832
rect 191196 467780 191248 467832
rect 62028 467100 62080 467152
rect 95240 467100 95292 467152
rect 104900 466420 104952 466472
rect 105544 466420 105596 466472
rect 60464 465672 60516 465724
rect 78772 465672 78824 465724
rect 124956 465060 125008 465112
rect 171048 465060 171100 465112
rect 197360 465060 197412 465112
rect 356336 465060 356388 465112
rect 356796 465060 356848 465112
rect 582380 465060 582432 465112
rect 358084 464992 358136 465044
rect 365720 464992 365772 465044
rect 106188 464312 106240 464364
rect 120816 464312 120868 464364
rect 64788 463700 64840 463752
rect 180248 463700 180300 463752
rect 93768 462952 93820 463004
rect 107660 462952 107712 463004
rect 3516 462340 3568 462392
rect 14556 462340 14608 462392
rect 127624 462340 127676 462392
rect 197360 462340 197412 462392
rect 358728 462340 358780 462392
rect 385132 462340 385184 462392
rect 59084 461660 59136 461712
rect 72424 461660 72476 461712
rect 52276 461592 52328 461644
rect 78036 461592 78088 461644
rect 76012 461456 76064 461508
rect 76564 461456 76616 461508
rect 76564 460912 76616 460964
rect 173900 460912 173952 460964
rect 65984 460164 66036 460216
rect 77944 460164 77996 460216
rect 143448 460164 143500 460216
rect 197360 460164 197412 460216
rect 370044 460164 370096 460216
rect 582564 460164 582616 460216
rect 142804 459552 142856 459604
rect 143448 459552 143500 459604
rect 358452 459552 358504 459604
rect 370044 459552 370096 459604
rect 4804 459484 4856 459536
rect 112536 459484 112588 459536
rect 64788 458804 64840 458856
rect 73252 458804 73304 458856
rect 131764 458192 131816 458244
rect 197360 458192 197412 458244
rect 108304 458124 108356 458176
rect 115296 458124 115348 458176
rect 52276 456764 52328 456816
rect 67640 456764 67692 456816
rect 68836 456764 68888 456816
rect 63316 456016 63368 456068
rect 67640 456016 67692 456068
rect 68652 456016 68704 456068
rect 68836 456016 68888 456068
rect 81440 456016 81492 456068
rect 68652 455404 68704 455456
rect 185676 455404 185728 455456
rect 358728 455404 358780 455456
rect 387800 455404 387852 455456
rect 582840 455404 582892 455456
rect 55036 455336 55088 455388
rect 56416 455336 56468 455388
rect 63316 454656 63368 454708
rect 75920 454656 75972 454708
rect 102784 454656 102836 454708
rect 125600 454656 125652 454708
rect 56416 454044 56468 454096
rect 87052 454044 87104 454096
rect 17224 453976 17276 454028
rect 17868 453976 17920 454028
rect 65616 453296 65668 453348
rect 75184 453296 75236 453348
rect 17224 452616 17276 452668
rect 124220 452616 124272 452668
rect 358728 452616 358780 452668
rect 376760 452616 376812 452668
rect 3424 451868 3476 451920
rect 121552 451868 121604 451920
rect 124956 451868 125008 451920
rect 116124 451256 116176 451308
rect 156604 451256 156656 451308
rect 66076 450576 66128 450628
rect 91100 450576 91152 450628
rect 48136 450508 48188 450560
rect 80888 450508 80940 450560
rect 96252 450508 96304 450560
rect 128452 450508 128504 450560
rect 91100 449896 91152 449948
rect 91560 449896 91612 449948
rect 159456 449896 159508 449948
rect 358728 449896 358780 449948
rect 364340 449896 364392 449948
rect 106924 449828 106976 449880
rect 131764 449828 131816 449880
rect 115204 449352 115256 449404
rect 120632 449352 120684 449404
rect 57704 449216 57756 449268
rect 78680 449216 78732 449268
rect 14556 449148 14608 449200
rect 68836 449148 68888 449200
rect 368388 449148 368440 449200
rect 582472 449148 582524 449200
rect 3148 448536 3200 448588
rect 14464 448536 14516 448588
rect 68836 448536 68888 448588
rect 103520 448536 103572 448588
rect 103704 448536 103756 448588
rect 168288 448536 168340 448588
rect 197360 448536 197412 448588
rect 358728 448536 358780 448588
rect 367284 448536 367336 448588
rect 368388 448536 368440 448588
rect 57888 447788 57940 447840
rect 83832 447788 83884 447840
rect 94780 447788 94832 447840
rect 127624 447788 127676 447840
rect 164884 447788 164936 447840
rect 192576 447788 192628 447840
rect 65892 447108 65944 447160
rect 71044 447108 71096 447160
rect 88892 447108 88944 447160
rect 132592 447108 132644 447160
rect 68928 447040 68980 447092
rect 73160 447040 73212 447092
rect 79324 447040 79376 447092
rect 130476 447040 130528 447092
rect 48044 446360 48096 446412
rect 71872 446360 71924 446412
rect 74816 446360 74868 446412
rect 90364 445748 90416 445800
rect 96528 445748 96580 445800
rect 100852 445748 100904 445800
rect 102232 445748 102284 445800
rect 112536 445748 112588 445800
rect 112904 445748 112956 445800
rect 142896 445748 142948 445800
rect 144276 445748 144328 445800
rect 197360 445748 197412 445800
rect 60556 444456 60608 444508
rect 93032 444456 93084 444508
rect 100760 444456 100812 444508
rect 127624 444456 127676 444508
rect 4804 444388 4856 444440
rect 118700 444388 118752 444440
rect 119160 444388 119212 444440
rect 121644 444388 121696 444440
rect 147496 444320 147548 444372
rect 148324 444320 148376 444372
rect 168380 443640 168432 443692
rect 184296 443640 184348 443692
rect 184388 443640 184440 443692
rect 197360 443640 197412 443692
rect 125508 442960 125560 443012
rect 168380 442960 168432 443012
rect 358728 442960 358780 443012
rect 383660 442960 383712 443012
rect 67364 442892 67416 442944
rect 67824 442892 67876 442944
rect 124128 442008 124180 442060
rect 131764 442008 131816 442060
rect 185676 441532 185728 441584
rect 197360 441532 197412 441584
rect 358728 440240 358780 440292
rect 368480 440240 368532 440292
rect 67364 438880 67416 438932
rect 67640 438880 67692 438932
rect 358728 438880 358780 438932
rect 361764 438880 361816 438932
rect 64696 438812 64748 438864
rect 66812 438812 66864 438864
rect 124128 438200 124180 438252
rect 132500 438200 132552 438252
rect 133144 438200 133196 438252
rect 126244 438132 126296 438184
rect 152556 438132 152608 438184
rect 50804 436092 50856 436144
rect 358728 436092 358780 436144
rect 379520 436092 379572 436144
rect 53104 436024 53156 436076
rect 66720 436024 66772 436076
rect 192576 433304 192628 433356
rect 197360 433304 197412 433356
rect 358728 433304 358780 433356
rect 380992 433304 381044 433356
rect 50896 433236 50948 433288
rect 54944 433236 54996 433288
rect 124128 432556 124180 432608
rect 142804 432556 142856 432608
rect 54944 431944 54996 431996
rect 66812 431944 66864 431996
rect 124128 431876 124180 431928
rect 124312 431876 124364 431928
rect 169116 431876 169168 431928
rect 50988 431196 51040 431248
rect 64696 431196 64748 431248
rect 66812 431196 66864 431248
rect 358728 430584 358780 430636
rect 376852 430584 376904 430636
rect 51080 429088 51132 429140
rect 52368 429088 52420 429140
rect 66812 429088 66864 429140
rect 122748 429088 122800 429140
rect 173164 429088 173216 429140
rect 22744 428408 22796 428460
rect 51080 428408 51132 428460
rect 178684 427796 178736 427848
rect 197360 427796 197412 427848
rect 358728 427796 358780 427848
rect 372712 427796 372764 427848
rect 356704 426776 356756 426828
rect 357532 426776 357584 426828
rect 152464 426436 152516 426488
rect 197360 426436 197412 426488
rect 41328 425688 41380 425740
rect 60740 425688 60792 425740
rect 60740 425076 60792 425128
rect 61844 425076 61896 425128
rect 66720 425076 66772 425128
rect 58900 423648 58952 423700
rect 63408 423648 63460 423700
rect 66812 423648 66864 423700
rect 178868 423648 178920 423700
rect 197360 423648 197412 423700
rect 358728 423648 358780 423700
rect 364616 423648 364668 423700
rect 374000 423648 374052 423700
rect 3424 423580 3476 423632
rect 17224 423580 17276 423632
rect 50988 421540 51040 421592
rect 59176 421540 59228 421592
rect 66260 421540 66312 421592
rect 122932 421540 122984 421592
rect 148968 421540 149020 421592
rect 178776 421540 178828 421592
rect 358728 420928 358780 420980
rect 370136 420928 370188 420980
rect 124128 420860 124180 420912
rect 159364 420860 159416 420912
rect 358728 418208 358780 418260
rect 365812 418208 365864 418260
rect 177304 418140 177356 418192
rect 197360 418140 197412 418192
rect 121184 415352 121236 415404
rect 126980 415352 127032 415404
rect 49608 415284 49660 415336
rect 53656 415284 53708 415336
rect 53656 413992 53708 414044
rect 66812 413992 66864 414044
rect 185676 413992 185728 414044
rect 197360 413992 197412 414044
rect 358728 413992 358780 414044
rect 367376 413992 367428 414044
rect 123852 413244 123904 413296
rect 136640 413244 136692 413296
rect 58992 411272 59044 411324
rect 66904 411272 66956 411324
rect 123576 411272 123628 411324
rect 151084 411272 151136 411324
rect 164148 411272 164200 411324
rect 197360 411272 197412 411324
rect 358728 411272 358780 411324
rect 389180 411272 389232 411324
rect 124864 409776 124916 409828
rect 197360 409776 197412 409828
rect 358728 408552 358780 408604
rect 365904 408552 365956 408604
rect 124128 407872 124180 407924
rect 133880 407872 133932 407924
rect 134616 407872 134668 407924
rect 122104 407056 122156 407108
rect 123024 407056 123076 407108
rect 124128 406172 124180 406224
rect 125508 406172 125560 406224
rect 59268 405764 59320 405816
rect 64604 405764 64656 405816
rect 66260 405764 66312 405816
rect 133236 405696 133288 405748
rect 197360 405696 197412 405748
rect 57888 403588 57940 403640
rect 66260 403588 66312 403640
rect 142896 403588 142948 403640
rect 167000 403588 167052 403640
rect 358728 403520 358780 403572
rect 363236 403520 363288 403572
rect 123760 403384 123812 403436
rect 124864 403384 124916 403436
rect 194048 401616 194100 401668
rect 197360 401616 197412 401668
rect 358728 401616 358780 401668
rect 378140 401616 378192 401668
rect 44088 401548 44140 401600
rect 48228 401548 48280 401600
rect 66260 401548 66312 401600
rect 124128 400868 124180 400920
rect 193220 400868 193272 400920
rect 193220 400188 193272 400240
rect 194140 400188 194192 400240
rect 60004 399440 60056 399492
rect 66260 399440 66312 399492
rect 124128 399440 124180 399492
rect 189908 399440 189960 399492
rect 187056 398828 187108 398880
rect 197360 398828 197412 398880
rect 357992 398828 358044 398880
rect 360476 398828 360528 398880
rect 2780 398692 2832 398744
rect 4804 398692 4856 398744
rect 48228 398080 48280 398132
rect 55128 398080 55180 398132
rect 60004 398080 60056 398132
rect 130476 397468 130528 397520
rect 187056 397468 187108 397520
rect 37188 396720 37240 396772
rect 66996 396720 67048 396772
rect 67272 396720 67324 396772
rect 133144 396720 133196 396772
rect 171140 396720 171192 396772
rect 169668 396040 169720 396092
rect 197360 396040 197412 396092
rect 358728 396040 358780 396092
rect 361856 396040 361908 396092
rect 124128 395292 124180 395344
rect 188528 395292 188580 395344
rect 191656 394680 191708 394732
rect 197360 394680 197412 394732
rect 134524 393320 134576 393372
rect 198464 393320 198516 393372
rect 61936 392028 61988 392080
rect 66168 392028 66220 392080
rect 66628 392028 66680 392080
rect 121460 392028 121512 392080
rect 153200 392028 153252 392080
rect 140136 391960 140188 392012
rect 197360 391960 197412 392012
rect 3424 391212 3476 391264
rect 81440 391008 81492 391060
rect 85856 391008 85908 391060
rect 140044 391212 140096 391264
rect 157984 391212 158036 391264
rect 175280 391212 175332 391264
rect 120448 390260 120500 390312
rect 120816 390260 120868 390312
rect 113088 389784 113140 389836
rect 120724 389784 120776 389836
rect 57704 389240 57756 389292
rect 85580 389240 85632 389292
rect 25504 389172 25556 389224
rect 110420 389172 110472 389224
rect 111432 389172 111484 389224
rect 43996 389104 44048 389156
rect 70308 389104 70360 389156
rect 76656 389104 76708 389156
rect 91652 389104 91704 389156
rect 93216 389104 93268 389156
rect 96252 389104 96304 389156
rect 130476 389104 130528 389156
rect 76380 389036 76432 389088
rect 79508 388492 79560 388544
rect 86224 388492 86276 388544
rect 77852 388424 77904 388476
rect 171784 388424 171836 388476
rect 191104 388424 191156 388476
rect 88524 387812 88576 387864
rect 90364 387812 90416 387864
rect 57796 387744 57848 387796
rect 82084 387744 82136 387796
rect 104164 387744 104216 387796
rect 128360 387744 128412 387796
rect 11704 387064 11756 387116
rect 123668 387064 123720 387116
rect 185768 387064 185820 387116
rect 187240 386384 187292 386436
rect 197360 386384 197412 386436
rect 60464 386316 60516 386368
rect 86960 386316 87012 386368
rect 3424 385636 3476 385688
rect 95240 385636 95292 385688
rect 107200 385636 107252 385688
rect 167092 385636 167144 385688
rect 171048 385636 171100 385688
rect 191104 385636 191156 385688
rect 117596 384276 117648 384328
rect 196624 384276 196676 384328
rect 111800 383664 111852 383716
rect 113088 383664 113140 383716
rect 184296 383664 184348 383716
rect 65984 383596 66036 383648
rect 82820 383596 82872 383648
rect 61844 382916 61896 382968
rect 165620 382916 165672 382968
rect 123484 382236 123536 382288
rect 192668 382236 192720 382288
rect 79968 381488 80020 381540
rect 169852 381488 169904 381540
rect 50896 380876 50948 380928
rect 173164 380876 173216 380928
rect 59084 380808 59136 380860
rect 74540 380808 74592 380860
rect 49608 380128 49660 380180
rect 59084 380128 59136 380180
rect 73160 380128 73212 380180
rect 140136 380128 140188 380180
rect 188528 379516 188580 379568
rect 189816 379516 189868 379568
rect 197360 379516 197412 379568
rect 357900 379516 357952 379568
rect 382280 379516 382332 379568
rect 101404 378768 101456 378820
rect 152556 378768 152608 378820
rect 67272 378156 67324 378208
rect 195244 378156 195296 378208
rect 358360 378088 358412 378140
rect 360384 378088 360436 378140
rect 361488 377952 361540 378004
rect 364524 377952 364576 378004
rect 355324 377544 355376 377596
rect 356244 377544 356296 377596
rect 197084 377476 197136 377528
rect 201592 377476 201644 377528
rect 140688 376796 140740 376848
rect 198740 376796 198792 376848
rect 199108 376796 199160 376848
rect 72424 376728 72476 376780
rect 73068 376728 73120 376780
rect 187056 376728 187108 376780
rect 189908 376660 189960 376712
rect 218060 376660 218112 376712
rect 218244 376660 218296 376712
rect 92388 376048 92440 376100
rect 115664 376048 115716 376100
rect 352656 376048 352708 376100
rect 358820 376048 358872 376100
rect 48228 375980 48280 376032
rect 184388 375980 184440 376032
rect 198740 375980 198792 376032
rect 242164 375980 242216 376032
rect 353944 375980 353996 376032
rect 363236 375980 363288 376032
rect 50988 375300 51040 375352
rect 202236 375300 202288 375352
rect 203524 375300 203576 375352
rect 204996 375300 205048 375352
rect 236644 375300 236696 375352
rect 238116 375300 238168 375352
rect 260104 375300 260156 375352
rect 261484 375300 261536 375352
rect 262496 375300 262548 375352
rect 273076 375300 273128 375352
rect 273996 375300 274048 375352
rect 274732 375300 274784 375352
rect 278044 375300 278096 375352
rect 279700 375300 279752 375352
rect 320180 375300 320232 375352
rect 321284 375300 321336 375352
rect 339500 375300 339552 375352
rect 342352 375300 342404 375352
rect 344468 375300 344520 375352
rect 582380 375300 582432 375352
rect 194600 375232 194652 375284
rect 196808 375232 196860 375284
rect 233884 375232 233936 375284
rect 236460 375232 236512 375284
rect 348424 375232 348476 375284
rect 352748 375232 352800 375284
rect 50804 375096 50856 375148
rect 50988 375096 51040 375148
rect 304264 374824 304316 374876
rect 306196 374824 306248 374876
rect 327724 374824 327776 374876
rect 331220 374824 331272 374876
rect 198924 374620 198976 374672
rect 204352 374620 204404 374672
rect 246396 374620 246448 374672
rect 253204 374620 253256 374672
rect 258724 374620 258776 374672
rect 281356 374620 281408 374672
rect 282184 374620 282236 374672
rect 296260 374620 296312 374672
rect 309876 374620 309928 374672
rect 327908 374620 327960 374672
rect 198740 374280 198792 374332
rect 200028 374280 200080 374332
rect 206468 374280 206520 374332
rect 208308 374280 208360 374332
rect 119988 374008 120040 374060
rect 195336 374008 195388 374060
rect 226984 374008 227036 374060
rect 229836 374008 229888 374060
rect 250444 374008 250496 374060
rect 255964 374008 256016 374060
rect 276664 374008 276716 374060
rect 277676 374008 277728 374060
rect 294604 374008 294656 374060
rect 297916 374008 297968 374060
rect 308404 374008 308456 374060
rect 313924 374008 313976 374060
rect 354036 374008 354088 374060
rect 356060 374008 356112 374060
rect 199016 373328 199068 373380
rect 207020 373328 207072 373380
rect 355416 373328 355468 373380
rect 364432 373328 364484 373380
rect 101404 373260 101456 373312
rect 133236 373260 133288 373312
rect 184296 373260 184348 373312
rect 251824 373260 251876 373312
rect 286324 373260 286376 373312
rect 293960 373260 294012 373312
rect 340144 373260 340196 373312
rect 357624 373260 357676 373312
rect 136824 372648 136876 372700
rect 175924 372648 175976 372700
rect 67548 372580 67600 372632
rect 191196 372580 191248 372632
rect 334624 372580 334676 372632
rect 336740 372580 336792 372632
rect 180248 372512 180300 372564
rect 197268 372512 197320 372564
rect 582932 372512 582984 372564
rect 56416 371832 56468 371884
rect 76564 371832 76616 371884
rect 341524 371832 341576 371884
rect 357532 371832 357584 371884
rect 358084 371832 358136 371884
rect 365904 371832 365956 371884
rect 66904 371220 66956 371272
rect 67364 371220 67416 371272
rect 213184 371220 213236 371272
rect 195336 371152 195388 371204
rect 234620 371152 234672 371204
rect 267648 370540 267700 370592
rect 357716 370540 357768 370592
rect 84844 370472 84896 370524
rect 120724 370472 120776 370524
rect 124864 370472 124916 370524
rect 162768 370472 162820 370524
rect 387800 370472 387852 370524
rect 234620 369860 234672 369912
rect 235264 369860 235316 369912
rect 345664 369180 345716 369232
rect 361672 369180 361724 369232
rect 56508 369112 56560 369164
rect 144276 369112 144328 369164
rect 190368 369112 190420 369164
rect 211804 369112 211856 369164
rect 347044 369112 347096 369164
rect 365812 369112 365864 369164
rect 134616 368908 134668 368960
rect 135168 368908 135220 368960
rect 147680 368568 147732 368620
rect 148324 368568 148376 368620
rect 184296 368568 184348 368620
rect 135168 368500 135220 368552
rect 195244 368500 195296 368552
rect 125416 368432 125468 368484
rect 127716 368432 127768 368484
rect 86224 367820 86276 367872
rect 124772 367820 124824 367872
rect 67732 367752 67784 367804
rect 124864 367752 124916 367804
rect 144828 367752 144880 367804
rect 202880 367752 202932 367804
rect 209136 367752 209188 367804
rect 242256 367752 242308 367804
rect 359096 367752 359148 367804
rect 124220 367072 124272 367124
rect 124772 367072 124824 367124
rect 196624 367072 196676 367124
rect 71688 366936 71740 366988
rect 73804 366936 73856 366988
rect 231860 366800 231912 366852
rect 232596 366800 232648 366852
rect 77944 366392 77996 366444
rect 130384 366392 130436 366444
rect 331956 366392 332008 366444
rect 360292 366392 360344 366444
rect 99012 366324 99064 366376
rect 157432 366324 157484 366376
rect 159364 366324 159416 366376
rect 166816 366324 166868 366376
rect 203616 366324 203668 366376
rect 209044 366324 209096 366376
rect 218060 366324 218112 366376
rect 273260 366324 273312 366376
rect 349252 366324 349304 366376
rect 349804 366324 349856 366376
rect 368572 366324 368624 366376
rect 139492 365712 139544 365764
rect 232596 365712 232648 365764
rect 197176 365644 197228 365696
rect 198832 365644 198884 365696
rect 338948 365032 339000 365084
rect 363052 365032 363104 365084
rect 71596 364964 71648 365016
rect 136824 364964 136876 365016
rect 137284 364964 137336 365016
rect 185400 364964 185452 365016
rect 206376 364964 206428 365016
rect 212540 364964 212592 365016
rect 213276 364964 213328 365016
rect 356336 364964 356388 365016
rect 134708 364352 134760 364404
rect 200120 364352 200172 364404
rect 206284 364352 206336 364404
rect 206468 364352 206520 364404
rect 209228 364352 209280 364404
rect 58900 363604 58952 363656
rect 130384 363604 130436 363656
rect 325608 363604 325660 363656
rect 363144 363604 363196 363656
rect 137284 362992 137336 363044
rect 188344 362992 188396 363044
rect 188712 362992 188764 363044
rect 103428 362924 103480 362976
rect 149704 362924 149756 362976
rect 151728 362924 151780 362976
rect 325608 362924 325660 362976
rect 322296 362244 322348 362296
rect 347780 362244 347832 362296
rect 82084 362176 82136 362228
rect 259552 362176 259604 362228
rect 260104 362176 260156 362228
rect 338856 362176 338908 362228
rect 374092 362176 374144 362228
rect 81624 361564 81676 361616
rect 82084 361564 82136 361616
rect 90548 361564 90600 361616
rect 186136 361496 186188 361548
rect 367284 361496 367336 361548
rect 175096 361428 175148 361480
rect 211160 361428 211212 361480
rect 103336 360816 103388 360868
rect 155316 360816 155368 360868
rect 173348 360272 173400 360324
rect 173900 360272 173952 360324
rect 90456 360204 90508 360256
rect 181536 360204 181588 360256
rect 202144 359524 202196 359576
rect 228364 359524 228416 359576
rect 80152 359456 80204 359508
rect 81348 359456 81400 359508
rect 273260 359456 273312 359508
rect 99104 358776 99156 358828
rect 192484 358776 192536 358828
rect 3332 358708 3384 358760
rect 15844 358708 15896 358760
rect 47584 358708 47636 358760
rect 48044 358708 48096 358760
rect 79324 358096 79376 358148
rect 93860 358096 93912 358148
rect 206468 358096 206520 358148
rect 253940 358096 253992 358148
rect 273904 358096 273956 358148
rect 285680 358096 285732 358148
rect 47584 358028 47636 358080
rect 139492 358028 139544 358080
rect 235540 358028 235592 358080
rect 356152 358028 356204 358080
rect 142988 357484 143040 357536
rect 190092 357484 190144 357536
rect 103520 357416 103572 357468
rect 170404 357416 170456 357468
rect 180064 357348 180116 357400
rect 180340 357348 180392 357400
rect 75736 356736 75788 356788
rect 98828 356736 98880 356788
rect 129832 356736 129884 356788
rect 160008 356736 160060 356788
rect 202144 356736 202196 356788
rect 64604 356668 64656 356720
rect 107752 356668 107804 356720
rect 110328 356668 110380 356720
rect 164240 356668 164292 356720
rect 164700 356668 164752 356720
rect 180340 356668 180392 356720
rect 201408 356668 201460 356720
rect 240232 356668 240284 356720
rect 132592 355988 132644 356040
rect 244280 355988 244332 356040
rect 244924 355988 244976 356040
rect 81348 355308 81400 355360
rect 132592 355308 132644 355360
rect 195888 355308 195940 355360
rect 230480 355308 230532 355360
rect 94504 354696 94556 354748
rect 195888 354696 195940 354748
rect 93216 353948 93268 354000
rect 120724 353948 120776 354000
rect 305644 353948 305696 354000
rect 340880 353948 340932 354000
rect 104900 353336 104952 353388
rect 199384 353336 199436 353388
rect 120632 353268 120684 353320
rect 220084 353268 220136 353320
rect 235264 352588 235316 352640
rect 249800 352588 249852 352640
rect 76656 352520 76708 352572
rect 158720 352520 158772 352572
rect 161296 352520 161348 352572
rect 222200 352520 222252 352572
rect 240784 352520 240836 352572
rect 580172 352520 580224 352572
rect 240232 352180 240284 352232
rect 240784 352180 240836 352232
rect 101496 351908 101548 351960
rect 180064 351908 180116 351960
rect 96436 351228 96488 351280
rect 120632 351228 120684 351280
rect 64696 351160 64748 351212
rect 66996 351160 67048 351212
rect 195244 351160 195296 351212
rect 255320 351160 255372 351212
rect 273996 351160 274048 351212
rect 124128 350548 124180 350600
rect 255320 350548 255372 350600
rect 233148 350480 233200 350532
rect 240140 350480 240192 350532
rect 86868 349868 86920 349920
rect 100024 349868 100076 349920
rect 110420 349868 110472 349920
rect 158904 349868 158956 349920
rect 25504 349800 25556 349852
rect 67824 349800 67876 349852
rect 125692 349800 125744 349852
rect 142988 349800 143040 349852
rect 169208 349800 169260 349852
rect 309140 349800 309192 349852
rect 155316 349596 155368 349648
rect 155868 349596 155920 349648
rect 155868 349120 155920 349172
rect 233148 349120 233200 349172
rect 105544 348372 105596 348424
rect 157984 348372 158036 348424
rect 196808 348372 196860 348424
rect 231124 348372 231176 348424
rect 130384 347828 130436 347880
rect 133880 347828 133932 347880
rect 129096 347760 129148 347812
rect 201592 347760 201644 347812
rect 202236 347760 202288 347812
rect 93768 347012 93820 347064
rect 137284 347012 137336 347064
rect 139308 347012 139360 347064
rect 191656 347012 191708 347064
rect 121552 346400 121604 346452
rect 122748 346400 122800 346452
rect 221464 346400 221516 346452
rect 135168 346332 135220 346384
rect 139400 346332 139452 346384
rect 2780 346264 2832 346316
rect 4804 346264 4856 346316
rect 84108 345720 84160 345772
rect 108488 345720 108540 345772
rect 119344 345720 119396 345772
rect 157340 345720 157392 345772
rect 58900 345652 58952 345704
rect 134524 345652 134576 345704
rect 146116 345040 146168 345092
rect 242256 345040 242308 345092
rect 156604 344496 156656 344548
rect 162952 344496 163004 344548
rect 110328 344360 110380 344412
rect 116676 344360 116728 344412
rect 79692 344292 79744 344344
rect 111064 344292 111116 344344
rect 120724 344292 120776 344344
rect 235540 344292 235592 344344
rect 114468 343680 114520 343732
rect 124036 343680 124088 343732
rect 63408 343612 63460 343664
rect 66904 343612 66956 343664
rect 120080 343612 120132 343664
rect 120724 343612 120776 343664
rect 144644 343612 144696 343664
rect 156604 343612 156656 343664
rect 155776 343544 155828 343596
rect 207112 343544 207164 343596
rect 97908 342932 97960 342984
rect 129004 342932 129056 342984
rect 73804 342864 73856 342916
rect 144644 342864 144696 342916
rect 148968 342864 149020 342916
rect 158904 342864 158956 342916
rect 207112 342320 207164 342372
rect 207664 342320 207716 342372
rect 85396 342252 85448 342304
rect 90548 342252 90600 342304
rect 141424 342252 141476 342304
rect 142068 342252 142120 342304
rect 155132 342252 155184 342304
rect 158812 342252 158864 342304
rect 227076 342252 227128 342304
rect 55036 341504 55088 341556
rect 86960 341504 87012 341556
rect 155224 341504 155276 341556
rect 195244 341504 195296 341556
rect 304264 341504 304316 341556
rect 372712 341504 372764 341556
rect 125048 340960 125100 341012
rect 140780 340960 140832 341012
rect 95148 340892 95200 340944
rect 254032 340892 254084 340944
rect 140780 340824 140832 340876
rect 153200 340824 153252 340876
rect 153844 340824 153896 340876
rect 229744 340212 229796 340264
rect 309784 340212 309836 340264
rect 52368 340144 52420 340196
rect 125048 340144 125100 340196
rect 156696 340144 156748 340196
rect 337384 340144 337436 340196
rect 61844 339464 61896 339516
rect 162308 339464 162360 339516
rect 156604 338784 156656 338836
rect 207756 338784 207808 338836
rect 64788 338716 64840 338768
rect 116584 338716 116636 338768
rect 201408 338716 201460 338768
rect 335360 338716 335412 338768
rect 118516 338172 118568 338224
rect 131120 338172 131172 338224
rect 147680 338172 147732 338224
rect 156880 338172 156932 338224
rect 117228 338104 117280 338156
rect 196808 338104 196860 338156
rect 77300 337424 77352 337476
rect 85580 337424 85632 337476
rect 52184 337356 52236 337408
rect 82820 337356 82872 337408
rect 107384 337356 107436 337408
rect 129096 337356 129148 337408
rect 139216 337356 139268 337408
rect 147680 337356 147732 337408
rect 170404 337356 170456 337408
rect 249064 337356 249116 337408
rect 275284 337356 275336 337408
rect 371332 337356 371384 337408
rect 149612 336812 149664 336864
rect 174544 336812 174596 336864
rect 136548 336744 136600 336796
rect 169852 336744 169904 336796
rect 155776 335996 155828 336048
rect 224408 335996 224460 336048
rect 148140 335384 148192 335436
rect 155132 335384 155184 335436
rect 60648 335316 60700 335368
rect 84660 335316 84712 335368
rect 134892 335316 134944 335368
rect 163504 335316 163556 335368
rect 155132 334772 155184 334824
rect 160744 334772 160796 334824
rect 129280 334636 129332 334688
rect 136548 334636 136600 334688
rect 149060 334636 149112 334688
rect 155868 334636 155920 334688
rect 189908 334636 189960 334688
rect 243636 334636 243688 334688
rect 135168 334568 135220 334620
rect 149612 334568 149664 334620
rect 173164 334568 173216 334620
rect 192668 334568 192720 334620
rect 223028 334568 223080 334620
rect 582380 334568 582432 334620
rect 3424 333956 3476 334008
rect 124220 333956 124272 334008
rect 124956 333956 125008 334008
rect 137100 333956 137152 334008
rect 139492 333956 139544 334008
rect 140780 333956 140832 334008
rect 172704 333956 172756 334008
rect 52276 333888 52328 333940
rect 94320 333888 94372 333940
rect 20 333208 72 333260
rect 52276 333208 52328 333260
rect 83372 333208 83424 333260
rect 106924 333208 106976 333260
rect 132132 333208 132184 333260
rect 140780 333208 140832 333260
rect 240876 333208 240928 333260
rect 349804 333208 349856 333260
rect 143080 332664 143132 332716
rect 252560 332664 252612 332716
rect 67824 332596 67876 332648
rect 72424 332596 72476 332648
rect 106648 332596 106700 332648
rect 229192 332596 229244 332648
rect 59084 332528 59136 332580
rect 101496 332528 101548 332580
rect 142896 332528 142948 332580
rect 146944 332528 146996 332580
rect 74264 332460 74316 332512
rect 76748 332460 76800 332512
rect 70768 332120 70820 332172
rect 71504 332120 71556 332172
rect 78588 332120 78640 332172
rect 79324 332120 79376 332172
rect 88248 332120 88300 332172
rect 90456 332120 90508 332172
rect 110880 332120 110932 332172
rect 111616 332120 111668 332172
rect 113824 332120 113876 332172
rect 114468 332120 114520 332172
rect 115296 332120 115348 332172
rect 115848 332120 115900 332172
rect 116768 332120 116820 332172
rect 117228 332120 117280 332172
rect 118516 332120 118568 332172
rect 119068 332120 119120 332172
rect 123300 332120 123352 332172
rect 124128 332120 124180 332172
rect 125600 332120 125652 332172
rect 126428 332120 126480 332172
rect 129924 332120 129976 332172
rect 130384 332120 130436 332172
rect 138664 332120 138716 332172
rect 139308 332120 139360 332172
rect 143816 332120 143868 332172
rect 144736 332120 144788 332172
rect 145288 332120 145340 332172
rect 146024 332120 146076 332172
rect 149704 332120 149756 332172
rect 150348 332120 150400 332172
rect 98552 331984 98604 332036
rect 99288 331984 99340 332036
rect 162216 331984 162268 332036
rect 164976 331984 165028 332036
rect 232596 331916 232648 331968
rect 244280 331916 244332 331968
rect 33784 331848 33836 331900
rect 59084 331848 59136 331900
rect 107844 331848 107896 331900
rect 135168 331848 135220 331900
rect 188620 331848 188672 331900
rect 202880 331848 202932 331900
rect 215392 331848 215444 331900
rect 292580 331848 292632 331900
rect 80244 331576 80296 331628
rect 81348 331576 81400 331628
rect 135720 331576 135772 331628
rect 141424 331576 141476 331628
rect 95608 331508 95660 331560
rect 96528 331508 96580 331560
rect 109408 331508 109460 331560
rect 110328 331508 110380 331560
rect 90456 331440 90508 331492
rect 93124 331440 93176 331492
rect 94136 331440 94188 331492
rect 95148 331440 95200 331492
rect 100024 331440 100076 331492
rect 100668 331440 100720 331492
rect 134248 331440 134300 331492
rect 139216 331440 139268 331492
rect 83096 331304 83148 331356
rect 84108 331304 84160 331356
rect 88984 331304 89036 331356
rect 89628 331304 89680 331356
rect 97080 331304 97132 331356
rect 97908 331304 97960 331356
rect 118976 331304 119028 331356
rect 119896 331304 119948 331356
rect 119988 331304 120040 331356
rect 120540 331304 120592 331356
rect 132776 331304 132828 331356
rect 133788 331304 133840 331356
rect 150348 331304 150400 331356
rect 158076 331304 158128 331356
rect 50988 331236 51040 331288
rect 69388 331236 69440 331288
rect 151176 331236 151228 331288
rect 187148 331236 187200 331288
rect 184296 331100 184348 331152
rect 188344 331100 188396 331152
rect 204904 330624 204956 330676
rect 224224 330624 224276 330676
rect 175924 330556 175976 330608
rect 209320 330556 209372 330608
rect 289084 330556 289136 330608
rect 355416 330556 355468 330608
rect 67272 330488 67324 330540
rect 73804 330488 73856 330540
rect 131764 330488 131816 330540
rect 184480 330488 184532 330540
rect 209228 330488 209280 330540
rect 306380 330488 306432 330540
rect 67732 329808 67784 329860
rect 77300 329808 77352 329860
rect 162216 329808 162268 329860
rect 174544 329740 174596 329792
rect 180340 329740 180392 329792
rect 114560 329672 114612 329724
rect 115710 329672 115762 329724
rect 154120 329128 154172 329180
rect 157248 329128 157300 329180
rect 169852 329128 169904 329180
rect 174544 329128 174596 329180
rect 32404 329060 32456 329112
rect 47584 329060 47636 329112
rect 59084 328516 59136 328568
rect 66628 328516 66680 328568
rect 7564 328448 7616 328500
rect 114560 329060 114612 329112
rect 136456 329060 136508 329112
rect 139308 329060 139360 329112
rect 156328 329060 156380 329112
rect 172704 329060 172756 329112
rect 231216 329060 231268 329112
rect 253296 329060 253348 329112
rect 317420 329060 317472 329112
rect 186228 328924 186280 328976
rect 192576 328924 192628 328976
rect 156696 328788 156748 328840
rect 158168 328584 158220 328636
rect 158904 328516 158956 328568
rect 172520 328516 172572 328568
rect 156788 328448 156840 328500
rect 170404 328448 170456 328500
rect 180156 327768 180208 327820
rect 209228 327768 209280 327820
rect 222936 327768 222988 327820
rect 263600 327768 263652 327820
rect 236736 327700 236788 327752
rect 57796 327088 57848 327140
rect 169852 327088 169904 327140
rect 162308 327020 162360 327072
rect 170496 327020 170548 327072
rect 178040 326408 178092 326460
rect 245016 326408 245068 326460
rect 185584 326340 185636 326392
rect 204904 326340 204956 326392
rect 215944 326340 215996 326392
rect 348424 326340 348476 326392
rect 158996 325660 159048 325712
rect 181628 325660 181680 325712
rect 159088 325592 159140 325644
rect 167092 325592 167144 325644
rect 177396 324980 177448 325032
rect 187240 324980 187292 325032
rect 195244 324980 195296 325032
rect 235908 324980 235960 325032
rect 295984 324980 296036 325032
rect 170404 324912 170456 324964
rect 236644 324912 236696 324964
rect 158720 324368 158772 324420
rect 159088 324368 159140 324420
rect 167092 324300 167144 324352
rect 171876 324300 171928 324352
rect 158720 324232 158772 324284
rect 178776 324232 178828 324284
rect 220084 323552 220136 323604
rect 251364 323552 251416 323604
rect 305736 323552 305788 323604
rect 336004 323552 336056 323604
rect 158904 322940 158956 322992
rect 243728 322940 243780 322992
rect 158996 322328 159048 322380
rect 258172 322328 258224 322380
rect 158720 322260 158772 322312
rect 162952 322260 163004 322312
rect 185584 322260 185636 322312
rect 251824 322192 251876 322244
rect 260932 322192 260984 322244
rect 344284 322192 344336 322244
rect 3516 321512 3568 321564
rect 66904 321512 66956 321564
rect 176108 320900 176160 320952
rect 193864 320900 193916 320952
rect 156696 320832 156748 320884
rect 169300 320832 169352 320884
rect 178040 320832 178092 320884
rect 237380 320832 237432 320884
rect 281448 320832 281500 320884
rect 331956 320832 332008 320884
rect 55128 320152 55180 320204
rect 66812 320152 66864 320204
rect 237380 320152 237432 320204
rect 238024 320152 238076 320204
rect 281448 320152 281500 320204
rect 159272 319472 159324 319524
rect 159916 319472 159968 319524
rect 169116 319472 169168 319524
rect 174544 319472 174596 319524
rect 195244 319472 195296 319524
rect 231124 319472 231176 319524
rect 267832 319472 267884 319524
rect 4068 319404 4120 319456
rect 11704 319404 11756 319456
rect 163504 319404 163556 319456
rect 247132 319404 247184 319456
rect 281356 319404 281408 319456
rect 355324 319404 355376 319456
rect 34428 318724 34480 318776
rect 55864 318792 55916 318844
rect 66904 318792 66956 318844
rect 236736 318724 236788 318776
rect 237288 318724 237340 318776
rect 64696 318112 64748 318164
rect 66812 318112 66864 318164
rect 189080 318112 189132 318164
rect 246120 318112 246172 318164
rect 156880 318044 156932 318096
rect 233884 318044 233936 318096
rect 298008 318044 298060 318096
rect 345664 318044 345716 318096
rect 158720 317568 158772 317620
rect 163596 317568 163648 317620
rect 50804 317432 50856 317484
rect 52276 317432 52328 317484
rect 237288 317432 237340 317484
rect 296904 317432 296956 317484
rect 298008 317432 298060 317484
rect 158720 317364 158772 317416
rect 159088 317364 159140 317416
rect 169208 317364 169260 317416
rect 177488 316752 177540 316804
rect 258264 316752 258316 316804
rect 15844 316684 15896 316736
rect 67364 316684 67416 316736
rect 199476 316684 199528 316736
rect 352656 316684 352708 316736
rect 199384 315324 199436 315376
rect 220084 315324 220136 315376
rect 181628 315256 181680 315308
rect 210424 315256 210476 315308
rect 210516 315256 210568 315308
rect 240784 315256 240836 315308
rect 321560 315256 321612 315308
rect 357440 315256 357492 315308
rect 251824 314644 251876 314696
rect 321560 314644 321612 314696
rect 58900 314576 58952 314628
rect 66812 314576 66864 314628
rect 184388 313964 184440 314016
rect 238116 313964 238168 314016
rect 228456 313896 228508 313948
rect 380992 313896 381044 313948
rect 158720 313352 158772 313404
rect 163504 313352 163556 313404
rect 61844 313216 61896 313268
rect 66444 313216 66496 313268
rect 206468 313216 206520 313268
rect 209872 313216 209924 313268
rect 166448 312604 166500 312656
rect 200764 312604 200816 312656
rect 185584 312536 185636 312588
rect 225972 312536 226024 312588
rect 227076 312536 227128 312588
rect 253940 312536 253992 312588
rect 160836 311856 160888 311908
rect 166264 311856 166316 311908
rect 224408 311856 224460 311908
rect 224868 311856 224920 311908
rect 260840 311856 260892 311908
rect 161388 311788 161440 311840
rect 162860 311788 162912 311840
rect 244924 311788 244976 311840
rect 248420 311788 248472 311840
rect 170496 311176 170548 311228
rect 222936 311176 222988 311228
rect 18604 311108 18656 311160
rect 67456 311108 67508 311160
rect 169300 311108 169352 311160
rect 192484 311108 192536 311160
rect 202236 311108 202288 311160
rect 207020 311108 207072 311160
rect 287060 311108 287112 311160
rect 158720 310496 158772 310548
rect 170404 310496 170456 310548
rect 184480 310428 184532 310480
rect 226432 310428 226484 310480
rect 36544 309748 36596 309800
rect 63408 309748 63460 309800
rect 66812 309748 66864 309800
rect 158812 309748 158864 309800
rect 174636 309748 174688 309800
rect 317328 309748 317380 309800
rect 338948 309748 339000 309800
rect 177488 309136 177540 309188
rect 218152 309136 218204 309188
rect 239496 309136 239548 309188
rect 316132 309136 316184 309188
rect 317328 309136 317380 309188
rect 158720 308456 158772 308508
rect 165620 308456 165672 308508
rect 202144 308456 202196 308508
rect 231124 308456 231176 308508
rect 232504 308456 232556 308508
rect 259644 308456 259696 308508
rect 157984 308388 158036 308440
rect 240876 308388 240928 308440
rect 57612 307708 57664 307760
rect 66904 307708 66956 307760
rect 231216 307708 231268 307760
rect 232228 307708 232280 307760
rect 232228 307096 232280 307148
rect 281356 307096 281408 307148
rect 189724 307028 189776 307080
rect 197176 307028 197228 307080
rect 262864 307028 262916 307080
rect 322296 307028 322348 307080
rect 158720 306348 158772 306400
rect 167644 306348 167696 306400
rect 169116 306348 169168 306400
rect 252744 306348 252796 306400
rect 3516 306280 3568 306332
rect 32404 306280 32456 306332
rect 61936 306280 61988 306332
rect 66812 306280 66864 306332
rect 233884 305940 233936 305992
rect 234252 305940 234304 305992
rect 158720 305056 158772 305108
rect 231216 305056 231268 305108
rect 234252 305056 234304 305108
rect 274640 305056 274692 305108
rect 165068 304988 165120 305040
rect 165528 304988 165580 305040
rect 262312 304988 262364 305040
rect 63224 304920 63276 304972
rect 66812 304920 66864 304972
rect 158812 304920 158864 304972
rect 168196 304920 168248 304972
rect 168196 304240 168248 304292
rect 175924 304240 175976 304292
rect 182088 304240 182140 304292
rect 206376 304240 206428 304292
rect 206652 303696 206704 303748
rect 282276 303696 282328 303748
rect 211804 303628 211856 303680
rect 305000 303628 305052 303680
rect 165620 302880 165672 302932
rect 180156 302880 180208 302932
rect 329104 302880 329156 302932
rect 357440 302880 357492 302932
rect 184388 302268 184440 302320
rect 209964 302268 210016 302320
rect 210516 302268 210568 302320
rect 229836 302268 229888 302320
rect 270592 302268 270644 302320
rect 208492 302200 208544 302252
rect 209320 302200 209372 302252
rect 269856 302200 269908 302252
rect 59268 302132 59320 302184
rect 66904 302132 66956 302184
rect 194140 301520 194192 301572
rect 203524 301520 203576 301572
rect 207664 301520 207716 301572
rect 221648 301520 221700 301572
rect 158720 301452 158772 301504
rect 244556 301452 244608 301504
rect 274640 301452 274692 301504
rect 302424 301452 302476 301504
rect 340236 301452 340288 301504
rect 57612 300840 57664 300892
rect 66812 300840 66864 300892
rect 233148 300772 233200 300824
rect 233700 300772 233752 300824
rect 159640 300092 159692 300144
rect 180248 300092 180300 300144
rect 215300 299616 215352 299668
rect 216036 299616 216088 299668
rect 256792 299548 256844 299600
rect 197176 299480 197228 299532
rect 231308 299480 231360 299532
rect 233700 299480 233752 299532
rect 582472 299480 582524 299532
rect 195796 298800 195848 298852
rect 204352 298800 204404 298852
rect 159640 298732 159692 298784
rect 174544 298732 174596 298784
rect 180616 298732 180668 298784
rect 201500 298732 201552 298784
rect 221556 298732 221608 298784
rect 241428 298732 241480 298784
rect 243728 298732 243780 298784
rect 251180 298732 251232 298784
rect 292580 298732 292632 298784
rect 361580 298732 361632 298784
rect 59268 298120 59320 298172
rect 66628 298120 66680 298172
rect 243636 298120 243688 298172
rect 292580 298120 292632 298172
rect 50896 298052 50948 298104
rect 66812 298052 66864 298104
rect 158720 298052 158772 298104
rect 175280 298052 175332 298104
rect 175740 298052 175792 298104
rect 201408 298052 201460 298104
rect 202788 298052 202840 298104
rect 158628 297372 158680 297424
rect 171140 297372 171192 297424
rect 188988 297372 189040 297424
rect 194048 297372 194100 297424
rect 253204 297372 253256 297424
rect 259460 297372 259512 297424
rect 206284 296760 206336 296812
rect 211436 296760 211488 296812
rect 198372 296692 198424 296744
rect 282920 296692 282972 296744
rect 164884 295944 164936 295996
rect 184388 295944 184440 295996
rect 208032 295944 208084 295996
rect 226340 295944 226392 295996
rect 231308 295944 231360 295996
rect 272524 295944 272576 295996
rect 40684 295332 40736 295384
rect 67732 295332 67784 295384
rect 158720 295332 158772 295384
rect 169852 295332 169904 295384
rect 191288 295332 191340 295384
rect 211068 295332 211120 295384
rect 211436 295332 211488 295384
rect 278136 295332 278188 295384
rect 57796 295264 57848 295316
rect 66812 295264 66864 295316
rect 162216 294652 162268 294704
rect 213828 294652 213880 294704
rect 224224 294652 224276 294704
rect 227444 294652 227496 294704
rect 160836 294584 160888 294636
rect 164240 294584 164292 294636
rect 253204 294584 253256 294636
rect 221464 293972 221516 294024
rect 223948 293972 224000 294024
rect 241980 293972 242032 294024
rect 242256 293972 242308 294024
rect 283012 293972 283064 294024
rect 14464 293904 14516 293956
rect 52368 293904 52420 293956
rect 66812 293904 66864 293956
rect 219716 292680 219768 292732
rect 280804 292680 280856 292732
rect 158720 292612 158772 292664
rect 220176 292612 220228 292664
rect 3516 292544 3568 292596
rect 14556 292544 14608 292596
rect 183100 292544 183152 292596
rect 254584 292544 254636 292596
rect 54944 292476 54996 292528
rect 66812 292476 66864 292528
rect 158076 291796 158128 291848
rect 194048 291796 194100 291848
rect 200028 291796 200080 291848
rect 358084 291796 358136 291848
rect 158720 291184 158772 291236
rect 247316 291184 247368 291236
rect 41328 290436 41380 290488
rect 63500 290436 63552 290488
rect 166448 290436 166500 290488
rect 177488 290436 177540 290488
rect 240508 290436 240560 290488
rect 259552 290436 259604 290488
rect 313372 290436 313424 290488
rect 358912 290436 358964 290488
rect 63500 289892 63552 289944
rect 64696 289892 64748 289944
rect 66812 289892 66864 289944
rect 184020 289892 184072 289944
rect 244648 289892 244700 289944
rect 158720 289824 158772 289876
rect 223580 289824 223632 289876
rect 245016 289824 245068 289876
rect 245936 289824 245988 289876
rect 313372 289824 313424 289876
rect 169852 289756 169904 289808
rect 209044 289756 209096 289808
rect 50804 289076 50856 289128
rect 66720 289076 66772 289128
rect 217324 288464 217376 288516
rect 248512 288464 248564 288516
rect 50896 288396 50948 288448
rect 66812 288396 66864 288448
rect 158812 288396 158864 288448
rect 231308 288396 231360 288448
rect 239404 288396 239456 288448
rect 582564 288396 582616 288448
rect 231216 288328 231268 288380
rect 237012 288328 237064 288380
rect 238116 287648 238168 287700
rect 242900 287648 242952 287700
rect 158720 287104 158772 287156
rect 171968 287104 172020 287156
rect 184204 287104 184256 287156
rect 216772 287104 216824 287156
rect 218060 287104 218112 287156
rect 255412 287104 255464 287156
rect 63408 287036 63460 287088
rect 64788 287036 64840 287088
rect 66628 287036 66680 287088
rect 170496 287036 170548 287088
rect 223672 287036 223724 287088
rect 45468 286968 45520 287020
rect 52460 286968 52512 287020
rect 57704 286968 57756 287020
rect 66812 286968 66864 287020
rect 158720 286968 158772 287020
rect 169116 286968 169168 287020
rect 210424 286968 210476 287020
rect 218060 286968 218112 287020
rect 52460 286288 52512 286340
rect 53564 286288 53616 286340
rect 66352 286288 66404 286340
rect 158720 286288 158772 286340
rect 165068 286288 165120 286340
rect 166356 286288 166408 286340
rect 188528 286288 188580 286340
rect 282276 286288 282328 286340
rect 582840 286288 582892 286340
rect 223580 286084 223632 286136
rect 224500 286084 224552 286136
rect 231124 285812 231176 285864
rect 231676 285812 231728 285864
rect 190368 285744 190420 285796
rect 210884 285744 210936 285796
rect 222108 285744 222160 285796
rect 222844 285744 222896 285796
rect 225420 285744 225472 285796
rect 226432 285744 226484 285796
rect 236092 285744 236144 285796
rect 237288 285744 237340 285796
rect 258724 285744 258776 285796
rect 269028 285744 269080 285796
rect 275284 285744 275336 285796
rect 198832 285676 198884 285728
rect 204628 285676 204680 285728
rect 207572 285676 207624 285728
rect 300952 285676 301004 285728
rect 56508 285608 56560 285660
rect 66720 285608 66772 285660
rect 200120 285268 200172 285320
rect 200948 285268 201000 285320
rect 240140 285268 240192 285320
rect 241060 285268 241112 285320
rect 243176 285268 243228 285320
rect 244096 285268 244148 285320
rect 240784 285132 240836 285184
rect 243820 285132 243872 285184
rect 48228 284928 48280 284980
rect 56508 284928 56560 284980
rect 169116 284928 169168 284980
rect 198832 284928 198884 284980
rect 187608 284384 187660 284436
rect 217692 284384 217744 284436
rect 158812 284248 158864 284300
rect 244464 284316 244516 284368
rect 245660 283908 245712 283960
rect 245936 283908 245988 283960
rect 245936 283772 245988 283824
rect 248420 283772 248472 283824
rect 56508 283568 56560 283620
rect 66996 283568 67048 283620
rect 158720 283568 158772 283620
rect 178132 283568 178184 283620
rect 64604 282888 64656 282940
rect 66812 282888 66864 282940
rect 178132 282888 178184 282940
rect 179328 282888 179380 282940
rect 158720 282820 158772 282872
rect 197268 282888 197320 282940
rect 199476 282888 199528 282940
rect 195888 282820 195940 282872
rect 198004 282820 198056 282872
rect 254584 282820 254636 282872
rect 255136 282820 255188 282872
rect 383660 282820 383712 282872
rect 197360 282752 197412 282804
rect 245752 282752 245804 282804
rect 260932 282752 260984 282804
rect 183100 282684 183152 282736
rect 182916 282140 182968 282192
rect 192576 282140 192628 282192
rect 272616 282140 272668 282192
rect 282184 282140 282236 282192
rect 282276 282140 282328 282192
rect 302332 282140 302384 282192
rect 302884 282140 302936 282192
rect 327724 282140 327776 282192
rect 192760 282072 192812 282124
rect 194140 282072 194192 282124
rect 245936 281528 245988 281580
rect 249892 281528 249944 281580
rect 180156 281460 180208 281512
rect 197360 281460 197412 281512
rect 173256 280780 173308 280832
rect 176016 280780 176068 280832
rect 245660 280780 245712 280832
rect 250076 280780 250128 280832
rect 298284 280780 298336 280832
rect 378232 280780 378284 280832
rect 196716 280440 196768 280492
rect 197268 280440 197320 280492
rect 198280 280440 198332 280492
rect 21364 280168 21416 280220
rect 61844 280168 61896 280220
rect 67180 280168 67232 280220
rect 158720 280100 158772 280152
rect 169300 280100 169352 280152
rect 196624 280100 196676 280152
rect 199384 280100 199436 280152
rect 245752 279488 245804 279540
rect 249984 279488 250036 279540
rect 54944 279420 54996 279472
rect 67088 279420 67140 279472
rect 167644 279420 167696 279472
rect 193220 279420 193272 279472
rect 245936 279420 245988 279472
rect 255596 279420 255648 279472
rect 158720 278740 158772 278792
rect 165068 278740 165120 278792
rect 193220 278740 193272 278792
rect 197360 278740 197412 278792
rect 255596 278740 255648 278792
rect 583116 278740 583168 278792
rect 196808 278672 196860 278724
rect 197268 278672 197320 278724
rect 245752 278672 245804 278724
rect 249984 278672 250036 278724
rect 389180 278672 389232 278724
rect 266268 278604 266320 278656
rect 289084 278604 289136 278656
rect 180156 278060 180208 278112
rect 198832 278060 198884 278112
rect 158812 277992 158864 278044
rect 189080 277992 189132 278044
rect 389180 277992 389232 278044
rect 583392 277992 583444 278044
rect 63224 277380 63276 277432
rect 66812 277380 66864 277432
rect 158720 277312 158772 277364
rect 165160 277312 165212 277364
rect 186044 277312 186096 277364
rect 197360 277312 197412 277364
rect 49608 276632 49660 276684
rect 60464 276632 60516 276684
rect 66812 276632 66864 276684
rect 189080 276632 189132 276684
rect 190276 276632 190328 276684
rect 197360 276632 197412 276684
rect 246120 276632 246172 276684
rect 318800 276632 318852 276684
rect 367192 276632 367244 276684
rect 244096 276020 244148 276072
rect 245752 276020 245804 276072
rect 159364 275272 159416 275324
rect 172060 275272 172112 275324
rect 262956 275272 263008 275324
rect 278044 275272 278096 275324
rect 280988 275272 281040 275324
rect 583300 275272 583352 275324
rect 175280 274728 175332 274780
rect 178040 274728 178092 274780
rect 185676 274728 185728 274780
rect 197452 274728 197504 274780
rect 35808 274592 35860 274644
rect 57244 274592 57296 274644
rect 66628 274660 66680 274712
rect 158812 274660 158864 274712
rect 167644 274660 167696 274712
rect 169300 274660 169352 274712
rect 197360 274660 197412 274712
rect 158720 274592 158772 274644
rect 191196 274592 191248 274644
rect 194048 274524 194100 274576
rect 197084 274524 197136 274576
rect 197360 274524 197412 274576
rect 245936 273912 245988 273964
rect 289820 273912 289872 273964
rect 369952 273912 370004 273964
rect 264336 273572 264388 273624
rect 269120 273572 269172 273624
rect 180064 273300 180116 273352
rect 197360 273300 197412 273352
rect 184848 273164 184900 273216
rect 197360 273164 197412 273216
rect 245844 273164 245896 273216
rect 251180 273164 251232 273216
rect 252468 273164 252520 273216
rect 192668 273096 192720 273148
rect 197452 273096 197504 273148
rect 168288 272484 168340 272536
rect 183560 272484 183612 272536
rect 252468 272484 252520 272536
rect 288440 272484 288492 272536
rect 365720 272484 365772 272536
rect 52092 271872 52144 271924
rect 66260 271872 66312 271924
rect 574744 271872 574796 271924
rect 579804 271872 579856 271924
rect 191104 271804 191156 271856
rect 191840 271804 191892 271856
rect 191196 271192 191248 271244
rect 198740 271192 198792 271244
rect 158720 271124 158772 271176
rect 181536 271124 181588 271176
rect 245936 271124 245988 271176
rect 256976 271124 257028 271176
rect 286048 271124 286100 271176
rect 372620 271124 372672 271176
rect 195152 270512 195204 270564
rect 197360 270512 197412 270564
rect 245752 270444 245804 270496
rect 254032 270444 254084 270496
rect 166908 269832 166960 269884
rect 180248 269832 180300 269884
rect 180340 269832 180392 269884
rect 196716 269832 196768 269884
rect 260104 269832 260156 269884
rect 295340 269832 295392 269884
rect 4068 269764 4120 269816
rect 11704 269764 11756 269816
rect 158536 269764 158588 269816
rect 195152 269764 195204 269816
rect 245844 269764 245896 269816
rect 287152 269764 287204 269816
rect 256884 269084 256936 269136
rect 169208 269016 169260 269068
rect 197360 269016 197412 269068
rect 249064 269016 249116 269068
rect 250076 269016 250128 269068
rect 254400 269016 254452 269068
rect 583024 269016 583076 269068
rect 158720 268948 158772 269000
rect 170496 268948 170548 269000
rect 189080 268948 189132 269000
rect 189816 268948 189868 269000
rect 197452 268948 197504 269000
rect 178776 268336 178828 268388
rect 189080 268336 189132 268388
rect 246764 268336 246816 268388
rect 254400 268336 254452 268388
rect 158720 267928 158772 267980
rect 162124 267928 162176 267980
rect 63316 267792 63368 267844
rect 66812 267792 66864 267844
rect 3332 267724 3384 267776
rect 22744 267724 22796 267776
rect 61936 267724 61988 267776
rect 67180 267724 67232 267776
rect 170496 267656 170548 267708
rect 182824 267656 182876 267708
rect 188344 267656 188396 267708
rect 197360 267656 197412 267708
rect 246948 267520 247000 267572
rect 248420 267520 248472 267572
rect 270408 266976 270460 267028
rect 362960 266976 363012 267028
rect 189080 266364 189132 266416
rect 195336 266364 195388 266416
rect 162216 265616 162268 265668
rect 178868 265616 178920 265668
rect 245936 265616 245988 265668
rect 248604 265616 248656 265668
rect 251272 265616 251324 265668
rect 53564 264936 53616 264988
rect 66812 264936 66864 264988
rect 195336 264936 195388 264988
rect 197452 264936 197504 264988
rect 187056 264868 187108 264920
rect 197360 264868 197412 264920
rect 245844 264868 245896 264920
rect 273260 264868 273312 264920
rect 167828 264188 167880 264240
rect 183008 264188 183060 264240
rect 162768 263644 162820 263696
rect 164240 263644 164292 263696
rect 182824 263644 182876 263696
rect 197360 263644 197412 263696
rect 53748 263576 53800 263628
rect 57704 263576 57756 263628
rect 66812 263576 66864 263628
rect 158720 263576 158772 263628
rect 186964 263576 187016 263628
rect 253204 263508 253256 263560
rect 385132 263508 385184 263560
rect 158076 262896 158128 262948
rect 166448 262896 166500 262948
rect 169208 262896 169260 262948
rect 191288 262896 191340 262948
rect 39856 262828 39908 262880
rect 49608 262828 49660 262880
rect 159364 262828 159416 262880
rect 196624 262828 196676 262880
rect 166540 262488 166592 262540
rect 168656 262488 168708 262540
rect 49608 262216 49660 262268
rect 66812 262216 66864 262268
rect 245936 262216 245988 262268
rect 252652 262216 252704 262268
rect 11704 262148 11756 262200
rect 66444 262148 66496 262200
rect 191380 262148 191432 262200
rect 193220 262148 193272 262200
rect 175096 261536 175148 261588
rect 184480 261536 184532 261588
rect 157984 261468 158036 261520
rect 191840 261468 191892 261520
rect 197360 261468 197412 261520
rect 246396 261468 246448 261520
rect 247316 261468 247368 261520
rect 251180 261468 251232 261520
rect 264244 261468 264296 261520
rect 323584 261468 323636 261520
rect 245844 260788 245896 260840
rect 253204 260788 253256 260840
rect 163504 260108 163556 260160
rect 188344 260108 188396 260160
rect 260104 260108 260156 260160
rect 282276 260108 282328 260160
rect 314660 260108 314712 260160
rect 364340 260108 364392 260160
rect 64788 259428 64840 259480
rect 66812 259428 66864 259480
rect 193128 259428 193180 259480
rect 197360 259428 197412 259480
rect 245936 259428 245988 259480
rect 314660 259428 314712 259480
rect 175188 259360 175240 259412
rect 177396 259360 177448 259412
rect 191748 259360 191800 259412
rect 197452 259360 197504 259412
rect 245844 259360 245896 259412
rect 254124 259360 254176 259412
rect 381544 259360 381596 259412
rect 580172 259360 580224 259412
rect 245936 259292 245988 259344
rect 252744 259292 252796 259344
rect 253020 259292 253072 259344
rect 254124 258748 254176 258800
rect 255136 258748 255188 258800
rect 278044 258748 278096 258800
rect 158720 258680 158772 258732
rect 184204 258680 184256 258732
rect 187240 258680 187292 258732
rect 194416 258680 194468 258732
rect 197360 258680 197412 258732
rect 253020 258680 253072 258732
rect 294052 258680 294104 258732
rect 356704 258680 356756 258732
rect 159456 257320 159508 257372
rect 177396 257320 177448 257372
rect 307668 257320 307720 257372
rect 376852 257320 376904 257372
rect 187608 257048 187660 257100
rect 188436 257048 188488 257100
rect 177948 256776 178000 256828
rect 180800 256776 180852 256828
rect 196624 256776 196676 256828
rect 197176 256776 197228 256828
rect 198096 256776 198148 256828
rect 160100 256708 160152 256760
rect 186136 256708 186188 256760
rect 197452 256708 197504 256760
rect 246028 256708 246080 256760
rect 262128 256708 262180 256760
rect 269028 256708 269080 256760
rect 306564 256708 306616 256760
rect 307668 256708 307720 256760
rect 173164 256640 173216 256692
rect 197360 256640 197412 256692
rect 245936 256640 245988 256692
rect 259552 256640 259604 256692
rect 260748 256640 260800 256692
rect 61752 255960 61804 256012
rect 66996 255960 67048 256012
rect 260748 255960 260800 256012
rect 310612 255960 310664 256012
rect 379520 255960 379572 256012
rect 173716 255348 173768 255400
rect 176660 255348 176712 255400
rect 58992 255280 59044 255332
rect 66812 255280 66864 255332
rect 158812 255280 158864 255332
rect 173808 255280 173860 255332
rect 3148 255212 3200 255264
rect 18604 255212 18656 255264
rect 158720 255212 158772 255264
rect 167000 255212 167052 255264
rect 186228 255280 186280 255332
rect 187792 255280 187844 255332
rect 197452 255280 197504 255332
rect 197360 255212 197412 255264
rect 245936 255212 245988 255264
rect 258172 255212 258224 255264
rect 167000 254532 167052 254584
rect 191288 254532 191340 254584
rect 246948 254532 247000 254584
rect 582932 254532 582984 254584
rect 245476 253852 245528 253904
rect 269028 253852 269080 253904
rect 60372 253240 60424 253292
rect 66904 253240 66956 253292
rect 160836 253172 160888 253224
rect 164884 253172 164936 253224
rect 300768 253172 300820 253224
rect 341524 253172 341576 253224
rect 60556 252968 60608 253020
rect 66996 252968 67048 253020
rect 67364 252968 67416 253020
rect 158720 252560 158772 252612
rect 176016 252560 176068 252612
rect 193036 252560 193088 252612
rect 197360 252560 197412 252612
rect 245476 252560 245528 252612
rect 299664 252560 299716 252612
rect 300768 252560 300820 252612
rect 165160 252492 165212 252544
rect 166540 252492 166592 252544
rect 176568 252492 176620 252544
rect 178040 252492 178092 252544
rect 245936 252492 245988 252544
rect 251364 252492 251416 252544
rect 252468 252492 252520 252544
rect 187148 251880 187200 251932
rect 194048 251880 194100 251932
rect 173808 251812 173860 251864
rect 191656 251812 191708 251864
rect 195796 251812 195848 251864
rect 197360 251812 197412 251864
rect 252468 251812 252520 251864
rect 566464 251812 566516 251864
rect 168288 251132 168340 251184
rect 169300 251132 169352 251184
rect 179328 250520 179380 250572
rect 187056 250520 187108 250572
rect 160744 250452 160796 250504
rect 184848 250452 184900 250504
rect 309048 250452 309100 250504
rect 340144 250452 340196 250504
rect 60556 249840 60608 249892
rect 66904 249840 66956 249892
rect 195704 249840 195756 249892
rect 197912 249840 197964 249892
rect 63132 249772 63184 249824
rect 66812 249772 66864 249824
rect 187240 249772 187292 249824
rect 197360 249772 197412 249824
rect 245752 249772 245804 249824
rect 248604 249772 248656 249824
rect 307852 249772 307904 249824
rect 309048 249772 309100 249824
rect 181536 249704 181588 249756
rect 183468 249704 183520 249756
rect 193864 249704 193916 249756
rect 194508 249704 194560 249756
rect 245936 249500 245988 249552
rect 249800 249500 249852 249552
rect 295984 249024 296036 249076
rect 300860 249024 300912 249076
rect 194508 248684 194560 248736
rect 197452 248684 197504 248736
rect 245936 248616 245988 248668
rect 249984 248616 250036 248668
rect 158812 248480 158864 248532
rect 176568 248480 176620 248532
rect 158720 248412 158772 248464
rect 180708 248412 180760 248464
rect 182824 248412 182876 248464
rect 183468 248412 183520 248464
rect 197360 248412 197412 248464
rect 169760 248344 169812 248396
rect 185676 248344 185728 248396
rect 246948 247732 247000 247784
rect 251364 247732 251416 247784
rect 329748 247732 329800 247784
rect 354036 247732 354088 247784
rect 189724 247664 189776 247716
rect 195704 247664 195756 247716
rect 244556 247664 244608 247716
rect 264336 247664 264388 247716
rect 326344 247664 326396 247716
rect 353300 247664 353352 247716
rect 162124 247460 162176 247512
rect 168380 247460 168432 247512
rect 191748 247120 191800 247172
rect 192760 247120 192812 247172
rect 52368 247052 52420 247104
rect 66904 247052 66956 247104
rect 167736 247052 167788 247104
rect 169760 247052 169812 247104
rect 192668 247052 192720 247104
rect 197452 247052 197504 247104
rect 260196 247052 260248 247104
rect 328460 247052 328512 247104
rect 329748 247052 329800 247104
rect 59176 246984 59228 247036
rect 66812 246984 66864 247036
rect 184480 246984 184532 247036
rect 197360 246984 197412 247036
rect 320640 246304 320692 246356
rect 353944 246304 353996 246356
rect 197084 246100 197136 246152
rect 199384 246100 199436 246152
rect 177856 245828 177908 245880
rect 178684 245828 178736 245880
rect 162308 245692 162360 245744
rect 166356 245692 166408 245744
rect 158812 245624 158864 245676
rect 177856 245624 177908 245676
rect 245752 245624 245804 245676
rect 266452 245624 266504 245676
rect 320272 245624 320324 245676
rect 320640 245624 320692 245676
rect 165068 244876 165120 244928
rect 177488 244876 177540 244928
rect 184848 244876 184900 244928
rect 197360 244876 197412 244928
rect 278136 244876 278188 244928
rect 291844 244876 291896 244928
rect 303804 244876 303856 244928
rect 342260 244876 342312 244928
rect 57888 244264 57940 244316
rect 64512 244264 64564 244316
rect 66352 244264 66404 244316
rect 158720 244264 158772 244316
rect 195612 244264 195664 244316
rect 250444 244264 250496 244316
rect 303804 244264 303856 244316
rect 381544 244264 381596 244316
rect 580172 244264 580224 244316
rect 182272 244196 182324 244248
rect 197360 244196 197412 244248
rect 266360 244196 266412 244248
rect 267648 244196 267700 244248
rect 267832 244196 267884 244248
rect 171968 243584 172020 243636
rect 181628 243584 181680 243636
rect 156972 243516 157024 243568
rect 168288 243516 168340 243568
rect 177396 243516 177448 243568
rect 181720 243516 181772 243568
rect 197084 243516 197136 243568
rect 249064 243312 249116 243364
rect 250076 243312 250128 243364
rect 158720 242904 158772 242956
rect 164976 242904 165028 242956
rect 190276 242836 190328 242888
rect 191104 242836 191156 242888
rect 300860 242156 300912 242208
rect 352564 242156 352616 242208
rect 69756 241816 69808 241868
rect 71044 241816 71096 241868
rect 156880 241544 156932 241596
rect 184756 241544 184808 241596
rect 155316 241476 155368 241528
rect 195980 241544 196032 241596
rect 196624 241544 196676 241596
rect 195520 241476 195572 241528
rect 197820 241476 197872 241528
rect 246396 241476 246448 241528
rect 247316 241476 247368 241528
rect 300860 241476 300912 241528
rect 3516 241408 3568 241460
rect 25504 241408 25556 241460
rect 67824 241408 67876 241460
rect 180064 241408 180116 241460
rect 180248 241408 180300 241460
rect 193956 241408 194008 241460
rect 196992 241408 197044 241460
rect 288532 241408 288584 241460
rect 291200 241408 291252 241460
rect 67456 240728 67508 240780
rect 97908 240728 97960 240780
rect 111432 240728 111484 240780
rect 136364 240728 136416 240780
rect 154488 240728 154540 240780
rect 158536 240728 158588 240780
rect 164884 240728 164936 240780
rect 177856 240728 177908 240780
rect 194324 240728 194376 240780
rect 200120 240320 200172 240372
rect 192484 240252 192536 240304
rect 114560 240116 114612 240168
rect 115204 240116 115256 240168
rect 126980 240116 127032 240168
rect 127532 240116 127584 240168
rect 138020 240116 138072 240168
rect 138572 240116 138624 240168
rect 195980 240116 196032 240168
rect 200304 240116 200356 240168
rect 201040 240116 201092 240168
rect 202144 240116 202196 240168
rect 202788 240116 202840 240168
rect 207296 240116 207348 240168
rect 213920 240116 213972 240168
rect 221832 240116 221884 240168
rect 225328 240116 225380 240168
rect 231952 240116 232004 240168
rect 233148 240116 233200 240168
rect 245660 240184 245712 240236
rect 248604 240184 248656 240236
rect 288532 240116 288584 240168
rect 44088 240048 44140 240100
rect 75920 240048 75972 240100
rect 76564 240048 76616 240100
rect 93216 240048 93268 240100
rect 93768 240048 93820 240100
rect 96712 240048 96764 240100
rect 97540 240048 97592 240100
rect 99656 240048 99708 240100
rect 100668 240048 100720 240100
rect 102600 240048 102652 240100
rect 103336 240048 103388 240100
rect 104072 240048 104124 240100
rect 104808 240048 104860 240100
rect 110696 240048 110748 240100
rect 218980 240048 219032 240100
rect 219900 240048 219952 240100
rect 72608 239980 72660 240032
rect 73068 239980 73120 240032
rect 119344 239980 119396 240032
rect 119988 239980 120040 240032
rect 125968 239980 126020 240032
rect 126796 239980 126848 240032
rect 131856 239980 131908 240032
rect 132408 239980 132460 240032
rect 133328 239980 133380 240032
rect 133788 239980 133840 240032
rect 149336 239980 149388 240032
rect 150256 239980 150308 240032
rect 152004 239980 152056 240032
rect 157340 239980 157392 240032
rect 197452 239980 197504 240032
rect 201500 239980 201552 240032
rect 244556 239980 244608 240032
rect 79232 239912 79284 239964
rect 79876 239912 79928 239964
rect 82176 239912 82228 239964
rect 82728 239912 82780 239964
rect 117320 239912 117372 239964
rect 117964 239912 118016 239964
rect 129832 239912 129884 239964
rect 130476 239912 130528 239964
rect 132592 239912 132644 239964
rect 133420 239912 133472 239964
rect 150808 239912 150860 239964
rect 154488 239912 154540 239964
rect 85856 239844 85908 239896
rect 86868 239844 86920 239896
rect 130384 239776 130436 239828
rect 131028 239776 131080 239828
rect 112168 239640 112220 239692
rect 112996 239640 113048 239692
rect 201500 239640 201552 239692
rect 202420 239640 202472 239692
rect 116584 239504 116636 239556
rect 117136 239504 117188 239556
rect 120816 239504 120868 239556
rect 121368 239504 121420 239556
rect 108948 239436 109000 239488
rect 129556 239436 129608 239488
rect 74080 239368 74132 239420
rect 111064 239368 111116 239420
rect 141424 239368 141476 239420
rect 141976 239368 142028 239420
rect 144184 239368 144236 239420
rect 144828 239368 144880 239420
rect 145012 239368 145064 239420
rect 145748 239368 145800 239420
rect 311992 239368 312044 239420
rect 334072 239368 334124 239420
rect 95976 239232 96028 239284
rect 96528 239232 96580 239284
rect 105544 239232 105596 239284
rect 106188 239232 106240 239284
rect 128728 239232 128780 239284
rect 129648 239232 129700 239284
rect 135536 239232 135588 239284
rect 136456 239232 136508 239284
rect 143540 239232 143592 239284
rect 144276 239232 144328 239284
rect 153752 239232 153804 239284
rect 154488 239232 154540 239284
rect 82636 238756 82688 238808
rect 84844 238756 84896 238808
rect 214564 238756 214616 238808
rect 221464 238756 221516 238808
rect 224868 238756 224920 238808
rect 67916 238688 67968 238740
rect 190184 238688 190236 238740
rect 200212 238688 200264 238740
rect 205548 238688 205600 238740
rect 222292 238688 222344 238740
rect 223304 238688 223356 238740
rect 237380 238756 237432 238808
rect 311992 238756 312044 238808
rect 258080 238688 258132 238740
rect 259644 238688 259696 238740
rect 361488 238688 361540 238740
rect 381544 238688 381596 238740
rect 129556 238620 129608 238672
rect 219900 238620 219952 238672
rect 225788 238620 225840 238672
rect 233148 238620 233200 238672
rect 240324 238620 240376 238672
rect 240784 238620 240836 238672
rect 250444 238620 250496 238672
rect 151912 238552 151964 238604
rect 157984 238552 158036 238604
rect 215668 238212 215720 238264
rect 216496 238212 216548 238264
rect 63316 238008 63368 238060
rect 69756 238008 69808 238060
rect 195244 238008 195296 238060
rect 202328 238008 202380 238060
rect 202328 237668 202380 237720
rect 204076 237668 204128 237720
rect 200212 237396 200264 237448
rect 200764 237396 200816 237448
rect 201500 237396 201552 237448
rect 202604 237396 202656 237448
rect 223396 237396 223448 237448
rect 229652 237396 229704 237448
rect 14556 237328 14608 237380
rect 55036 237328 55088 237380
rect 138020 237328 138072 237380
rect 138112 237328 138164 237380
rect 156972 237328 157024 237380
rect 197084 237328 197136 237380
rect 207664 237328 207716 237380
rect 241796 237328 241848 237380
rect 242256 237328 242308 237380
rect 249064 237328 249116 237380
rect 242164 237260 242216 237312
rect 252560 237260 252612 237312
rect 239404 237192 239456 237244
rect 246304 237192 246356 237244
rect 157340 237124 157392 237176
rect 162216 237124 162268 237176
rect 207020 236716 207072 236768
rect 240692 236716 240744 236768
rect 64604 236648 64656 236700
rect 73804 236648 73856 236700
rect 78496 236648 78548 236700
rect 88340 236648 88392 236700
rect 97908 236648 97960 236700
rect 239220 236648 239272 236700
rect 88340 235968 88392 236020
rect 88984 235968 89036 236020
rect 162124 235968 162176 236020
rect 164148 235968 164200 236020
rect 76104 235900 76156 235952
rect 121644 235900 121696 235952
rect 147220 235900 147272 235952
rect 136364 235832 136416 235884
rect 155316 235832 155368 235884
rect 195612 235900 195664 235952
rect 241244 235900 241296 235952
rect 182088 235832 182140 235884
rect 203616 235832 203668 235884
rect 240876 235560 240928 235612
rect 243268 235560 243320 235612
rect 11704 235220 11756 235272
rect 52184 235220 52236 235272
rect 60372 235220 60424 235272
rect 146208 235220 146260 235272
rect 157432 235220 157484 235272
rect 166908 235220 166960 235272
rect 171876 235220 171928 235272
rect 227720 235220 227772 235272
rect 228732 235220 228784 235272
rect 295984 235220 296036 235272
rect 207388 235084 207440 235136
rect 209044 235084 209096 235136
rect 211804 234608 211856 234660
rect 212540 234608 212592 234660
rect 295524 234608 295576 234660
rect 295984 234608 296036 234660
rect 22744 234540 22796 234592
rect 92480 234540 92532 234592
rect 145012 234540 145064 234592
rect 237380 234540 237432 234592
rect 96712 234472 96764 234524
rect 150440 234472 150492 234524
rect 200304 234472 200356 234524
rect 270500 234472 270552 234524
rect 271236 234472 271288 234524
rect 92480 234132 92532 234184
rect 93124 234132 93176 234184
rect 163504 233860 163556 233912
rect 187240 233860 187292 233912
rect 127072 233180 127124 233232
rect 227720 233180 227772 233232
rect 235356 233180 235408 233232
rect 253940 233180 253992 233232
rect 143356 233112 143408 233164
rect 157340 233112 157392 233164
rect 65892 232568 65944 232620
rect 129004 232568 129056 232620
rect 224316 232568 224368 232620
rect 273904 232568 273956 232620
rect 61752 232500 61804 232552
rect 126244 232500 126296 232552
rect 208400 232500 208452 232552
rect 223396 232500 223448 232552
rect 253940 232500 253992 232552
rect 582748 232500 582800 232552
rect 126796 231752 126848 231804
rect 175188 231752 175240 231804
rect 176016 231752 176068 231804
rect 247316 231752 247368 231804
rect 140688 231684 140740 231736
rect 167736 231684 167788 231736
rect 200580 231684 200632 231736
rect 202144 231684 202196 231736
rect 218980 231684 219032 231736
rect 267740 231684 267792 231736
rect 269028 231684 269080 231736
rect 74540 231072 74592 231124
rect 138388 231072 138440 231124
rect 269028 231072 269080 231124
rect 288624 231072 288676 231124
rect 204168 230936 204220 230988
rect 210424 230936 210476 230988
rect 142160 230392 142212 230444
rect 234068 230392 234120 230444
rect 275928 230392 275980 230444
rect 276664 230392 276716 230444
rect 293960 230392 294012 230444
rect 294604 230392 294656 230444
rect 150256 230324 150308 230376
rect 157432 230324 157484 230376
rect 188344 230324 188396 230376
rect 206284 230324 206336 230376
rect 206836 230324 206888 230376
rect 66076 229712 66128 229764
rect 147496 229712 147548 229764
rect 167644 229712 167696 229764
rect 184204 229712 184256 229764
rect 208492 229712 208544 229764
rect 275928 229712 275980 229764
rect 287704 229712 287756 229764
rect 306472 229712 306524 229764
rect 262956 229100 263008 229152
rect 293960 229100 294012 229152
rect 86224 229032 86276 229084
rect 158168 229032 158220 229084
rect 181628 229032 181680 229084
rect 223764 229032 223816 229084
rect 110328 228964 110380 229016
rect 156788 228964 156840 229016
rect 156604 228352 156656 228404
rect 166448 228352 166500 228404
rect 234068 228352 234120 228404
rect 277584 228352 277636 228404
rect 223764 227740 223816 227792
rect 226984 227740 227036 227792
rect 229100 227740 229152 227792
rect 231952 227740 232004 227792
rect 259368 227740 259420 227792
rect 260104 227740 260156 227792
rect 60556 227672 60608 227724
rect 156604 227672 156656 227724
rect 187148 227672 187200 227724
rect 243544 227672 243596 227724
rect 126244 227604 126296 227656
rect 187700 227604 187752 227656
rect 302148 227060 302200 227112
rect 302884 227060 302936 227112
rect 196624 226992 196676 227044
rect 245844 226992 245896 227044
rect 302332 226992 302384 227044
rect 316040 226992 316092 227044
rect 156604 226584 156656 226636
rect 162308 226584 162360 226636
rect 187700 226312 187752 226364
rect 188528 226312 188580 226364
rect 279608 226312 279660 226364
rect 302332 226312 302384 226364
rect 103336 226244 103388 226296
rect 184756 226244 184808 226296
rect 221004 226244 221056 226296
rect 276020 226244 276072 226296
rect 142804 226176 142856 226228
rect 156880 226176 156932 226228
rect 194048 226176 194100 226228
rect 222844 226176 222896 226228
rect 276020 225564 276072 225616
rect 287244 225564 287296 225616
rect 184756 224952 184808 225004
rect 195152 224952 195204 225004
rect 84844 224884 84896 224936
rect 189724 224884 189776 224936
rect 195244 224884 195296 224936
rect 249800 224884 249852 224936
rect 126980 224816 127032 224868
rect 227260 224816 227312 224868
rect 277584 224204 277636 224256
rect 309140 224204 309192 224256
rect 322940 224204 322992 224256
rect 69020 223524 69072 223576
rect 231124 223524 231176 223576
rect 233240 223524 233292 223576
rect 138388 223456 138440 223508
rect 155224 223456 155276 223508
rect 155776 223456 155828 223508
rect 215116 223456 215168 223508
rect 238300 223456 238352 223508
rect 269948 223592 270000 223644
rect 279424 222844 279476 222896
rect 295432 222844 295484 222896
rect 69664 222096 69716 222148
rect 182916 222096 182968 222148
rect 184204 222096 184256 222148
rect 244372 222096 244424 222148
rect 100760 221416 100812 221468
rect 195888 221416 195940 221468
rect 202420 221416 202472 221468
rect 276664 221416 276716 221468
rect 91192 220736 91244 220788
rect 211344 220736 211396 220788
rect 227260 220736 227312 220788
rect 262956 220736 263008 220788
rect 104900 220668 104952 220720
rect 193128 220668 193180 220720
rect 193128 220056 193180 220108
rect 227076 220056 227128 220108
rect 215208 219444 215260 219496
rect 228364 219444 228416 219496
rect 124220 219376 124272 219428
rect 227720 219376 227772 219428
rect 231860 219376 231912 219428
rect 279608 219376 279660 219428
rect 73068 219308 73120 219360
rect 156604 219308 156656 219360
rect 170404 219308 170456 219360
rect 215208 219308 215260 219360
rect 95240 217948 95292 218000
rect 244280 217948 244332 218000
rect 132316 217880 132368 217932
rect 192668 217880 192720 217932
rect 195888 217880 195940 217932
rect 212540 217880 212592 217932
rect 192484 216656 192536 216708
rect 192668 216656 192720 216708
rect 212540 216656 212592 216708
rect 213184 216656 213236 216708
rect 117320 216588 117372 216640
rect 224224 216588 224276 216640
rect 177488 216520 177540 216572
rect 220176 216520 220228 216572
rect 220452 216520 220504 216572
rect 91100 215908 91152 215960
rect 92388 215908 92440 215960
rect 175280 215908 175332 215960
rect 164976 215228 165028 215280
rect 249892 215228 249944 215280
rect 114468 214616 114520 214668
rect 187148 214616 187200 214668
rect 35164 214548 35216 214600
rect 159364 214548 159416 214600
rect 197176 214548 197228 214600
rect 233332 214548 233384 214600
rect 260748 214548 260800 214600
rect 291292 214548 291344 214600
rect 100576 213868 100628 213920
rect 183284 213868 183336 213920
rect 184480 213868 184532 213920
rect 198648 213868 198700 213920
rect 199476 213868 199528 213920
rect 124312 213188 124364 213240
rect 198648 213188 198700 213240
rect 189080 212576 189132 212628
rect 190368 212576 190420 212628
rect 232136 212576 232188 212628
rect 207756 212508 207808 212560
rect 208216 212508 208268 212560
rect 278136 212508 278188 212560
rect 86960 212440 87012 212492
rect 209688 212440 209740 212492
rect 144828 211760 144880 211812
rect 237380 211760 237432 211812
rect 209688 211148 209740 211200
rect 214656 211148 214708 211200
rect 184848 210468 184900 210520
rect 244464 210468 244516 210520
rect 71044 210400 71096 210452
rect 188344 210400 188396 210452
rect 216496 209788 216548 209840
rect 245936 209788 245988 209840
rect 67732 209720 67784 209772
rect 206376 209720 206428 209772
rect 132408 209652 132460 209704
rect 248512 209652 248564 209704
rect 216680 208360 216732 208412
rect 217968 208360 218020 208412
rect 307852 208360 307904 208412
rect 70400 208292 70452 208344
rect 216496 208292 216548 208344
rect 187148 208224 187200 208276
rect 245752 208224 245804 208276
rect 133788 206932 133840 206984
rect 248696 206932 248748 206984
rect 122840 206864 122892 206916
rect 225604 206864 225656 206916
rect 82728 205572 82780 205624
rect 253940 205572 253992 205624
rect 106188 205504 106240 205556
rect 216680 205504 216732 205556
rect 218060 204280 218112 204332
rect 218244 204280 218296 204332
rect 229376 204280 229428 204332
rect 73804 204212 73856 204264
rect 217140 204212 217192 204264
rect 188344 204144 188396 204196
rect 234620 204144 234672 204196
rect 173164 203532 173216 203584
rect 184204 203532 184256 203584
rect 225696 203532 225748 203584
rect 284392 203532 284444 203584
rect 3424 202784 3476 202836
rect 137284 202784 137336 202836
rect 147588 202784 147640 202836
rect 247132 202784 247184 202836
rect 168288 202716 168340 202768
rect 169116 202716 169168 202768
rect 141976 202104 142028 202156
rect 168288 202104 168340 202156
rect 194416 202104 194468 202156
rect 245660 202104 245712 202156
rect 117228 200812 117280 200864
rect 190460 200812 190512 200864
rect 236828 200812 236880 200864
rect 245752 200812 245804 200864
rect 272524 200812 272576 200864
rect 290004 200812 290056 200864
rect 3424 200744 3476 200796
rect 169024 200744 169076 200796
rect 209044 200744 209096 200796
rect 238116 200744 238168 200796
rect 262864 200744 262916 200796
rect 281540 200744 281592 200796
rect 49608 200064 49660 200116
rect 177304 200064 177356 200116
rect 129004 199996 129056 200048
rect 195520 199996 195572 200048
rect 215208 199452 215260 199504
rect 242348 199452 242400 199504
rect 202328 199384 202380 199436
rect 238760 199384 238812 199436
rect 284300 198704 284352 198756
rect 294604 198704 294656 198756
rect 76564 198636 76616 198688
rect 238944 198636 238996 198688
rect 126888 198568 126940 198620
rect 252560 198568 252612 198620
rect 260196 198024 260248 198076
rect 270592 198024 270644 198076
rect 241428 197956 241480 198008
rect 306656 197956 306708 198008
rect 103428 197276 103480 197328
rect 163504 197276 163556 197328
rect 201408 196664 201460 196716
rect 232596 196664 232648 196716
rect 50896 196596 50948 196648
rect 204260 196596 204312 196648
rect 206468 196596 206520 196648
rect 284300 196596 284352 196648
rect 106280 195916 106332 195968
rect 162768 195916 162820 195968
rect 162768 195304 162820 195356
rect 192668 195304 192720 195356
rect 119988 195236 120040 195288
rect 177304 195236 177356 195288
rect 191380 195236 191432 195288
rect 200856 195236 200908 195288
rect 206284 195236 206336 195288
rect 245844 195236 245896 195288
rect 207664 193944 207716 193996
rect 227720 193944 227772 193996
rect 188528 193876 188580 193928
rect 217416 193876 217468 193928
rect 113088 193808 113140 193860
rect 191196 193808 191248 193860
rect 220268 193808 220320 193860
rect 276848 193808 276900 193860
rect 291844 193808 291896 193860
rect 301136 193808 301188 193860
rect 214656 192516 214708 192568
rect 233884 192516 233936 192568
rect 177396 192448 177448 192500
rect 247132 192448 247184 192500
rect 267004 192448 267056 192500
rect 292672 192448 292724 192500
rect 115204 191836 115256 191888
rect 196808 191836 196860 191888
rect 227720 191224 227772 191276
rect 253204 191224 253256 191276
rect 90364 191156 90416 191208
rect 192576 191156 192628 191208
rect 202144 191156 202196 191208
rect 232504 191156 232556 191208
rect 259368 191156 259420 191208
rect 305092 191156 305144 191208
rect 52092 191088 52144 191140
rect 167000 191088 167052 191140
rect 192484 191088 192536 191140
rect 228456 191088 228508 191140
rect 238116 191088 238168 191140
rect 303896 191088 303948 191140
rect 136640 190408 136692 190460
rect 243912 190408 243964 190460
rect 217324 189728 217376 189780
rect 238852 189728 238904 189780
rect 125508 189048 125560 189100
rect 174636 189048 174688 189100
rect 3516 188980 3568 189032
rect 15844 188980 15896 189032
rect 164884 188368 164936 188420
rect 241612 188368 241664 188420
rect 275928 188368 275980 188420
rect 295616 188368 295668 188420
rect 89628 188300 89680 188352
rect 220268 188300 220320 188352
rect 262128 188300 262180 188352
rect 299480 188300 299532 188352
rect 302148 188300 302200 188352
rect 314752 188300 314804 188352
rect 133144 187688 133196 187740
rect 164976 187688 165028 187740
rect 255964 187620 256016 187672
rect 258080 187620 258132 187672
rect 198648 186940 198700 186992
rect 242992 186940 243044 186992
rect 223488 186668 223540 186720
rect 227168 186668 227220 186720
rect 113088 186396 113140 186448
rect 177396 186396 177448 186448
rect 133788 186328 133840 186380
rect 210516 186328 210568 186380
rect 53472 186260 53524 186312
rect 169392 186260 169444 186312
rect 202236 186260 202288 186312
rect 292856 186328 292908 186380
rect 232596 185716 232648 185768
rect 242900 185716 242952 185768
rect 230204 185648 230256 185700
rect 233056 185648 233108 185700
rect 213184 185580 213236 185632
rect 238944 185580 238996 185632
rect 269764 185580 269816 185632
rect 285956 185580 286008 185632
rect 118608 184900 118660 184952
rect 185584 184900 185636 184952
rect 227076 184220 227128 184272
rect 244556 184220 244608 184272
rect 191104 184152 191156 184204
rect 230572 184152 230624 184204
rect 244188 184152 244240 184204
rect 283564 184152 283616 184204
rect 316776 184152 316828 184204
rect 326344 184152 326396 184204
rect 129004 183608 129056 183660
rect 167828 183608 167880 183660
rect 107568 183540 107620 183592
rect 166356 183540 166408 183592
rect 180708 182860 180760 182912
rect 229468 182860 229520 182912
rect 199384 182792 199436 182844
rect 248604 182792 248656 182844
rect 280896 182792 280948 182844
rect 291384 182792 291436 182844
rect 134800 182248 134852 182300
rect 162860 182248 162912 182300
rect 121920 182180 121972 182232
rect 173256 182180 173308 182232
rect 271236 181500 271288 181552
rect 283196 181500 283248 181552
rect 184296 181432 184348 181484
rect 237472 181432 237524 181484
rect 273904 181432 273956 181484
rect 288716 181432 288768 181484
rect 105912 180888 105964 180940
rect 170404 180888 170456 180940
rect 132408 180820 132460 180872
rect 214932 180820 214984 180872
rect 226248 180820 226300 180872
rect 251364 180820 251416 180872
rect 220268 180140 220320 180192
rect 232228 180140 232280 180192
rect 278136 180140 278188 180192
rect 280252 180140 280304 180192
rect 187056 180072 187108 180124
rect 226432 180072 226484 180124
rect 233884 180072 233936 180124
rect 241520 180072 241572 180124
rect 253204 180072 253256 180124
rect 276020 180072 276072 180124
rect 284944 180072 284996 180124
rect 298376 180072 298428 180124
rect 119896 179460 119948 179512
rect 167736 179460 167788 179512
rect 126796 179392 126848 179444
rect 206284 179392 206336 179444
rect 227168 179392 227220 179444
rect 229284 179392 229336 179444
rect 276848 179392 276900 179444
rect 279148 179392 279200 179444
rect 281448 179392 281500 179444
rect 284484 179392 284536 179444
rect 220176 178712 220228 178764
rect 233240 178712 233292 178764
rect 279424 178712 279476 178764
rect 296996 178712 297048 178764
rect 200856 178644 200908 178696
rect 231952 178644 232004 178696
rect 232504 178644 232556 178696
rect 292764 178644 292816 178696
rect 123300 178100 123352 178152
rect 169116 178100 169168 178152
rect 148232 178032 148284 178084
rect 203616 178032 203668 178084
rect 129464 177964 129516 178016
rect 133144 177964 133196 178016
rect 203524 177964 203576 178016
rect 226340 177964 226392 178016
rect 114192 177556 114244 177608
rect 115204 177556 115256 177608
rect 127992 177556 128044 177608
rect 129004 177556 129056 177608
rect 278044 177352 278096 177404
rect 287336 177352 287388 177404
rect 228364 177284 228416 177336
rect 233424 177284 233476 177336
rect 268384 177284 268436 177336
rect 281816 177284 281868 177336
rect 158996 176740 159048 176792
rect 173164 176740 173216 176792
rect 128176 176672 128228 176724
rect 207020 176672 207072 176724
rect 135720 176604 135772 176656
rect 213920 176604 213972 176656
rect 197268 176536 197320 176588
rect 229100 176672 229152 176724
rect 269948 176604 270000 176656
rect 281724 176604 281776 176656
rect 334624 176604 334676 176656
rect 283564 175992 283616 176044
rect 284576 175992 284628 176044
rect 130752 175924 130804 175976
rect 165528 175924 165580 175976
rect 226432 175924 226484 175976
rect 233516 175924 233568 175976
rect 276664 175924 276716 175976
rect 226524 175788 226576 175840
rect 228456 175788 228508 175840
rect 231860 175788 231912 175840
rect 283012 175924 283064 175976
rect 283196 175924 283248 175976
rect 283196 175788 283248 175840
rect 210516 175176 210568 175228
rect 214012 175176 214064 175228
rect 214564 175176 214616 175228
rect 239588 175244 239640 175296
rect 264980 175244 265032 175296
rect 230664 175176 230716 175228
rect 232228 175176 232280 175228
rect 256976 175176 257028 175228
rect 280988 175176 281040 175228
rect 281908 175176 281960 175228
rect 282184 175176 282236 175228
rect 285772 175176 285824 175228
rect 229376 175108 229428 175160
rect 162860 175040 162912 175092
rect 213920 175040 213972 175092
rect 280804 175040 280856 175092
rect 285772 175040 285824 175092
rect 229008 174972 229060 175024
rect 231952 174972 232004 175024
rect 260288 173952 260340 174004
rect 265072 173952 265124 174004
rect 236644 173884 236696 173936
rect 264980 173884 265032 173936
rect 165528 173816 165580 173868
rect 213920 173816 213972 173868
rect 282460 173816 282512 173868
rect 302424 173816 302476 173868
rect 230756 173136 230808 173188
rect 247224 173136 247276 173188
rect 230388 172524 230440 172576
rect 233332 172524 233384 172576
rect 249248 172524 249300 172576
rect 264980 172524 265032 172576
rect 164976 172456 165028 172508
rect 213920 172456 213972 172508
rect 231400 172456 231452 172508
rect 252560 172456 252612 172508
rect 207020 172388 207072 172440
rect 214012 172388 214064 172440
rect 231308 172388 231360 172440
rect 240140 172388 240192 172440
rect 254676 171164 254728 171216
rect 264980 171164 265032 171216
rect 167920 171096 167972 171148
rect 182916 171096 182968 171148
rect 247684 171096 247736 171148
rect 265072 171096 265124 171148
rect 167828 171028 167880 171080
rect 213920 171028 213972 171080
rect 206284 170960 206336 171012
rect 214012 170960 214064 171012
rect 282276 170892 282328 170944
rect 285772 170892 285824 170944
rect 246672 170348 246724 170400
rect 256792 170348 256844 170400
rect 261484 169804 261536 169856
rect 265072 169804 265124 169856
rect 231216 169736 231268 169788
rect 234620 169736 234672 169788
rect 234896 169736 234948 169788
rect 238024 169736 238076 169788
rect 238300 169736 238352 169788
rect 264980 169736 265032 169788
rect 169116 169668 169168 169720
rect 214012 169668 214064 169720
rect 282828 169668 282880 169720
rect 292856 169668 292908 169720
rect 174636 169600 174688 169652
rect 213920 169600 213972 169652
rect 230572 169464 230624 169516
rect 233240 169464 233292 169516
rect 231124 169396 231176 169448
rect 234804 169396 234856 169448
rect 233884 168512 233936 168564
rect 238760 168512 238812 168564
rect 243544 168444 243596 168496
rect 264980 168444 265032 168496
rect 238024 168376 238076 168428
rect 265072 168376 265124 168428
rect 166540 168308 166592 168360
rect 214012 168308 214064 168360
rect 282276 168308 282328 168360
rect 290096 168308 290148 168360
rect 173256 168240 173308 168292
rect 213920 168240 213972 168292
rect 231400 168036 231452 168088
rect 237472 168036 237524 168088
rect 231400 167084 231452 167136
rect 236828 167084 236880 167136
rect 239772 167084 239824 167136
rect 264980 167084 265032 167136
rect 236736 167016 236788 167068
rect 265072 167016 265124 167068
rect 167736 166948 167788 167000
rect 213920 166948 213972 167000
rect 566464 166948 566516 167000
rect 580172 166948 580224 167000
rect 171784 166880 171836 166932
rect 214012 166880 214064 166932
rect 231768 166676 231820 166728
rect 234896 166676 234948 166728
rect 234068 166064 234120 166116
rect 238944 166064 238996 166116
rect 245108 165656 245160 165708
rect 265072 165656 265124 165708
rect 235264 165588 235316 165640
rect 264980 165588 265032 165640
rect 166448 165520 166500 165572
rect 214012 165520 214064 165572
rect 180156 165452 180208 165504
rect 213920 165452 213972 165504
rect 281908 165316 281960 165368
rect 284576 165316 284628 165368
rect 231492 165180 231544 165232
rect 235448 165180 235500 165232
rect 253388 164296 253440 164348
rect 264980 164296 265032 164348
rect 240784 164228 240836 164280
rect 265072 164228 265124 164280
rect 3240 164160 3292 164212
rect 40684 164160 40736 164212
rect 177396 164160 177448 164212
rect 214012 164160 214064 164212
rect 230020 164160 230072 164212
rect 230664 164160 230716 164212
rect 231032 164160 231084 164212
rect 255412 164160 255464 164212
rect 196808 164092 196860 164144
rect 213920 164092 213972 164144
rect 231676 164092 231728 164144
rect 244372 164092 244424 164144
rect 282828 163276 282880 163328
rect 288716 163276 288768 163328
rect 258908 162936 258960 162988
rect 265072 162936 265124 162988
rect 245016 162868 245068 162920
rect 264980 162868 265032 162920
rect 164884 162800 164936 162852
rect 213920 162800 213972 162852
rect 230388 162800 230440 162852
rect 230848 162800 230900 162852
rect 230940 162800 230992 162852
rect 233516 162800 233568 162852
rect 282828 162800 282880 162852
rect 296904 162800 296956 162852
rect 207756 162732 207808 162784
rect 214012 162732 214064 162784
rect 184480 162120 184532 162172
rect 207664 162120 207716 162172
rect 231124 162120 231176 162172
rect 260288 162120 260340 162172
rect 262864 161644 262916 161696
rect 265072 161644 265124 161696
rect 243912 161440 243964 161492
rect 264980 161440 265032 161492
rect 166356 161372 166408 161424
rect 214012 161372 214064 161424
rect 282828 161372 282880 161424
rect 303804 161372 303856 161424
rect 170496 161304 170548 161356
rect 213920 161304 213972 161356
rect 231676 160692 231728 160744
rect 242992 160692 243044 160744
rect 281724 160556 281776 160608
rect 284484 160556 284536 160608
rect 257436 160148 257488 160200
rect 264980 160148 265032 160200
rect 234160 160080 234212 160132
rect 265072 160080 265124 160132
rect 170404 160012 170456 160064
rect 213920 160012 213972 160064
rect 231768 160012 231820 160064
rect 248420 160012 248472 160064
rect 281908 160012 281960 160064
rect 318800 160012 318852 160064
rect 231400 159944 231452 159996
rect 240968 159944 241020 159996
rect 282368 159944 282420 159996
rect 292764 159944 292816 159996
rect 254584 158788 254636 158840
rect 264980 158788 265032 158840
rect 240876 158720 240928 158772
rect 265072 158720 265124 158772
rect 169024 158652 169076 158704
rect 214012 158652 214064 158704
rect 192484 158584 192536 158636
rect 213920 158584 213972 158636
rect 231216 158584 231268 158636
rect 236000 158584 236052 158636
rect 282828 157564 282880 157616
rect 287336 157564 287388 157616
rect 249340 157428 249392 157480
rect 264980 157428 265032 157480
rect 240968 157360 241020 157412
rect 265072 157360 265124 157412
rect 167644 157292 167696 157344
rect 214012 157292 214064 157344
rect 188528 157224 188580 157276
rect 213920 157224 213972 157276
rect 231768 157224 231820 157276
rect 244280 157224 244332 157276
rect 280068 156612 280120 156664
rect 285864 156612 285916 156664
rect 247868 156000 247920 156052
rect 264980 156000 265032 156052
rect 235540 155932 235592 155984
rect 265072 155932 265124 155984
rect 166264 155864 166316 155916
rect 214012 155864 214064 155916
rect 281632 155864 281684 155916
rect 321560 155864 321612 155916
rect 184572 155796 184624 155848
rect 213920 155796 213972 155848
rect 231492 155796 231544 155848
rect 234068 155796 234120 155848
rect 231676 155184 231728 155236
rect 240416 155184 240468 155236
rect 250536 154640 250588 154692
rect 264980 154640 265032 154692
rect 238116 154572 238168 154624
rect 265164 154572 265216 154624
rect 231492 154504 231544 154556
rect 242900 154504 242952 154556
rect 231768 154436 231820 154488
rect 241612 154436 241664 154488
rect 281632 154436 281684 154488
rect 295616 154436 295668 154488
rect 206376 153280 206428 153332
rect 213920 153280 213972 153332
rect 249064 153280 249116 153332
rect 264980 153280 265032 153332
rect 198188 153212 198240 153264
rect 214012 153212 214064 153264
rect 243728 153212 243780 153264
rect 265072 153212 265124 153264
rect 281632 153144 281684 153196
rect 296996 153144 297048 153196
rect 231492 152940 231544 152992
rect 237380 152940 237432 152992
rect 236920 152464 236972 152516
rect 265348 152464 265400 152516
rect 281632 152464 281684 152516
rect 295524 152464 295576 152516
rect 211804 152192 211856 152244
rect 214012 152192 214064 152244
rect 252008 151784 252060 151836
rect 264980 151784 265032 151836
rect 231492 151716 231544 151768
rect 245936 151716 245988 151768
rect 281816 151036 281868 151088
rect 300860 151036 300912 151088
rect 231676 150900 231728 150952
rect 234712 150900 234764 150952
rect 187148 150492 187200 150544
rect 213920 150492 213972 150544
rect 247776 150492 247828 150544
rect 264980 150492 265032 150544
rect 169116 150424 169168 150476
rect 214012 150424 214064 150476
rect 235448 150424 235500 150476
rect 265072 150424 265124 150476
rect 3516 150356 3568 150408
rect 11704 150356 11756 150408
rect 182916 150356 182968 150408
rect 214104 150356 214156 150408
rect 281632 150356 281684 150408
rect 294144 150356 294196 150408
rect 281724 150288 281776 150340
rect 292672 150288 292724 150340
rect 173164 149676 173216 149728
rect 213920 149676 213972 149728
rect 232688 149676 232740 149728
rect 265624 149676 265676 149728
rect 244924 149064 244976 149116
rect 264980 149064 265032 149116
rect 281632 148996 281684 149048
rect 294052 148996 294104 149048
rect 231492 148792 231544 148844
rect 233884 148792 233936 148844
rect 232872 148316 232924 148368
rect 265164 148316 265216 148368
rect 173256 147636 173308 147688
rect 213920 147636 213972 147688
rect 229928 147636 229980 147688
rect 232136 147636 232188 147688
rect 238208 147636 238260 147688
rect 264980 147636 265032 147688
rect 282828 147568 282880 147620
rect 306656 147568 306708 147620
rect 181444 146888 181496 146940
rect 192484 146888 192536 146940
rect 192576 146888 192628 146940
rect 204996 146888 205048 146940
rect 206284 146888 206336 146940
rect 214564 146888 214616 146940
rect 262772 146344 262824 146396
rect 265072 146344 265124 146396
rect 166264 146276 166316 146328
rect 213920 146276 213972 146328
rect 256056 146276 256108 146328
rect 264980 146276 265032 146328
rect 231676 146208 231728 146260
rect 245844 146208 245896 146260
rect 282368 146208 282420 146260
rect 291476 146208 291528 146260
rect 184296 145528 184348 145580
rect 214012 145528 214064 145580
rect 262588 144984 262640 145036
rect 265072 144984 265124 145036
rect 201408 144916 201460 144968
rect 213920 144916 213972 144968
rect 246580 144916 246632 144968
rect 264980 144916 265032 144968
rect 231216 144848 231268 144900
rect 238300 144848 238352 144900
rect 167644 144168 167696 144220
rect 201408 144168 201460 144220
rect 236828 144168 236880 144220
rect 262772 144168 262824 144220
rect 209044 143624 209096 143676
rect 213920 143624 213972 143676
rect 184388 143556 184440 143608
rect 214012 143556 214064 143608
rect 252100 143556 252152 143608
rect 264980 143556 265032 143608
rect 282828 143488 282880 143540
rect 290004 143488 290056 143540
rect 231676 143420 231728 143472
rect 234252 143420 234304 143472
rect 231308 142876 231360 142928
rect 254676 142876 254728 142928
rect 238392 142808 238444 142860
rect 262588 142808 262640 142860
rect 258816 142740 258868 142792
rect 264980 142740 265032 142792
rect 177488 142128 177540 142180
rect 213920 142128 213972 142180
rect 282092 142060 282144 142112
rect 299480 142060 299532 142112
rect 282828 141992 282880 142044
rect 298284 141992 298336 142044
rect 180064 141380 180116 141432
rect 200764 141380 200816 141432
rect 250812 141380 250864 141432
rect 265716 141380 265768 141432
rect 231124 141312 231176 141364
rect 233884 141312 233936 141364
rect 203524 140768 203576 140820
rect 213920 140768 213972 140820
rect 231768 140700 231820 140752
rect 247132 140700 247184 140752
rect 282828 140700 282880 140752
rect 313372 140700 313424 140752
rect 231676 140020 231728 140072
rect 247684 140020 247736 140072
rect 189724 139408 189776 139460
rect 213920 139408 213972 139460
rect 263048 139408 263100 139460
rect 265348 139408 265400 139460
rect 282828 139340 282880 139392
rect 302516 139340 302568 139392
rect 231492 138864 231544 138916
rect 235356 138864 235408 138916
rect 176016 138660 176068 138712
rect 214012 138660 214064 138712
rect 202144 137980 202196 138032
rect 213920 137980 213972 138032
rect 233884 137980 233936 138032
rect 264980 137980 265032 138032
rect 265716 137980 265768 138032
rect 267096 137980 267148 138032
rect 3516 137912 3568 137964
rect 17224 137912 17276 137964
rect 231584 137912 231636 137964
rect 251364 137912 251416 137964
rect 282828 137912 282880 137964
rect 299664 137912 299716 137964
rect 198096 136688 198148 136740
rect 213920 136688 213972 136740
rect 171784 136620 171836 136672
rect 214012 136620 214064 136672
rect 247684 136620 247736 136672
rect 264980 136620 265032 136672
rect 230572 136552 230624 136604
rect 232688 136552 232740 136604
rect 282828 136552 282880 136604
rect 303896 136552 303948 136604
rect 167828 135872 167880 135924
rect 213184 135872 213236 135924
rect 231492 135872 231544 135924
rect 236644 135872 236696 135924
rect 243636 135328 243688 135380
rect 264980 135328 265032 135380
rect 180064 135260 180116 135312
rect 213920 135260 213972 135312
rect 235356 135260 235408 135312
rect 265072 135260 265124 135312
rect 231584 135192 231636 135244
rect 264244 135192 264296 135244
rect 282460 135124 282512 135176
rect 285956 135124 286008 135176
rect 192576 134512 192628 134564
rect 214104 134512 214156 134564
rect 230756 134512 230808 134564
rect 239772 134512 239824 134564
rect 173164 133900 173216 133952
rect 213920 133900 213972 133952
rect 239496 133900 239548 133952
rect 264980 133900 265032 133952
rect 230848 133832 230900 133884
rect 257620 133832 257672 133884
rect 282736 133832 282788 133884
rect 311992 133832 312044 133884
rect 231768 133764 231820 133816
rect 249248 133764 249300 133816
rect 282828 133764 282880 133816
rect 300952 133764 301004 133816
rect 174636 133152 174688 133204
rect 206376 133152 206428 133204
rect 249432 133152 249484 133204
rect 265808 133152 265860 133204
rect 209136 132540 209188 132592
rect 213920 132540 213972 132592
rect 181444 132472 181496 132524
rect 214012 132472 214064 132524
rect 257344 132472 257396 132524
rect 264980 132472 265032 132524
rect 231676 132404 231728 132456
rect 261484 132404 261536 132456
rect 282828 132404 282880 132456
rect 316132 132404 316184 132456
rect 231124 131724 231176 131776
rect 253480 131724 253532 131776
rect 210516 131180 210568 131232
rect 214012 131180 214064 131232
rect 195520 131112 195572 131164
rect 213920 131112 213972 131164
rect 260472 131112 260524 131164
rect 264980 131112 265032 131164
rect 230572 131044 230624 131096
rect 243544 131044 243596 131096
rect 282828 131044 282880 131096
rect 307760 131044 307812 131096
rect 282736 130976 282788 131028
rect 307852 130976 307904 131028
rect 231676 129888 231728 129940
rect 238024 129888 238076 129940
rect 180156 129752 180208 129804
rect 213920 129752 213972 129804
rect 254676 129752 254728 129804
rect 264980 129752 265032 129804
rect 231768 129684 231820 129736
rect 239680 129684 239732 129736
rect 281816 129684 281868 129736
rect 284300 129684 284352 129736
rect 178776 129004 178828 129056
rect 214840 129004 214892 129056
rect 230940 129004 230992 129056
rect 258908 129004 258960 129056
rect 283564 129004 283616 129056
rect 301136 129004 301188 129056
rect 207756 128324 207808 128376
rect 213920 128324 213972 128376
rect 243820 128324 243872 128376
rect 247684 128324 247736 128376
rect 261484 128324 261536 128376
rect 265164 128324 265216 128376
rect 282828 128256 282880 128308
rect 314752 128256 314804 128308
rect 282736 128188 282788 128240
rect 305092 128188 305144 128240
rect 231768 127916 231820 127968
rect 236736 127916 236788 127968
rect 230572 127644 230624 127696
rect 245108 127644 245160 127696
rect 241060 127576 241112 127628
rect 264980 127576 265032 127628
rect 203616 127032 203668 127084
rect 213920 127032 213972 127084
rect 170404 126964 170456 127016
rect 214012 126964 214064 127016
rect 247684 126964 247736 127016
rect 264980 126964 265032 127016
rect 231768 126896 231820 126948
rect 260104 126896 260156 126948
rect 282368 126896 282420 126948
rect 287152 126896 287204 126948
rect 230848 126828 230900 126880
rect 235264 126828 235316 126880
rect 282092 126216 282144 126268
rect 306564 126216 306616 126268
rect 193864 125672 193916 125724
rect 213920 125672 213972 125724
rect 182916 125604 182968 125656
rect 214012 125604 214064 125656
rect 261576 125604 261628 125656
rect 264980 125604 265032 125656
rect 231492 125536 231544 125588
rect 253388 125536 253440 125588
rect 282828 125536 282880 125588
rect 320272 125536 320324 125588
rect 231768 125468 231820 125520
rect 240784 125468 240836 125520
rect 282736 125468 282788 125520
rect 292580 125468 292632 125520
rect 177580 124856 177632 124908
rect 214748 124856 214800 124908
rect 253480 124856 253532 124908
rect 265624 124856 265676 124908
rect 167736 124176 167788 124228
rect 213920 124176 213972 124228
rect 260196 124176 260248 124228
rect 264980 124176 265032 124228
rect 231768 124108 231820 124160
rect 260380 124108 260432 124160
rect 231676 124040 231728 124092
rect 245016 124040 245068 124092
rect 282828 123632 282880 123684
rect 288440 123632 288492 123684
rect 188528 123428 188580 123480
rect 214012 123428 214064 123480
rect 282184 123428 282236 123480
rect 314660 123428 314712 123480
rect 170496 122816 170548 122868
rect 213920 122816 213972 122868
rect 250720 122816 250772 122868
rect 264980 122816 265032 122868
rect 231768 122748 231820 122800
rect 242256 122748 242308 122800
rect 282828 122748 282880 122800
rect 298192 122748 298244 122800
rect 230756 122068 230808 122120
rect 253204 122068 253256 122120
rect 282644 122068 282696 122120
rect 303712 122068 303764 122120
rect 199476 121524 199528 121576
rect 214012 121524 214064 121576
rect 260104 121524 260156 121576
rect 265072 121524 265124 121576
rect 178684 121456 178736 121508
rect 213920 121456 213972 121508
rect 255964 121456 256016 121508
rect 264980 121456 265032 121508
rect 282828 121388 282880 121440
rect 289912 121388 289964 121440
rect 230572 121184 230624 121236
rect 234160 121184 234212 121236
rect 282092 120912 282144 120964
rect 285680 120912 285732 120964
rect 231584 120708 231636 120760
rect 252008 120708 252060 120760
rect 174728 120164 174780 120216
rect 213920 120164 213972 120216
rect 261668 120164 261720 120216
rect 265072 120164 265124 120216
rect 169208 120096 169260 120148
rect 214012 120096 214064 120148
rect 238300 120096 238352 120148
rect 264980 120096 265032 120148
rect 231492 120028 231544 120080
rect 240876 120028 240928 120080
rect 282828 120028 282880 120080
rect 298376 120028 298428 120080
rect 241152 119348 241204 119400
rect 264612 119348 264664 119400
rect 284944 119348 284996 119400
rect 305000 119348 305052 119400
rect 210424 118736 210476 118788
rect 214012 118736 214064 118788
rect 205180 118668 205232 118720
rect 213920 118668 213972 118720
rect 231492 118668 231544 118720
rect 238392 118668 238444 118720
rect 247960 118668 248012 118720
rect 264980 118668 265032 118720
rect 231400 118600 231452 118652
rect 254584 118600 254636 118652
rect 282828 118600 282880 118652
rect 293960 118600 294012 118652
rect 231768 118532 231820 118584
rect 240968 118532 241020 118584
rect 282828 117920 282880 117972
rect 288624 117920 288676 117972
rect 184480 117376 184532 117428
rect 214012 117376 214064 117428
rect 170588 117308 170640 117360
rect 213920 117308 213972 117360
rect 252008 117308 252060 117360
rect 264980 117308 265032 117360
rect 230940 117240 230992 117292
rect 236920 117240 236972 117292
rect 290648 117240 290700 117292
rect 360200 117240 360252 117292
rect 230756 116696 230808 116748
rect 235540 116696 235592 116748
rect 177396 116560 177448 116612
rect 195520 116560 195572 116612
rect 282828 116560 282880 116612
rect 290648 116560 290700 116612
rect 195428 116016 195480 116068
rect 213920 116016 213972 116068
rect 254584 116016 254636 116068
rect 265072 116016 265124 116068
rect 187056 115948 187108 116000
rect 214012 115948 214064 116000
rect 236736 115948 236788 116000
rect 264980 115948 265032 116000
rect 231768 115880 231820 115932
rect 251916 115880 251968 115932
rect 282828 115880 282880 115932
rect 301044 115880 301096 115932
rect 382280 115880 382332 115932
rect 231032 115812 231084 115864
rect 238116 115812 238168 115864
rect 187240 114588 187292 114640
rect 213920 114588 213972 114640
rect 257436 114588 257488 114640
rect 265072 114588 265124 114640
rect 171876 114520 171928 114572
rect 214012 114520 214064 114572
rect 242256 114520 242308 114572
rect 264980 114520 265032 114572
rect 230572 114452 230624 114504
rect 250536 114452 250588 114504
rect 231584 114316 231636 114368
rect 233976 114316 234028 114368
rect 282828 114112 282880 114164
rect 287244 114112 287296 114164
rect 173440 113772 173492 113824
rect 214104 113772 214156 113824
rect 281724 113772 281776 113824
rect 299572 113772 299624 113824
rect 257620 113228 257672 113280
rect 265072 113228 265124 113280
rect 193956 113160 194008 113212
rect 213920 113160 213972 113212
rect 250444 113160 250496 113212
rect 264980 113160 265032 113212
rect 231768 113092 231820 113144
rect 250812 113092 250864 113144
rect 282828 113092 282880 113144
rect 317512 113092 317564 113144
rect 368480 113092 368532 113144
rect 231676 113024 231728 113076
rect 243728 113024 243780 113076
rect 169024 112412 169076 112464
rect 211804 112412 211856 112464
rect 211896 111868 211948 111920
rect 214012 111868 214064 111920
rect 260380 111868 260432 111920
rect 265900 111868 265952 111920
rect 172152 111800 172204 111852
rect 213920 111800 213972 111852
rect 247868 111800 247920 111852
rect 264980 111800 265032 111852
rect 3148 111732 3200 111784
rect 35164 111732 35216 111784
rect 167828 111732 167880 111784
rect 187148 111732 187200 111784
rect 282828 111732 282880 111784
rect 295432 111732 295484 111784
rect 282092 111596 282144 111648
rect 284944 111596 284996 111648
rect 230940 111052 230992 111104
rect 256056 111052 256108 111104
rect 230572 110848 230624 110900
rect 232872 110848 232924 110900
rect 196808 110508 196860 110560
rect 213920 110508 213972 110560
rect 176200 110440 176252 110492
rect 214012 110440 214064 110492
rect 245016 110440 245068 110492
rect 264980 110440 265032 110492
rect 168196 110372 168248 110424
rect 169116 110372 169168 110424
rect 231768 110372 231820 110424
rect 247776 110372 247828 110424
rect 282644 110372 282696 110424
rect 295340 110372 295392 110424
rect 230756 109964 230808 110016
rect 235448 109964 235500 110016
rect 199384 109080 199436 109132
rect 214012 109080 214064 109132
rect 170680 109012 170732 109064
rect 213920 109012 213972 109064
rect 235540 109012 235592 109064
rect 265072 109012 265124 109064
rect 231768 108944 231820 108996
rect 257528 108944 257580 108996
rect 281724 108944 281776 108996
rect 328460 108944 328512 108996
rect 231492 108876 231544 108928
rect 244924 108876 244976 108928
rect 282828 108876 282880 108928
rect 309140 108876 309192 108928
rect 167920 107720 167972 107772
rect 213920 107720 213972 107772
rect 262956 107720 263008 107772
rect 265348 107720 265400 107772
rect 166356 107652 166408 107704
rect 214012 107652 214064 107704
rect 256148 107652 256200 107704
rect 264980 107652 265032 107704
rect 231768 107584 231820 107636
rect 265716 107584 265768 107636
rect 231492 107516 231544 107568
rect 249432 107516 249484 107568
rect 282828 106904 282880 106956
rect 287060 106904 287112 106956
rect 202328 106360 202380 106412
rect 214012 106360 214064 106412
rect 167828 106292 167880 106344
rect 213920 106292 213972 106344
rect 249248 106292 249300 106344
rect 264980 106292 265032 106344
rect 282828 106224 282880 106276
rect 291200 106224 291252 106276
rect 231768 106020 231820 106072
rect 238208 106020 238260 106072
rect 245200 105612 245252 105664
rect 262128 105612 262180 105664
rect 230756 105544 230808 105596
rect 264428 105544 264480 105596
rect 282828 105272 282880 105324
rect 288532 105272 288584 105324
rect 191288 104932 191340 104984
rect 214012 104932 214064 104984
rect 169116 104864 169168 104916
rect 213920 104864 213972 104916
rect 263140 104864 263192 104916
rect 264980 104864 265032 104916
rect 230940 104796 230992 104848
rect 236828 104796 236880 104848
rect 282828 104796 282880 104848
rect 291384 104796 291436 104848
rect 281540 104728 281592 104780
rect 284392 104728 284444 104780
rect 250628 104184 250680 104236
rect 263048 104184 263100 104236
rect 164884 104116 164936 104168
rect 177488 104116 177540 104168
rect 230572 104116 230624 104168
rect 252100 104116 252152 104168
rect 261760 103912 261812 103964
rect 264980 103912 265032 103964
rect 178868 103504 178920 103556
rect 213920 103504 213972 103556
rect 231768 103436 231820 103488
rect 246580 103436 246632 103488
rect 282092 103436 282144 103488
rect 291292 103436 291344 103488
rect 231492 103368 231544 103420
rect 241152 103368 241204 103420
rect 181628 102756 181680 102808
rect 209044 102756 209096 102808
rect 212448 102212 212500 102264
rect 214012 102212 214064 102264
rect 258908 102212 258960 102264
rect 265072 102212 265124 102264
rect 185584 102144 185636 102196
rect 213920 102144 213972 102196
rect 240876 102144 240928 102196
rect 264980 102144 265032 102196
rect 231676 102076 231728 102128
rect 258816 102076 258868 102128
rect 282276 102076 282328 102128
rect 296812 102076 296864 102128
rect 230664 102008 230716 102060
rect 242348 102008 242400 102060
rect 196716 101396 196768 101448
rect 217232 101396 217284 101448
rect 258724 100784 258776 100836
rect 264980 100784 265032 100836
rect 177488 100716 177540 100768
rect 213920 100716 213972 100768
rect 263048 100716 263100 100768
rect 265072 100716 265124 100768
rect 230664 100648 230716 100700
rect 254768 100648 254820 100700
rect 231768 100580 231820 100632
rect 253480 100580 253532 100632
rect 169300 99968 169352 100020
rect 202144 99968 202196 100020
rect 205088 99968 205140 100020
rect 214840 99968 214892 100020
rect 282000 99968 282052 100020
rect 310612 99968 310664 100020
rect 166448 99356 166500 99408
rect 213920 99356 213972 99408
rect 264428 99356 264480 99408
rect 265992 99356 266044 99408
rect 281632 99288 281684 99340
rect 283564 99288 283616 99340
rect 173348 98608 173400 98660
rect 214104 98608 214156 98660
rect 242348 98064 242400 98116
rect 265072 98064 265124 98116
rect 166540 97996 166592 98048
rect 213920 97996 213972 98048
rect 231216 97996 231268 98048
rect 264980 97996 265032 98048
rect 3516 97928 3568 97980
rect 33784 97928 33836 97980
rect 204904 97928 204956 97980
rect 229100 97928 229152 97980
rect 229192 97316 229244 97368
rect 264980 97316 265032 97368
rect 165528 96636 165580 96688
rect 213920 96636 213972 96688
rect 265072 97248 265124 97300
rect 282184 97248 282236 97300
rect 310520 97248 310572 97300
rect 219348 96024 219400 96076
rect 165436 95888 165488 95940
rect 216036 95888 216088 95940
rect 255872 95888 255924 95940
rect 267832 95888 267884 95940
rect 230480 95276 230532 95328
rect 232596 95276 232648 95328
rect 206376 95208 206428 95260
rect 213920 95208 213972 95260
rect 225696 95208 225748 95260
rect 264980 95208 265032 95260
rect 267648 95208 267700 95260
rect 269212 95208 269264 95260
rect 259368 95140 259420 95192
rect 279332 95140 279384 95192
rect 176108 94528 176160 94580
rect 214564 94528 214616 94580
rect 209044 94460 209096 94512
rect 260380 94460 260432 94512
rect 117136 93916 117188 93968
rect 169208 93916 169260 93968
rect 107752 93848 107804 93900
rect 195428 93848 195480 93900
rect 224224 93848 224276 93900
rect 230020 93848 230072 93900
rect 264888 93848 264940 93900
rect 267924 93848 267976 93900
rect 267832 93780 267884 93832
rect 273996 93780 274048 93832
rect 115848 93168 115900 93220
rect 174728 93168 174780 93220
rect 216036 93168 216088 93220
rect 234160 93168 234212 93220
rect 60648 93100 60700 93152
rect 90364 93100 90416 93152
rect 95056 93100 95108 93152
rect 166356 93100 166408 93152
rect 211804 93100 211856 93152
rect 243820 93100 243872 93152
rect 276756 93100 276808 93152
rect 305644 93100 305696 93152
rect 86776 92488 86828 92540
rect 115296 92488 115348 92540
rect 136088 92420 136140 92472
rect 173256 92420 173308 92472
rect 217324 91808 217376 91860
rect 245200 91808 245252 91860
rect 62028 91740 62080 91792
rect 88984 91740 89036 91792
rect 160744 91740 160796 91792
rect 171784 91740 171836 91792
rect 202144 91740 202196 91792
rect 231308 91740 231360 91792
rect 102048 91128 102100 91180
rect 115204 91128 115256 91180
rect 152096 91128 152148 91180
rect 158720 91128 158772 91180
rect 89076 91060 89128 91112
rect 122104 91060 122156 91112
rect 132408 91060 132460 91112
rect 134524 91060 134576 91112
rect 134708 91060 134760 91112
rect 153108 91060 153160 91112
rect 112352 90992 112404 91044
rect 210424 90992 210476 91044
rect 110328 90924 110380 90976
rect 170588 90924 170640 90976
rect 222844 90380 222896 90432
rect 235356 90380 235408 90432
rect 65984 90312 66036 90364
rect 111064 90312 111116 90364
rect 220084 90312 220136 90364
rect 263140 90312 263192 90364
rect 119712 89632 119764 89684
rect 199476 89632 199528 89684
rect 121736 89564 121788 89616
rect 170496 89564 170548 89616
rect 218704 89020 218756 89072
rect 239680 89020 239732 89072
rect 103336 88952 103388 89004
rect 120080 88952 120132 89004
rect 171784 88952 171836 89004
rect 209228 88952 209280 89004
rect 214564 88952 214616 89004
rect 261760 88952 261812 89004
rect 120816 88272 120868 88324
rect 216128 88272 216180 88324
rect 114376 88204 114428 88256
rect 205180 88204 205232 88256
rect 209136 87660 209188 87712
rect 232780 87660 232832 87712
rect 67732 87592 67784 87644
rect 105544 87592 105596 87644
rect 227076 87592 227128 87644
rect 253388 87592 253440 87644
rect 111248 86912 111300 86964
rect 184480 86912 184532 86964
rect 158720 86844 158772 86896
rect 206284 86844 206336 86896
rect 3240 86232 3292 86284
rect 21364 86232 21416 86284
rect 66076 86232 66128 86284
rect 111156 86232 111208 86284
rect 184296 86232 184348 86284
rect 261668 86232 261720 86284
rect 104256 85484 104308 85536
rect 193956 85484 194008 85536
rect 151544 85416 151596 85468
rect 174636 85416 174688 85468
rect 206284 84872 206336 84924
rect 231216 84872 231268 84924
rect 67364 84804 67416 84856
rect 120724 84804 120776 84856
rect 204996 84804 205048 84856
rect 264428 84804 264480 84856
rect 93768 84124 93820 84176
rect 202328 84124 202380 84176
rect 126704 84056 126756 84108
rect 182916 84056 182968 84108
rect 207664 83444 207716 83496
rect 284944 83444 284996 83496
rect 85488 82764 85540 82816
rect 177488 82764 177540 82816
rect 126796 82696 126848 82748
rect 162216 82696 162268 82748
rect 204904 82084 204956 82136
rect 238300 82084 238352 82136
rect 99196 81336 99248 81388
rect 196808 81336 196860 81388
rect 126888 81268 126940 81320
rect 164884 81268 164936 81320
rect 115848 79976 115900 80028
rect 173440 79976 173492 80028
rect 133788 79908 133840 79960
rect 166264 79908 166316 79960
rect 151636 78616 151688 78668
rect 198188 78616 198240 78668
rect 129004 78548 129056 78600
rect 157984 78548 158036 78600
rect 159364 77936 159416 77988
rect 254768 77936 254820 77988
rect 64788 77188 64840 77240
rect 171968 77188 172020 77240
rect 117228 77120 117280 77172
rect 160744 77120 160796 77172
rect 115296 75828 115348 75880
rect 200856 75828 200908 75880
rect 111156 75760 111208 75812
rect 185584 75760 185636 75812
rect 106096 74468 106148 74520
rect 177396 74468 177448 74520
rect 124036 74400 124088 74452
rect 167736 74400 167788 74452
rect 111708 73108 111760 73160
rect 173164 73108 173216 73160
rect 123484 73040 123536 73092
rect 178868 73040 178920 73092
rect 3516 71680 3568 71732
rect 36544 71680 36596 71732
rect 101956 71680 102008 71732
rect 164976 71680 165028 71732
rect 128268 71612 128320 71664
rect 181628 71612 181680 71664
rect 120724 70320 120776 70372
rect 196716 70320 196768 70372
rect 112996 70252 113048 70304
rect 180064 70252 180116 70304
rect 115204 68960 115256 69012
rect 205088 68960 205140 69012
rect 110236 68892 110288 68944
rect 187056 68892 187108 68944
rect 105544 67532 105596 67584
rect 214656 67532 214708 67584
rect 151728 67464 151780 67516
rect 169024 67464 169076 67516
rect 101864 66172 101916 66224
rect 176108 66172 176160 66224
rect 307760 66172 307812 66224
rect 338764 66172 338816 66224
rect 125416 66104 125468 66156
rect 193864 66104 193916 66156
rect 110144 64812 110196 64864
rect 213276 64812 213328 64864
rect 86868 64132 86920 64184
rect 249156 64132 249208 64184
rect 97908 63452 97960 63504
rect 199384 63452 199436 63504
rect 122104 63384 122156 63436
rect 173348 63384 173400 63436
rect 134524 62024 134576 62076
rect 215944 62024 215996 62076
rect 119896 61956 119948 62008
rect 178776 61956 178828 62008
rect 125508 60664 125560 60716
rect 203524 60664 203576 60716
rect 244280 60052 244332 60104
rect 302240 60052 302292 60104
rect 97908 59984 97960 60036
rect 245108 59984 245160 60036
rect 99288 59304 99340 59356
rect 170404 59304 170456 59356
rect 3332 58828 3384 58880
rect 7564 58828 7616 58880
rect 102048 58624 102100 58676
rect 264336 58624 264388 58676
rect 106924 57876 106976 57928
rect 207756 57876 207808 57928
rect 111708 57196 111760 57248
rect 267740 57196 267792 57248
rect 91008 56516 91060 56568
rect 191288 56516 191340 56568
rect 115848 55836 115900 55888
rect 245016 55836 245068 55888
rect 75736 55156 75788 55208
rect 206376 55156 206428 55208
rect 123484 54476 123536 54528
rect 209136 54476 209188 54528
rect 118608 53728 118660 53780
rect 178684 53728 178736 53780
rect 88984 53116 89036 53168
rect 112444 53116 112496 53168
rect 84108 53048 84160 53100
rect 217324 53048 217376 53100
rect 103428 52368 103480 52420
rect 202236 52368 202288 52420
rect 121368 51688 121420 51740
rect 246396 51688 246448 51740
rect 114468 51008 114520 51060
rect 198096 51008 198148 51060
rect 34428 50328 34480 50380
rect 258724 50328 258776 50380
rect 123944 49648 123996 49700
rect 188528 49648 188580 49700
rect 37188 48968 37240 49020
rect 246488 48968 246540 49020
rect 90364 47608 90416 47660
rect 274640 47608 274692 47660
rect 12348 47540 12400 47592
rect 251916 47540 251968 47592
rect 98644 46248 98696 46300
rect 270592 46248 270644 46300
rect 49608 46180 49660 46232
rect 254584 46180 254636 46232
rect 3516 45500 3568 45552
rect 43444 45500 43496 45552
rect 86776 44820 86828 44872
rect 250536 44820 250588 44872
rect 87604 43460 87656 43512
rect 210424 43460 210476 43512
rect 9588 43392 9640 43444
rect 253204 43392 253256 43444
rect 91008 42032 91060 42084
rect 262956 42032 263008 42084
rect 77208 40740 77260 40792
rect 256056 40740 256108 40792
rect 28908 40672 28960 40724
rect 270500 40672 270552 40724
rect 103428 39380 103480 39432
rect 239404 39380 239456 39432
rect 59268 39312 59320 39364
rect 238208 39312 238260 39364
rect 71044 37884 71096 37936
rect 228364 37884 228416 37936
rect 125508 36592 125560 36644
rect 151084 36592 151136 36644
rect 26148 36524 26200 36576
rect 206284 36524 206336 36576
rect 206376 36524 206428 36576
rect 224224 36524 224276 36576
rect 116584 35232 116636 35284
rect 184296 35232 184348 35284
rect 192484 35232 192536 35284
rect 220176 35232 220228 35284
rect 182916 35164 182968 35216
rect 269120 35164 269172 35216
rect 2872 33056 2924 33108
rect 32404 33056 32456 33108
rect 583392 33056 583444 33108
rect 583668 33056 583720 33108
rect 110328 32444 110380 32496
rect 260196 32444 260248 32496
rect 52368 32376 52420 32428
rect 250536 32376 250588 32428
rect 61936 31084 61988 31136
rect 220084 31084 220136 31136
rect 74448 31016 74500 31068
rect 251824 31016 251876 31068
rect 13728 29656 13780 29708
rect 250444 29656 250496 29708
rect 63408 29588 63460 29640
rect 310520 29588 310572 29640
rect 85488 28296 85540 28348
rect 260104 28296 260156 28348
rect 1400 28228 1452 28280
rect 231124 28228 231176 28280
rect 48228 26868 48280 26920
rect 251180 26868 251232 26920
rect 92388 25576 92440 25628
rect 240784 25576 240836 25628
rect 73068 25508 73120 25560
rect 267832 25508 267884 25560
rect 322204 25508 322256 25560
rect 328460 25508 328512 25560
rect 20628 24148 20680 24200
rect 247684 24148 247736 24200
rect 57244 24080 57296 24132
rect 324412 24080 324464 24132
rect 56508 22788 56560 22840
rect 216036 22788 216088 22840
rect 88248 22720 88300 22772
rect 255964 22720 256016 22772
rect 37096 21428 37148 21480
rect 225604 21428 225656 21480
rect 46848 21360 46900 21412
rect 238116 21360 238168 21412
rect 114468 20000 114520 20052
rect 182916 20000 182968 20052
rect 187056 20000 187108 20052
rect 209044 20000 209096 20052
rect 24768 19932 24820 19984
rect 159364 19932 159416 19984
rect 184204 19932 184256 19984
rect 291844 19932 291896 19984
rect 319444 19932 319496 19984
rect 378140 19932 378192 19984
rect 6828 18640 6880 18692
rect 98644 18640 98696 18692
rect 99288 18640 99340 18692
rect 206376 18640 206428 18692
rect 65524 18572 65576 18624
rect 262864 18572 262916 18624
rect 119896 17212 119948 17264
rect 204996 17212 205048 17264
rect 259552 17212 259604 17264
rect 276020 17212 276072 17264
rect 96252 15920 96304 15972
rect 222844 15920 222896 15972
rect 309784 15920 309836 15972
rect 322112 15920 322164 15972
rect 50988 15852 51040 15904
rect 297272 15852 297324 15904
rect 313924 15852 313976 15904
rect 345296 15852 345348 15904
rect 118608 14492 118660 14544
rect 233884 14492 233936 14544
rect 27528 14424 27580 14476
rect 227076 14424 227128 14476
rect 331220 14424 331272 14476
rect 374000 14424 374052 14476
rect 300124 13744 300176 13796
rect 349160 13744 349212 13796
rect 100668 13132 100720 13184
rect 242164 13132 242216 13184
rect 28816 13064 28868 13116
rect 242256 13064 242308 13116
rect 299664 12452 299716 12504
rect 300124 12452 300176 12504
rect 81348 11772 81400 11824
rect 204904 11772 204956 11824
rect 340972 11772 341024 11824
rect 342168 11772 342220 11824
rect 53656 11704 53708 11756
rect 238024 11704 238076 11756
rect 257068 11704 257120 11756
rect 358820 11704 358872 11756
rect 67548 10344 67600 10396
rect 264244 10344 264296 10396
rect 42708 10276 42760 10328
rect 243544 10276 243596 10328
rect 249984 9596 250036 9648
rect 250536 9596 250588 9648
rect 376760 9596 376812 9648
rect 106924 8916 106976 8968
rect 211804 8916 211856 8968
rect 71504 7624 71556 7676
rect 226984 7624 227036 7676
rect 55128 7556 55180 7608
rect 262956 7556 263008 7608
rect 375380 7556 375432 7608
rect 302884 6808 302936 6860
rect 369860 6808 369912 6860
rect 574744 6808 574796 6860
rect 580172 6808 580224 6860
rect 102232 6196 102284 6248
rect 202144 6196 202196 6248
rect 17040 6128 17092 6180
rect 249064 6128 249116 6180
rect 284944 6128 284996 6180
rect 301964 6128 302016 6180
rect 325608 6128 325660 6180
rect 332692 6128 332744 6180
rect 241704 5516 241756 5568
rect 246304 5516 246356 5568
rect 305736 5516 305788 5568
rect 307944 5516 307996 5568
rect 338672 5448 338724 5500
rect 367100 5448 367152 5500
rect 54944 4836 54996 4888
rect 214564 4836 214616 4888
rect 60832 4768 60884 4820
rect 232504 4768 232556 4820
rect 232596 4156 232648 4208
rect 235816 4156 235868 4208
rect 177304 4088 177356 4140
rect 257068 4088 257120 4140
rect 296076 4088 296128 4140
rect 298100 4088 298152 4140
rect 316684 4088 316736 4140
rect 319720 4088 319772 4140
rect 116400 4020 116452 4072
rect 123484 4020 123536 4072
rect 255872 4020 255924 4072
rect 282184 4020 282236 4072
rect 310244 4020 310296 4072
rect 317420 4020 317472 4072
rect 63224 3816 63276 3868
rect 65524 3816 65576 3868
rect 305552 3748 305604 3800
rect 306472 3748 306524 3800
rect 2872 3544 2924 3596
rect 3976 3544 4028 3596
rect 8760 3476 8812 3528
rect 9588 3476 9640 3528
rect 9956 3476 10008 3528
rect 10968 3476 11020 3528
rect 15936 3476 15988 3528
rect 16488 3476 16540 3528
rect 18236 3476 18288 3528
rect 19248 3476 19300 3528
rect 24216 3476 24268 3528
rect 24768 3476 24820 3528
rect 25320 3476 25372 3528
rect 26148 3476 26200 3528
rect 26516 3476 26568 3528
rect 27528 3476 27580 3528
rect 27712 3476 27764 3528
rect 28816 3476 28868 3528
rect 32404 3476 32456 3528
rect 33048 3476 33100 3528
rect 33600 3476 33652 3528
rect 34428 3476 34480 3528
rect 34796 3476 34848 3528
rect 35808 3476 35860 3528
rect 35992 3476 36044 3528
rect 37096 3476 37148 3528
rect 40684 3476 40736 3528
rect 41328 3476 41380 3528
rect 41880 3476 41932 3528
rect 42708 3476 42760 3528
rect 43076 3476 43128 3528
rect 44088 3476 44140 3528
rect 44272 3476 44324 3528
rect 71044 3612 71096 3664
rect 70216 3544 70268 3596
rect 87604 3612 87656 3664
rect 85672 3544 85724 3596
rect 86776 3544 86828 3596
rect 95056 3544 95108 3596
rect 66720 3476 66772 3528
rect 67548 3476 67600 3528
rect 67916 3476 67968 3528
rect 68928 3476 68980 3528
rect 69112 3476 69164 3528
rect 70308 3476 70360 3528
rect 72608 3476 72660 3528
rect 73068 3476 73120 3528
rect 73804 3476 73856 3528
rect 74448 3476 74500 3528
rect 76196 3476 76248 3528
rect 77208 3476 77260 3528
rect 80888 3476 80940 3528
rect 81348 3476 81400 3528
rect 84476 3476 84528 3528
rect 85488 3476 85540 3528
rect 89168 3476 89220 3528
rect 89628 3476 89680 3528
rect 90364 3476 90416 3528
rect 91008 3476 91060 3528
rect 91560 3476 91612 3528
rect 92388 3476 92440 3528
rect 92756 3476 92808 3528
rect 93768 3476 93820 3528
rect 93952 3476 94004 3528
rect 95148 3476 95200 3528
rect 97448 3476 97500 3528
rect 97908 3476 97960 3528
rect 98644 3476 98696 3528
rect 99288 3476 99340 3528
rect 99840 3476 99892 3528
rect 100668 3476 100720 3528
rect 101036 3476 101088 3528
rect 102048 3476 102100 3528
rect 126244 3544 126296 3596
rect 124680 3476 124732 3528
rect 125508 3476 125560 3528
rect 129372 3476 129424 3528
rect 130384 3476 130436 3528
rect 291844 3476 291896 3528
rect 292580 3476 292632 3528
rect 307760 3476 307812 3528
rect 309048 3476 309100 3528
rect 324320 3476 324372 3528
rect 325608 3476 325660 3528
rect 336004 3476 336056 3528
rect 337476 3476 337528 3528
rect 349252 3476 349304 3528
rect 357440 3476 357492 3528
rect 581000 3476 581052 3528
rect 583484 3476 583536 3528
rect 20536 3408 20588 3460
rect 48964 3408 49016 3460
rect 49608 3408 49660 3460
rect 52552 3408 52604 3460
rect 53656 3408 53708 3460
rect 56048 3408 56100 3460
rect 56508 3408 56560 3460
rect 57244 3408 57296 3460
rect 57888 3408 57940 3460
rect 58440 3408 58492 3460
rect 59268 3408 59320 3460
rect 59636 3408 59688 3460
rect 60648 3408 60700 3460
rect 64328 3408 64380 3460
rect 64788 3408 64840 3460
rect 83280 3408 83332 3460
rect 84108 3408 84160 3460
rect 61384 3340 61436 3392
rect 77392 3340 77444 3392
rect 105728 3408 105780 3460
rect 106188 3408 106240 3460
rect 108120 3408 108172 3460
rect 108948 3408 109000 3460
rect 109316 3408 109368 3460
rect 110328 3408 110380 3460
rect 114008 3408 114060 3460
rect 114468 3408 114520 3460
rect 115204 3408 115256 3460
rect 115848 3408 115900 3460
rect 117596 3408 117648 3460
rect 118608 3408 118660 3460
rect 118792 3408 118844 3460
rect 119804 3408 119856 3460
rect 122288 3408 122340 3460
rect 122748 3408 122800 3460
rect 123484 3408 123536 3460
rect 187056 3408 187108 3460
rect 195244 3408 195296 3460
rect 246396 3408 246448 3460
rect 288992 3408 289044 3460
rect 296720 3408 296772 3460
rect 323584 3408 323636 3460
rect 348056 3408 348108 3460
rect 350448 3408 350500 3460
rect 360292 3408 360344 3460
rect 116584 3340 116636 3392
rect 582196 3272 582248 3324
rect 583576 3272 583628 3324
rect 75000 3204 75052 3256
rect 75828 3204 75880 3256
rect 268384 3136 268436 3188
rect 276020 3136 276072 3188
rect 280804 3136 280856 3188
rect 283104 3136 283156 3188
rect 337384 3136 337436 3188
rect 339868 3136 339920 3188
rect 11152 3000 11204 3052
rect 15844 3000 15896 3052
rect 50160 3000 50212 3052
rect 50896 3000 50948 3052
rect 82084 3000 82136 3052
rect 82728 3000 82780 3052
rect 110512 3000 110564 3052
rect 111524 3000 111576 3052
rect 19432 2932 19484 2984
rect 20628 2932 20680 2984
rect 309876 2932 309928 2984
rect 315028 2932 315080 2984
rect 112812 2116 112864 2168
rect 218704 2116 218756 2168
rect 220176 2116 220228 2168
rect 240508 2116 240560 2168
rect 51356 2048 51408 2100
rect 58624 2048 58676 2100
rect 65524 2048 65576 2100
rect 233976 2048 234028 2100
rect 253204 2048 253256 2100
rect 272432 2048 272484 2100
rect 331864 2048 331916 2100
rect 340972 2048 341024 2100
rect 332600 552 332652 604
rect 333888 552 333940 604
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40052 703582 40356 703610
rect 8128 702506 8156 703520
rect 8116 702500 8168 702506
rect 8116 702442 8168 702448
rect 24320 699718 24348 703520
rect 24308 699712 24360 699718
rect 24308 699654 24360 699660
rect 25504 699712 25556 699718
rect 25504 699654 25556 699660
rect 3422 684312 3478 684321
rect 3422 684247 3478 684256
rect 3436 683194 3464 684247
rect 3424 683188 3476 683194
rect 3424 683130 3476 683136
rect 11704 683188 11756 683194
rect 11704 683130 11756 683136
rect 3514 671256 3570 671265
rect 3514 671191 3570 671200
rect 3528 670750 3556 671191
rect 3516 670744 3568 670750
rect 3516 670686 3568 670692
rect 3422 658200 3478 658209
rect 3422 658135 3424 658144
rect 3476 658135 3478 658144
rect 7564 658164 7616 658170
rect 3424 658106 3476 658112
rect 7564 658106 7616 658112
rect 3424 632120 3476 632126
rect 3422 632088 3424 632097
rect 3476 632088 3478 632097
rect 3422 632023 3478 632032
rect 3146 619168 3202 619177
rect 3146 619103 3202 619112
rect 3160 618322 3188 619103
rect 3148 618316 3200 618322
rect 3148 618258 3200 618264
rect 3238 606112 3294 606121
rect 3238 606047 3294 606056
rect 3252 605878 3280 606047
rect 3240 605872 3292 605878
rect 3240 605814 3292 605820
rect 7576 591326 7604 658106
rect 7564 591320 7616 591326
rect 7564 591262 7616 591268
rect 3424 589348 3476 589354
rect 3424 589290 3476 589296
rect 3436 580009 3464 589290
rect 3422 580000 3478 580009
rect 3422 579935 3478 579944
rect 3422 566944 3478 566953
rect 3422 566879 3478 566888
rect 3436 565894 3464 566879
rect 3424 565888 3476 565894
rect 3424 565830 3476 565836
rect 3422 553888 3478 553897
rect 3422 553823 3478 553832
rect 3436 540258 3464 553823
rect 11716 543046 11744 683130
rect 14464 670744 14516 670750
rect 14464 670686 14516 670692
rect 11704 543040 11756 543046
rect 11704 542982 11756 542988
rect 14476 541686 14504 670686
rect 17224 632120 17276 632126
rect 17224 632062 17276 632068
rect 15844 618316 15896 618322
rect 15844 618258 15896 618264
rect 14464 541680 14516 541686
rect 14464 541622 14516 541628
rect 3424 540252 3476 540258
rect 3424 540194 3476 540200
rect 3424 538892 3476 538898
rect 3424 538834 3476 538840
rect 3436 527921 3464 538834
rect 8208 537532 8260 537538
rect 8208 537474 8260 537480
rect 3422 527912 3478 527921
rect 3422 527847 3478 527856
rect 2778 514856 2834 514865
rect 2778 514791 2780 514800
rect 2832 514791 2834 514800
rect 2780 514762 2832 514768
rect 3330 475688 3386 475697
rect 3330 475623 3386 475632
rect 3344 475386 3372 475623
rect 3332 475380 3384 475386
rect 3332 475322 3384 475328
rect 3436 451926 3464 527847
rect 4804 514820 4856 514826
rect 4804 514762 4856 514768
rect 3516 502308 3568 502314
rect 3516 502250 3568 502256
rect 3528 501809 3556 502250
rect 3514 501800 3570 501809
rect 3514 501735 3570 501744
rect 3514 462632 3570 462641
rect 3514 462567 3570 462576
rect 3528 462398 3556 462567
rect 3516 462392 3568 462398
rect 3516 462334 3568 462340
rect 4816 459542 4844 514762
rect 8220 475386 8248 537474
rect 15856 536110 15884 618258
rect 17236 576162 17264 632062
rect 25516 592686 25544 699654
rect 40052 594114 40080 703582
rect 40328 703474 40356 703582
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 412652 703582 413508 703610
rect 40512 703474 40540 703520
rect 40328 703446 40540 703474
rect 62028 702908 62080 702914
rect 62028 702850 62080 702856
rect 40040 594108 40092 594114
rect 40040 594050 40092 594056
rect 25504 592680 25556 592686
rect 25504 592622 25556 592628
rect 55036 587920 55088 587926
rect 55036 587862 55088 587868
rect 48136 582412 48188 582418
rect 48136 582354 48188 582360
rect 17224 576156 17276 576162
rect 17224 576098 17276 576104
rect 43444 565888 43496 565894
rect 43444 565830 43496 565836
rect 41328 560312 41380 560318
rect 41328 560254 41380 560260
rect 36544 543040 36596 543046
rect 36544 542982 36596 542988
rect 36556 542434 36584 542982
rect 36544 542428 36596 542434
rect 36544 542370 36596 542376
rect 37188 542428 37240 542434
rect 37188 542370 37240 542376
rect 15844 536104 15896 536110
rect 15844 536046 15896 536052
rect 11704 534744 11756 534750
rect 11704 534686 11756 534692
rect 11716 502314 11744 534686
rect 17868 532024 17920 532030
rect 17868 531966 17920 531972
rect 11704 502308 11756 502314
rect 11704 502250 11756 502256
rect 8208 475380 8260 475386
rect 8208 475322 8260 475328
rect 14556 462392 14608 462398
rect 14556 462334 14608 462340
rect 4804 459536 4856 459542
rect 4804 459478 4856 459484
rect 3424 451920 3476 451926
rect 3424 451862 3476 451868
rect 3146 449576 3202 449585
rect 3146 449511 3202 449520
rect 3160 448594 3188 449511
rect 14568 449206 14596 462334
rect 17880 454034 17908 531966
rect 35806 526416 35862 526425
rect 35806 526351 35862 526360
rect 34428 525088 34480 525094
rect 34428 525030 34480 525036
rect 25504 475380 25556 475386
rect 25504 475322 25556 475328
rect 17224 454028 17276 454034
rect 17224 453970 17276 453976
rect 17868 454028 17920 454034
rect 17868 453970 17920 453976
rect 17236 452674 17264 453970
rect 17224 452668 17276 452674
rect 17224 452610 17276 452616
rect 14556 449200 14608 449206
rect 14556 449142 14608 449148
rect 3148 448588 3200 448594
rect 3148 448530 3200 448536
rect 14464 448588 14516 448594
rect 14464 448530 14516 448536
rect 4804 444440 4856 444446
rect 4804 444382 4856 444388
rect 3424 423632 3476 423638
rect 3422 423600 3424 423609
rect 3476 423600 3478 423609
rect 3422 423535 3478 423544
rect 3422 410544 3478 410553
rect 3422 410479 3478 410488
rect 2780 398744 2832 398750
rect 2780 398686 2832 398692
rect 2792 397497 2820 398686
rect 2778 397488 2834 397497
rect 2778 397423 2834 397432
rect 3436 391270 3464 410479
rect 4816 398750 4844 444382
rect 4804 398744 4856 398750
rect 4804 398686 4856 398692
rect 3424 391264 3476 391270
rect 3424 391206 3476 391212
rect 11704 387116 11756 387122
rect 11704 387058 11756 387064
rect 3424 385688 3476 385694
rect 3424 385630 3476 385636
rect 3436 383654 3464 385630
rect 3436 383626 3556 383654
rect 3528 371385 3556 383626
rect 4802 381032 4858 381041
rect 4802 380967 4858 380976
rect 3514 371376 3570 371385
rect 3514 371311 3570 371320
rect 3332 358760 3384 358766
rect 3332 358702 3384 358708
rect 3344 358465 3372 358702
rect 3330 358456 3386 358465
rect 3330 358391 3386 358400
rect 2780 346316 2832 346322
rect 2780 346258 2832 346264
rect 2792 345409 2820 346258
rect 2778 345400 2834 345409
rect 2778 345335 2834 345344
rect 3424 334008 3476 334014
rect 3424 333950 3476 333956
rect 20 333260 72 333266
rect 20 333202 72 333208
rect 32 6905 60 333202
rect 3332 267776 3384 267782
rect 3332 267718 3384 267724
rect 3344 267209 3372 267718
rect 3330 267200 3386 267209
rect 3330 267135 3386 267144
rect 3148 255264 3200 255270
rect 3148 255206 3200 255212
rect 3160 254153 3188 255206
rect 3146 254144 3202 254153
rect 3146 254079 3202 254088
rect 3436 214985 3464 333950
rect 3528 321570 3556 371311
rect 4816 346322 4844 380967
rect 4804 346316 4856 346322
rect 4804 346258 4856 346264
rect 7564 328500 7616 328506
rect 7564 328442 7616 328448
rect 3516 321564 3568 321570
rect 3516 321506 3568 321512
rect 4068 319456 4120 319462
rect 4068 319398 4120 319404
rect 4080 319297 4108 319398
rect 4066 319288 4122 319297
rect 4066 319223 4122 319232
rect 3516 306332 3568 306338
rect 3516 306274 3568 306280
rect 3528 306241 3556 306274
rect 3514 306232 3570 306241
rect 3514 306167 3570 306176
rect 3514 293176 3570 293185
rect 3514 293111 3570 293120
rect 3528 292602 3556 293111
rect 3516 292596 3568 292602
rect 3516 292538 3568 292544
rect 4080 269822 4108 319223
rect 4068 269816 4120 269822
rect 4068 269758 4120 269764
rect 3516 241460 3568 241466
rect 3516 241402 3568 241408
rect 3528 241097 3556 241402
rect 3514 241088 3570 241097
rect 3514 241023 3570 241032
rect 3422 214976 3478 214985
rect 3422 214911 3478 214920
rect 3424 202836 3476 202842
rect 3424 202778 3476 202784
rect 3436 201929 3464 202778
rect 3422 201920 3478 201929
rect 3422 201855 3478 201864
rect 3424 200796 3476 200802
rect 3424 200738 3476 200744
rect 3240 164212 3292 164218
rect 3240 164154 3292 164160
rect 3252 162897 3280 164154
rect 3238 162888 3294 162897
rect 3238 162823 3294 162832
rect 3148 111784 3200 111790
rect 3148 111726 3200 111732
rect 3160 110673 3188 111726
rect 3146 110664 3202 110673
rect 3146 110599 3202 110608
rect 3240 86284 3292 86290
rect 3240 86226 3292 86232
rect 3252 84697 3280 86226
rect 3238 84688 3294 84697
rect 3238 84623 3294 84632
rect 3332 58880 3384 58886
rect 3332 58822 3384 58828
rect 3344 58585 3372 58822
rect 3330 58576 3386 58585
rect 3330 58511 3386 58520
rect 2872 33108 2924 33114
rect 2872 33050 2924 33056
rect 2884 32473 2912 33050
rect 2870 32464 2926 32473
rect 2870 32399 2926 32408
rect 1400 28280 1452 28286
rect 1400 28222 1452 28228
rect 1412 16574 1440 28222
rect 3436 19417 3464 200738
rect 3516 189032 3568 189038
rect 3516 188974 3568 188980
rect 3528 188873 3556 188974
rect 3514 188864 3570 188873
rect 3514 188799 3570 188808
rect 3516 150408 3568 150414
rect 3516 150350 3568 150356
rect 3528 149841 3556 150350
rect 3514 149832 3570 149841
rect 3514 149767 3570 149776
rect 3516 137964 3568 137970
rect 3516 137906 3568 137912
rect 3528 136785 3556 137906
rect 3514 136776 3570 136785
rect 3514 136711 3570 136720
rect 3516 97980 3568 97986
rect 3516 97922 3568 97928
rect 3528 97617 3556 97922
rect 3514 97608 3570 97617
rect 3514 97543 3570 97552
rect 5446 79384 5502 79393
rect 5446 79319 5502 79328
rect 3516 71732 3568 71738
rect 3516 71674 3568 71680
rect 3528 71641 3556 71674
rect 3514 71632 3570 71641
rect 3514 71567 3570 71576
rect 3516 45552 3568 45558
rect 3514 45520 3516 45529
rect 3568 45520 3570 45529
rect 3514 45455 3570 45464
rect 4066 35184 4122 35193
rect 4066 35119 4122 35128
rect 3422 19408 3478 19417
rect 3422 19343 3478 19352
rect 3974 17232 4030 17241
rect 3974 17167 4030 17176
rect 3988 16574 4016 17167
rect 1412 16546 1716 16574
rect 570 8936 626 8945
rect 570 8871 626 8880
rect 18 6896 74 6905
rect 18 6831 74 6840
rect 584 480 612 8871
rect 1688 480 1716 16546
rect 3896 16546 4016 16574
rect 2872 3596 2924 3602
rect 2872 3538 2924 3544
rect 2884 480 2912 3538
rect 3896 3482 3924 16546
rect 4080 6914 4108 35119
rect 5460 6914 5488 79319
rect 7576 58886 7604 328442
rect 11716 319462 11744 387058
rect 11704 319456 11756 319462
rect 11704 319398 11756 319404
rect 14476 293962 14504 448530
rect 17236 423638 17264 452610
rect 22744 428460 22796 428466
rect 22744 428402 22796 428408
rect 17224 423632 17276 423638
rect 17224 423574 17276 423580
rect 15842 383752 15898 383761
rect 15842 383687 15898 383696
rect 15856 358766 15884 383687
rect 15844 358760 15896 358766
rect 15844 358702 15896 358708
rect 17222 330032 17278 330041
rect 17222 329967 17278 329976
rect 15844 316736 15896 316742
rect 15844 316678 15896 316684
rect 14464 293956 14516 293962
rect 14464 293898 14516 293904
rect 14556 292596 14608 292602
rect 14556 292538 14608 292544
rect 11704 269816 11756 269822
rect 11704 269758 11756 269764
rect 11716 262206 11744 269758
rect 11704 262200 11756 262206
rect 11704 262142 11756 262148
rect 14568 237386 14596 292538
rect 14556 237380 14608 237386
rect 14556 237322 14608 237328
rect 11704 235272 11756 235278
rect 11704 235214 11756 235220
rect 11716 150414 11744 235214
rect 15856 189038 15884 316678
rect 15844 189032 15896 189038
rect 15844 188974 15896 188980
rect 11704 150408 11756 150414
rect 11704 150350 11756 150356
rect 17236 137970 17264 329967
rect 18604 311160 18656 311166
rect 18604 311102 18656 311108
rect 18616 255270 18644 311102
rect 21364 280220 21416 280226
rect 21364 280162 21416 280168
rect 18604 255264 18656 255270
rect 18604 255206 18656 255212
rect 17224 137964 17276 137970
rect 17224 137906 17276 137912
rect 21376 86290 21404 280162
rect 22756 267782 22784 428402
rect 25516 389230 25544 475322
rect 25504 389224 25556 389230
rect 25504 389166 25556 389172
rect 25504 349852 25556 349858
rect 25504 349794 25556 349800
rect 22744 267776 22796 267782
rect 22744 267718 22796 267724
rect 22756 234598 22784 267718
rect 25516 241466 25544 349794
rect 33784 331900 33836 331906
rect 33784 331842 33836 331848
rect 32404 329112 32456 329118
rect 32404 329054 32456 329060
rect 32416 306338 32444 329054
rect 32404 306332 32456 306338
rect 32404 306274 32456 306280
rect 25504 241460 25556 241466
rect 25504 241402 25556 241408
rect 22744 234592 22796 234598
rect 22744 234534 22796 234540
rect 32402 222864 32458 222873
rect 32402 222799 32458 222808
rect 21364 86284 21416 86290
rect 21364 86226 21416 86232
rect 30286 83464 30342 83473
rect 30286 83399 30342 83408
rect 15842 80744 15898 80753
rect 15842 80679 15898 80688
rect 15106 61432 15162 61441
rect 15106 61367 15162 61376
rect 7564 58880 7616 58886
rect 7564 58822 7616 58828
rect 12348 47592 12400 47598
rect 12348 47534 12400 47540
rect 9588 43444 9640 43450
rect 9588 43386 9640 43392
rect 6828 18692 6880 18698
rect 6828 18634 6880 18640
rect 6840 6914 6868 18634
rect 3988 6886 4108 6914
rect 5276 6886 5488 6914
rect 6472 6886 6868 6914
rect 3988 3602 4016 6886
rect 3976 3596 4028 3602
rect 3976 3538 4028 3544
rect 3896 3454 4108 3482
rect 4080 480 4108 3454
rect 5276 480 5304 6886
rect 6472 480 6500 6886
rect 9600 3534 9628 43386
rect 10966 42120 11022 42129
rect 10966 42055 11022 42064
rect 10980 3534 11008 42055
rect 8760 3528 8812 3534
rect 8760 3470 8812 3476
rect 9588 3528 9640 3534
rect 9588 3470 9640 3476
rect 9956 3528 10008 3534
rect 9956 3470 10008 3476
rect 10968 3528 11020 3534
rect 10968 3470 11020 3476
rect 7654 3360 7710 3369
rect 7654 3295 7710 3304
rect 7668 480 7696 3295
rect 8772 480 8800 3470
rect 9968 480 9996 3470
rect 11152 3052 11204 3058
rect 11152 2994 11204 3000
rect 11164 480 11192 2994
rect 12360 480 12388 47534
rect 13728 29708 13780 29714
rect 13728 29650 13780 29656
rect 13740 6914 13768 29650
rect 15120 6914 15148 61367
rect 13556 6886 13768 6914
rect 14752 6886 15148 6914
rect 13556 480 13584 6886
rect 14752 480 14780 6886
rect 15856 3058 15884 80679
rect 19246 75304 19302 75313
rect 19246 75239 19302 75248
rect 16486 33824 16542 33833
rect 16486 33759 16542 33768
rect 16500 3534 16528 33759
rect 17040 6180 17092 6186
rect 17040 6122 17092 6128
rect 15936 3528 15988 3534
rect 15936 3470 15988 3476
rect 16488 3528 16540 3534
rect 16488 3470 16540 3476
rect 15844 3052 15896 3058
rect 15844 2994 15896 3000
rect 15948 480 15976 3470
rect 17052 480 17080 6122
rect 19260 3534 19288 75239
rect 23386 54496 23442 54505
rect 23386 54431 23442 54440
rect 22006 51776 22062 51785
rect 22006 51711 22062 51720
rect 20628 24200 20680 24206
rect 20628 24142 20680 24148
rect 18236 3528 18288 3534
rect 18236 3470 18288 3476
rect 19248 3528 19300 3534
rect 19248 3470 19300 3476
rect 18248 480 18276 3470
rect 20536 3460 20588 3466
rect 20536 3402 20588 3408
rect 19432 2984 19484 2990
rect 19432 2926 19484 2932
rect 19444 480 19472 2926
rect 20548 1714 20576 3402
rect 20640 2990 20668 24142
rect 22020 6914 22048 51711
rect 23400 6914 23428 54431
rect 28908 40724 28960 40730
rect 28908 40666 28960 40672
rect 26148 36576 26200 36582
rect 26148 36518 26200 36524
rect 24768 19984 24820 19990
rect 24768 19926 24820 19932
rect 21836 6886 22048 6914
rect 23032 6886 23428 6914
rect 20628 2984 20680 2990
rect 20628 2926 20680 2932
rect 20548 1686 20668 1714
rect 20640 480 20668 1686
rect 21836 480 21864 6886
rect 23032 480 23060 6886
rect 24780 3534 24808 19926
rect 26160 3534 26188 36518
rect 27528 14476 27580 14482
rect 27528 14418 27580 14424
rect 27540 3534 27568 14418
rect 28816 13116 28868 13122
rect 28816 13058 28868 13064
rect 28828 3534 28856 13058
rect 24216 3528 24268 3534
rect 24216 3470 24268 3476
rect 24768 3528 24820 3534
rect 24768 3470 24820 3476
rect 25320 3528 25372 3534
rect 25320 3470 25372 3476
rect 26148 3528 26200 3534
rect 26148 3470 26200 3476
rect 26516 3528 26568 3534
rect 26516 3470 26568 3476
rect 27528 3528 27580 3534
rect 27528 3470 27580 3476
rect 27712 3528 27764 3534
rect 27712 3470 27764 3476
rect 28816 3528 28868 3534
rect 28816 3470 28868 3476
rect 24228 480 24256 3470
rect 25332 480 25360 3470
rect 26528 480 26556 3470
rect 27724 480 27752 3470
rect 28920 480 28948 40666
rect 30300 6914 30328 83399
rect 31666 55856 31722 55865
rect 31666 55791 31722 55800
rect 31680 6914 31708 55791
rect 32416 33114 32444 222799
rect 33796 97986 33824 331842
rect 34440 318782 34468 525030
rect 34428 318776 34480 318782
rect 34428 318718 34480 318724
rect 35820 274650 35848 526351
rect 37200 396778 37228 542370
rect 41340 531282 41368 560254
rect 43456 536790 43484 565830
rect 43444 536784 43496 536790
rect 43444 536726 43496 536732
rect 43996 536104 44048 536110
rect 43996 536046 44048 536052
rect 41328 531276 41380 531282
rect 41328 531218 41380 531224
rect 39948 518220 40000 518226
rect 39948 518162 40000 518168
rect 37188 396772 37240 396778
rect 37188 396714 37240 396720
rect 39854 384296 39910 384305
rect 39854 384231 39910 384240
rect 36544 309800 36596 309806
rect 36544 309742 36596 309748
rect 35808 274644 35860 274650
rect 35808 274586 35860 274592
rect 35164 214600 35216 214606
rect 35164 214542 35216 214548
rect 35176 111790 35204 214542
rect 35164 111784 35216 111790
rect 35164 111726 35216 111732
rect 33784 97980 33836 97986
rect 33784 97922 33836 97928
rect 36556 71738 36584 309742
rect 39868 262886 39896 384231
rect 39856 262880 39908 262886
rect 39856 262822 39908 262828
rect 39960 238649 39988 518162
rect 41340 425746 41368 531218
rect 41328 425740 41380 425746
rect 41328 425682 41380 425688
rect 41326 415440 41382 415449
rect 41326 415375 41382 415384
rect 40684 295384 40736 295390
rect 40684 295326 40736 295332
rect 39946 238640 40002 238649
rect 39946 238575 40002 238584
rect 40696 164218 40724 295326
rect 41340 290494 41368 415375
rect 44008 389162 44036 536046
rect 48148 532778 48176 582354
rect 52276 579692 52328 579698
rect 52276 579634 52328 579640
rect 50896 564460 50948 564466
rect 50896 564402 50948 564408
rect 49608 554056 49660 554062
rect 49608 553998 49660 554004
rect 48228 545148 48280 545154
rect 48228 545090 48280 545096
rect 48136 532772 48188 532778
rect 48136 532714 48188 532720
rect 46848 520940 46900 520946
rect 46848 520882 46900 520888
rect 45468 514072 45520 514078
rect 45468 514014 45520 514020
rect 44088 401600 44140 401606
rect 44088 401542 44140 401548
rect 43996 389156 44048 389162
rect 43996 389098 44048 389104
rect 41328 290488 41380 290494
rect 41328 290430 41380 290436
rect 44100 240106 44128 401542
rect 45480 287026 45508 514014
rect 45468 287020 45520 287026
rect 45468 286962 45520 286968
rect 46860 257961 46888 520882
rect 48148 450566 48176 532714
rect 48136 450560 48188 450566
rect 48136 450502 48188 450508
rect 48044 446412 48096 446418
rect 48044 446354 48096 446360
rect 48056 358766 48084 446354
rect 48240 401606 48268 545090
rect 49620 415342 49648 553998
rect 50804 436144 50856 436150
rect 50804 436086 50856 436092
rect 49608 415336 49660 415342
rect 49608 415278 49660 415284
rect 48228 401600 48280 401606
rect 48228 401542 48280 401548
rect 48228 398132 48280 398138
rect 48228 398074 48280 398080
rect 48240 376038 48268 398074
rect 50816 383654 50844 436086
rect 50908 433294 50936 564402
rect 50988 563100 51040 563106
rect 50988 563042 51040 563048
rect 50896 433288 50948 433294
rect 50896 433230 50948 433236
rect 51000 431254 51028 563042
rect 52288 461650 52316 579634
rect 53104 566500 53156 566506
rect 53104 566442 53156 566448
rect 52368 561740 52420 561746
rect 52368 561682 52420 561688
rect 52276 461644 52328 461650
rect 52276 461586 52328 461592
rect 52276 456816 52328 456822
rect 52276 456758 52328 456764
rect 50988 431248 51040 431254
rect 50988 431190 51040 431196
rect 51080 429140 51132 429146
rect 51080 429082 51132 429088
rect 51092 428466 51120 429082
rect 51080 428460 51132 428466
rect 51080 428402 51132 428408
rect 50988 421592 51040 421598
rect 50988 421534 51040 421540
rect 50816 383626 50936 383654
rect 50908 380934 50936 383626
rect 50896 380928 50948 380934
rect 50896 380870 50948 380876
rect 49608 380180 49660 380186
rect 49608 380122 49660 380128
rect 48228 376032 48280 376038
rect 48228 375974 48280 375980
rect 48240 373994 48268 375974
rect 48148 373966 48268 373994
rect 47584 358760 47636 358766
rect 47584 358702 47636 358708
rect 48044 358760 48096 358766
rect 48044 358702 48096 358708
rect 47596 358086 47624 358702
rect 47584 358080 47636 358086
rect 47584 358022 47636 358028
rect 47596 329118 47624 358022
rect 47584 329112 47636 329118
rect 47584 329054 47636 329060
rect 46846 257952 46902 257961
rect 46846 257887 46902 257896
rect 48148 240145 48176 373966
rect 48228 284980 48280 284986
rect 48228 284922 48280 284928
rect 48134 240136 48190 240145
rect 44088 240100 44140 240106
rect 48134 240071 48190 240080
rect 44088 240042 44140 240048
rect 43442 221504 43498 221513
rect 43442 221439 43498 221448
rect 40684 164212 40736 164218
rect 40684 164154 40736 164160
rect 41326 77888 41382 77897
rect 41326 77823 41382 77832
rect 36544 71732 36596 71738
rect 36544 71674 36596 71680
rect 38566 58576 38622 58585
rect 38566 58511 38622 58520
rect 35806 57216 35862 57225
rect 35806 57151 35862 57160
rect 34428 50380 34480 50386
rect 34428 50322 34480 50328
rect 33046 36544 33102 36553
rect 33046 36479 33102 36488
rect 32404 33108 32456 33114
rect 32404 33050 32456 33056
rect 30116 6886 30328 6914
rect 31312 6886 31708 6914
rect 30116 480 30144 6886
rect 31312 480 31340 6886
rect 33060 3534 33088 36479
rect 34440 3534 34468 50322
rect 35820 3534 35848 57151
rect 37188 49020 37240 49026
rect 37188 48962 37240 48968
rect 37096 21480 37148 21486
rect 37096 21422 37148 21428
rect 37108 3534 37136 21422
rect 32404 3528 32456 3534
rect 32404 3470 32456 3476
rect 33048 3528 33100 3534
rect 33048 3470 33100 3476
rect 33600 3528 33652 3534
rect 33600 3470 33652 3476
rect 34428 3528 34480 3534
rect 34428 3470 34480 3476
rect 34796 3528 34848 3534
rect 34796 3470 34848 3476
rect 35808 3528 35860 3534
rect 35808 3470 35860 3476
rect 35992 3528 36044 3534
rect 35992 3470 36044 3476
rect 37096 3528 37148 3534
rect 37096 3470 37148 3476
rect 32416 480 32444 3470
rect 33612 480 33640 3470
rect 34808 480 34836 3470
rect 36004 480 36032 3470
rect 37200 480 37228 48962
rect 38580 6914 38608 58511
rect 39946 48920 40002 48929
rect 39946 48855 40002 48864
rect 39960 6914 39988 48855
rect 38396 6886 38608 6914
rect 39592 6886 39988 6914
rect 38396 480 38424 6886
rect 39592 480 39620 6886
rect 41340 3534 41368 77823
rect 43456 45558 43484 221439
rect 48134 65512 48190 65521
rect 48134 65447 48190 65456
rect 45466 59936 45522 59945
rect 45466 59871 45522 59880
rect 44086 50280 44142 50289
rect 44086 50215 44142 50224
rect 43444 45552 43496 45558
rect 43444 45494 43496 45500
rect 42708 10328 42760 10334
rect 42708 10270 42760 10276
rect 42720 3534 42748 10270
rect 44100 3534 44128 50215
rect 40684 3528 40736 3534
rect 40684 3470 40736 3476
rect 41328 3528 41380 3534
rect 41328 3470 41380 3476
rect 41880 3528 41932 3534
rect 41880 3470 41932 3476
rect 42708 3528 42760 3534
rect 42708 3470 42760 3476
rect 43076 3528 43128 3534
rect 43076 3470 43128 3476
rect 44088 3528 44140 3534
rect 44088 3470 44140 3476
rect 44272 3528 44324 3534
rect 44272 3470 44324 3476
rect 40696 480 40724 3470
rect 41892 480 41920 3470
rect 43088 480 43116 3470
rect 44284 480 44312 3470
rect 45480 480 45508 59871
rect 46848 21412 46900 21418
rect 46848 21354 46900 21360
rect 46860 6914 46888 21354
rect 48148 6914 48176 65447
rect 48240 26926 48268 284922
rect 49620 276690 49648 380122
rect 50804 375148 50856 375154
rect 50804 375090 50856 375096
rect 50816 317490 50844 375090
rect 50804 317484 50856 317490
rect 50804 317426 50856 317432
rect 50908 298110 50936 380870
rect 51000 375358 51028 421534
rect 50988 375352 51040 375358
rect 50988 375294 51040 375300
rect 51000 375154 51028 375294
rect 50988 375148 51040 375154
rect 50988 375090 51040 375096
rect 52184 337408 52236 337414
rect 52184 337350 52236 337356
rect 50988 331288 51040 331294
rect 50988 331230 51040 331236
rect 50896 298104 50948 298110
rect 50896 298046 50948 298052
rect 50804 289128 50856 289134
rect 50804 289070 50856 289076
rect 49608 276684 49660 276690
rect 49608 276626 49660 276632
rect 49608 262880 49660 262886
rect 49608 262822 49660 262828
rect 49620 262274 49648 262822
rect 49608 262268 49660 262274
rect 49608 262210 49660 262216
rect 49620 200122 49648 262210
rect 50816 213625 50844 289070
rect 50896 288448 50948 288454
rect 50896 288390 50948 288396
rect 50802 213616 50858 213625
rect 50802 213551 50858 213560
rect 49608 200116 49660 200122
rect 49608 200058 49660 200064
rect 50908 196654 50936 288390
rect 50896 196648 50948 196654
rect 50896 196590 50948 196596
rect 50894 73808 50950 73817
rect 50894 73743 50950 73752
rect 49608 46232 49660 46238
rect 49608 46174 49660 46180
rect 48228 26920 48280 26926
rect 48228 26862 48280 26868
rect 46676 6886 46888 6914
rect 47872 6886 48176 6914
rect 46676 480 46704 6886
rect 47872 480 47900 6886
rect 49620 3466 49648 46174
rect 48964 3460 49016 3466
rect 48964 3402 49016 3408
rect 49608 3460 49660 3466
rect 49608 3402 49660 3408
rect 48976 480 49004 3402
rect 50908 3058 50936 73743
rect 51000 15910 51028 331230
rect 52092 271924 52144 271930
rect 52092 271866 52144 271872
rect 52104 191146 52132 271866
rect 52196 235929 52224 337350
rect 52288 333946 52316 456758
rect 52380 429146 52408 561682
rect 53116 436082 53144 566442
rect 53656 554804 53708 554810
rect 53656 554746 53708 554752
rect 53104 436076 53156 436082
rect 53104 436018 53156 436024
rect 52368 429140 52420 429146
rect 52368 429082 52420 429088
rect 53668 415449 53696 554746
rect 55048 455394 55076 587862
rect 59084 586560 59136 586566
rect 59084 586502 59136 586508
rect 57888 585200 57940 585206
rect 57888 585142 57940 585148
rect 56508 549296 56560 549302
rect 56508 549238 56560 549244
rect 55128 543788 55180 543794
rect 55128 543730 55180 543736
rect 55036 455388 55088 455394
rect 55036 455330 55088 455336
rect 55034 445768 55090 445777
rect 55034 445703 55090 445712
rect 53746 444544 53802 444553
rect 53746 444479 53802 444488
rect 53654 415440 53710 415449
rect 53654 415375 53710 415384
rect 53656 415336 53708 415342
rect 53656 415278 53708 415284
rect 53668 414050 53696 415278
rect 53656 414044 53708 414050
rect 53656 413986 53708 413992
rect 52368 340196 52420 340202
rect 52368 340138 52420 340144
rect 52276 333940 52328 333946
rect 52276 333882 52328 333888
rect 52288 333266 52316 333882
rect 52276 333260 52328 333266
rect 52276 333202 52328 333208
rect 52276 317484 52328 317490
rect 52276 317426 52328 317432
rect 52288 314945 52316 317426
rect 52274 314936 52330 314945
rect 52274 314871 52330 314880
rect 52182 235920 52238 235929
rect 52182 235855 52238 235864
rect 52196 235278 52224 235855
rect 52184 235272 52236 235278
rect 52184 235214 52236 235220
rect 52288 226001 52316 314871
rect 52380 293962 52408 340138
rect 52368 293956 52420 293962
rect 52368 293898 52420 293904
rect 52460 287020 52512 287026
rect 52460 286962 52512 286968
rect 52472 286346 52500 286962
rect 52460 286340 52512 286346
rect 52460 286282 52512 286288
rect 53564 286340 53616 286346
rect 53564 286282 53616 286288
rect 53576 285705 53604 286282
rect 53562 285696 53618 285705
rect 53562 285631 53618 285640
rect 53470 268424 53526 268433
rect 53470 268359 53526 268368
rect 52368 247104 52420 247110
rect 52368 247046 52420 247052
rect 52274 225992 52330 226001
rect 52274 225927 52330 225936
rect 52092 191140 52144 191146
rect 52092 191082 52144 191088
rect 52380 32434 52408 247046
rect 53484 186318 53512 268359
rect 53564 264988 53616 264994
rect 53564 264930 53616 264936
rect 53576 217841 53604 264930
rect 53668 241505 53696 413986
rect 53760 263634 53788 444479
rect 54944 433288 54996 433294
rect 54944 433230 54996 433236
rect 54956 432002 54984 433230
rect 54944 431996 54996 432002
rect 54944 431938 54996 431944
rect 54956 373289 54984 431938
rect 54942 373280 54998 373289
rect 54942 373215 54998 373224
rect 55048 368393 55076 445703
rect 55140 398138 55168 543730
rect 56520 520266 56548 549238
rect 57796 538960 57848 538966
rect 57796 538902 57848 538908
rect 56508 520260 56560 520266
rect 56508 520202 56560 520208
rect 56416 455388 56468 455394
rect 56416 455330 56468 455336
rect 56428 454102 56456 455330
rect 56416 454096 56468 454102
rect 56416 454038 56468 454044
rect 55128 398132 55180 398138
rect 55128 398074 55180 398080
rect 56428 371890 56456 454038
rect 56520 407153 56548 520202
rect 57704 449268 57756 449274
rect 57704 449210 57756 449216
rect 56506 407144 56562 407153
rect 56506 407079 56562 407088
rect 57716 389298 57744 449210
rect 57704 389292 57756 389298
rect 57704 389234 57756 389240
rect 57808 387802 57836 538902
rect 57900 447846 57928 585142
rect 59096 529310 59124 586502
rect 61844 574116 61896 574122
rect 61844 574058 61896 574064
rect 60648 571396 60700 571402
rect 60648 571338 60700 571344
rect 59176 558476 59228 558482
rect 59176 558418 59228 558424
rect 59084 529304 59136 529310
rect 59084 529246 59136 529252
rect 59084 461712 59136 461718
rect 59084 461654 59136 461660
rect 57888 447840 57940 447846
rect 57888 447782 57940 447788
rect 58900 423700 58952 423706
rect 58900 423642 58952 423648
rect 57888 403640 57940 403646
rect 57888 403582 57940 403588
rect 57796 387796 57848 387802
rect 57796 387738 57848 387744
rect 56416 371884 56468 371890
rect 56416 371826 56468 371832
rect 56508 369164 56560 369170
rect 56508 369106 56560 369112
rect 55034 368384 55090 368393
rect 55034 368319 55090 368328
rect 55048 354674 55076 368319
rect 54956 354646 55076 354674
rect 54956 292534 54984 354646
rect 55036 341556 55088 341562
rect 55036 341498 55088 341504
rect 54944 292528 54996 292534
rect 54944 292470 54996 292476
rect 54944 279472 54996 279478
rect 54944 279414 54996 279420
rect 53748 263628 53800 263634
rect 53748 263570 53800 263576
rect 53654 241496 53710 241505
rect 53654 241431 53710 241440
rect 53562 217832 53618 217841
rect 53562 217767 53618 217776
rect 54956 204241 54984 279414
rect 55048 237386 55076 341498
rect 55128 320204 55180 320210
rect 55128 320146 55180 320152
rect 55036 237380 55088 237386
rect 55036 237322 55088 237328
rect 54942 204232 54998 204241
rect 54942 204167 54998 204176
rect 53472 186312 53524 186318
rect 53472 186254 53524 186260
rect 53746 71088 53802 71097
rect 53746 71023 53802 71032
rect 52368 32428 52420 32434
rect 52368 32370 52420 32376
rect 50988 15904 51040 15910
rect 50988 15846 51040 15852
rect 53656 11756 53708 11762
rect 53656 11698 53708 11704
rect 53668 3466 53696 11698
rect 52552 3460 52604 3466
rect 52552 3402 52604 3408
rect 53656 3460 53708 3466
rect 53656 3402 53708 3408
rect 50160 3052 50212 3058
rect 50160 2994 50212 3000
rect 50896 3052 50948 3058
rect 50896 2994 50948 3000
rect 50172 480 50200 2994
rect 51356 2100 51408 2106
rect 51356 2042 51408 2048
rect 51368 480 51396 2042
rect 52564 480 52592 3402
rect 53760 480 53788 71023
rect 55140 7614 55168 320146
rect 55864 318844 55916 318850
rect 55864 318786 55916 318792
rect 55876 71233 55904 318786
rect 56520 285666 56548 369106
rect 57702 338736 57758 338745
rect 57702 338671 57758 338680
rect 57610 335608 57666 335617
rect 57610 335543 57666 335552
rect 57624 307766 57652 335543
rect 57612 307760 57664 307766
rect 57612 307702 57664 307708
rect 57612 300892 57664 300898
rect 57612 300834 57664 300840
rect 56508 285660 56560 285666
rect 56508 285602 56560 285608
rect 56520 284986 56548 285602
rect 56508 284980 56560 284986
rect 56508 284922 56560 284928
rect 56508 283620 56560 283626
rect 56508 283562 56560 283568
rect 56520 215937 56548 283562
rect 57244 274644 57296 274650
rect 57244 274586 57296 274592
rect 56506 215928 56562 215937
rect 56506 215863 56562 215872
rect 55862 71224 55918 71233
rect 55862 71159 55918 71168
rect 57256 24138 57284 274586
rect 57624 232801 57652 300834
rect 57716 287026 57744 338671
rect 57796 327140 57848 327146
rect 57796 327082 57848 327088
rect 57808 295322 57836 327082
rect 57796 295316 57848 295322
rect 57796 295258 57848 295264
rect 57704 287020 57756 287026
rect 57704 286962 57756 286968
rect 57704 263628 57756 263634
rect 57704 263570 57756 263576
rect 57610 232792 57666 232801
rect 57610 232727 57666 232736
rect 57716 230217 57744 263570
rect 57900 244322 57928 403582
rect 58912 363662 58940 423642
rect 58992 411324 59044 411330
rect 58992 411266 59044 411272
rect 58900 363656 58952 363662
rect 58900 363598 58952 363604
rect 58900 345704 58952 345710
rect 58900 345646 58952 345652
rect 58912 314634 58940 345646
rect 59004 345014 59032 411266
rect 59096 380866 59124 461654
rect 59188 421598 59216 558418
rect 59268 547936 59320 547942
rect 59268 547878 59320 547884
rect 59176 421592 59228 421598
rect 59176 421534 59228 421540
rect 59280 405822 59308 547878
rect 60464 465724 60516 465730
rect 60464 465666 60516 465672
rect 59268 405816 59320 405822
rect 59268 405758 59320 405764
rect 60004 399492 60056 399498
rect 60004 399434 60056 399440
rect 60016 398138 60044 399434
rect 60004 398132 60056 398138
rect 60004 398074 60056 398080
rect 60476 386374 60504 465666
rect 60660 445913 60688 571338
rect 61856 462913 61884 574058
rect 62040 558482 62068 702850
rect 68284 700324 68336 700330
rect 68284 700266 68336 700272
rect 65800 699712 65852 699718
rect 65800 699654 65852 699660
rect 64696 581052 64748 581058
rect 64696 580994 64748 581000
rect 63316 568608 63368 568614
rect 63316 568550 63368 568556
rect 62028 558476 62080 558482
rect 62028 558418 62080 558424
rect 62040 557598 62068 558418
rect 62028 557592 62080 557598
rect 62028 557534 62080 557540
rect 61936 539640 61988 539646
rect 61936 539582 61988 539588
rect 61842 462904 61898 462913
rect 61842 462839 61898 462848
rect 60646 445904 60702 445913
rect 60646 445839 60702 445848
rect 60556 444508 60608 444514
rect 60556 444450 60608 444456
rect 60464 386368 60516 386374
rect 60464 386310 60516 386316
rect 59084 380860 59136 380866
rect 59084 380802 59136 380808
rect 59096 380186 59124 380802
rect 59084 380180 59136 380186
rect 59084 380122 59136 380128
rect 59174 374096 59230 374105
rect 59174 374031 59230 374040
rect 59004 344986 59124 345014
rect 59096 332586 59124 344986
rect 59084 332580 59136 332586
rect 59084 332522 59136 332528
rect 59096 331906 59124 332522
rect 59084 331900 59136 331906
rect 59084 331842 59136 331848
rect 59084 328568 59136 328574
rect 59084 328510 59136 328516
rect 58900 314628 58952 314634
rect 58900 314570 58952 314576
rect 58992 255332 59044 255338
rect 58992 255274 59044 255280
rect 57888 244316 57940 244322
rect 57888 244258 57940 244264
rect 57702 230208 57758 230217
rect 57702 230143 57758 230152
rect 59004 224913 59032 255274
rect 59096 231441 59124 328510
rect 59188 247042 59216 374031
rect 59266 334384 59322 334393
rect 59266 334319 59322 334328
rect 59280 302190 59308 334319
rect 59268 302184 59320 302190
rect 59268 302126 59320 302132
rect 59268 298172 59320 298178
rect 59268 298114 59320 298120
rect 59176 247036 59228 247042
rect 59176 246978 59228 246984
rect 59082 231432 59138 231441
rect 59082 231367 59138 231376
rect 58990 224904 59046 224913
rect 58990 224839 59046 224848
rect 57886 72584 57942 72593
rect 57886 72519 57942 72528
rect 57244 24132 57296 24138
rect 57244 24074 57296 24080
rect 56508 22840 56560 22846
rect 56508 22782 56560 22788
rect 55128 7608 55180 7614
rect 55128 7550 55180 7556
rect 54944 4888 54996 4894
rect 54944 4830 54996 4836
rect 54956 480 54984 4830
rect 56520 3466 56548 22782
rect 57900 3466 57928 72519
rect 59280 72457 59308 298114
rect 60464 276684 60516 276690
rect 60464 276626 60516 276632
rect 60372 253292 60424 253298
rect 60372 253234 60424 253240
rect 60384 235278 60412 253234
rect 60372 235272 60424 235278
rect 60372 235214 60424 235220
rect 60476 194585 60504 276626
rect 60568 253026 60596 444450
rect 60740 425740 60792 425746
rect 60740 425682 60792 425688
rect 60752 425134 60780 425682
rect 60740 425128 60792 425134
rect 60740 425070 60792 425076
rect 61844 425128 61896 425134
rect 61844 425070 61896 425076
rect 61856 382974 61884 425070
rect 61948 392086 61976 539582
rect 62028 467152 62080 467158
rect 62028 467094 62080 467100
rect 61936 392080 61988 392086
rect 61936 392022 61988 392028
rect 61844 382968 61896 382974
rect 61844 382910 61896 382916
rect 61934 363080 61990 363089
rect 61934 363015 61990 363024
rect 61844 339516 61896 339522
rect 61844 339458 61896 339464
rect 60648 335368 60700 335374
rect 60648 335310 60700 335316
rect 60556 253020 60608 253026
rect 60556 252962 60608 252968
rect 60556 249892 60608 249898
rect 60556 249834 60608 249840
rect 60568 227730 60596 249834
rect 60556 227724 60608 227730
rect 60556 227666 60608 227672
rect 60462 194576 60518 194585
rect 60462 194511 60518 194520
rect 60660 93158 60688 335310
rect 61856 313274 61884 339458
rect 61844 313268 61896 313274
rect 61844 313210 61896 313216
rect 61948 306338 61976 363015
rect 61936 306332 61988 306338
rect 61936 306274 61988 306280
rect 61844 280220 61896 280226
rect 61844 280162 61896 280168
rect 61752 256012 61804 256018
rect 61752 255954 61804 255960
rect 61764 232558 61792 255954
rect 61752 232552 61804 232558
rect 61752 232494 61804 232500
rect 61856 220833 61884 280162
rect 61936 267776 61988 267782
rect 61936 267718 61988 267724
rect 61842 220824 61898 220833
rect 61842 220759 61898 220768
rect 61948 187649 61976 267718
rect 61934 187640 61990 187649
rect 61934 187575 61990 187584
rect 60648 93152 60700 93158
rect 60648 93094 60700 93100
rect 62040 91798 62068 467094
rect 63328 456074 63356 568550
rect 63408 558952 63460 558958
rect 63408 558894 63460 558900
rect 63316 456068 63368 456074
rect 63316 456010 63368 456016
rect 63316 454708 63368 454714
rect 63316 454650 63368 454656
rect 62854 416664 62910 416673
rect 62854 416599 62910 416608
rect 62868 415449 62896 416599
rect 62854 415440 62910 415449
rect 62854 415375 62910 415384
rect 63328 387025 63356 454650
rect 63420 423706 63448 558894
rect 64708 530602 64736 580994
rect 64788 567248 64840 567254
rect 64788 567190 64840 567196
rect 64696 530596 64748 530602
rect 64696 530538 64748 530544
rect 64800 463758 64828 567190
rect 65812 538966 65840 699654
rect 67456 596828 67508 596834
rect 67456 596770 67508 596776
rect 65984 594856 66036 594862
rect 65984 594798 66036 594804
rect 65890 573472 65946 573481
rect 65890 573407 65946 573416
rect 65904 542337 65932 573407
rect 65996 554062 66024 594798
rect 66074 590744 66130 590753
rect 66074 590679 66130 590688
rect 65984 554056 66036 554062
rect 65984 553998 66036 554004
rect 65890 542328 65946 542337
rect 65890 542263 65946 542272
rect 65800 538960 65852 538966
rect 65800 538902 65852 538908
rect 65984 538960 66036 538966
rect 65984 538902 66036 538908
rect 65996 538286 66024 538902
rect 65984 538280 66036 538286
rect 65984 538222 66036 538228
rect 64788 463752 64840 463758
rect 64788 463694 64840 463700
rect 64800 460934 64828 463694
rect 64708 460906 64828 460934
rect 64708 438870 64736 460906
rect 65984 460216 66036 460222
rect 65984 460158 66036 460164
rect 64788 458856 64840 458862
rect 64788 458798 64840 458804
rect 64696 438864 64748 438870
rect 64696 438806 64748 438812
rect 64696 431248 64748 431254
rect 64696 431190 64748 431196
rect 63408 423700 63460 423706
rect 63408 423642 63460 423648
rect 63406 415440 63462 415449
rect 63406 415375 63462 415384
rect 63420 389201 63448 415375
rect 64604 405816 64656 405822
rect 64604 405758 64656 405764
rect 63406 389192 63462 389201
rect 63406 389127 63462 389136
rect 63314 387016 63370 387025
rect 63314 386951 63370 386960
rect 63314 378720 63370 378729
rect 63314 378655 63370 378664
rect 63222 332752 63278 332761
rect 63222 332687 63278 332696
rect 63236 304978 63264 332687
rect 63224 304972 63276 304978
rect 63224 304914 63276 304920
rect 63224 277432 63276 277438
rect 63224 277374 63276 277380
rect 63132 249824 63184 249830
rect 63132 249766 63184 249772
rect 63144 226953 63172 249766
rect 63236 230353 63264 277374
rect 63328 267850 63356 378655
rect 64616 356726 64644 405758
rect 64708 376689 64736 431190
rect 64800 391241 64828 458798
rect 65616 453348 65668 453354
rect 65616 453290 65668 453296
rect 64786 391232 64842 391241
rect 64786 391167 64842 391176
rect 65628 388793 65656 453290
rect 65892 447160 65944 447166
rect 65892 447102 65944 447108
rect 65798 389056 65854 389065
rect 65798 388991 65854 389000
rect 65614 388784 65670 388793
rect 65614 388719 65670 388728
rect 64694 376680 64750 376689
rect 64694 376615 64750 376624
rect 64604 356720 64656 356726
rect 64604 356662 64656 356668
rect 64696 351212 64748 351218
rect 64696 351154 64748 351160
rect 63408 343664 63460 343670
rect 63408 343606 63460 343612
rect 63420 309806 63448 343606
rect 64708 318170 64736 351154
rect 64788 338768 64840 338774
rect 64788 338710 64840 338716
rect 64696 318164 64748 318170
rect 64696 318106 64748 318112
rect 63408 309800 63460 309806
rect 63408 309742 63460 309748
rect 63500 290488 63552 290494
rect 63500 290430 63552 290436
rect 63512 289950 63540 290430
rect 63500 289944 63552 289950
rect 63500 289886 63552 289892
rect 64696 289944 64748 289950
rect 64696 289886 64748 289892
rect 63408 287088 63460 287094
rect 63408 287030 63460 287036
rect 63316 267844 63368 267850
rect 63316 267786 63368 267792
rect 63328 238066 63356 267786
rect 63316 238060 63368 238066
rect 63316 238002 63368 238008
rect 63222 230344 63278 230353
rect 63222 230279 63278 230288
rect 63130 226944 63186 226953
rect 63130 226879 63186 226888
rect 62028 91792 62080 91798
rect 62028 91734 62080 91740
rect 61382 79520 61438 79529
rect 61382 79455 61438 79464
rect 59266 72448 59322 72457
rect 59266 72383 59322 72392
rect 60646 69592 60702 69601
rect 60646 69527 60702 69536
rect 58622 64152 58678 64161
rect 58622 64087 58678 64096
rect 56048 3460 56100 3466
rect 56048 3402 56100 3408
rect 56508 3460 56560 3466
rect 56508 3402 56560 3408
rect 57244 3460 57296 3466
rect 57244 3402 57296 3408
rect 57888 3460 57940 3466
rect 57888 3402 57940 3408
rect 58440 3460 58492 3466
rect 58440 3402 58492 3408
rect 56060 480 56088 3402
rect 57256 480 57284 3402
rect 58452 480 58480 3402
rect 58636 2106 58664 64087
rect 59268 39364 59320 39370
rect 59268 39306 59320 39312
rect 59280 3466 59308 39306
rect 60660 3466 60688 69527
rect 60832 4820 60884 4826
rect 60832 4762 60884 4768
rect 59268 3460 59320 3466
rect 59268 3402 59320 3408
rect 59636 3460 59688 3466
rect 59636 3402 59688 3408
rect 60648 3460 60700 3466
rect 60648 3402 60700 3408
rect 58624 2100 58676 2106
rect 58624 2042 58676 2048
rect 59648 480 59676 3402
rect 60844 480 60872 4762
rect 61396 3398 61424 79455
rect 61936 31136 61988 31142
rect 61936 31078 61988 31084
rect 61948 16574 61976 31078
rect 63420 29646 63448 287030
rect 64604 282940 64656 282946
rect 64604 282882 64656 282888
rect 64512 244316 64564 244322
rect 64512 244258 64564 244264
rect 64524 219201 64552 244258
rect 64616 236706 64644 282882
rect 64604 236700 64656 236706
rect 64604 236642 64656 236648
rect 64708 231713 64736 289886
rect 64800 287094 64828 338710
rect 65812 322425 65840 388991
rect 65904 388929 65932 447102
rect 65890 388920 65946 388929
rect 65890 388855 65946 388864
rect 65996 383654 66024 460158
rect 66088 450634 66116 590679
rect 66810 588432 66866 588441
rect 66810 588367 66866 588376
rect 66824 587926 66852 588367
rect 66812 587920 66864 587926
rect 66812 587862 66864 587868
rect 66260 586560 66312 586566
rect 66258 586528 66260 586537
rect 66312 586528 66314 586537
rect 66258 586463 66314 586472
rect 66810 585712 66866 585721
rect 66810 585647 66866 585656
rect 66824 585206 66852 585647
rect 66812 585200 66864 585206
rect 66812 585142 66864 585148
rect 66810 582992 66866 583001
rect 66810 582927 66866 582936
rect 66824 582418 66852 582927
rect 66812 582412 66864 582418
rect 66812 582354 66864 582360
rect 66442 581768 66498 581777
rect 66442 581703 66498 581712
rect 66456 581058 66484 581703
rect 66444 581052 66496 581058
rect 66444 580994 66496 581000
rect 66810 580272 66866 580281
rect 66810 580207 66866 580216
rect 66824 579698 66852 580207
rect 66812 579692 66864 579698
rect 66812 579634 66864 579640
rect 67270 577552 67326 577561
rect 67270 577487 67326 577496
rect 67086 574832 67142 574841
rect 67086 574767 67142 574776
rect 67100 574122 67128 574767
rect 67088 574116 67140 574122
rect 67088 574058 67140 574064
rect 66810 572112 66866 572121
rect 66810 572047 66866 572056
rect 66824 571402 66852 572047
rect 66812 571396 66864 571402
rect 66812 571338 66864 571344
rect 67178 570752 67234 570761
rect 67178 570687 67234 570696
rect 66810 569392 66866 569401
rect 66810 569327 66866 569336
rect 66824 568614 66852 569327
rect 66812 568608 66864 568614
rect 66812 568550 66864 568556
rect 66718 568032 66774 568041
rect 66718 567967 66774 567976
rect 66732 567254 66760 567967
rect 66720 567248 66772 567254
rect 66720 567190 66772 567196
rect 66810 565040 66866 565049
rect 66810 564975 66866 564984
rect 66824 564466 66852 564975
rect 66812 564460 66864 564466
rect 66812 564402 66864 564408
rect 66810 563680 66866 563689
rect 66810 563615 66866 563624
rect 66824 563106 66852 563615
rect 66812 563100 66864 563106
rect 66812 563042 66864 563048
rect 66810 562320 66866 562329
rect 66810 562255 66866 562264
rect 66824 561746 66852 562255
rect 66812 561740 66864 561746
rect 66812 561682 66864 561688
rect 66810 560960 66866 560969
rect 66810 560895 66866 560904
rect 66824 560318 66852 560895
rect 66812 560312 66864 560318
rect 66812 560254 66864 560260
rect 66810 559600 66866 559609
rect 66810 559535 66866 559544
rect 66824 558958 66852 559535
rect 66812 558952 66864 558958
rect 66812 558894 66864 558900
rect 66810 558240 66866 558249
rect 66810 558175 66866 558184
rect 66824 557598 66852 558175
rect 66812 557592 66864 557598
rect 66812 557534 66864 557540
rect 66810 555520 66866 555529
rect 66810 555455 66866 555464
rect 66824 554810 66852 555455
rect 66812 554804 66864 554810
rect 66812 554746 66864 554752
rect 66534 554160 66590 554169
rect 66534 554095 66590 554104
rect 66548 554062 66576 554095
rect 66536 554056 66588 554062
rect 66536 553998 66588 554004
rect 66442 550080 66498 550089
rect 66442 550015 66498 550024
rect 66456 549302 66484 550015
rect 66444 549296 66496 549302
rect 66444 549238 66496 549244
rect 66442 548720 66498 548729
rect 66442 548655 66498 548664
rect 66456 547942 66484 548655
rect 66444 547936 66496 547942
rect 66444 547878 66496 547884
rect 66166 547360 66222 547369
rect 66166 547295 66222 547304
rect 66180 517478 66208 547295
rect 66810 545184 66866 545193
rect 66810 545119 66812 545128
rect 66864 545119 66866 545128
rect 66812 545090 66864 545096
rect 66810 544640 66866 544649
rect 66810 544575 66866 544584
rect 66824 543794 66852 544575
rect 66812 543788 66864 543794
rect 66812 543730 66864 543736
rect 66810 543280 66866 543289
rect 66810 543215 66866 543224
rect 66824 542434 66852 543215
rect 66812 542428 66864 542434
rect 66812 542370 66864 542376
rect 67086 541920 67142 541929
rect 67086 541855 67142 541864
rect 67100 541686 67128 541855
rect 67088 541680 67140 541686
rect 67088 541622 67140 541628
rect 67192 538214 67220 570687
rect 67284 539782 67312 577487
rect 67362 576192 67418 576201
rect 67362 576127 67364 576136
rect 67416 576127 67418 576136
rect 67364 576098 67416 576104
rect 67376 569906 67404 576098
rect 67364 569900 67416 569906
rect 67364 569842 67416 569848
rect 67468 566817 67496 596770
rect 68296 585206 68324 700266
rect 72988 699718 73016 703520
rect 86868 702568 86920 702574
rect 86868 702510 86920 702516
rect 72976 699712 73028 699718
rect 72976 699654 73028 699660
rect 74632 599004 74684 599010
rect 74632 598946 74684 598952
rect 70308 597576 70360 597582
rect 70308 597518 70360 597524
rect 69112 591320 69164 591326
rect 69112 591262 69164 591268
rect 69124 590714 69152 591262
rect 70124 590776 70176 590782
rect 70320 590753 70348 597518
rect 74644 596174 74672 598946
rect 74644 596146 75040 596174
rect 72882 595504 72938 595513
rect 72882 595439 72938 595448
rect 70124 590718 70176 590724
rect 70306 590744 70362 590753
rect 69112 590708 69164 590714
rect 69112 590650 69164 590656
rect 69124 589084 69152 590650
rect 70136 589084 70164 590718
rect 71134 590744 71190 590753
rect 70306 590679 70362 590688
rect 70400 590708 70452 590714
rect 71134 590679 71190 590688
rect 70400 590650 70452 590656
rect 70412 589966 70440 590650
rect 70400 589960 70452 589966
rect 70400 589902 70452 589908
rect 71148 589084 71176 590679
rect 72174 588526 72464 588554
rect 72436 588470 72464 588526
rect 72896 588470 72924 595439
rect 73988 593428 74040 593434
rect 73988 593370 74040 593376
rect 73160 590776 73212 590782
rect 73160 590718 73212 590724
rect 73068 590708 73120 590714
rect 73068 590650 73120 590656
rect 73080 589084 73108 590650
rect 73172 589937 73200 590718
rect 73158 589928 73214 589937
rect 73158 589863 73214 589872
rect 74000 589084 74028 593370
rect 74908 589348 74960 589354
rect 74908 589290 74960 589296
rect 74920 589084 74948 589290
rect 75012 589098 75040 596146
rect 86880 594930 86908 702510
rect 88800 702500 88852 702506
rect 88800 702442 88852 702448
rect 87604 699712 87656 699718
rect 87604 699654 87656 699660
rect 87616 595513 87644 699654
rect 88812 596174 88840 702442
rect 89180 699718 89208 703520
rect 95148 702636 95200 702642
rect 95148 702578 95200 702584
rect 89168 699712 89220 699718
rect 89168 699654 89220 699660
rect 90364 605872 90416 605878
rect 90364 605814 90416 605820
rect 88812 596146 89024 596174
rect 87602 595504 87658 595513
rect 87602 595439 87658 595448
rect 86868 594924 86920 594930
rect 86868 594866 86920 594872
rect 80336 592680 80388 592686
rect 80336 592622 80388 592628
rect 75644 592136 75696 592142
rect 75644 592078 75696 592084
rect 78586 592104 78642 592113
rect 75656 589354 75684 592078
rect 78586 592039 78642 592048
rect 77666 589520 77722 589529
rect 77666 589455 77722 589464
rect 75644 589348 75696 589354
rect 75644 589290 75696 589296
rect 76748 589348 76800 589354
rect 76748 589290 76800 589296
rect 75012 589070 75762 589098
rect 76760 589084 76788 589290
rect 77680 589084 77708 589455
rect 78600 589084 78628 592039
rect 80348 588554 80376 592622
rect 84108 592068 84160 592074
rect 84108 592010 84160 592016
rect 83186 591016 83242 591025
rect 83186 590951 83242 590960
rect 82266 590744 82322 590753
rect 81716 590708 81768 590714
rect 82266 590679 82322 590688
rect 81716 590650 81768 590656
rect 81346 589384 81402 589393
rect 81346 589319 81402 589328
rect 81360 589084 81388 589319
rect 81728 588713 81756 590650
rect 82280 589084 82308 590679
rect 83200 589084 83228 590951
rect 84120 589084 84148 592010
rect 86776 590776 86828 590782
rect 86776 590718 86828 590724
rect 85028 590708 85080 590714
rect 85028 590650 85080 590656
rect 85040 589084 85068 590650
rect 86224 590640 86276 590646
rect 86224 590582 86276 590588
rect 86236 589098 86264 590582
rect 85974 589070 86264 589098
rect 86788 589084 86816 590718
rect 86880 590714 86908 594866
rect 86868 590708 86920 590714
rect 86868 590650 86920 590656
rect 81714 588704 81770 588713
rect 81714 588639 81770 588648
rect 88062 588568 88118 588577
rect 79534 588538 79824 588554
rect 80348 588540 80744 588554
rect 79534 588532 79836 588538
rect 79534 588526 79784 588532
rect 80362 588526 80744 588540
rect 87814 588526 88062 588554
rect 79784 588474 79836 588480
rect 80716 588470 80744 588526
rect 88062 588503 88118 588512
rect 72424 588464 72476 588470
rect 72424 588406 72476 588412
rect 72884 588464 72936 588470
rect 72884 588406 72936 588412
rect 80704 588464 80756 588470
rect 80704 588406 80756 588412
rect 88734 588390 88932 588418
rect 88904 587450 88932 588390
rect 88892 587444 88944 587450
rect 88892 587386 88944 587392
rect 88996 587330 89024 596146
rect 90376 594454 90404 605814
rect 90364 594448 90416 594454
rect 90364 594390 90416 594396
rect 91100 594448 91152 594454
rect 91100 594390 91152 594396
rect 89812 594108 89864 594114
rect 89812 594050 89864 594056
rect 89076 589960 89128 589966
rect 89076 589902 89128 589908
rect 88812 587302 89024 587330
rect 67548 585200 67600 585206
rect 67548 585142 67600 585148
rect 68284 585200 68336 585206
rect 68284 585142 68336 585148
rect 67560 574841 67588 585142
rect 67638 584352 67694 584361
rect 67638 584287 67694 584296
rect 67546 574832 67602 574841
rect 67546 574767 67602 574776
rect 67454 566808 67510 566817
rect 67454 566743 67510 566752
rect 67468 566506 67496 566743
rect 67456 566500 67508 566506
rect 67456 566442 67508 566448
rect 67454 552800 67510 552809
rect 67454 552735 67510 552744
rect 67364 541680 67416 541686
rect 67364 541622 67416 541628
rect 67272 539776 67324 539782
rect 67272 539718 67324 539724
rect 67376 539458 67404 541622
rect 67468 539578 67496 552735
rect 67548 539640 67600 539646
rect 67546 539608 67548 539617
rect 67600 539608 67602 539617
rect 67456 539572 67508 539578
rect 67546 539543 67602 539552
rect 67456 539514 67508 539520
rect 67376 539430 67588 539458
rect 67456 539368 67508 539374
rect 67456 539310 67508 539316
rect 67192 538186 67404 538214
rect 67376 538121 67404 538186
rect 67362 538112 67418 538121
rect 67362 538047 67418 538056
rect 67086 537432 67142 537441
rect 67086 537367 67142 537376
rect 66902 523832 66958 523841
rect 66902 523767 66958 523776
rect 66916 523734 66944 523767
rect 66904 523728 66956 523734
rect 67100 523705 67128 537367
rect 66904 523670 66956 523676
rect 67086 523696 67142 523705
rect 66168 517472 66220 517478
rect 66168 517414 66220 517420
rect 66076 450628 66128 450634
rect 66076 450570 66128 450576
rect 66180 403730 66208 517414
rect 66812 438864 66864 438870
rect 66812 438806 66864 438812
rect 66824 437889 66852 438806
rect 66810 437880 66866 437889
rect 66810 437815 66866 437824
rect 66720 436076 66772 436082
rect 66720 436018 66772 436024
rect 66732 435441 66760 436018
rect 66718 435432 66774 435441
rect 66718 435367 66774 435376
rect 66810 433120 66866 433129
rect 66810 433055 66866 433064
rect 66824 432002 66852 433055
rect 66812 431996 66864 432002
rect 66812 431938 66864 431944
rect 66812 431248 66864 431254
rect 66812 431190 66864 431196
rect 66824 431089 66852 431190
rect 66810 431080 66866 431089
rect 66810 431015 66866 431024
rect 66812 429140 66864 429146
rect 66812 429082 66864 429088
rect 66824 428641 66852 429082
rect 66810 428632 66866 428641
rect 66810 428567 66866 428576
rect 66718 426320 66774 426329
rect 66718 426255 66774 426264
rect 66732 425134 66760 426255
rect 66720 425128 66772 425134
rect 66720 425070 66772 425076
rect 66810 424144 66866 424153
rect 66810 424079 66866 424088
rect 66824 423706 66852 424079
rect 66812 423700 66864 423706
rect 66812 423642 66864 423648
rect 66258 421968 66314 421977
rect 66258 421903 66314 421912
rect 66272 421598 66300 421903
rect 66260 421592 66312 421598
rect 66260 421534 66312 421540
rect 66810 415168 66866 415177
rect 66810 415103 66866 415112
rect 66824 414050 66852 415103
rect 66812 414044 66864 414050
rect 66812 413986 66864 413992
rect 66916 411330 66944 523670
rect 67086 523631 67142 523640
rect 67376 442950 67404 538047
rect 67364 442944 67416 442950
rect 67364 442886 67416 442892
rect 67364 438932 67416 438938
rect 67364 438874 67416 438880
rect 66904 411324 66956 411330
rect 66904 411266 66956 411272
rect 66916 410689 66944 411266
rect 66902 410680 66958 410689
rect 66902 410615 66958 410624
rect 66258 406192 66314 406201
rect 66258 406127 66314 406136
rect 66272 405822 66300 406127
rect 66260 405816 66312 405822
rect 66260 405758 66312 405764
rect 66258 403744 66314 403753
rect 66180 403702 66258 403730
rect 66258 403679 66314 403688
rect 66272 403646 66300 403679
rect 66260 403640 66312 403646
rect 66260 403582 66312 403588
rect 66260 401600 66312 401606
rect 66258 401568 66260 401577
rect 66312 401568 66314 401577
rect 66258 401503 66314 401512
rect 66258 399528 66314 399537
rect 66258 399463 66260 399472
rect 66312 399463 66314 399472
rect 66260 399434 66312 399440
rect 66994 396944 67050 396953
rect 66994 396879 67050 396888
rect 67008 396778 67036 396879
rect 66996 396772 67048 396778
rect 66996 396714 67048 396720
rect 67272 396772 67324 396778
rect 67272 396714 67324 396720
rect 66626 392592 66682 392601
rect 66626 392527 66682 392536
rect 66640 392086 66668 392527
rect 66168 392080 66220 392086
rect 66168 392022 66220 392028
rect 66628 392080 66680 392086
rect 66628 392022 66680 392028
rect 65984 383648 66036 383654
rect 65984 383590 66036 383596
rect 66074 360904 66130 360913
rect 66074 360839 66130 360848
rect 65890 336832 65946 336841
rect 65890 336767 65946 336776
rect 65798 322416 65854 322425
rect 65798 322351 65854 322360
rect 65904 303113 65932 336767
rect 65982 322416 66038 322425
rect 65982 322351 66038 322360
rect 65890 303104 65946 303113
rect 65890 303039 65946 303048
rect 64788 287088 64840 287094
rect 64788 287030 64840 287036
rect 65890 281344 65946 281353
rect 65890 281279 65946 281288
rect 64788 259480 64840 259486
rect 64788 259422 64840 259428
rect 64694 231704 64750 231713
rect 64694 231639 64750 231648
rect 64510 219192 64566 219201
rect 64510 219127 64566 219136
rect 64800 190369 64828 259422
rect 65904 232626 65932 281279
rect 65996 234569 66024 322351
rect 66088 271833 66116 360839
rect 66180 315874 66208 392022
rect 67284 378214 67312 396714
rect 67272 378208 67324 378214
rect 67272 378150 67324 378156
rect 67284 373994 67312 378150
rect 67008 373966 67312 373994
rect 66904 371272 66956 371278
rect 66904 371214 66956 371220
rect 66916 343670 66944 371214
rect 67008 351218 67036 373966
rect 67376 371278 67404 438874
rect 67468 412865 67496 539310
rect 67454 412856 67510 412865
rect 67454 412791 67510 412800
rect 67364 371272 67416 371278
rect 67364 371214 67416 371220
rect 66996 351212 67048 351218
rect 66996 351154 67048 351160
rect 67362 345672 67418 345681
rect 67362 345607 67418 345616
rect 66904 343664 66956 343670
rect 66904 343606 66956 343612
rect 67272 330540 67324 330546
rect 67272 330482 67324 330488
rect 66626 328944 66682 328953
rect 66626 328879 66682 328888
rect 66640 328574 66668 328879
rect 66628 328568 66680 328574
rect 66628 328510 66680 328516
rect 67284 324601 67312 330482
rect 67270 324592 67326 324601
rect 67270 324527 67326 324536
rect 66904 321564 66956 321570
rect 66904 321506 66956 321512
rect 66810 321328 66866 321337
rect 66810 321263 66866 321272
rect 66824 320210 66852 321263
rect 66916 320249 66944 321506
rect 66902 320240 66958 320249
rect 66812 320204 66864 320210
rect 66902 320175 66958 320184
rect 66812 320146 66864 320152
rect 66902 319152 66958 319161
rect 66902 319087 66958 319096
rect 66916 318850 66944 319087
rect 66904 318844 66956 318850
rect 66904 318786 66956 318792
rect 66812 318164 66864 318170
rect 66812 318106 66864 318112
rect 66824 318073 66852 318106
rect 66810 318064 66866 318073
rect 66810 317999 66866 318008
rect 67376 316985 67404 345607
rect 67362 316976 67418 316985
rect 67362 316911 67418 316920
rect 67376 316742 67404 316911
rect 67364 316736 67416 316742
rect 67364 316678 67416 316684
rect 66258 315888 66314 315897
rect 66180 315846 66258 315874
rect 66074 271824 66130 271833
rect 66074 271759 66130 271768
rect 66074 260944 66130 260953
rect 66074 260879 66130 260888
rect 65982 234560 66038 234569
rect 65982 234495 66038 234504
rect 65892 232620 65944 232626
rect 65892 232562 65944 232568
rect 66088 229770 66116 260879
rect 66076 229764 66128 229770
rect 66076 229706 66128 229712
rect 66180 224777 66208 315846
rect 66258 315823 66314 315832
rect 66812 314628 66864 314634
rect 66812 314570 66864 314576
rect 66824 313993 66852 314570
rect 66810 313984 66866 313993
rect 66810 313919 66866 313928
rect 66444 313268 66496 313274
rect 66444 313210 66496 313216
rect 66456 312905 66484 313210
rect 66442 312896 66498 312905
rect 66442 312831 66498 312840
rect 66994 311808 67050 311817
rect 66994 311743 67050 311752
rect 66812 309800 66864 309806
rect 66812 309742 66864 309748
rect 66824 309641 66852 309742
rect 66810 309632 66866 309641
rect 66810 309567 66866 309576
rect 66904 307760 66956 307766
rect 66904 307702 66956 307708
rect 66916 307465 66944 307702
rect 66902 307456 66958 307465
rect 66902 307391 66958 307400
rect 66812 306332 66864 306338
rect 66812 306274 66864 306280
rect 66824 305289 66852 306274
rect 66810 305280 66866 305289
rect 66810 305215 66866 305224
rect 66812 304972 66864 304978
rect 66812 304914 66864 304920
rect 66824 304201 66852 304914
rect 66810 304192 66866 304201
rect 66810 304127 66866 304136
rect 66904 302184 66956 302190
rect 66904 302126 66956 302132
rect 66810 302016 66866 302025
rect 66810 301951 66866 301960
rect 66824 300898 66852 301951
rect 66916 300937 66944 302126
rect 66902 300928 66958 300937
rect 66812 300892 66864 300898
rect 66902 300863 66958 300872
rect 66812 300834 66864 300840
rect 66626 298752 66682 298761
rect 66626 298687 66682 298696
rect 66640 298178 66668 298687
rect 66628 298172 66680 298178
rect 66628 298114 66680 298120
rect 66812 298104 66864 298110
rect 66812 298046 66864 298052
rect 66824 297673 66852 298046
rect 66810 297664 66866 297673
rect 66810 297599 66866 297608
rect 66718 295488 66774 295497
rect 66718 295423 66774 295432
rect 66732 289134 66760 295423
rect 66812 295316 66864 295322
rect 66812 295258 66864 295264
rect 66824 294409 66852 295258
rect 66810 294400 66866 294409
rect 66810 294335 66866 294344
rect 66812 293956 66864 293962
rect 66812 293898 66864 293904
rect 66824 293321 66852 293898
rect 66810 293312 66866 293321
rect 66810 293247 66866 293256
rect 66812 292528 66864 292534
rect 66812 292470 66864 292476
rect 66824 292233 66852 292470
rect 66810 292224 66866 292233
rect 66810 292159 66866 292168
rect 66810 291136 66866 291145
rect 66810 291071 66866 291080
rect 66824 289950 66852 291071
rect 66902 290048 66958 290057
rect 66902 289983 66958 289992
rect 66812 289944 66864 289950
rect 66812 289886 66864 289892
rect 66720 289128 66772 289134
rect 66720 289070 66772 289076
rect 66810 288960 66866 288969
rect 66810 288895 66866 288904
rect 66824 288454 66852 288895
rect 66812 288448 66864 288454
rect 66812 288390 66864 288396
rect 66626 287872 66682 287881
rect 66626 287807 66682 287816
rect 66640 287094 66668 287807
rect 66628 287088 66680 287094
rect 66628 287030 66680 287036
rect 66812 287020 66864 287026
rect 66812 286962 66864 286968
rect 66350 286784 66406 286793
rect 66350 286719 66406 286728
rect 66364 286346 66392 286719
rect 66352 286340 66404 286346
rect 66352 286282 66404 286288
rect 66824 285705 66852 286962
rect 66810 285696 66866 285705
rect 66720 285660 66772 285666
rect 66810 285631 66866 285640
rect 66720 285602 66772 285608
rect 66732 284617 66760 285602
rect 66718 284608 66774 284617
rect 66718 284543 66774 284552
rect 66810 283520 66866 283529
rect 66810 283455 66866 283464
rect 66824 282946 66852 283455
rect 66812 282940 66864 282946
rect 66812 282882 66864 282888
rect 66810 278080 66866 278089
rect 66810 278015 66866 278024
rect 66824 277438 66852 278015
rect 66812 277432 66864 277438
rect 66812 277374 66864 277380
rect 66810 277264 66866 277273
rect 66810 277199 66866 277208
rect 66824 276690 66852 277199
rect 66812 276684 66864 276690
rect 66812 276626 66864 276632
rect 66626 275088 66682 275097
rect 66626 275023 66682 275032
rect 66640 274718 66668 275023
rect 66628 274712 66680 274718
rect 66628 274654 66680 274660
rect 66258 272912 66314 272921
rect 66258 272847 66314 272856
rect 66272 271930 66300 272847
rect 66260 271924 66312 271930
rect 66260 271866 66312 271872
rect 66810 268560 66866 268569
rect 66810 268495 66866 268504
rect 66824 267850 66852 268495
rect 66812 267844 66864 267850
rect 66812 267786 66864 267792
rect 66810 265296 66866 265305
rect 66810 265231 66866 265240
rect 66824 264994 66852 265231
rect 66812 264988 66864 264994
rect 66812 264930 66864 264936
rect 66810 264208 66866 264217
rect 66810 264143 66866 264152
rect 66824 263634 66852 264143
rect 66812 263628 66864 263634
rect 66812 263570 66864 263576
rect 66810 263120 66866 263129
rect 66810 263055 66866 263064
rect 66824 262274 66852 263055
rect 66812 262268 66864 262274
rect 66812 262210 66864 262216
rect 66444 262200 66496 262206
rect 66444 262142 66496 262148
rect 66456 262041 66484 262142
rect 66442 262032 66498 262041
rect 66442 261967 66498 261976
rect 66810 259856 66866 259865
rect 66810 259791 66866 259800
rect 66824 259486 66852 259791
rect 66812 259480 66864 259486
rect 66812 259422 66864 259428
rect 66810 256592 66866 256601
rect 66810 256527 66866 256536
rect 66824 255338 66852 256527
rect 66812 255332 66864 255338
rect 66812 255274 66864 255280
rect 66916 253298 66944 289983
rect 67008 283626 67036 311743
rect 67468 311166 67496 412791
rect 67560 394913 67588 539430
rect 67652 456822 67680 584287
rect 67730 578912 67786 578921
rect 67730 578847 67786 578856
rect 67744 534070 67772 578847
rect 88812 576854 88840 587302
rect 88892 587172 88944 587178
rect 88892 587114 88944 587120
rect 88904 577561 88932 587114
rect 89088 582374 89116 589902
rect 89168 588464 89220 588470
rect 89168 588406 89220 588412
rect 89180 586634 89208 588406
rect 89168 586628 89220 586634
rect 89168 586570 89220 586576
rect 89718 586256 89774 586265
rect 89718 586191 89774 586200
rect 88996 582346 89116 582374
rect 88890 577552 88946 577561
rect 88890 577487 88946 577496
rect 88812 576826 88932 576854
rect 68284 569900 68336 569906
rect 68284 569842 68336 569848
rect 67732 534064 67784 534070
rect 67732 534006 67784 534012
rect 68296 476134 68324 569842
rect 88904 560153 88932 576826
rect 88890 560144 88946 560153
rect 88890 560079 88946 560088
rect 70400 539640 70452 539646
rect 71872 539640 71924 539646
rect 70452 539588 70610 539594
rect 70400 539582 70610 539588
rect 71872 539582 71924 539588
rect 88156 539640 88208 539646
rect 88156 539582 88208 539588
rect 70412 539566 70610 539582
rect 68664 539294 68770 539322
rect 69584 539294 69690 539322
rect 68664 536625 68692 539294
rect 69584 536790 69612 539294
rect 69572 536784 69624 536790
rect 69572 536726 69624 536732
rect 68650 536616 68706 536625
rect 68650 536551 68706 536560
rect 68664 535537 68692 536551
rect 69584 535537 69612 536726
rect 68650 535528 68706 535537
rect 68650 535463 68706 535472
rect 69570 535528 69626 535537
rect 69570 535463 69626 535472
rect 68284 476128 68336 476134
rect 68284 476070 68336 476076
rect 68928 476128 68980 476134
rect 68928 476070 68980 476076
rect 67640 456816 67692 456822
rect 67640 456758 67692 456764
rect 68836 456816 68888 456822
rect 68836 456758 68888 456764
rect 68848 456074 68876 456758
rect 67640 456068 67692 456074
rect 67640 456010 67692 456016
rect 68652 456068 68704 456074
rect 68652 456010 68704 456016
rect 68836 456068 68888 456074
rect 68836 456010 68888 456016
rect 67652 439929 67680 456010
rect 68664 455462 68692 456010
rect 68652 455456 68704 455462
rect 68652 455398 68704 455404
rect 68836 449200 68888 449206
rect 68836 449142 68888 449148
rect 68848 448594 68876 449142
rect 68836 448588 68888 448594
rect 68836 448530 68888 448536
rect 68848 446434 68876 448530
rect 68940 447098 68968 476070
rect 70214 447128 70270 447137
rect 68928 447092 68980 447098
rect 70214 447063 70270 447072
rect 68928 447034 68980 447040
rect 68664 446406 68876 446434
rect 67824 442944 67876 442950
rect 67824 442886 67876 442892
rect 67836 442241 67864 442886
rect 67822 442232 67878 442241
rect 67822 442167 67878 442176
rect 67638 439920 67694 439929
rect 67638 439855 67694 439864
rect 67652 438938 67680 439855
rect 67640 438932 67692 438938
rect 67640 438874 67692 438880
rect 67730 419656 67786 419665
rect 67730 419591 67786 419600
rect 67546 394904 67602 394913
rect 67546 394839 67602 394848
rect 67560 372638 67588 394839
rect 67548 372632 67600 372638
rect 67548 372574 67600 372580
rect 67456 311160 67508 311166
rect 67456 311102 67508 311108
rect 67468 310729 67496 311102
rect 67454 310720 67510 310729
rect 67454 310655 67510 310664
rect 67086 306368 67142 306377
rect 67086 306303 67142 306312
rect 66996 283620 67048 283626
rect 66996 283562 67048 283568
rect 67100 279478 67128 306303
rect 67560 299849 67588 372574
rect 67744 367810 67772 419591
rect 67732 367804 67784 367810
rect 67732 367746 67784 367752
rect 67836 349858 67864 442167
rect 68664 389337 68692 446406
rect 68742 445904 68798 445913
rect 68742 445839 68798 445848
rect 68756 444380 68784 445839
rect 70228 444380 70256 447063
rect 70412 446457 70440 539566
rect 70780 539294 71530 539322
rect 70780 528554 70808 539294
rect 70504 528526 70808 528554
rect 70504 527542 70532 528526
rect 70492 527536 70544 527542
rect 70492 527478 70544 527484
rect 71044 527536 71096 527542
rect 71044 527478 71096 527484
rect 71056 527202 71084 527478
rect 71044 527196 71096 527202
rect 71044 527138 71096 527144
rect 71056 447166 71084 527138
rect 71044 447160 71096 447166
rect 71044 447102 71096 447108
rect 70398 446448 70454 446457
rect 71884 446418 71912 539582
rect 72344 539294 72450 539322
rect 73172 539294 73370 539322
rect 73540 539294 74290 539322
rect 75104 539294 75210 539322
rect 75932 539294 76130 539322
rect 76760 539294 77050 539322
rect 77864 539294 77970 539322
rect 78692 539294 78890 539322
rect 79060 539294 79810 539322
rect 80072 539294 80730 539322
rect 81544 539294 81650 539322
rect 81820 539294 82570 539322
rect 82832 539294 83490 539322
rect 84304 539294 84410 539322
rect 84580 539294 85330 539322
rect 86342 539294 86632 539322
rect 72344 538214 72372 539294
rect 72344 538186 72464 538214
rect 72436 536761 72464 538186
rect 72422 536752 72478 536761
rect 72422 536687 72478 536696
rect 72436 461718 72464 536687
rect 73172 536110 73200 539294
rect 73160 536104 73212 536110
rect 73160 536046 73212 536052
rect 73540 528554 73568 539294
rect 75104 538214 75132 539294
rect 75104 538186 75224 538214
rect 75196 536790 75224 538186
rect 75184 536784 75236 536790
rect 75184 536726 75236 536732
rect 73264 528526 73568 528554
rect 72424 461712 72476 461718
rect 72424 461654 72476 461660
rect 73264 458862 73292 528526
rect 73252 458856 73304 458862
rect 73252 458798 73304 458804
rect 75196 453354 75224 536726
rect 75932 454714 75960 539294
rect 76760 538286 76788 539294
rect 76748 538280 76800 538286
rect 76748 538222 76800 538228
rect 76564 534064 76616 534070
rect 76564 534006 76616 534012
rect 76576 461514 76604 534006
rect 77864 532846 77892 539294
rect 77852 532840 77904 532846
rect 77852 532782 77904 532788
rect 77864 528554 77892 532782
rect 77864 528526 77984 528554
rect 76012 461508 76064 461514
rect 76012 461450 76064 461456
rect 76564 461508 76616 461514
rect 76564 461450 76616 461456
rect 75920 454708 75972 454714
rect 75920 454650 75972 454656
rect 75184 453348 75236 453354
rect 75184 453290 75236 453296
rect 73160 447092 73212 447098
rect 73160 447034 73212 447040
rect 70398 446383 70454 446392
rect 71872 446412 71924 446418
rect 71872 446354 71924 446360
rect 71778 445904 71834 445913
rect 71778 445839 71834 445848
rect 71792 444380 71820 445839
rect 73172 444380 73200 447034
rect 74816 446412 74868 446418
rect 74816 446354 74868 446360
rect 74828 444380 74856 446354
rect 76024 444394 76052 461450
rect 76576 460970 76604 461450
rect 76564 460964 76616 460970
rect 76564 460906 76616 460912
rect 77956 460222 77984 528526
rect 78036 461644 78088 461650
rect 78036 461586 78088 461592
rect 77944 460216 77996 460222
rect 77944 460158 77996 460164
rect 78048 448633 78076 461586
rect 78692 449274 78720 539294
rect 79060 528554 79088 539294
rect 79324 530596 79376 530602
rect 79324 530538 79376 530544
rect 78784 528526 79088 528554
rect 78784 465730 78812 528526
rect 78772 465724 78824 465730
rect 78772 465666 78824 465672
rect 78680 449268 78732 449274
rect 78680 449210 78732 449216
rect 78034 448624 78090 448633
rect 78034 448559 78090 448568
rect 78048 444394 78076 448559
rect 79336 447098 79364 530538
rect 80072 529242 80100 539294
rect 81544 535634 81572 539294
rect 81532 535628 81584 535634
rect 81532 535570 81584 535576
rect 80060 529236 80112 529242
rect 80060 529178 80112 529184
rect 81820 528554 81848 539294
rect 81452 528526 81848 528554
rect 81452 456249 81480 528526
rect 82832 462913 82860 539294
rect 84304 536518 84332 539294
rect 84292 536512 84344 536518
rect 84292 536454 84344 536460
rect 83464 535628 83516 535634
rect 83464 535570 83516 535576
rect 82818 462904 82874 462913
rect 82818 462839 82874 462848
rect 83476 460193 83504 535570
rect 84580 528554 84608 539294
rect 86604 538214 86632 539294
rect 86972 539294 87354 539322
rect 86604 538186 86908 538214
rect 86880 538150 86908 538186
rect 86868 538144 86920 538150
rect 86868 538086 86920 538092
rect 85580 529304 85632 529310
rect 85580 529246 85632 529252
rect 84212 528526 84608 528554
rect 83462 460184 83518 460193
rect 83462 460119 83518 460128
rect 81438 456240 81494 456249
rect 81438 456175 81494 456184
rect 81440 456068 81492 456074
rect 81440 456010 81492 456016
rect 80888 450560 80940 450566
rect 80888 450502 80940 450508
rect 79324 447092 79376 447098
rect 79324 447034 79376 447040
rect 76024 444366 76314 444394
rect 77878 444366 78076 444394
rect 79336 444394 79364 447034
rect 79414 444544 79470 444553
rect 79414 444479 79470 444488
rect 79428 444394 79456 444479
rect 79336 444380 79456 444394
rect 80900 444380 80928 450502
rect 81452 444394 81480 456010
rect 83832 447840 83884 447846
rect 83832 447782 83884 447788
rect 83844 444553 83872 447782
rect 84212 447273 84240 528526
rect 84198 447264 84254 447273
rect 84198 447199 84254 447208
rect 85592 445777 85620 529246
rect 86880 457473 86908 538086
rect 86866 457464 86922 457473
rect 86866 457399 86922 457408
rect 86972 454753 87000 539294
rect 88168 536625 88196 539582
rect 88366 539294 88656 539322
rect 88628 538218 88656 539294
rect 88616 538212 88668 538218
rect 88616 538154 88668 538160
rect 88154 536616 88210 536625
rect 88154 536551 88210 536560
rect 86958 454744 87014 454753
rect 86958 454679 87014 454688
rect 87052 454096 87104 454102
rect 87052 454038 87104 454044
rect 85578 445768 85634 445777
rect 85578 445703 85634 445712
rect 83830 444544 83886 444553
rect 83830 444479 83886 444488
rect 79336 444366 79442 444380
rect 81452 444366 82386 444394
rect 83844 444380 83872 444479
rect 85592 444380 85620 445703
rect 87064 444689 87092 454038
rect 88996 451274 89024 582346
rect 89626 560144 89682 560153
rect 89626 560079 89682 560088
rect 89640 558958 89668 560079
rect 89628 558952 89680 558958
rect 89628 558894 89680 558900
rect 89626 543824 89682 543833
rect 89626 543759 89682 543768
rect 89640 538218 89668 543759
rect 89732 538898 89760 586191
rect 89824 567361 89852 594050
rect 90362 589928 90418 589937
rect 90362 589863 90418 589872
rect 89810 567352 89866 567361
rect 89810 567287 89866 567296
rect 89824 567254 89852 567287
rect 89812 567248 89864 567254
rect 89812 567190 89864 567196
rect 89720 538892 89772 538898
rect 89720 538834 89772 538840
rect 89628 538212 89680 538218
rect 89628 538154 89680 538160
rect 89076 536512 89128 536518
rect 89076 536454 89128 536460
rect 89088 459649 89116 536454
rect 89640 535498 89668 538154
rect 89628 535492 89680 535498
rect 89628 535434 89680 535440
rect 89074 459640 89130 459649
rect 89074 459575 89130 459584
rect 88904 451246 89024 451274
rect 88904 447166 88932 451246
rect 88892 447160 88944 447166
rect 88892 447102 88944 447108
rect 87050 444680 87106 444689
rect 87050 444615 87106 444624
rect 87064 444380 87092 444615
rect 88904 444394 88932 447102
rect 90376 445806 90404 589863
rect 91112 576745 91140 594390
rect 93766 589384 93822 589393
rect 93766 589319 93822 589328
rect 93124 587716 93176 587722
rect 93124 587658 93176 587664
rect 91742 587616 91798 587625
rect 91742 587551 91798 587560
rect 91756 586566 91784 587551
rect 91744 586560 91796 586566
rect 91744 586502 91796 586508
rect 91374 584896 91430 584905
rect 91374 584831 91430 584840
rect 91388 584458 91416 584831
rect 91376 584452 91428 584458
rect 91376 584394 91428 584400
rect 91192 583704 91244 583710
rect 91190 583672 91192 583681
rect 91244 583672 91246 583681
rect 91190 583607 91246 583616
rect 91742 582176 91798 582185
rect 91742 582111 91798 582120
rect 91756 581058 91784 582111
rect 91744 581052 91796 581058
rect 91744 580994 91796 581000
rect 91742 580816 91798 580825
rect 91742 580751 91798 580760
rect 91756 579698 91784 580751
rect 91744 579692 91796 579698
rect 91744 579634 91796 579640
rect 91742 579456 91798 579465
rect 91742 579391 91798 579400
rect 91756 578270 91784 579391
rect 91744 578264 91796 578270
rect 91744 578206 91796 578212
rect 91098 576736 91154 576745
rect 91098 576671 91154 576680
rect 91112 576162 91140 576671
rect 91100 576156 91152 576162
rect 91100 576098 91152 576104
rect 91098 575376 91154 575385
rect 91098 575311 91154 575320
rect 91112 574122 91140 575311
rect 91100 574116 91152 574122
rect 91100 574058 91152 574064
rect 91098 572656 91154 572665
rect 91098 572591 91154 572600
rect 91112 571402 91140 572591
rect 91190 571432 91246 571441
rect 91100 571396 91152 571402
rect 91190 571367 91246 571376
rect 91100 571338 91152 571344
rect 91098 570072 91154 570081
rect 91098 570007 91100 570016
rect 91152 570007 91154 570016
rect 91100 569978 91152 569984
rect 91204 569226 91232 571367
rect 93136 569974 93164 587658
rect 93124 569968 93176 569974
rect 93124 569910 93176 569916
rect 91192 569220 91244 569226
rect 91192 569162 91244 569168
rect 91098 568712 91154 568721
rect 91098 568647 91154 568656
rect 91112 568614 91140 568647
rect 91100 568608 91152 568614
rect 91100 568550 91152 568556
rect 91376 565888 91428 565894
rect 91374 565856 91376 565865
rect 91428 565856 91430 565865
rect 91374 565791 91430 565800
rect 91374 564496 91430 564505
rect 91374 564431 91376 564440
rect 91428 564431 91430 564440
rect 91376 564402 91428 564408
rect 91374 563136 91430 563145
rect 91374 563071 91376 563080
rect 91428 563071 91430 563080
rect 91376 563042 91428 563048
rect 91098 561504 91154 561513
rect 91098 561439 91154 561448
rect 90456 535492 90508 535498
rect 90456 535434 90508 535440
rect 90468 456113 90496 535434
rect 91112 532030 91140 561439
rect 92386 558784 92442 558793
rect 92386 558719 92442 558728
rect 91190 557424 91246 557433
rect 91190 557359 91246 557368
rect 91204 556238 91232 557359
rect 92400 556850 92428 558719
rect 92388 556844 92440 556850
rect 92388 556786 92440 556792
rect 91192 556232 91244 556238
rect 91192 556174 91244 556180
rect 91742 556064 91798 556073
rect 91742 555999 91798 556008
rect 91756 554810 91784 555999
rect 91744 554804 91796 554810
rect 91744 554746 91796 554752
rect 91742 554704 91798 554713
rect 91742 554639 91798 554648
rect 91756 553450 91784 554639
rect 91744 553444 91796 553450
rect 91744 553386 91796 553392
rect 91742 553344 91798 553353
rect 91742 553279 91798 553288
rect 91756 552158 91784 553279
rect 91744 552152 91796 552158
rect 91190 552120 91246 552129
rect 91744 552094 91796 552100
rect 91190 552055 91192 552064
rect 91244 552055 91246 552064
rect 91192 552026 91244 552032
rect 91190 550760 91246 550769
rect 91190 550695 91246 550704
rect 91204 550662 91232 550695
rect 91192 550656 91244 550662
rect 91192 550598 91244 550604
rect 91480 547942 91508 547973
rect 91468 547936 91520 547942
rect 91466 547904 91468 547913
rect 91520 547904 91522 547913
rect 91466 547839 91522 547848
rect 91190 546544 91246 546553
rect 91190 546479 91192 546488
rect 91244 546479 91246 546488
rect 91192 546450 91244 546456
rect 91204 545306 91232 546450
rect 91204 545278 91324 545306
rect 91190 545184 91246 545193
rect 91190 545119 91192 545128
rect 91244 545119 91246 545128
rect 91192 545090 91244 545096
rect 91190 542464 91246 542473
rect 91190 542399 91192 542408
rect 91244 542399 91246 542408
rect 91192 542370 91244 542376
rect 91192 541680 91244 541686
rect 91192 541622 91244 541628
rect 91204 541249 91232 541622
rect 91190 541240 91246 541249
rect 91190 541175 91246 541184
rect 91296 541090 91324 545278
rect 91204 541062 91324 541090
rect 91204 534750 91232 541062
rect 91480 540954 91508 547839
rect 91834 543960 91890 543969
rect 91834 543895 91890 543904
rect 91848 543794 91876 543895
rect 91836 543788 91888 543794
rect 91836 543730 91888 543736
rect 91296 540926 91508 540954
rect 91296 537538 91324 540926
rect 92386 539744 92442 539753
rect 92386 539679 92442 539688
rect 92400 539646 92428 539679
rect 92388 539640 92440 539646
rect 92388 539582 92440 539588
rect 91284 537532 91336 537538
rect 91284 537474 91336 537480
rect 91192 534744 91244 534750
rect 91192 534686 91244 534692
rect 91100 532024 91152 532030
rect 91100 531966 91152 531972
rect 90454 456104 90510 456113
rect 90454 456039 90510 456048
rect 91100 450628 91152 450634
rect 91100 450570 91152 450576
rect 91112 449954 91140 450570
rect 91100 449948 91152 449954
rect 91100 449890 91152 449896
rect 91560 449948 91612 449954
rect 91560 449890 91612 449896
rect 90364 445800 90416 445806
rect 90364 445742 90416 445748
rect 90376 444394 90404 445742
rect 88550 444366 88932 444394
rect 90206 444366 90404 444394
rect 91572 444380 91600 449890
rect 93032 444508 93084 444514
rect 93032 444450 93084 444456
rect 93044 444394 93072 444450
rect 93136 444394 93164 569910
rect 93676 543788 93728 543794
rect 93676 543730 93728 543736
rect 93216 539640 93268 539646
rect 93216 539582 93268 539588
rect 93228 464409 93256 539582
rect 93688 534721 93716 543730
rect 93674 534712 93730 534721
rect 93674 534647 93730 534656
rect 93214 464400 93270 464409
rect 93214 464335 93270 464344
rect 93780 463010 93808 589319
rect 95160 584458 95188 702578
rect 99288 702500 99340 702506
rect 99288 702442 99340 702448
rect 98644 599004 98696 599010
rect 98644 598946 98696 598952
rect 96620 592136 96672 592142
rect 96620 592078 96672 592084
rect 95240 586560 95292 586566
rect 95240 586502 95292 586508
rect 95148 584452 95200 584458
rect 95148 584394 95200 584400
rect 94504 570036 94556 570042
rect 94504 569978 94556 569984
rect 94516 566506 94544 569978
rect 94504 566500 94556 566506
rect 94504 566442 94556 566448
rect 95146 549400 95202 549409
rect 95146 549335 95202 549344
rect 94504 545148 94556 545154
rect 94504 545090 94556 545096
rect 94516 467129 94544 545090
rect 94502 467120 94558 467129
rect 94502 467055 94558 467064
rect 93768 463004 93820 463010
rect 93768 462946 93820 462952
rect 95160 460193 95188 549335
rect 95252 467158 95280 586502
rect 95332 547936 95384 547942
rect 95332 547878 95384 547884
rect 95344 547194 95372 547878
rect 95332 547188 95384 547194
rect 95332 547130 95384 547136
rect 95240 467152 95292 467158
rect 95240 467094 95292 467100
rect 95146 460184 95202 460193
rect 95146 460119 95202 460128
rect 96252 450560 96304 450566
rect 96252 450502 96304 450508
rect 94780 447840 94832 447846
rect 94780 447782 94832 447788
rect 94792 445777 94820 447782
rect 94778 445768 94834 445777
rect 94778 445703 94834 445712
rect 93044 444380 93164 444394
rect 94792 444380 94820 445703
rect 96264 444380 96292 450502
rect 96528 445800 96580 445806
rect 96632 445777 96660 592078
rect 97264 574116 97316 574122
rect 97264 574058 97316 574064
rect 97276 558210 97304 574058
rect 97264 558204 97316 558210
rect 97264 558146 97316 558152
rect 97356 552152 97408 552158
rect 97356 552094 97408 552100
rect 97264 546508 97316 546514
rect 97264 546450 97316 546456
rect 97276 457473 97304 546450
rect 97368 469849 97396 552094
rect 97354 469840 97410 469849
rect 97354 469775 97410 469784
rect 97262 457464 97318 457473
rect 97262 457399 97318 457408
rect 98656 456929 98684 598946
rect 99300 583710 99328 702442
rect 105464 700330 105492 703520
rect 137848 700398 137876 703520
rect 154132 702545 154160 703520
rect 170324 702982 170352 703520
rect 170312 702976 170364 702982
rect 170312 702918 170364 702924
rect 154118 702536 154174 702545
rect 154118 702471 154174 702480
rect 170324 702434 170352 702918
rect 202800 702846 202828 703520
rect 202788 702840 202840 702846
rect 202788 702782 202840 702788
rect 197268 702704 197320 702710
rect 197268 702646 197320 702652
rect 170324 702406 170444 702434
rect 129648 700392 129700 700398
rect 129648 700334 129700 700340
rect 137836 700392 137888 700398
rect 137836 700334 137888 700340
rect 105452 700324 105504 700330
rect 105452 700266 105504 700272
rect 113180 594924 113232 594930
rect 113180 594866 113232 594872
rect 103518 592104 103574 592113
rect 103518 592039 103574 592048
rect 112536 592068 112588 592074
rect 100758 591016 100814 591025
rect 100758 590951 100814 590960
rect 100772 589966 100800 590951
rect 100760 589960 100812 589966
rect 100760 589902 100812 589908
rect 100850 589520 100906 589529
rect 100850 589455 100906 589464
rect 100760 589348 100812 589354
rect 100760 589290 100812 589296
rect 99288 583704 99340 583710
rect 99288 583646 99340 583652
rect 100024 568608 100076 568614
rect 100024 568550 100076 568556
rect 98736 542428 98788 542434
rect 98736 542370 98788 542376
rect 98748 470665 98776 542370
rect 98734 470656 98790 470665
rect 98734 470591 98790 470600
rect 97998 456920 98054 456929
rect 97998 456855 98054 456864
rect 98642 456920 98698 456929
rect 98642 456855 98698 456864
rect 96528 445742 96580 445748
rect 96618 445768 96674 445777
rect 96540 444961 96568 445742
rect 96618 445703 96674 445712
rect 97630 445768 97686 445777
rect 97630 445703 97686 445712
rect 96526 444952 96582 444961
rect 96526 444887 96582 444896
rect 97644 444380 97672 445703
rect 98012 444394 98040 456855
rect 100036 451897 100064 568550
rect 100116 552084 100168 552090
rect 100116 552026 100168 552032
rect 100128 474065 100156 552026
rect 100114 474056 100170 474065
rect 100114 473991 100170 474000
rect 100022 451888 100078 451897
rect 100022 451823 100078 451832
rect 100772 444514 100800 589290
rect 100864 445806 100892 589455
rect 102784 565888 102836 565894
rect 102784 565830 102836 565836
rect 100944 532840 100996 532846
rect 100944 532782 100996 532788
rect 100956 532710 100984 532782
rect 100944 532704 100996 532710
rect 100944 532646 100996 532652
rect 102796 454714 102824 565830
rect 102784 454708 102836 454714
rect 102784 454650 102836 454656
rect 103532 448594 103560 592039
rect 112536 592010 112588 592016
rect 111064 589960 111116 589966
rect 111064 589902 111116 589908
rect 105544 587920 105596 587926
rect 105544 587862 105596 587868
rect 104164 583704 104216 583710
rect 104164 583646 104216 583652
rect 104176 453257 104204 583646
rect 105556 467838 105584 587862
rect 106924 586628 106976 586634
rect 106924 586570 106976 586576
rect 106188 554804 106240 554810
rect 106188 554746 106240 554752
rect 105544 467832 105596 467838
rect 105544 467774 105596 467780
rect 105556 466478 105584 467774
rect 104900 466472 104952 466478
rect 104900 466414 104952 466420
rect 105544 466472 105596 466478
rect 105544 466414 105596 466420
rect 104162 453248 104218 453257
rect 104162 453183 104218 453192
rect 103520 448588 103572 448594
rect 103520 448530 103572 448536
rect 103704 448588 103756 448594
rect 103704 448530 103756 448536
rect 100852 445800 100904 445806
rect 100850 445768 100852 445777
rect 102232 445800 102284 445806
rect 100904 445768 100906 445777
rect 102232 445742 102284 445748
rect 100850 445703 100906 445712
rect 100760 444508 100812 444514
rect 100760 444450 100812 444456
rect 93058 444366 93150 444380
rect 98012 444366 99130 444394
rect 100772 444380 100800 444450
rect 102244 444380 102272 445742
rect 103716 444380 103744 448530
rect 104912 444394 104940 466414
rect 106200 464370 106228 554746
rect 106188 464364 106240 464370
rect 106188 464306 106240 464312
rect 106936 449886 106964 586570
rect 109038 582992 109094 583001
rect 109038 582927 109094 582936
rect 108304 579692 108356 579698
rect 108304 579634 108356 579640
rect 107016 564460 107068 564466
rect 107016 564402 107068 564408
rect 107028 479505 107056 564402
rect 107014 479496 107070 479505
rect 107014 479431 107070 479440
rect 107660 463004 107712 463010
rect 107660 462946 107712 462952
rect 106924 449880 106976 449886
rect 106924 449822 106976 449828
rect 104912 444366 105386 444394
rect 106936 444380 106964 449822
rect 107672 444394 107700 462946
rect 108316 458182 108344 579634
rect 108948 550656 109000 550662
rect 108948 550598 109000 550604
rect 108960 467809 108988 550598
rect 108946 467800 109002 467809
rect 108946 467735 109002 467744
rect 108304 458176 108356 458182
rect 108304 458118 108356 458124
rect 109052 447137 109080 582927
rect 111076 561746 111104 589902
rect 111064 561740 111116 561746
rect 111064 561682 111116 561688
rect 111708 561740 111760 561746
rect 111708 561682 111760 561688
rect 109038 447128 109094 447137
rect 109038 447063 109094 447072
rect 109052 444689 109080 447063
rect 111720 444689 111748 561682
rect 112444 553444 112496 553450
rect 112444 553386 112496 553392
rect 112456 458833 112484 553386
rect 112548 552090 112576 592010
rect 112536 552084 112588 552090
rect 112536 552026 112588 552032
rect 112548 459542 112576 552026
rect 112536 459536 112588 459542
rect 112536 459478 112588 459484
rect 112442 458824 112498 458833
rect 112442 458759 112498 458768
rect 112548 445806 112576 459478
rect 112536 445800 112588 445806
rect 112536 445742 112588 445748
rect 112904 445800 112956 445806
rect 113192 445777 113220 594866
rect 116584 593428 116636 593434
rect 116584 593370 116636 593376
rect 115296 590776 115348 590782
rect 115296 590718 115348 590724
rect 115204 571396 115256 571402
rect 115204 571338 115256 571344
rect 115216 449410 115244 571338
rect 115308 564466 115336 590718
rect 115296 564460 115348 564466
rect 115296 564402 115348 564408
rect 116596 478174 116624 593370
rect 118698 585712 118754 585721
rect 118698 585647 118754 585656
rect 117964 564460 118016 564466
rect 117964 564402 118016 564408
rect 117976 553489 118004 564402
rect 117962 553480 118018 553489
rect 117962 553415 118018 553424
rect 118606 553480 118662 553489
rect 118606 553415 118662 553424
rect 116584 478168 116636 478174
rect 116584 478110 116636 478116
rect 115296 458176 115348 458182
rect 115296 458118 115348 458124
rect 115204 449404 115256 449410
rect 115204 449346 115256 449352
rect 115308 447273 115336 458118
rect 116124 451308 116176 451314
rect 116124 451250 116176 451256
rect 115294 447264 115350 447273
rect 115294 447199 115350 447208
rect 112904 445742 112956 445748
rect 113178 445768 113234 445777
rect 109038 444680 109094 444689
rect 109038 444615 109094 444624
rect 111706 444680 111762 444689
rect 111706 444615 111762 444624
rect 109052 444394 109080 444615
rect 111720 444394 111748 444615
rect 107672 444366 108330 444394
rect 109052 444366 109802 444394
rect 111550 444366 111748 444394
rect 112916 444380 112944 445742
rect 113178 445703 113234 445712
rect 114374 445768 114430 445777
rect 114374 445703 114430 445712
rect 114388 444380 114416 445703
rect 116136 444380 116164 451250
rect 118620 445777 118648 553415
rect 117594 445768 117650 445777
rect 117594 445703 117650 445712
rect 118606 445768 118662 445777
rect 118606 445703 118662 445712
rect 117608 444380 117636 445703
rect 118712 444446 118740 585647
rect 120724 578264 120776 578270
rect 120724 578206 120776 578212
rect 120632 449404 120684 449410
rect 120632 449346 120684 449352
rect 118700 444440 118752 444446
rect 119160 444440 119212 444446
rect 118700 444382 118752 444388
rect 119094 444388 119160 444394
rect 119094 444382 119212 444388
rect 119094 444366 119200 444382
rect 120644 422294 120672 449346
rect 120736 429321 120764 578206
rect 123024 576156 123076 576162
rect 123024 576098 123076 576104
rect 122104 558952 122156 558958
rect 122104 558894 122156 558900
rect 121460 556232 121512 556238
rect 121460 556174 121512 556180
rect 120816 464364 120868 464370
rect 120816 464306 120868 464312
rect 120722 429312 120778 429321
rect 120722 429247 120778 429256
rect 120644 422266 120764 422294
rect 120736 417081 120764 422266
rect 120722 417072 120778 417081
rect 120722 417007 120778 417016
rect 120630 414624 120686 414633
rect 120630 414559 120686 414568
rect 77666 391096 77722 391105
rect 92938 391096 92994 391105
rect 85606 391068 85896 391082
rect 85592 391066 85896 391068
rect 77666 391031 77722 391040
rect 81440 391060 81492 391066
rect 69938 390416 69994 390425
rect 68650 389328 68706 389337
rect 68650 389263 68706 389272
rect 68756 389065 68784 390388
rect 77680 390402 77708 391031
rect 81440 391002 81492 391008
rect 85592 391060 85908 391066
rect 85592 391054 85856 391060
rect 69994 390388 70334 390402
rect 69994 390374 70348 390388
rect 69938 390351 69994 390360
rect 70320 389162 70348 390374
rect 70308 389156 70360 389162
rect 70308 389098 70360 389104
rect 71792 389065 71820 390388
rect 68742 389056 68798 389065
rect 68742 388991 68798 389000
rect 71778 389056 71834 389065
rect 71778 388991 71834 389000
rect 73066 389056 73122 389065
rect 73066 388991 73122 389000
rect 69662 380216 69718 380225
rect 69662 380151 69718 380160
rect 67824 349852 67876 349858
rect 67824 349794 67876 349800
rect 69676 335354 69704 380151
rect 73080 376786 73108 388991
rect 73172 388929 73200 390388
rect 74552 390374 74842 390402
rect 77680 390388 77878 390402
rect 73158 388920 73214 388929
rect 73158 388855 73214 388864
rect 73802 388920 73858 388929
rect 73802 388855 73858 388864
rect 73160 380180 73212 380186
rect 73160 380122 73212 380128
rect 72424 376780 72476 376786
rect 72424 376722 72476 376728
rect 73068 376780 73120 376786
rect 73068 376722 73120 376728
rect 71688 366988 71740 366994
rect 71688 366930 71740 366936
rect 71596 365016 71648 365022
rect 71596 364958 71648 364964
rect 71608 345014 71636 364958
rect 71516 344986 71636 345014
rect 69846 344312 69902 344321
rect 69846 344247 69902 344256
rect 69400 335326 69704 335354
rect 67824 332648 67876 332654
rect 67824 332590 67876 332596
rect 67732 329860 67784 329866
rect 67732 329802 67784 329808
rect 67638 310720 67694 310729
rect 67638 310655 67694 310664
rect 67546 299840 67602 299849
rect 67546 299775 67602 299784
rect 67454 282432 67510 282441
rect 67454 282367 67510 282376
rect 67178 280256 67234 280265
rect 67178 280191 67180 280200
rect 67232 280191 67234 280200
rect 67180 280162 67232 280168
rect 67088 279472 67140 279478
rect 67088 279414 67140 279420
rect 67178 279168 67234 279177
rect 67178 279103 67234 279112
rect 66994 274000 67050 274009
rect 66994 273935 67050 273944
rect 67008 256018 67036 273935
rect 67192 267782 67220 279103
rect 67180 267776 67232 267782
rect 67180 267718 67232 267724
rect 66996 256012 67048 256018
rect 66996 255954 67048 255960
rect 67270 255504 67326 255513
rect 67270 255439 67326 255448
rect 66994 253328 67050 253337
rect 66904 253292 66956 253298
rect 66994 253263 67050 253272
rect 66904 253234 66956 253240
rect 67008 253026 67036 253263
rect 66996 253020 67048 253026
rect 66996 252962 67048 252968
rect 66902 251152 66958 251161
rect 66902 251087 66958 251096
rect 66810 250064 66866 250073
rect 66810 249999 66866 250008
rect 66824 249830 66852 249999
rect 66916 249898 66944 251087
rect 66904 249892 66956 249898
rect 66904 249834 66956 249840
rect 66812 249824 66864 249830
rect 66812 249766 66864 249772
rect 66902 247888 66958 247897
rect 66902 247823 66958 247832
rect 66916 247110 66944 247823
rect 66904 247104 66956 247110
rect 66904 247046 66956 247052
rect 66812 247036 66864 247042
rect 66812 246978 66864 246984
rect 66824 246809 66852 246978
rect 66810 246800 66866 246809
rect 66810 246735 66866 246744
rect 66350 244624 66406 244633
rect 66350 244559 66406 244568
rect 66364 244322 66392 244559
rect 66352 244316 66404 244322
rect 66352 244258 66404 244264
rect 67086 242856 67142 242865
rect 67086 242791 67142 242800
rect 66166 224768 66222 224777
rect 66166 224703 66222 224712
rect 67100 204921 67128 242791
rect 67284 236609 67312 255439
rect 67364 253020 67416 253026
rect 67364 252962 67416 252968
rect 67376 241777 67404 252962
rect 67362 241768 67418 241777
rect 67362 241703 67418 241712
rect 67468 240786 67496 282367
rect 67546 266384 67602 266393
rect 67546 266319 67602 266328
rect 67456 240780 67508 240786
rect 67456 240722 67508 240728
rect 67270 236600 67326 236609
rect 67270 236535 67326 236544
rect 67086 204912 67142 204921
rect 67086 204847 67142 204856
rect 64786 190360 64842 190369
rect 64786 190295 64842 190304
rect 66166 129296 66222 129305
rect 66166 129231 66222 129240
rect 65982 125216 66038 125225
rect 65982 125151 66038 125160
rect 64970 122632 65026 122641
rect 64970 122567 65026 122576
rect 64984 121553 65012 122567
rect 64786 121544 64842 121553
rect 64786 121479 64842 121488
rect 64970 121544 65026 121553
rect 64970 121479 65026 121488
rect 64800 77246 64828 121479
rect 65890 102368 65946 102377
rect 65890 102303 65946 102312
rect 65904 95033 65932 102303
rect 65890 95024 65946 95033
rect 65890 94959 65946 94968
rect 65996 90370 66024 125151
rect 66074 123584 66130 123593
rect 66074 123519 66130 123528
rect 65984 90364 66036 90370
rect 65984 90306 66036 90312
rect 66088 86290 66116 123519
rect 66076 86284 66128 86290
rect 66076 86226 66128 86232
rect 66180 81433 66208 129231
rect 67454 126304 67510 126313
rect 67454 126239 67510 126248
rect 67362 120864 67418 120873
rect 67362 120799 67418 120808
rect 67376 84862 67404 120799
rect 67468 89049 67496 126239
rect 67454 89040 67510 89049
rect 67454 88975 67510 88984
rect 67364 84856 67416 84862
rect 67364 84798 67416 84804
rect 66166 81424 66222 81433
rect 66166 81359 66222 81368
rect 64788 77240 64840 77246
rect 64788 77182 64840 77188
rect 64786 68368 64842 68377
rect 64786 68303 64842 68312
rect 63408 29640 63460 29646
rect 63408 29582 63460 29588
rect 61948 16546 62068 16574
rect 61384 3392 61436 3398
rect 61384 3334 61436 3340
rect 62040 480 62068 16546
rect 63224 3868 63276 3874
rect 63224 3810 63276 3816
rect 63236 480 63264 3810
rect 64800 3466 64828 68303
rect 67560 68241 67588 266319
rect 67652 228993 67680 310655
rect 67744 296585 67772 329802
rect 67836 308553 67864 332590
rect 69400 331294 69428 335326
rect 69388 331288 69440 331294
rect 69388 331230 69440 331236
rect 69400 329474 69428 331230
rect 69860 329633 69888 344247
rect 71516 332178 71544 344986
rect 71700 335354 71728 366930
rect 71608 335326 71728 335354
rect 70768 332172 70820 332178
rect 70768 332114 70820 332120
rect 71504 332172 71556 332178
rect 71504 332114 71556 332120
rect 70030 331800 70086 331809
rect 70030 331735 70086 331744
rect 69846 329624 69902 329633
rect 69846 329559 69902 329568
rect 70044 329474 70072 331735
rect 70780 329474 70808 332114
rect 71608 329474 71636 335326
rect 72238 334112 72294 334121
rect 72238 334047 72294 334056
rect 72252 329474 72280 334047
rect 72436 332654 72464 376722
rect 73066 365800 73122 365809
rect 73066 365735 73122 365744
rect 72424 332648 72476 332654
rect 72424 332590 72476 332596
rect 73080 329474 73108 365735
rect 69000 329446 69428 329474
rect 69736 329446 70072 329474
rect 70472 329446 70808 329474
rect 71208 329446 71636 329474
rect 71944 329446 72280 329474
rect 72680 329446 73108 329474
rect 73172 329474 73200 380122
rect 73816 379545 73844 388855
rect 74552 380866 74580 390374
rect 76392 389094 76420 390388
rect 77680 390374 77892 390388
rect 76656 389156 76708 389162
rect 76656 389098 76708 389104
rect 76380 389088 76432 389094
rect 76380 389030 76432 389036
rect 76392 385665 76420 389030
rect 76378 385656 76434 385665
rect 76378 385591 76434 385600
rect 75826 382936 75882 382945
rect 75826 382871 75882 382880
rect 74540 380860 74592 380866
rect 74540 380802 74592 380808
rect 73802 379536 73858 379545
rect 73802 379471 73858 379480
rect 73816 366994 73844 379471
rect 73804 366988 73856 366994
rect 73804 366930 73856 366936
rect 75736 356788 75788 356794
rect 75736 356730 75788 356736
rect 73804 342916 73856 342922
rect 73804 342858 73856 342864
rect 73816 330546 73844 342858
rect 74264 332512 74316 332518
rect 74264 332454 74316 332460
rect 73804 330540 73856 330546
rect 73804 330482 73856 330488
rect 74276 329474 74304 332454
rect 75182 331256 75238 331265
rect 75182 331191 75238 331200
rect 75196 329474 75224 331191
rect 75748 329474 75776 356730
rect 75840 331265 75868 382871
rect 76564 371884 76616 371890
rect 76564 371826 76616 371832
rect 76576 345014 76604 371826
rect 76668 352578 76696 389098
rect 77864 388482 77892 390374
rect 79520 388793 79548 390388
rect 79506 388784 79562 388793
rect 79506 388719 79562 388728
rect 79520 388550 79548 388719
rect 79508 388544 79560 388550
rect 79508 388486 79560 388492
rect 77852 388476 77904 388482
rect 77852 388418 77904 388424
rect 80900 387025 80928 390388
rect 81452 389065 81480 391002
rect 82096 390374 82386 390402
rect 82832 390374 83858 390402
rect 81438 389056 81494 389065
rect 81438 388991 81494 389000
rect 82096 387802 82124 390374
rect 82084 387796 82136 387802
rect 82084 387738 82136 387744
rect 79966 387016 80022 387025
rect 79966 386951 80022 386960
rect 80886 387016 80942 387025
rect 80886 386951 80942 386960
rect 79980 381546 80008 386951
rect 79968 381540 80020 381546
rect 79968 381482 80020 381488
rect 81346 373416 81402 373425
rect 81346 373351 81402 373360
rect 77944 366444 77996 366450
rect 77944 366386 77996 366392
rect 76746 353424 76802 353433
rect 76746 353359 76802 353368
rect 76656 352572 76708 352578
rect 76656 352514 76708 352520
rect 76576 344986 76696 345014
rect 75826 331256 75882 331265
rect 75826 331191 75882 331200
rect 76668 329905 76696 344986
rect 76760 332518 76788 353359
rect 77300 337476 77352 337482
rect 77300 337418 77352 337424
rect 77114 337376 77170 337385
rect 77114 337311 77170 337320
rect 76748 332512 76800 332518
rect 76748 332454 76800 332460
rect 76654 329896 76710 329905
rect 76654 329831 76710 329840
rect 76668 329474 76696 329831
rect 77128 329746 77156 337311
rect 77312 329866 77340 337418
rect 77300 329860 77352 329866
rect 77300 329802 77352 329808
rect 73172 329446 73416 329474
rect 74152 329446 74304 329474
rect 74888 329446 75224 329474
rect 75624 329446 75776 329474
rect 76360 329446 76696 329474
rect 77082 329718 77156 329746
rect 77082 329460 77110 329718
rect 77482 329216 77538 329225
rect 77956 329202 77984 366386
rect 81360 359514 81388 373351
rect 82096 362234 82124 387738
rect 82832 383654 82860 390374
rect 85592 389298 85620 391054
rect 92994 391068 93058 391082
rect 92994 391054 93072 391068
rect 92938 391031 92994 391040
rect 85856 391002 85908 391008
rect 89810 390416 89866 390425
rect 85580 389292 85632 389298
rect 85580 389234 85632 389240
rect 82820 383648 82872 383654
rect 82820 383590 82872 383596
rect 82084 362228 82136 362234
rect 82084 362170 82136 362176
rect 82096 361622 82124 362170
rect 81624 361616 81676 361622
rect 81624 361558 81676 361564
rect 82084 361616 82136 361622
rect 82084 361558 82136 361564
rect 80152 359508 80204 359514
rect 80152 359450 80204 359456
rect 81348 359508 81400 359514
rect 81348 359450 81400 359456
rect 79324 358148 79376 358154
rect 79324 358090 79376 358096
rect 79336 332178 79364 358090
rect 80164 345014 80192 359450
rect 81348 355360 81400 355366
rect 81348 355302 81400 355308
rect 80164 344986 80376 345014
rect 79692 344344 79744 344350
rect 79692 344286 79744 344292
rect 78588 332172 78640 332178
rect 78588 332114 78640 332120
rect 79324 332172 79376 332178
rect 79324 332114 79376 332120
rect 78600 329746 78628 332114
rect 78554 329718 78628 329746
rect 78554 329460 78582 329718
rect 79704 329474 79732 344286
rect 80244 331628 80296 331634
rect 80244 331570 80296 331576
rect 80256 329474 80284 331570
rect 79304 329446 79732 329474
rect 80040 329446 80284 329474
rect 80348 329474 80376 344986
rect 81360 331634 81388 355302
rect 81636 345014 81664 361558
rect 81636 344986 81848 345014
rect 81438 339552 81494 339561
rect 81438 339487 81494 339496
rect 81348 331628 81400 331634
rect 81348 331570 81400 331576
rect 81452 329746 81480 339487
rect 81452 329718 81526 329746
rect 80348 329446 80776 329474
rect 81498 329460 81526 329718
rect 81820 329474 81848 344986
rect 82832 337414 82860 383590
rect 84844 370524 84896 370530
rect 84844 370466 84896 370472
rect 84108 345772 84160 345778
rect 84108 345714 84160 345720
rect 82820 337408 82872 337414
rect 82820 337350 82872 337356
rect 83372 333260 83424 333266
rect 83372 333202 83424 333208
rect 83096 331356 83148 331362
rect 83096 331298 83148 331304
rect 83108 329474 83136 331298
rect 81820 329446 82248 329474
rect 82800 329446 83136 329474
rect 77538 329174 77984 329202
rect 83186 329216 83242 329225
rect 77482 329151 77538 329160
rect 83384 329202 83412 333202
rect 84120 331362 84148 345714
rect 84660 335368 84712 335374
rect 84856 335354 84884 370466
rect 85396 342304 85448 342310
rect 85396 342246 85448 342252
rect 84712 335326 84884 335354
rect 84660 335310 84712 335316
rect 84108 331356 84160 331362
rect 84108 331298 84160 331304
rect 84672 329474 84700 335310
rect 85408 329474 85436 342246
rect 85592 337482 85620 389234
rect 86224 388544 86276 388550
rect 86224 388486 86276 388492
rect 86236 367878 86264 388486
rect 86972 386374 87000 390388
rect 88536 387870 88564 390388
rect 89866 390374 90496 390402
rect 89810 390351 89866 390360
rect 90468 388929 90496 390374
rect 91664 389162 91692 390388
rect 91652 389156 91704 389162
rect 91652 389098 91704 389104
rect 91664 389065 91692 389098
rect 91650 389056 91706 389065
rect 91650 388991 91706 389000
rect 90454 388920 90510 388929
rect 90454 388855 90510 388864
rect 88524 387864 88576 387870
rect 88524 387806 88576 387812
rect 90364 387864 90416 387870
rect 90364 387806 90416 387812
rect 86960 386368 87012 386374
rect 86960 386310 87012 386316
rect 86224 367872 86276 367878
rect 86224 367814 86276 367820
rect 86868 349920 86920 349926
rect 86868 349862 86920 349868
rect 85670 338192 85726 338201
rect 85670 338127 85726 338136
rect 85580 337476 85632 337482
rect 85580 337418 85632 337424
rect 85684 329746 85712 338127
rect 85684 329718 85758 329746
rect 84272 329446 84700 329474
rect 85008 329446 85436 329474
rect 85730 329460 85758 329718
rect 86880 329474 86908 349862
rect 86972 341562 87000 386310
rect 89626 371376 89682 371385
rect 89626 371311 89682 371320
rect 87602 370560 87658 370569
rect 87602 370495 87658 370504
rect 87616 345014 87644 370495
rect 87156 344986 87644 345014
rect 87156 342281 87184 344986
rect 87142 342272 87198 342281
rect 87142 342207 87198 342216
rect 86960 341556 87012 341562
rect 86960 341498 87012 341504
rect 87156 329746 87184 342207
rect 89534 341048 89590 341057
rect 89534 340983 89590 340992
rect 88248 332172 88300 332178
rect 88248 332114 88300 332120
rect 87156 329718 87230 329746
rect 86480 329446 86908 329474
rect 87202 329460 87230 329718
rect 88260 329474 88288 332114
rect 88984 331356 89036 331362
rect 88984 331298 89036 331304
rect 88996 329474 89024 331298
rect 89548 329474 89576 340983
rect 89640 331362 89668 371311
rect 90376 353297 90404 387806
rect 90468 383654 90496 388855
rect 93044 388793 93072 391054
rect 115754 390688 115810 390697
rect 115754 390623 115810 390632
rect 94226 390416 94282 390425
rect 97354 390416 97410 390425
rect 94282 390374 95004 390402
rect 94226 390351 94282 390360
rect 93216 389156 93268 389162
rect 93216 389098 93268 389104
rect 93030 388784 93086 388793
rect 93030 388719 93086 388728
rect 90468 383626 90588 383654
rect 90560 361622 90588 383626
rect 92388 376100 92440 376106
rect 92388 376042 92440 376048
rect 90548 361616 90600 361622
rect 90548 361558 90600 361564
rect 90456 360256 90508 360262
rect 90456 360198 90508 360204
rect 90362 353288 90418 353297
rect 90362 353223 90418 353232
rect 90468 332178 90496 360198
rect 90560 342310 90588 361558
rect 91006 351112 91062 351121
rect 91006 351047 91062 351056
rect 90548 342304 90600 342310
rect 90548 342246 90600 342252
rect 90456 332172 90508 332178
rect 90456 332114 90508 332120
rect 90456 331492 90508 331498
rect 90456 331434 90508 331440
rect 89628 331356 89680 331362
rect 89628 331298 89680 331304
rect 90468 329474 90496 331434
rect 91020 329474 91048 351047
rect 91926 330168 91982 330177
rect 91926 330103 91982 330112
rect 91940 329474 91968 330103
rect 92400 329746 92428 376042
rect 93122 369880 93178 369889
rect 93122 369815 93178 369824
rect 93136 331498 93164 369815
rect 93228 354006 93256 389098
rect 94976 383654 95004 390374
rect 96264 389162 96292 390388
rect 98826 390416 98882 390425
rect 97410 390374 97856 390402
rect 97354 390351 97410 390360
rect 96252 389156 96304 389162
rect 96252 389098 96304 389104
rect 96264 389065 96292 389098
rect 95238 389056 95294 389065
rect 95238 388991 95294 389000
rect 96250 389056 96306 389065
rect 96250 388991 96306 389000
rect 95252 385694 95280 388991
rect 95240 385688 95292 385694
rect 95240 385630 95292 385636
rect 94976 383626 95188 383654
rect 95160 364449 95188 383626
rect 97262 374640 97318 374649
rect 97262 374575 97318 374584
rect 93858 364440 93914 364449
rect 93858 364375 93914 364384
rect 95146 364440 95202 364449
rect 95146 364375 95202 364384
rect 93872 358154 93900 364375
rect 93860 358148 93912 358154
rect 93860 358090 93912 358096
rect 96526 356144 96582 356153
rect 96526 356079 96582 356088
rect 94504 354748 94556 354754
rect 94504 354690 94556 354696
rect 93216 354000 93268 354006
rect 93216 353942 93268 353948
rect 93768 347064 93820 347070
rect 93768 347006 93820 347012
rect 93780 335354 93808 347006
rect 94516 335354 94544 354690
rect 96436 351280 96488 351286
rect 96436 351222 96488 351228
rect 95148 340944 95200 340950
rect 95148 340886 95200 340892
rect 93504 335326 93808 335354
rect 94332 335326 94544 335354
rect 93124 331492 93176 331498
rect 93124 331434 93176 331440
rect 87952 329446 88288 329474
rect 88688 329446 89024 329474
rect 89424 329446 89576 329474
rect 90160 329446 90496 329474
rect 90896 329446 91048 329474
rect 91632 329446 91968 329474
rect 92354 329718 92428 329746
rect 92354 329460 92382 329718
rect 93504 329474 93532 335326
rect 94332 333946 94360 335326
rect 94320 333940 94372 333946
rect 94320 333882 94372 333888
rect 94136 331492 94188 331498
rect 94136 331434 94188 331440
rect 94148 329474 94176 331434
rect 93104 329446 93532 329474
rect 93840 329446 94176 329474
rect 94332 329474 94360 333882
rect 95160 331498 95188 340886
rect 95608 331560 95660 331566
rect 95608 331502 95660 331508
rect 95148 331492 95200 331498
rect 95148 331434 95200 331440
rect 95620 329474 95648 331502
rect 96448 329474 96476 351222
rect 96540 331566 96568 356079
rect 97276 341465 97304 374575
rect 97828 360097 97856 390374
rect 102138 390416 102194 390425
rect 98882 390374 99130 390402
rect 98826 390351 98882 390360
rect 99024 366382 99052 390374
rect 100772 390289 100800 390388
rect 104990 390416 105046 390425
rect 102194 390388 102350 390402
rect 102194 390374 102364 390388
rect 103822 390374 104204 390402
rect 102138 390351 102194 390360
rect 100758 390280 100814 390289
rect 100758 390215 100814 390224
rect 100772 389065 100800 390215
rect 102336 389065 102364 390374
rect 99194 389056 99250 389065
rect 99194 388991 99250 389000
rect 100758 389056 100814 389065
rect 100758 388991 100814 389000
rect 102322 389056 102378 389065
rect 102322 388991 102378 389000
rect 103334 389056 103390 389065
rect 103334 388991 103390 389000
rect 99012 366376 99064 366382
rect 99012 366318 99064 366324
rect 97814 360088 97870 360097
rect 97814 360023 97870 360032
rect 99104 358828 99156 358834
rect 99104 358770 99156 358776
rect 98826 356960 98882 356969
rect 98826 356895 98882 356904
rect 98840 356794 98868 356895
rect 98828 356788 98880 356794
rect 98828 356730 98880 356736
rect 97908 342984 97960 342990
rect 97908 342926 97960 342932
rect 97262 341456 97318 341465
rect 97262 341391 97318 341400
rect 97814 332888 97870 332897
rect 97814 332823 97870 332832
rect 96528 331560 96580 331566
rect 96528 331502 96580 331508
rect 97080 331356 97132 331362
rect 97080 331298 97132 331304
rect 97092 329474 97120 331298
rect 97828 329474 97856 332823
rect 97920 331362 97948 342926
rect 98552 332036 98604 332042
rect 98552 331978 98604 331984
rect 97908 331356 97960 331362
rect 97908 331298 97960 331304
rect 98564 329474 98592 331978
rect 99116 329474 99144 358770
rect 99208 356969 99236 388991
rect 101402 388784 101458 388793
rect 101402 388719 101458 388728
rect 101416 378826 101444 388719
rect 101404 378820 101456 378826
rect 101404 378762 101456 378768
rect 101404 373312 101456 373318
rect 101404 373254 101456 373260
rect 99286 371920 99342 371929
rect 99286 371855 99342 371864
rect 99194 356960 99250 356969
rect 99194 356895 99250 356904
rect 99300 332042 99328 371855
rect 100022 370016 100078 370025
rect 100022 369951 100078 369960
rect 100036 349926 100064 369951
rect 100024 349920 100076 349926
rect 100024 349862 100076 349868
rect 100666 349752 100722 349761
rect 100666 349687 100722 349696
rect 100574 346488 100630 346497
rect 100574 346423 100630 346432
rect 99288 332036 99340 332042
rect 99288 331978 99340 331984
rect 100024 331492 100076 331498
rect 100024 331434 100076 331440
rect 100036 329474 100064 331434
rect 100588 329474 100616 346423
rect 100680 331498 100708 349687
rect 101416 337521 101444 373254
rect 103348 360874 103376 388991
rect 104176 387802 104204 390374
rect 106554 390416 106610 390425
rect 105046 390374 105386 390402
rect 104990 390351 105046 390360
rect 108026 390416 108082 390425
rect 106610 390374 107240 390402
rect 106554 390351 106610 390360
rect 104164 387796 104216 387802
rect 104164 387738 104216 387744
rect 103428 362976 103480 362982
rect 103428 362918 103480 362924
rect 103336 360868 103388 360874
rect 103336 360810 103388 360816
rect 103334 355328 103390 355337
rect 103334 355263 103390 355272
rect 101496 351960 101548 351966
rect 101496 351902 101548 351908
rect 101402 337512 101458 337521
rect 101402 337447 101458 337456
rect 101508 332586 101536 351902
rect 102046 344040 102102 344049
rect 102046 343975 102102 343984
rect 101496 332580 101548 332586
rect 101496 332522 101548 332528
rect 100668 331492 100720 331498
rect 100668 331434 100720 331440
rect 101508 329474 101536 332522
rect 102060 329474 102088 343975
rect 103348 335354 103376 355263
rect 103072 335326 103376 335354
rect 103072 329474 103100 335326
rect 103440 329746 103468 362918
rect 103520 357468 103572 357474
rect 103520 357410 103572 357416
rect 103532 345014 103560 357410
rect 103532 344986 103744 345014
rect 94332 329446 94576 329474
rect 95312 329446 95648 329474
rect 96048 329446 96476 329474
rect 96784 329446 97120 329474
rect 97520 329446 97856 329474
rect 98256 329446 98592 329474
rect 98992 329446 99144 329474
rect 99728 329446 100064 329474
rect 100464 329446 100616 329474
rect 101200 329446 101536 329474
rect 101936 329446 102088 329474
rect 102672 329446 103100 329474
rect 103394 329718 103468 329746
rect 103394 329460 103422 329718
rect 103716 329474 103744 344986
rect 104176 340105 104204 387738
rect 105004 381041 105032 390351
rect 106922 388376 106978 388385
rect 106922 388311 106978 388320
rect 106186 381576 106242 381585
rect 106186 381511 106242 381520
rect 104990 381032 105046 381041
rect 104990 380967 105046 380976
rect 105542 381032 105598 381041
rect 105542 380967 105598 380976
rect 104900 353388 104952 353394
rect 104900 353330 104952 353336
rect 104162 340096 104218 340105
rect 104162 340031 104218 340040
rect 104912 329746 104940 353330
rect 105556 348430 105584 380967
rect 105544 348424 105596 348430
rect 105544 348366 105596 348372
rect 106200 346361 106228 381511
rect 104990 346352 105046 346361
rect 104990 346287 105046 346296
rect 106186 346352 106242 346361
rect 106186 346287 106242 346296
rect 105004 345014 105032 346287
rect 106200 345817 106228 346287
rect 106186 345808 106242 345817
rect 106186 345743 106242 345752
rect 105004 344986 105216 345014
rect 104866 329718 104940 329746
rect 103716 329446 104144 329474
rect 104866 329460 104894 329718
rect 105188 329474 105216 344986
rect 106936 333266 106964 388311
rect 107212 385694 107240 390374
rect 109498 390416 109554 390425
rect 108082 390388 108422 390402
rect 108082 390374 108436 390388
rect 108026 390351 108082 390360
rect 108408 389337 108436 390374
rect 109554 390374 110276 390402
rect 109498 390351 109554 390360
rect 108394 389328 108450 389337
rect 108394 389263 108450 389272
rect 107200 385688 107252 385694
rect 107200 385630 107252 385636
rect 110248 383654 110276 390374
rect 111444 389230 111472 390388
rect 110420 389224 110472 389230
rect 110420 389166 110472 389172
rect 111432 389224 111484 389230
rect 111432 389166 111484 389172
rect 110248 383626 110368 383654
rect 110234 357504 110290 357513
rect 110234 357439 110290 357448
rect 107752 356720 107804 356726
rect 107752 356662 107804 356668
rect 107764 351257 107792 356662
rect 107750 351248 107806 351257
rect 107750 351183 107806 351192
rect 107764 345014 107792 351183
rect 108486 349208 108542 349217
rect 108486 349143 108542 349152
rect 108500 345778 108528 349143
rect 108488 345772 108540 345778
rect 108488 345714 108540 345720
rect 107764 344986 107976 345014
rect 107384 337408 107436 337414
rect 107384 337350 107436 337356
rect 106924 333260 106976 333266
rect 106924 333202 106976 333208
rect 106648 332648 106700 332654
rect 106648 332590 106700 332596
rect 106660 329474 106688 332590
rect 107396 329474 107424 337350
rect 107844 331900 107896 331906
rect 107844 331842 107896 331848
rect 107856 329474 107884 331842
rect 105188 329446 105616 329474
rect 106352 329446 106688 329474
rect 107088 329446 107424 329474
rect 107640 329446 107884 329474
rect 107948 329474 107976 344986
rect 109408 331560 109460 331566
rect 109408 331502 109460 331508
rect 109420 329474 109448 331502
rect 110248 329474 110276 357439
rect 110340 356726 110368 383626
rect 110328 356720 110380 356726
rect 110328 356662 110380 356668
rect 110432 349926 110460 389166
rect 112916 389065 112944 390388
rect 113088 389836 113140 389842
rect 113088 389778 113140 389784
rect 112902 389056 112958 389065
rect 112902 388991 112958 389000
rect 113100 383722 113128 389778
rect 114388 389065 114416 390388
rect 113178 389056 113234 389065
rect 113178 388991 113234 389000
rect 114374 389056 114430 389065
rect 114374 388991 114430 389000
rect 111800 383716 111852 383722
rect 111800 383658 111852 383664
rect 113088 383716 113140 383722
rect 113088 383658 113140 383664
rect 111062 381032 111118 381041
rect 111062 380967 111118 380976
rect 110420 349920 110472 349926
rect 110420 349862 110472 349868
rect 110328 344412 110380 344418
rect 110328 344354 110380 344360
rect 110340 331566 110368 344354
rect 111076 344350 111104 380967
rect 111706 348392 111762 348401
rect 111706 348327 111762 348336
rect 111064 344344 111116 344350
rect 111064 344286 111116 344292
rect 111614 340912 111670 340921
rect 111614 340847 111670 340856
rect 111628 332178 111656 340847
rect 110880 332172 110932 332178
rect 110880 332114 110932 332120
rect 111616 332172 111668 332178
rect 111616 332114 111668 332120
rect 110328 331560 110380 331566
rect 110328 331502 110380 331508
rect 110892 329474 110920 332114
rect 111720 329474 111748 348327
rect 107948 329446 108376 329474
rect 109112 329446 109448 329474
rect 109848 329446 110276 329474
rect 110584 329446 110920 329474
rect 111320 329446 111748 329474
rect 111812 329474 111840 383658
rect 113192 353433 113220 388991
rect 115662 379264 115718 379273
rect 115662 379199 115718 379208
rect 115676 378321 115704 379199
rect 115662 378312 115718 378321
rect 115662 378247 115718 378256
rect 114558 376544 114614 376553
rect 114558 376479 114614 376488
rect 113178 353424 113234 353433
rect 113178 353359 113234 353368
rect 113822 353424 113878 353433
rect 113822 353359 113878 353368
rect 113836 343641 113864 353359
rect 114468 343732 114520 343738
rect 114468 343674 114520 343680
rect 113822 343632 113878 343641
rect 113822 343567 113878 343576
rect 112350 339688 112406 339697
rect 112350 339623 112406 339632
rect 112364 329474 112392 339623
rect 114480 332178 114508 343674
rect 113824 332172 113876 332178
rect 113824 332114 113876 332120
rect 114468 332172 114520 332178
rect 114468 332114 114520 332120
rect 113836 329474 113864 332114
rect 114466 331256 114522 331265
rect 114466 331191 114522 331200
rect 114480 329474 114508 331191
rect 114572 329730 114600 376479
rect 115676 376106 115704 378247
rect 115768 376553 115796 390623
rect 115938 390416 115994 390425
rect 117870 390416 117926 390425
rect 115994 390374 116532 390402
rect 117622 390388 117870 390402
rect 115938 390351 115994 390360
rect 116504 377505 116532 390374
rect 117608 390374 117870 390388
rect 117608 384334 117636 390374
rect 117870 390351 117926 390360
rect 118790 390416 118846 390425
rect 118846 390374 119384 390402
rect 118790 390351 118846 390360
rect 117596 384328 117648 384334
rect 117596 384270 117648 384276
rect 119356 383761 119384 390374
rect 120460 390318 120488 390388
rect 120448 390312 120500 390318
rect 120448 390254 120500 390260
rect 120460 388385 120488 390254
rect 120446 388376 120502 388385
rect 120446 388311 120502 388320
rect 119342 383752 119398 383761
rect 119342 383687 119398 383696
rect 116490 377496 116546 377505
rect 116490 377431 116546 377440
rect 115754 376544 115810 376553
rect 115754 376479 115810 376488
rect 115664 376100 115716 376106
rect 115664 376042 115716 376048
rect 115768 375465 115796 376479
rect 115754 375456 115810 375465
rect 115754 375391 115810 375400
rect 116582 367704 116638 367713
rect 116582 367639 116638 367648
rect 115846 361040 115902 361049
rect 115846 360975 115902 360984
rect 115860 332178 115888 360975
rect 116596 338774 116624 367639
rect 116674 364576 116730 364585
rect 116674 364511 116730 364520
rect 116688 344418 116716 364511
rect 118606 353424 118662 353433
rect 118606 353359 118662 353368
rect 116676 344412 116728 344418
rect 116676 344354 116728 344360
rect 118514 339416 118570 339425
rect 118514 339351 118570 339360
rect 116584 338768 116636 338774
rect 116584 338710 116636 338716
rect 118528 338230 118556 339351
rect 118516 338224 118568 338230
rect 118516 338166 118568 338172
rect 117228 338156 117280 338162
rect 117228 338098 117280 338104
rect 117042 332616 117098 332625
rect 117042 332551 117098 332560
rect 115296 332172 115348 332178
rect 115296 332114 115348 332120
rect 115848 332172 115900 332178
rect 115848 332114 115900 332120
rect 116768 332172 116820 332178
rect 116768 332114 116820 332120
rect 114560 329724 114612 329730
rect 114560 329666 114612 329672
rect 111812 329446 112056 329474
rect 112364 329446 112792 329474
rect 113528 329446 113864 329474
rect 114264 329446 114508 329474
rect 83242 329174 83536 329202
rect 83186 329151 83242 329160
rect 114572 329118 114600 329666
rect 115308 329474 115336 332114
rect 115710 329724 115762 329730
rect 115710 329666 115762 329672
rect 115000 329446 115336 329474
rect 115722 329460 115750 329666
rect 116780 329474 116808 332114
rect 116472 329446 116808 329474
rect 117056 329338 117084 332551
rect 117240 332178 117268 338098
rect 118528 332178 118556 338166
rect 117228 332172 117280 332178
rect 117228 332114 117280 332120
rect 118516 332172 118568 332178
rect 118516 332114 118568 332120
rect 118620 329746 118648 353359
rect 119356 345778 119384 383687
rect 119986 378176 120042 378185
rect 119986 378111 120042 378120
rect 120000 374066 120028 378111
rect 119988 374060 120040 374066
rect 119988 374002 120040 374008
rect 119344 345772 119396 345778
rect 119344 345714 119396 345720
rect 119894 343904 119950 343913
rect 119894 343839 119950 343848
rect 119068 332172 119120 332178
rect 119068 332114 119120 332120
rect 118976 331356 119028 331362
rect 118976 331298 119028 331304
rect 118344 329718 118648 329746
rect 118344 329474 118372 329718
rect 118988 329474 119016 331298
rect 117944 329446 118372 329474
rect 118680 329446 119016 329474
rect 119080 329474 119108 332114
rect 119908 331362 119936 343839
rect 120000 331362 120028 374002
rect 120644 353326 120672 414559
rect 120736 389842 120764 417007
rect 120828 390318 120856 464306
rect 121184 415404 121236 415410
rect 121184 415346 121236 415352
rect 121196 415313 121224 415346
rect 121182 415304 121238 415313
rect 121182 415239 121238 415248
rect 121472 392737 121500 556174
rect 121552 451920 121604 451926
rect 121552 451862 121604 451868
rect 121564 440065 121592 451862
rect 121644 444440 121696 444446
rect 121644 444382 121696 444388
rect 121656 442241 121684 444382
rect 121642 442232 121698 442241
rect 121642 442167 121698 442176
rect 121550 440056 121606 440065
rect 121550 439991 121606 440000
rect 121550 435432 121606 435441
rect 121550 435367 121606 435376
rect 121458 392728 121514 392737
rect 121458 392663 121514 392672
rect 121472 392086 121500 392663
rect 121460 392080 121512 392086
rect 121460 392022 121512 392028
rect 120816 390312 120868 390318
rect 120816 390254 120868 390260
rect 120724 389836 120776 389842
rect 120724 389778 120776 389784
rect 120722 387016 120778 387025
rect 120722 386951 120778 386960
rect 120736 370530 120764 386951
rect 121564 381585 121592 435367
rect 122116 407114 122144 558894
rect 122932 558204 122984 558210
rect 122932 558146 122984 558152
rect 122748 429140 122800 429146
rect 122748 429082 122800 429088
rect 122760 428505 122788 429082
rect 122746 428496 122802 428505
rect 122746 428431 122802 428440
rect 122104 407108 122156 407114
rect 122104 407050 122156 407056
rect 121550 381576 121606 381585
rect 121550 381511 121606 381520
rect 120724 370524 120776 370530
rect 120724 370466 120776 370472
rect 121458 358048 121514 358057
rect 121458 357983 121514 357992
rect 120724 354000 120776 354006
rect 120724 353942 120776 353948
rect 120632 353320 120684 353326
rect 120632 353262 120684 353268
rect 120644 351286 120672 353262
rect 120632 351280 120684 351286
rect 120632 351222 120684 351228
rect 120736 344350 120764 353942
rect 120724 344344 120776 344350
rect 120724 344286 120776 344292
rect 120736 343670 120764 344286
rect 120080 343664 120132 343670
rect 120080 343606 120132 343612
rect 120724 343664 120776 343670
rect 120724 343606 120776 343612
rect 119896 331356 119948 331362
rect 119896 331298 119948 331304
rect 119988 331356 120040 331362
rect 119988 331298 120040 331304
rect 120092 329746 120120 343606
rect 120540 331356 120592 331362
rect 120540 331298 120592 331304
rect 120092 329718 120166 329746
rect 119080 329446 119416 329474
rect 120138 329460 120166 329718
rect 120552 329474 120580 331298
rect 121472 329474 121500 357983
rect 121734 353968 121790 353977
rect 121734 353903 121790 353912
rect 121552 346452 121604 346458
rect 121552 346394 121604 346400
rect 121564 345681 121592 346394
rect 121550 345672 121606 345681
rect 121550 345607 121606 345616
rect 121748 345014 121776 353903
rect 122760 346458 122788 428431
rect 122944 421977 122972 558146
rect 123036 424153 123064 576098
rect 126980 569220 127032 569226
rect 126980 569162 127032 569168
rect 126992 568614 127020 569162
rect 126980 568608 127032 568614
rect 126980 568550 127032 568556
rect 124864 550656 124916 550662
rect 124864 550598 124916 550604
rect 124876 528562 124904 550598
rect 126888 546508 126940 546514
rect 126888 546450 126940 546456
rect 124864 528556 124916 528562
rect 124864 528498 124916 528504
rect 124956 527196 125008 527202
rect 124956 527138 125008 527144
rect 124968 510610 124996 527138
rect 124956 510604 125008 510610
rect 124956 510546 125008 510552
rect 124956 465112 125008 465118
rect 124956 465054 125008 465060
rect 124220 452668 124272 452674
rect 124220 452610 124272 452616
rect 123574 451888 123630 451897
rect 123574 451823 123630 451832
rect 123482 426048 123538 426057
rect 123482 425983 123538 425992
rect 123022 424144 123078 424153
rect 123022 424079 123078 424088
rect 122930 421968 122986 421977
rect 122930 421903 122986 421912
rect 122944 421598 122972 421903
rect 122932 421592 122984 421598
rect 122932 421534 122984 421540
rect 123036 412634 123064 424079
rect 122852 412606 123064 412634
rect 122852 348537 122880 412606
rect 123024 407108 123076 407114
rect 123024 407050 123076 407056
rect 123036 397361 123064 407050
rect 123022 397352 123078 397361
rect 123022 397287 123078 397296
rect 122930 394768 122986 394777
rect 122930 394703 122986 394712
rect 122944 384305 122972 394703
rect 122930 384296 122986 384305
rect 122930 384231 122986 384240
rect 123496 382294 123524 425983
rect 123588 411330 123616 451823
rect 124126 442096 124182 442105
rect 124126 442031 124128 442040
rect 124180 442031 124182 442040
rect 124128 442002 124180 442008
rect 124128 438252 124180 438258
rect 124128 438194 124180 438200
rect 124140 437889 124168 438194
rect 124126 437880 124182 437889
rect 124126 437815 124182 437824
rect 124126 433120 124182 433129
rect 124126 433055 124182 433064
rect 124140 432614 124168 433055
rect 124128 432608 124180 432614
rect 124128 432550 124180 432556
rect 124128 431928 124180 431934
rect 124128 431870 124180 431876
rect 124140 431089 124168 431870
rect 124126 431080 124182 431089
rect 124126 431015 124182 431024
rect 124128 420912 124180 420918
rect 124126 420880 124128 420889
rect 124180 420880 124182 420889
rect 124126 420815 124182 420824
rect 123852 413296 123904 413302
rect 123852 413238 123904 413244
rect 123864 412865 123892 413238
rect 123850 412856 123906 412865
rect 123850 412791 123906 412800
rect 123576 411324 123628 411330
rect 123576 411266 123628 411272
rect 123588 410689 123616 411266
rect 123574 410680 123630 410689
rect 123574 410615 123630 410624
rect 123758 403744 123814 403753
rect 123758 403679 123814 403688
rect 123772 403442 123800 403679
rect 123760 403436 123812 403442
rect 123760 403378 123812 403384
rect 123864 393314 123892 412791
rect 124126 408368 124182 408377
rect 124126 408303 124182 408312
rect 124140 407930 124168 408303
rect 124128 407924 124180 407930
rect 124128 407866 124180 407872
rect 124128 406224 124180 406230
rect 124126 406192 124128 406201
rect 124180 406192 124182 406201
rect 124126 406127 124182 406136
rect 124126 401568 124182 401577
rect 124126 401503 124182 401512
rect 124140 400926 124168 401503
rect 124128 400920 124180 400926
rect 124128 400862 124180 400868
rect 124126 399528 124182 399537
rect 124232 399514 124260 452610
rect 124968 451926 124996 465054
rect 125600 454708 125652 454714
rect 125600 454650 125652 454656
rect 124956 451920 125008 451926
rect 124956 451862 125008 451868
rect 124310 447264 124366 447273
rect 124310 447199 124366 447208
rect 124324 431934 124352 447199
rect 124862 444816 124918 444825
rect 124862 444751 124918 444760
rect 124312 431928 124364 431934
rect 124312 431870 124364 431876
rect 124876 409834 124904 444751
rect 125506 443864 125562 443873
rect 125506 443799 125562 443808
rect 125520 443018 125548 443799
rect 125508 443012 125560 443018
rect 125508 442954 125560 442960
rect 124864 409828 124916 409834
rect 124864 409770 124916 409776
rect 125612 406994 125640 454650
rect 126244 438184 126296 438190
rect 126244 438126 126296 438132
rect 125520 406966 125640 406994
rect 125520 406230 125548 406966
rect 125508 406224 125560 406230
rect 125508 406166 125560 406172
rect 124864 403436 124916 403442
rect 124864 403378 124916 403384
rect 124182 399486 124260 399514
rect 124126 399463 124128 399472
rect 124180 399463 124182 399472
rect 124128 399434 124180 399440
rect 124126 397352 124182 397361
rect 124126 397287 124182 397296
rect 124140 395350 124168 397287
rect 124128 395344 124180 395350
rect 124128 395286 124180 395292
rect 123680 393286 123892 393314
rect 123680 387122 123708 393286
rect 123668 387116 123720 387122
rect 123668 387058 123720 387064
rect 123484 382288 123536 382294
rect 123484 382230 123536 382236
rect 123206 349072 123262 349081
rect 123206 349007 123262 349016
rect 122838 348528 122894 348537
rect 122838 348463 122894 348472
rect 122748 346452 122800 346458
rect 122748 346394 122800 346400
rect 123220 345014 123248 349007
rect 121748 344986 121960 345014
rect 123220 344986 123432 345014
rect 121932 329474 121960 344986
rect 123300 332172 123352 332178
rect 123300 332114 123352 332120
rect 123312 329474 123340 332114
rect 120552 329446 120888 329474
rect 121472 329446 121624 329474
rect 121932 329446 122360 329474
rect 123096 329446 123340 329474
rect 123404 329474 123432 344986
rect 123496 344321 123524 382230
rect 124876 370530 124904 403378
rect 125520 373994 125548 406166
rect 126256 374649 126284 438126
rect 126242 374640 126298 374649
rect 126242 374575 126298 374584
rect 125428 373966 125548 373994
rect 124864 370524 124916 370530
rect 124864 370466 124916 370472
rect 125428 368490 125456 373966
rect 125506 368656 125562 368665
rect 125506 368591 125562 368600
rect 125416 368484 125468 368490
rect 125416 368426 125468 368432
rect 125520 368393 125548 368591
rect 125506 368384 125562 368393
rect 125506 368319 125562 368328
rect 126900 368257 126928 546450
rect 126992 415410 127020 568550
rect 128360 541680 128412 541686
rect 128360 541622 128412 541628
rect 128372 541006 128400 541622
rect 129660 541006 129688 700334
rect 130384 700324 130436 700330
rect 130384 700266 130436 700272
rect 128360 541000 128412 541006
rect 128360 540942 128412 540948
rect 129648 541000 129700 541006
rect 129648 540942 129700 540948
rect 127624 462392 127676 462398
rect 127624 462334 127676 462340
rect 127636 447846 127664 462334
rect 127624 447840 127676 447846
rect 127624 447782 127676 447788
rect 127624 444508 127676 444514
rect 127624 444450 127676 444456
rect 126980 415404 127032 415410
rect 126980 415346 127032 415352
rect 125598 368248 125654 368257
rect 125598 368183 125654 368192
rect 126886 368248 126942 368257
rect 126886 368183 126942 368192
rect 124772 367872 124824 367878
rect 124772 367814 124824 367820
rect 124784 367130 124812 367814
rect 124864 367804 124916 367810
rect 124864 367746 124916 367752
rect 124220 367124 124272 367130
rect 124220 367066 124272 367072
rect 124772 367124 124824 367130
rect 124772 367066 124824 367072
rect 124128 350600 124180 350606
rect 124128 350542 124180 350548
rect 124140 349081 124168 350542
rect 124126 349072 124182 349081
rect 124126 349007 124182 349016
rect 124126 347848 124182 347857
rect 124126 347783 124182 347792
rect 123482 344312 123538 344321
rect 123482 344247 123538 344256
rect 124034 343768 124090 343777
rect 124034 343703 124036 343712
rect 124088 343703 124090 343712
rect 124036 343674 124088 343680
rect 124140 332178 124168 347783
rect 124232 334014 124260 367066
rect 124876 350577 124904 367746
rect 124862 350568 124918 350577
rect 124862 350503 124918 350512
rect 124220 334008 124272 334014
rect 124220 333950 124272 333956
rect 124128 332172 124180 332178
rect 124128 332114 124180 332120
rect 124876 330041 124904 350503
rect 125048 341012 125100 341018
rect 125048 340954 125100 340960
rect 125060 340202 125088 340954
rect 125048 340196 125100 340202
rect 125048 340138 125100 340144
rect 124956 334008 125008 334014
rect 124956 333950 125008 333956
rect 124862 330032 124918 330041
rect 124862 329967 124918 329976
rect 124876 329474 124904 329967
rect 123404 329446 123832 329474
rect 124568 329446 124904 329474
rect 124968 329474 124996 333950
rect 125612 332178 125640 368183
rect 126900 367169 126928 368183
rect 126886 367160 126942 367169
rect 126886 367095 126942 367104
rect 127636 367033 127664 444450
rect 128372 387802 128400 540942
rect 129648 539708 129700 539714
rect 129648 539650 129700 539656
rect 129660 536790 129688 539650
rect 130396 538218 130424 700266
rect 170416 596834 170444 702406
rect 170404 596828 170456 596834
rect 170404 596770 170456 596776
rect 187606 589384 187662 589393
rect 187606 589319 187608 589328
rect 187660 589319 187662 589328
rect 187608 589290 187660 589296
rect 132500 584452 132552 584458
rect 132500 584394 132552 584400
rect 130384 538212 130436 538218
rect 130384 538154 130436 538160
rect 129648 536784 129700 536790
rect 129648 536726 129700 536732
rect 130476 535560 130528 535566
rect 130476 535502 130528 535508
rect 129740 529236 129792 529242
rect 129740 529178 129792 529184
rect 129752 528630 129780 529178
rect 129740 528624 129792 528630
rect 129740 528566 129792 528572
rect 128452 478168 128504 478174
rect 128452 478110 128504 478116
rect 128464 477562 128492 478110
rect 128452 477556 128504 477562
rect 128452 477498 128504 477504
rect 128464 450566 128492 477498
rect 128452 450560 128504 450566
rect 128452 450502 128504 450508
rect 129002 448624 129058 448633
rect 129002 448559 129058 448568
rect 128360 387796 128412 387802
rect 128360 387738 128412 387744
rect 127716 368484 127768 368490
rect 127716 368426 127768 368432
rect 126978 367024 127034 367033
rect 126978 366959 127034 366968
rect 127622 367024 127678 367033
rect 127622 366959 127678 366968
rect 126992 366353 127020 366959
rect 126978 366344 127034 366353
rect 126978 366279 127034 366288
rect 125692 349852 125744 349858
rect 125692 349794 125744 349800
rect 125600 332172 125652 332178
rect 125600 332114 125652 332120
rect 125704 329474 125732 349794
rect 126992 335354 127020 366279
rect 127728 351937 127756 368426
rect 127070 351928 127126 351937
rect 127070 351863 127126 351872
rect 127714 351928 127770 351937
rect 127714 351863 127770 351872
rect 127084 345014 127112 351863
rect 129016 345137 129044 448559
rect 129752 353297 129780 528566
rect 130384 492720 130436 492726
rect 130384 492662 130436 492668
rect 130396 366450 130424 492662
rect 130488 447098 130516 535502
rect 131764 458244 131816 458250
rect 131764 458186 131816 458192
rect 131776 449886 131804 458186
rect 131764 449880 131816 449886
rect 131764 449822 131816 449828
rect 130476 447092 130528 447098
rect 130476 447034 130528 447040
rect 131764 442060 131816 442066
rect 131764 442002 131816 442008
rect 131776 407833 131804 442002
rect 132512 438258 132540 584394
rect 142804 581052 142856 581058
rect 142804 580994 142856 581000
rect 133880 567316 133932 567322
rect 133880 567258 133932 567264
rect 133142 541104 133198 541113
rect 133142 541039 133198 541048
rect 133156 536761 133184 541039
rect 133142 536752 133198 536761
rect 133142 536687 133198 536696
rect 132592 447160 132644 447166
rect 132592 447102 132644 447108
rect 132500 438252 132552 438258
rect 132500 438194 132552 438200
rect 131762 407824 131818 407833
rect 131762 407759 131818 407768
rect 130476 397520 130528 397526
rect 130476 397462 130528 397468
rect 130488 389162 130516 397462
rect 130476 389156 130528 389162
rect 130476 389098 130528 389104
rect 130384 366444 130436 366450
rect 130384 366386 130436 366392
rect 130384 363656 130436 363662
rect 130384 363598 130436 363604
rect 129832 356788 129884 356794
rect 129832 356730 129884 356736
rect 129738 353288 129794 353297
rect 129738 353223 129794 353232
rect 129752 352073 129780 353223
rect 129738 352064 129794 352073
rect 129738 351999 129794 352008
rect 129096 347812 129148 347818
rect 129096 347754 129148 347760
rect 129002 345128 129058 345137
rect 129002 345063 129058 345072
rect 127084 344986 127848 345014
rect 126992 335326 127112 335354
rect 126428 332172 126480 332178
rect 126428 332114 126480 332120
rect 126440 329474 126468 332114
rect 127084 329474 127112 335326
rect 127820 329474 127848 344986
rect 129016 342990 129044 345063
rect 129004 342984 129056 342990
rect 129004 342926 129056 342932
rect 129108 337414 129136 347754
rect 129844 345014 129872 356730
rect 130396 347886 130424 363598
rect 132604 356046 132632 447102
rect 133144 438252 133196 438258
rect 133144 438194 133196 438200
rect 133156 396778 133184 438194
rect 133892 407930 133920 567258
rect 137100 566500 137152 566506
rect 137100 566442 137152 566448
rect 137112 565894 137140 566442
rect 136640 565888 136692 565894
rect 136640 565830 136692 565836
rect 137100 565888 137152 565894
rect 137100 565830 137152 565836
rect 134708 563100 134760 563106
rect 134708 563042 134760 563048
rect 134720 559609 134748 563042
rect 134706 559600 134762 559609
rect 134706 559535 134762 559544
rect 136652 413302 136680 565830
rect 137926 545184 137982 545193
rect 137926 545119 137982 545128
rect 136640 413296 136692 413302
rect 136640 413238 136692 413244
rect 133880 407924 133932 407930
rect 133880 407866 133932 407872
rect 134616 407924 134668 407930
rect 134616 407866 134668 407872
rect 133236 405748 133288 405754
rect 133236 405690 133288 405696
rect 133144 396772 133196 396778
rect 133144 396714 133196 396720
rect 133248 373318 133276 405690
rect 134524 393372 134576 393378
rect 134524 393314 134576 393320
rect 133236 373312 133288 373318
rect 133236 373254 133288 373260
rect 133786 361720 133842 361729
rect 133786 361655 133842 361664
rect 132592 356040 132644 356046
rect 132592 355982 132644 355988
rect 132604 355366 132632 355982
rect 132592 355360 132644 355366
rect 132592 355302 132644 355308
rect 133694 354784 133750 354793
rect 133694 354719 133750 354728
rect 130474 352064 130530 352073
rect 130474 351999 130530 352008
rect 130384 347880 130436 347886
rect 130384 347822 130436 347828
rect 129844 344986 130056 345014
rect 129096 337408 129148 337414
rect 129096 337350 129148 337356
rect 129280 334688 129332 334694
rect 129280 334630 129332 334636
rect 129292 329474 129320 334630
rect 129924 332172 129976 332178
rect 129924 332114 129976 332120
rect 129936 329474 129964 332114
rect 124968 329446 125304 329474
rect 125704 329446 126040 329474
rect 126440 329446 126776 329474
rect 127084 329446 127512 329474
rect 127820 329446 128248 329474
rect 128984 329446 129320 329474
rect 129720 329446 129964 329474
rect 130028 329474 130056 344986
rect 130396 332178 130424 347822
rect 130488 342417 130516 351999
rect 130474 342408 130530 342417
rect 130474 342343 130530 342352
rect 131210 342408 131266 342417
rect 131210 342343 131266 342352
rect 131118 338328 131174 338337
rect 131118 338263 131174 338272
rect 131132 338230 131160 338263
rect 131120 338224 131172 338230
rect 131120 338166 131172 338172
rect 131224 335354 131252 342343
rect 131762 338464 131818 338473
rect 131762 338399 131818 338408
rect 131132 335326 131252 335354
rect 130384 332172 130436 332178
rect 130384 332114 130436 332120
rect 131132 329746 131160 335326
rect 131776 330546 131804 338399
rect 133708 335354 133736 354719
rect 133616 335326 133736 335354
rect 132132 333260 132184 333266
rect 132132 333202 132184 333208
rect 131764 330540 131816 330546
rect 131764 330482 131816 330488
rect 131132 329718 131206 329746
rect 130028 329446 130456 329474
rect 131178 329460 131206 329718
rect 132144 329474 132172 333202
rect 132776 331356 132828 331362
rect 132776 331298 132828 331304
rect 132788 329474 132816 331298
rect 133616 329474 133644 335326
rect 133800 331362 133828 361655
rect 133878 352064 133934 352073
rect 133878 351999 133934 352008
rect 133892 347886 133920 351999
rect 133880 347880 133932 347886
rect 133880 347822 133932 347828
rect 134536 345710 134564 393314
rect 134628 368966 134656 407866
rect 136824 372700 136876 372706
rect 136824 372642 136876 372648
rect 134616 368960 134668 368966
rect 134616 368902 134668 368908
rect 135168 368960 135220 368966
rect 135168 368902 135220 368908
rect 135180 368558 135208 368902
rect 135168 368552 135220 368558
rect 135168 368494 135220 368500
rect 134708 364404 134760 364410
rect 134708 364346 134760 364352
rect 134720 351121 134748 364346
rect 134706 351112 134762 351121
rect 134706 351047 134762 351056
rect 135180 346390 135208 368494
rect 136836 365022 136864 372642
rect 136824 365016 136876 365022
rect 136824 364958 136876 364964
rect 137284 365016 137336 365022
rect 137284 364958 137336 364964
rect 137296 364721 137324 364958
rect 137282 364712 137338 364721
rect 137282 364647 137338 364656
rect 137284 363044 137336 363050
rect 137284 362986 137336 362992
rect 136638 358864 136694 358873
rect 136638 358799 136694 358808
rect 135168 346384 135220 346390
rect 135168 346326 135220 346332
rect 134524 345704 134576 345710
rect 134524 345646 134576 345652
rect 136652 345014 136680 358799
rect 137296 347070 137324 362986
rect 137940 358873 137968 545119
rect 142066 542464 142122 542473
rect 142066 542399 142122 542408
rect 140044 473408 140096 473414
rect 140044 473350 140096 473356
rect 140056 391270 140084 473350
rect 141422 444952 141478 444961
rect 141422 444887 141478 444896
rect 140136 392012 140188 392018
rect 140136 391954 140188 391960
rect 140044 391264 140096 391270
rect 140044 391206 140096 391212
rect 140148 380186 140176 391954
rect 140136 380180 140188 380186
rect 140136 380122 140188 380128
rect 140688 376848 140740 376854
rect 140688 376790 140740 376796
rect 139492 365764 139544 365770
rect 139492 365706 139544 365712
rect 137926 358864 137982 358873
rect 137926 358799 137982 358808
rect 139504 358086 139532 365706
rect 139492 358080 139544 358086
rect 139492 358022 139544 358028
rect 137284 347064 137336 347070
rect 137284 347006 137336 347012
rect 139308 347064 139360 347070
rect 139308 347006 139360 347012
rect 136652 344986 137232 345014
rect 136548 336796 136600 336802
rect 136548 336738 136600 336744
rect 134892 335368 134944 335374
rect 134892 335310 134944 335316
rect 134248 331492 134300 331498
rect 134248 331434 134300 331440
rect 133788 331356 133840 331362
rect 133788 331298 133840 331304
rect 134260 329474 134288 331434
rect 134904 329474 134932 335310
rect 136560 334694 136588 336738
rect 136548 334688 136600 334694
rect 136548 334630 136600 334636
rect 135168 334620 135220 334626
rect 135168 334562 135220 334568
rect 135180 331906 135208 334562
rect 137100 334008 137152 334014
rect 137100 333950 137152 333956
rect 135168 331900 135220 331906
rect 135168 331842 135220 331848
rect 135720 331628 135772 331634
rect 135720 331570 135772 331576
rect 135732 329474 135760 331570
rect 137112 329474 137140 333950
rect 131928 329446 132172 329474
rect 132480 329446 132816 329474
rect 133216 329446 133644 329474
rect 133952 329446 134288 329474
rect 134688 329446 134932 329474
rect 135424 329446 135760 329474
rect 136896 329446 137140 329474
rect 137204 329474 137232 344986
rect 139216 337408 139268 337414
rect 139216 337350 139268 337356
rect 138664 332172 138716 332178
rect 138664 332114 138716 332120
rect 138676 329474 138704 332114
rect 139228 331498 139256 337350
rect 139320 332178 139348 347006
rect 139400 346384 139452 346390
rect 139400 346326 139452 346332
rect 139308 332172 139360 332178
rect 139308 332114 139360 332120
rect 139216 331492 139268 331498
rect 139216 331434 139268 331440
rect 137204 329446 137632 329474
rect 138368 329446 138704 329474
rect 139412 329474 139440 346326
rect 139504 334014 139532 358022
rect 139492 334008 139544 334014
rect 139492 333950 139544 333956
rect 140700 329474 140728 376790
rect 141436 349353 141464 444887
rect 140778 349344 140834 349353
rect 140778 349279 140834 349288
rect 141422 349344 141478 349353
rect 141422 349279 141478 349288
rect 140792 345014 140820 349279
rect 140792 344986 140912 345014
rect 140780 341012 140832 341018
rect 140780 340954 140832 340960
rect 140792 340882 140820 340954
rect 140780 340876 140832 340882
rect 140780 340818 140832 340824
rect 140780 334008 140832 334014
rect 140780 333950 140832 333956
rect 140792 333266 140820 333950
rect 140780 333260 140832 333266
rect 140780 333202 140832 333208
rect 139412 329446 139840 329474
rect 140576 329446 140728 329474
rect 140884 329474 140912 344986
rect 142080 342310 142108 542399
rect 142816 533633 142844 580994
rect 149704 571396 149756 571402
rect 149704 571338 149756 571344
rect 146944 560312 146996 560318
rect 146944 560254 146996 560260
rect 146956 535401 146984 560254
rect 148322 537160 148378 537169
rect 148322 537095 148378 537104
rect 146942 535392 146998 535401
rect 146942 535327 146998 535336
rect 143446 534032 143502 534041
rect 143446 533967 143502 533976
rect 143460 533633 143488 533967
rect 142802 533624 142858 533633
rect 142802 533559 142858 533568
rect 143446 533624 143502 533633
rect 143446 533559 143502 533568
rect 143460 460222 143488 533559
rect 147588 521688 147640 521694
rect 147588 521630 147640 521636
rect 147128 476808 147180 476814
rect 147128 476750 147180 476756
rect 147140 476134 147168 476750
rect 147128 476128 147180 476134
rect 147128 476070 147180 476076
rect 147496 476128 147548 476134
rect 147496 476070 147548 476076
rect 144184 474768 144236 474774
rect 144184 474710 144236 474716
rect 143448 460216 143500 460222
rect 143448 460158 143500 460164
rect 143460 459610 143488 460158
rect 142804 459604 142856 459610
rect 142804 459546 142856 459552
rect 143448 459604 143500 459610
rect 143448 459546 143500 459552
rect 142816 432614 142844 459546
rect 142896 445800 142948 445806
rect 142896 445742 142948 445748
rect 142804 432608 142856 432614
rect 142804 432550 142856 432556
rect 141424 342304 141476 342310
rect 141424 342246 141476 342252
rect 142068 342304 142120 342310
rect 142068 342246 142120 342252
rect 141436 331634 141464 342246
rect 142816 341601 142844 432550
rect 142908 403646 142936 445742
rect 142896 403640 142948 403646
rect 142896 403582 142948 403588
rect 144196 391921 144224 474710
rect 144276 445800 144328 445806
rect 144276 445742 144328 445748
rect 144182 391912 144238 391921
rect 144182 391847 144238 391856
rect 142894 377360 142950 377369
rect 142894 377295 142950 377304
rect 142802 341592 142858 341601
rect 142802 341527 142858 341536
rect 142908 332586 142936 377295
rect 144288 369170 144316 445742
rect 147508 444378 147536 476070
rect 147496 444372 147548 444378
rect 147496 444314 147548 444320
rect 144276 369164 144328 369170
rect 144276 369106 144328 369112
rect 144828 367804 144880 367810
rect 144828 367746 144880 367752
rect 142988 357536 143040 357542
rect 142988 357478 143040 357484
rect 143000 349858 143028 357478
rect 142988 349852 143040 349858
rect 142988 349794 143040 349800
rect 144734 345672 144790 345681
rect 144734 345607 144790 345616
rect 144644 343664 144696 343670
rect 144644 343606 144696 343612
rect 144656 342922 144684 343606
rect 144644 342916 144696 342922
rect 144644 342858 144696 342864
rect 143080 332716 143132 332722
rect 143080 332658 143132 332664
rect 142896 332580 142948 332586
rect 142896 332522 142948 332528
rect 141424 331628 141476 331634
rect 141424 331570 141476 331576
rect 141882 331392 141938 331401
rect 141882 331327 141938 331336
rect 140884 329446 141312 329474
rect 117056 329310 117208 329338
rect 141896 329202 141924 331327
rect 143092 329474 143120 332658
rect 144748 332178 144776 345607
rect 143816 332172 143868 332178
rect 143816 332114 143868 332120
rect 144736 332172 144788 332178
rect 144736 332114 144788 332120
rect 143828 329474 143856 332114
rect 144840 329474 144868 367746
rect 147600 363225 147628 521630
rect 148336 447137 148364 537095
rect 148322 447128 148378 447137
rect 148322 447063 148378 447072
rect 148324 444372 148376 444378
rect 148324 444314 148376 444320
rect 148336 368626 148364 444314
rect 148968 421592 149020 421598
rect 148968 421534 149020 421540
rect 147680 368620 147732 368626
rect 147680 368562 147732 368568
rect 148324 368620 148376 368626
rect 148324 368562 148376 368568
rect 147586 363216 147642 363225
rect 147586 363151 147642 363160
rect 146206 362264 146262 362273
rect 146206 362199 146262 362208
rect 146116 345092 146168 345098
rect 146116 345034 146168 345040
rect 146128 340218 146156 345034
rect 146036 340190 146156 340218
rect 146036 332178 146064 340190
rect 146220 335354 146248 362199
rect 147600 355337 147628 363151
rect 147586 355328 147642 355337
rect 147586 355263 147642 355272
rect 146942 347984 146998 347993
rect 146942 347919 146998 347928
rect 146128 335326 146248 335354
rect 145288 332172 145340 332178
rect 145288 332114 145340 332120
rect 146024 332172 146076 332178
rect 146024 332114 146076 332120
rect 145300 329474 145328 332114
rect 146128 329474 146156 335326
rect 146758 334248 146814 334257
rect 146758 334183 146814 334192
rect 146772 329474 146800 334183
rect 146956 332586 146984 347919
rect 147034 345128 147090 345137
rect 147034 345063 147090 345072
rect 147048 337521 147076 345063
rect 147692 345014 147720 368562
rect 147692 344986 148272 345014
rect 147680 338224 147732 338230
rect 147680 338166 147732 338172
rect 147034 337512 147090 337521
rect 147034 337447 147090 337456
rect 147692 337414 147720 338166
rect 147680 337408 147732 337414
rect 147680 337350 147732 337356
rect 148140 335436 148192 335442
rect 148140 335378 148192 335384
rect 146944 332580 146996 332586
rect 146944 332522 146996 332528
rect 142784 329446 143120 329474
rect 143520 329446 143856 329474
rect 144256 329446 144868 329474
rect 144992 329446 145328 329474
rect 145728 329446 146156 329474
rect 146464 329446 146800 329474
rect 146956 329474 146984 332522
rect 148152 329474 148180 335378
rect 146956 329446 147200 329474
rect 147936 329446 148180 329474
rect 148244 329474 148272 344986
rect 148980 342922 149008 421534
rect 149716 362982 149744 571338
rect 177304 564528 177356 564534
rect 177304 564470 177356 564476
rect 166816 564460 166868 564466
rect 166816 564402 166868 564408
rect 160008 558952 160060 558958
rect 160008 558894 160060 558900
rect 152464 556844 152516 556850
rect 152464 556786 152516 556792
rect 152476 487830 152504 556786
rect 157984 538892 158036 538898
rect 157984 538834 158036 538840
rect 156604 512644 156656 512650
rect 156604 512586 156656 512592
rect 152556 489932 152608 489938
rect 152556 489874 152608 489880
rect 152464 487824 152516 487830
rect 152464 487766 152516 487772
rect 152568 438190 152596 489874
rect 155222 467936 155278 467945
rect 155222 467871 155278 467880
rect 152556 438184 152608 438190
rect 152556 438126 152608 438132
rect 152464 426488 152516 426494
rect 152464 426430 152516 426436
rect 151084 411324 151136 411330
rect 151084 411266 151136 411272
rect 149704 362976 149756 362982
rect 149704 362918 149756 362924
rect 149716 355337 149744 362918
rect 149702 355328 149758 355337
rect 149702 355263 149758 355272
rect 150346 353560 150402 353569
rect 150346 353495 150402 353504
rect 148968 342916 149020 342922
rect 148968 342858 149020 342864
rect 149612 336864 149664 336870
rect 149612 336806 149664 336812
rect 149060 334688 149112 334694
rect 149060 334630 149112 334636
rect 149072 334393 149100 334630
rect 149624 334626 149652 336806
rect 149612 334620 149664 334626
rect 149612 334562 149664 334568
rect 149058 334384 149114 334393
rect 149058 334319 149114 334328
rect 150360 332178 150388 353495
rect 151096 334665 151124 411266
rect 152476 367713 152504 426430
rect 153200 392080 153252 392086
rect 153200 392022 153252 392028
rect 152556 378820 152608 378826
rect 152556 378762 152608 378768
rect 152462 367704 152518 367713
rect 152462 367639 152518 367648
rect 151728 362976 151780 362982
rect 151728 362918 151780 362924
rect 151082 334656 151138 334665
rect 151082 334591 151138 334600
rect 149704 332172 149756 332178
rect 149704 332114 149756 332120
rect 150348 332172 150400 332178
rect 150348 332114 150400 332120
rect 149716 329474 149744 332114
rect 150348 331356 150400 331362
rect 150348 331298 150400 331304
rect 150360 329474 150388 331298
rect 151176 331288 151228 331294
rect 151176 331230 151228 331236
rect 151188 329474 151216 331230
rect 151740 329474 151768 362918
rect 152568 358737 152596 378762
rect 152554 358728 152610 358737
rect 152554 358663 152610 358672
rect 153106 358728 153162 358737
rect 153106 358663 153162 358672
rect 153120 357785 153148 358663
rect 153106 357776 153162 357785
rect 153106 357711 153162 357720
rect 153014 339824 153070 339833
rect 153014 339759 153070 339768
rect 153028 338745 153056 339759
rect 153014 338736 153070 338745
rect 153014 338671 153070 338680
rect 152646 330032 152702 330041
rect 152646 329967 152702 329976
rect 152660 329474 152688 329967
rect 153120 329746 153148 357711
rect 153212 340882 153240 392022
rect 155236 356017 155264 467871
rect 156616 451314 156644 512586
rect 156604 451308 156656 451314
rect 156604 451250 156656 451256
rect 155316 360868 155368 360874
rect 155316 360810 155368 360816
rect 155222 356008 155278 356017
rect 155222 355943 155278 355952
rect 155222 353424 155278 353433
rect 155222 353359 155278 353368
rect 155132 342304 155184 342310
rect 155132 342246 155184 342252
rect 155144 341465 155172 342246
rect 155236 341562 155264 353359
rect 155328 349654 155356 360810
rect 155316 349648 155368 349654
rect 155316 349590 155368 349596
rect 155868 349648 155920 349654
rect 155868 349590 155920 349596
rect 155880 349178 155908 349590
rect 155868 349172 155920 349178
rect 155868 349114 155920 349120
rect 155774 344040 155830 344049
rect 155774 343975 155830 343984
rect 155788 343602 155816 343975
rect 155776 343596 155828 343602
rect 155776 343538 155828 343544
rect 155224 341556 155276 341562
rect 155224 341498 155276 341504
rect 155130 341456 155186 341465
rect 155130 341391 155186 341400
rect 155498 341048 155554 341057
rect 155498 340983 155554 340992
rect 153200 340876 153252 340882
rect 153200 340818 153252 340824
rect 153844 340876 153896 340882
rect 153844 340818 153896 340824
rect 153856 339425 153884 340818
rect 153842 339416 153898 339425
rect 153842 339351 153898 339360
rect 155512 338065 155540 340983
rect 155498 338056 155554 338065
rect 155498 337991 155554 338000
rect 155774 336832 155830 336841
rect 155774 336767 155830 336776
rect 155788 336054 155816 336767
rect 155776 336048 155828 336054
rect 155776 335990 155828 335996
rect 155132 335436 155184 335442
rect 155132 335378 155184 335384
rect 155144 334830 155172 335378
rect 155880 335354 155908 349114
rect 156616 344554 156644 451250
rect 157996 444553 158024 538834
rect 159362 535800 159418 535809
rect 159362 535735 159418 535744
rect 157982 444544 158038 444553
rect 157982 444479 158038 444488
rect 157996 391270 158024 444479
rect 159376 420918 159404 535735
rect 159456 449948 159508 449954
rect 159456 449890 159508 449896
rect 159364 420912 159416 420918
rect 159364 420854 159416 420860
rect 157984 391264 158036 391270
rect 157984 391206 158036 391212
rect 156786 368656 156842 368665
rect 156786 368591 156842 368600
rect 156694 367160 156750 367169
rect 156694 367095 156750 367104
rect 156604 344548 156656 344554
rect 156604 344490 156656 344496
rect 156604 343664 156656 343670
rect 156604 343606 156656 343612
rect 156616 338842 156644 343606
rect 156708 340202 156736 367095
rect 156696 340196 156748 340202
rect 156696 340138 156748 340144
rect 156604 338836 156656 338842
rect 156604 338778 156656 338784
rect 155696 335326 155908 335354
rect 155132 334824 155184 334830
rect 155132 334766 155184 334772
rect 154854 331936 154910 331945
rect 154854 331871 154910 331880
rect 148244 329446 148672 329474
rect 149408 329446 149744 329474
rect 150144 329446 150388 329474
rect 150880 329446 151216 329474
rect 151616 329446 151768 329474
rect 152352 329446 152688 329474
rect 153074 329718 153148 329746
rect 153074 329460 153102 329718
rect 154868 329474 154896 331871
rect 155696 329474 155724 335326
rect 155868 334688 155920 334694
rect 155866 334656 155868 334665
rect 155920 334656 155922 334665
rect 155866 334591 155922 334600
rect 154560 329446 154896 329474
rect 155296 329446 155724 329474
rect 141896 329174 142048 329202
rect 153824 329186 154160 329202
rect 153824 329180 154172 329186
rect 153824 329174 154120 329180
rect 154120 329122 154172 329128
rect 114560 329112 114612 329118
rect 136456 329112 136508 329118
rect 114560 329054 114612 329060
rect 136160 329060 136456 329066
rect 139308 329112 139360 329118
rect 136160 329054 136508 329060
rect 139104 329060 139308 329066
rect 156328 329112 156380 329118
rect 139104 329054 139360 329060
rect 156032 329060 156328 329066
rect 156800 329089 156828 368591
rect 157432 366376 157484 366382
rect 157432 366318 157484 366324
rect 159364 366376 159416 366382
rect 159364 366318 159416 366324
rect 157340 345772 157392 345778
rect 157340 345714 157392 345720
rect 156880 338224 156932 338230
rect 156880 338166 156932 338172
rect 156032 329054 156380 329060
rect 156786 329080 156842 329089
rect 136160 329038 136496 329054
rect 139104 329038 139348 329054
rect 156032 329038 156368 329054
rect 156786 329015 156842 329024
rect 156584 328902 156828 328930
rect 156696 328840 156748 328846
rect 156696 328782 156748 328788
rect 156708 320890 156736 328782
rect 156800 328506 156828 328902
rect 156788 328500 156840 328506
rect 156788 328442 156840 328448
rect 156696 320884 156748 320890
rect 156696 320826 156748 320832
rect 156892 318102 156920 338166
rect 157248 329180 157300 329186
rect 157248 329122 157300 329128
rect 157260 328545 157288 329122
rect 157246 328536 157302 328545
rect 157246 328471 157302 328480
rect 156880 318096 156932 318102
rect 156880 318038 156932 318044
rect 67822 308544 67878 308553
rect 67822 308479 67878 308488
rect 157352 300393 157380 345714
rect 157444 331401 157472 366318
rect 159376 358057 159404 366318
rect 159362 358048 159418 358057
rect 159362 357983 159418 357992
rect 158720 352572 158772 352578
rect 158720 352514 158772 352520
rect 157984 348424 158036 348430
rect 157984 348366 158036 348372
rect 157430 331392 157486 331401
rect 157430 331327 157486 331336
rect 157996 308446 158024 348366
rect 158076 331356 158128 331362
rect 158076 331298 158128 331304
rect 157984 308440 158036 308446
rect 157984 308382 158036 308388
rect 157338 300384 157394 300393
rect 157338 300319 157394 300328
rect 67730 296576 67786 296585
rect 67730 296511 67786 296520
rect 67744 295390 67772 296511
rect 67732 295384 67784 295390
rect 67732 295326 67784 295332
rect 156786 271144 156842 271153
rect 156786 271079 156842 271088
rect 67822 270736 67878 270745
rect 67822 270671 67878 270680
rect 67730 245712 67786 245721
rect 67730 245647 67786 245656
rect 67638 228984 67694 228993
rect 67638 228919 67694 228928
rect 67744 209778 67772 245647
rect 67836 241466 67864 270671
rect 80978 242040 81034 242049
rect 69584 241998 70104 242026
rect 67928 241590 68816 241618
rect 69032 241590 69368 241618
rect 67824 241460 67876 241466
rect 67824 241402 67876 241408
rect 67928 238746 67956 241590
rect 67916 238740 67968 238746
rect 67916 238682 67968 238688
rect 69032 223582 69060 241590
rect 69584 238754 69612 241998
rect 154670 242040 154726 242049
rect 81034 241998 81388 242026
rect 80978 241975 81034 241984
rect 69754 241904 69810 241913
rect 69754 241839 69756 241848
rect 69808 241839 69810 241848
rect 71044 241868 71096 241874
rect 69756 241810 69808 241816
rect 71044 241810 71096 241816
rect 69662 241768 69718 241777
rect 69662 241703 69718 241712
rect 69124 238726 69612 238754
rect 69124 238513 69152 238726
rect 69110 238504 69166 238513
rect 69110 238439 69166 238448
rect 69020 223576 69072 223582
rect 69020 223518 69072 223524
rect 69676 222154 69704 241703
rect 70412 241590 70840 241618
rect 69756 238060 69808 238066
rect 69756 238002 69808 238008
rect 69664 222148 69716 222154
rect 69664 222090 69716 222096
rect 69768 217977 69796 238002
rect 69754 217968 69810 217977
rect 69754 217903 69810 217912
rect 67732 209772 67784 209778
rect 67732 209714 67784 209720
rect 70412 208350 70440 241590
rect 71056 210458 71084 241810
rect 71576 241590 71728 241618
rect 72312 241590 72648 241618
rect 71700 239465 71728 241590
rect 72620 240038 72648 241590
rect 72712 241590 73048 241618
rect 73784 241590 74120 241618
rect 74520 241590 74580 241618
rect 75256 241590 75868 241618
rect 72608 240032 72660 240038
rect 72608 239974 72660 239980
rect 71686 239456 71742 239465
rect 71686 239391 71742 239400
rect 72712 238754 72740 241590
rect 73068 240032 73120 240038
rect 73068 239974 73120 239980
rect 71792 238726 72740 238754
rect 71792 238649 71820 238726
rect 71778 238640 71834 238649
rect 71778 238575 71834 238584
rect 71792 237425 71820 238575
rect 71778 237416 71834 237425
rect 71778 237351 71834 237360
rect 72422 237416 72478 237425
rect 72422 237351 72478 237360
rect 71044 210452 71096 210458
rect 71044 210394 71096 210400
rect 70400 208344 70452 208350
rect 70400 208286 70452 208292
rect 72436 195265 72464 237351
rect 73080 219366 73108 239974
rect 74092 239426 74120 241590
rect 74080 239420 74132 239426
rect 74080 239362 74132 239368
rect 73804 236700 73856 236706
rect 73804 236642 73856 236648
rect 73068 219360 73120 219366
rect 73068 219302 73120 219308
rect 73816 204270 73844 236642
rect 74552 231130 74580 241590
rect 74540 231124 74592 231130
rect 74540 231066 74592 231072
rect 75840 210905 75868 241590
rect 75932 241590 75992 241618
rect 76116 241590 76728 241618
rect 77312 241590 77464 241618
rect 77588 241590 78200 241618
rect 78936 241590 79272 241618
rect 79672 241590 80008 241618
rect 80408 241590 80744 241618
rect 75932 240106 75960 241590
rect 75920 240100 75972 240106
rect 75920 240042 75972 240048
rect 76116 235958 76144 241590
rect 77312 240145 77340 241590
rect 77298 240136 77354 240145
rect 76564 240100 76616 240106
rect 77298 240071 77354 240080
rect 76564 240042 76616 240048
rect 76104 235952 76156 235958
rect 76104 235894 76156 235900
rect 75826 210896 75882 210905
rect 75826 210831 75882 210840
rect 73804 204264 73856 204270
rect 73804 204206 73856 204212
rect 76576 198694 76604 240042
rect 77588 238754 77616 241590
rect 79244 239970 79272 241590
rect 79232 239964 79284 239970
rect 79232 239906 79284 239912
rect 79876 239964 79928 239970
rect 79876 239906 79928 239912
rect 77312 238726 77616 238754
rect 77312 214577 77340 238726
rect 78494 237280 78550 237289
rect 78494 237215 78550 237224
rect 78508 236706 78536 237215
rect 78496 236700 78548 236706
rect 78496 236642 78548 236648
rect 77298 214568 77354 214577
rect 77298 214503 77354 214512
rect 76564 198688 76616 198694
rect 79888 198665 79916 239906
rect 76564 198630 76616 198636
rect 79874 198656 79930 198665
rect 79874 198591 79930 198600
rect 72422 195256 72478 195265
rect 72422 195191 72478 195200
rect 79980 192545 80008 241590
rect 80716 239601 80744 241590
rect 80702 239592 80758 239601
rect 80702 239527 80758 239536
rect 81360 206281 81388 241998
rect 154726 241998 155264 242026
rect 154670 241975 154726 241984
rect 81880 241590 82216 241618
rect 82616 241590 82676 241618
rect 82188 239970 82216 241590
rect 82176 239964 82228 239970
rect 82176 239906 82228 239912
rect 82648 238814 82676 241590
rect 83338 241505 83366 241604
rect 83476 241590 84088 241618
rect 84824 241590 85160 241618
rect 85560 241590 85896 241618
rect 86296 241590 86816 241618
rect 83324 241496 83380 241505
rect 83324 241431 83380 241440
rect 83476 240122 83504 241590
rect 83554 241496 83610 241505
rect 83554 241431 83610 241440
rect 82832 240094 83504 240122
rect 82728 239964 82780 239970
rect 82728 239906 82780 239912
rect 82636 238808 82688 238814
rect 82636 238750 82688 238756
rect 81346 206272 81402 206281
rect 81346 206207 81402 206216
rect 82740 205630 82768 239906
rect 82832 209681 82860 240094
rect 83568 238754 83596 241431
rect 85132 240009 85160 241590
rect 85118 240000 85174 240009
rect 85118 239935 85174 239944
rect 85868 239902 85896 241590
rect 85856 239896 85908 239902
rect 85856 239838 85908 239844
rect 86222 239456 86278 239465
rect 86222 239391 86278 239400
rect 83476 238726 83596 238754
rect 84844 238808 84896 238814
rect 84844 238750 84896 238756
rect 83476 230489 83504 238726
rect 83462 230480 83518 230489
rect 83462 230415 83518 230424
rect 84856 224942 84884 238750
rect 86236 229090 86264 239391
rect 86224 229084 86276 229090
rect 86224 229026 86276 229032
rect 84844 224936 84896 224942
rect 84844 224878 84896 224884
rect 82818 209672 82874 209681
rect 82818 209607 82874 209616
rect 86788 208321 86816 241590
rect 86972 241590 87032 241618
rect 87156 241590 87768 241618
rect 88352 241590 88504 241618
rect 89240 241590 89668 241618
rect 86868 239896 86920 239902
rect 86868 239838 86920 239844
rect 86774 208312 86830 208321
rect 86774 208247 86830 208256
rect 82728 205624 82780 205630
rect 82728 205566 82780 205572
rect 86880 197305 86908 239838
rect 86972 212498 87000 241590
rect 87156 212537 87184 241590
rect 87602 239592 87658 239601
rect 87602 239527 87658 239536
rect 87142 212528 87198 212537
rect 86960 212492 87012 212498
rect 87142 212463 87198 212472
rect 86960 212434 87012 212440
rect 87616 206825 87644 239527
rect 88352 236706 88380 241590
rect 88340 236700 88392 236706
rect 88340 236642 88392 236648
rect 88352 236026 88380 236642
rect 88340 236020 88392 236026
rect 88340 235962 88392 235968
rect 88984 236020 89036 236026
rect 88984 235962 89036 235968
rect 87602 206816 87658 206825
rect 87602 206751 87658 206760
rect 86866 197296 86922 197305
rect 86866 197231 86922 197240
rect 88996 193905 89024 235962
rect 88982 193896 89038 193905
rect 88982 193831 89038 193840
rect 79966 192536 80022 192545
rect 79966 192471 80022 192480
rect 89640 188358 89668 241590
rect 89732 241590 89976 241618
rect 90712 241590 91048 241618
rect 89732 237289 89760 241590
rect 89718 237280 89774 237289
rect 89718 237215 89774 237224
rect 89732 236065 89760 237215
rect 89718 236056 89774 236065
rect 89718 235991 89774 236000
rect 90362 236056 90418 236065
rect 90362 235991 90418 236000
rect 90376 191214 90404 235991
rect 91020 216481 91048 241590
rect 91112 241590 91448 241618
rect 91572 241590 92184 241618
rect 92920 241590 93256 241618
rect 91006 216472 91062 216481
rect 91006 216407 91062 216416
rect 91112 215966 91140 241590
rect 91572 238754 91600 241590
rect 93228 240106 93256 241590
rect 93320 241590 93472 241618
rect 93872 241590 94208 241618
rect 94424 241590 94944 241618
rect 95680 241590 96016 241618
rect 93216 240100 93268 240106
rect 93216 240042 93268 240048
rect 93320 238754 93348 241590
rect 93768 240100 93820 240106
rect 93768 240042 93820 240048
rect 91204 238726 91600 238754
rect 92492 238726 93348 238754
rect 91204 220794 91232 238726
rect 92492 234598 92520 238726
rect 92480 234592 92532 234598
rect 92480 234534 92532 234540
rect 92492 234190 92520 234534
rect 92480 234184 92532 234190
rect 92480 234126 92532 234132
rect 93124 234184 93176 234190
rect 93124 234126 93176 234132
rect 91192 220788 91244 220794
rect 91192 220730 91244 220736
rect 91100 215960 91152 215966
rect 91100 215902 91152 215908
rect 92388 215960 92440 215966
rect 92388 215902 92440 215908
rect 92400 199345 92428 215902
rect 92386 199336 92442 199345
rect 92386 199271 92442 199280
rect 93136 193225 93164 234126
rect 93780 209545 93808 240042
rect 93872 219337 93900 241590
rect 94424 238754 94452 241590
rect 95988 239290 96016 241590
rect 96080 241590 96416 241618
rect 96632 241590 97152 241618
rect 97552 241590 97888 241618
rect 98012 241590 98624 241618
rect 99360 241590 99696 241618
rect 100096 241590 100616 241618
rect 95976 239284 96028 239290
rect 95976 239226 96028 239232
rect 96080 238754 96108 241590
rect 96528 239284 96580 239290
rect 96528 239226 96580 239232
rect 93964 238726 94452 238754
rect 95252 238726 96108 238754
rect 93964 235929 93992 238726
rect 93950 235920 94006 235929
rect 93950 235855 94006 235864
rect 95146 235920 95202 235929
rect 95146 235855 95202 235864
rect 95160 235249 95188 235855
rect 95146 235240 95202 235249
rect 95146 235175 95202 235184
rect 93858 219328 93914 219337
rect 93858 219263 93914 219272
rect 95146 219328 95202 219337
rect 95146 219263 95202 219272
rect 93766 209536 93822 209545
rect 93766 209471 93822 209480
rect 93122 193216 93178 193225
rect 93122 193151 93178 193160
rect 90364 191208 90416 191214
rect 90364 191150 90416 191156
rect 89628 188352 89680 188358
rect 89628 188294 89680 188300
rect 95160 186289 95188 219263
rect 95252 218006 95280 238726
rect 95240 218000 95292 218006
rect 95240 217942 95292 217948
rect 96540 206961 96568 239226
rect 96632 238241 96660 241590
rect 97552 240106 97580 241590
rect 97908 240780 97960 240786
rect 97908 240722 97960 240728
rect 96712 240100 96764 240106
rect 96712 240042 96764 240048
rect 97540 240100 97592 240106
rect 97540 240042 97592 240048
rect 96618 238232 96674 238241
rect 96618 238167 96674 238176
rect 96724 234530 96752 240042
rect 97920 236706 97948 240722
rect 97908 236700 97960 236706
rect 97908 236642 97960 236648
rect 96712 234524 96764 234530
rect 96712 234466 96764 234472
rect 98012 211177 98040 241590
rect 99668 240106 99696 241590
rect 99656 240100 99708 240106
rect 99656 240042 99708 240048
rect 100588 213926 100616 241590
rect 100772 241590 100832 241618
rect 100956 241590 101568 241618
rect 102304 241590 102640 241618
rect 100668 240100 100720 240106
rect 100668 240042 100720 240048
rect 100576 213920 100628 213926
rect 100576 213862 100628 213868
rect 100680 212401 100708 240042
rect 100772 221474 100800 241590
rect 100956 224641 100984 241590
rect 102612 240106 102640 241590
rect 102796 241590 103040 241618
rect 103776 241590 104112 241618
rect 102600 240100 102652 240106
rect 102600 240042 102652 240048
rect 102796 228857 102824 241590
rect 104084 240106 104112 241590
rect 104176 241590 104512 241618
rect 105248 241590 105584 241618
rect 103336 240100 103388 240106
rect 103336 240042 103388 240048
rect 104072 240100 104124 240106
rect 104072 240042 104124 240048
rect 102782 228848 102838 228857
rect 102782 228783 102838 228792
rect 103348 226302 103376 240042
rect 104176 238754 104204 241590
rect 104808 240100 104860 240106
rect 104808 240042 104860 240048
rect 103532 238726 104204 238754
rect 103426 236736 103482 236745
rect 103532 236722 103560 238726
rect 103482 236694 103560 236722
rect 103426 236671 103482 236680
rect 103336 226296 103388 226302
rect 103336 226238 103388 226244
rect 100942 224632 100998 224641
rect 100942 224567 100998 224576
rect 102046 224632 102102 224641
rect 102046 224567 102102 224576
rect 100760 221468 100812 221474
rect 100760 221410 100812 221416
rect 100666 212392 100722 212401
rect 100666 212327 100722 212336
rect 97998 211168 98054 211177
rect 97998 211103 98054 211112
rect 99286 211168 99342 211177
rect 99286 211103 99342 211112
rect 99300 210769 99328 211103
rect 99286 210760 99342 210769
rect 99286 210695 99342 210704
rect 96526 206952 96582 206961
rect 96526 206887 96582 206896
rect 99300 186969 99328 210695
rect 102060 203561 102088 224567
rect 102046 203552 102102 203561
rect 102046 203487 102102 203496
rect 103440 197334 103468 236671
rect 103428 197328 103480 197334
rect 103428 197270 103480 197276
rect 104820 191049 104848 240042
rect 105556 239290 105584 241590
rect 105648 241590 105984 241618
rect 106292 241590 106720 241618
rect 107456 241590 107608 241618
rect 105544 239284 105596 239290
rect 105544 239226 105596 239232
rect 105648 238754 105676 241590
rect 106188 239284 106240 239290
rect 106188 239226 106240 239232
rect 104912 238726 105676 238754
rect 104912 220726 104940 238726
rect 104900 220720 104952 220726
rect 104900 220662 104952 220668
rect 106200 205562 106228 239226
rect 106188 205556 106240 205562
rect 106188 205498 106240 205504
rect 106292 195974 106320 241590
rect 106280 195968 106332 195974
rect 106280 195910 106332 195916
rect 104806 191040 104862 191049
rect 104806 190975 104862 190984
rect 107580 189689 107608 241590
rect 107672 241590 108192 241618
rect 108928 241590 108988 241618
rect 109664 241590 110092 241618
rect 110400 241590 110736 241618
rect 111136 241590 111472 241618
rect 111872 241590 112208 241618
rect 112608 241590 113128 241618
rect 113344 241590 113680 241618
rect 114080 241590 114508 241618
rect 107672 236745 107700 241590
rect 108960 239494 108988 241590
rect 108948 239488 109000 239494
rect 108948 239430 109000 239436
rect 110064 238754 110092 241590
rect 110708 240106 110736 241590
rect 111444 240786 111472 241590
rect 111432 240780 111484 240786
rect 111432 240722 111484 240728
rect 110696 240100 110748 240106
rect 110696 240042 110748 240048
rect 112180 239698 112208 241590
rect 112168 239692 112220 239698
rect 112168 239634 112220 239640
rect 112996 239692 113048 239698
rect 112996 239634 113048 239640
rect 111064 239420 111116 239426
rect 111064 239362 111116 239368
rect 110064 238726 110368 238754
rect 107658 236736 107714 236745
rect 107658 236671 107714 236680
rect 110340 229022 110368 238726
rect 110328 229016 110380 229022
rect 110328 228958 110380 228964
rect 111076 222057 111104 239362
rect 111062 222048 111118 222057
rect 111062 221983 111118 221992
rect 113008 217705 113036 239634
rect 112994 217696 113050 217705
rect 112994 217631 113050 217640
rect 113100 193866 113128 241590
rect 113652 239601 113680 241590
rect 113638 239592 113694 239601
rect 113638 239527 113694 239536
rect 114480 214674 114508 241590
rect 114664 241590 114816 241618
rect 115216 241590 115552 241618
rect 116288 241590 116624 241618
rect 117024 241590 117268 241618
rect 114560 240168 114612 240174
rect 114560 240110 114612 240116
rect 114572 238377 114600 240110
rect 114558 238368 114614 238377
rect 114558 238303 114614 238312
rect 114664 235929 114692 241590
rect 115216 240174 115244 241590
rect 115204 240168 115256 240174
rect 115204 240110 115256 240116
rect 116596 239562 116624 241590
rect 116584 239556 116636 239562
rect 116584 239498 116636 239504
rect 117136 239556 117188 239562
rect 117136 239498 117188 239504
rect 114650 235920 114706 235929
rect 114650 235855 114706 235864
rect 114468 214668 114520 214674
rect 114468 214610 114520 214616
rect 117148 207641 117176 239498
rect 117134 207632 117190 207641
rect 117134 207567 117190 207576
rect 117240 200870 117268 241590
rect 117424 241590 117760 241618
rect 117976 241590 118312 241618
rect 119048 241590 119384 241618
rect 117320 239964 117372 239970
rect 117320 239906 117372 239912
rect 117332 216646 117360 239906
rect 117424 233073 117452 241590
rect 117976 239970 118004 241590
rect 119356 240038 119384 241590
rect 119448 241590 119784 241618
rect 120520 241590 120856 241618
rect 121256 241590 121408 241618
rect 121992 241590 122328 241618
rect 122728 241590 122788 241618
rect 119344 240032 119396 240038
rect 119344 239974 119396 239980
rect 117964 239964 118016 239970
rect 117964 239906 118016 239912
rect 119448 238754 119476 241590
rect 119988 240032 120040 240038
rect 119988 239974 120040 239980
rect 118712 238726 119476 238754
rect 117410 233064 117466 233073
rect 117410 232999 117466 233008
rect 117320 216640 117372 216646
rect 117320 216582 117372 216588
rect 118712 209409 118740 238726
rect 118698 209400 118754 209409
rect 118698 209335 118754 209344
rect 117228 200864 117280 200870
rect 117228 200806 117280 200812
rect 120000 195294 120028 239974
rect 120828 239562 120856 241590
rect 121380 240825 121408 241590
rect 121366 240816 121422 240825
rect 121366 240751 121422 240760
rect 121642 240272 121698 240281
rect 121642 240207 121698 240216
rect 120816 239556 120868 239562
rect 120816 239498 120868 239504
rect 121368 239556 121420 239562
rect 121368 239498 121420 239504
rect 121380 202881 121408 239498
rect 121656 235958 121684 240207
rect 122300 239465 122328 241590
rect 122286 239456 122342 239465
rect 122286 239391 122342 239400
rect 121644 235952 121696 235958
rect 121644 235894 121696 235900
rect 121366 202872 121422 202881
rect 121366 202807 121422 202816
rect 122760 196625 122788 241590
rect 122852 241590 123464 241618
rect 124200 241590 124260 241618
rect 122852 206922 122880 241590
rect 124232 219434 124260 241590
rect 124324 241590 124936 241618
rect 125672 241590 126008 241618
rect 126408 241590 126928 241618
rect 124220 219428 124272 219434
rect 124220 219370 124272 219376
rect 124324 213246 124352 241590
rect 125980 240038 126008 241590
rect 125968 240032 126020 240038
rect 125968 239974 126020 239980
rect 126796 240032 126848 240038
rect 126796 239974 126848 239980
rect 126244 232552 126296 232558
rect 126244 232494 126296 232500
rect 126256 227662 126284 232494
rect 126808 231810 126836 239974
rect 126796 231804 126848 231810
rect 126796 231746 126848 231752
rect 126244 227656 126296 227662
rect 126244 227598 126296 227604
rect 124312 213240 124364 213246
rect 124312 213182 124364 213188
rect 122840 206916 122892 206922
rect 122840 206858 122892 206864
rect 126900 198626 126928 241590
rect 127084 241590 127144 241618
rect 127544 241590 127880 241618
rect 128616 241590 128768 241618
rect 126980 240168 127032 240174
rect 126980 240110 127032 240116
rect 126992 224874 127020 240110
rect 127084 233238 127112 241590
rect 127544 240174 127572 241590
rect 127532 240168 127584 240174
rect 127532 240110 127584 240116
rect 128740 239290 128768 241590
rect 128832 241590 129352 241618
rect 130088 241590 130424 241618
rect 128728 239284 128780 239290
rect 128728 239226 128780 239232
rect 128832 238754 128860 241590
rect 129832 239964 129884 239970
rect 129832 239906 129884 239912
rect 129556 239488 129608 239494
rect 129556 239430 129608 239436
rect 128372 238726 128860 238754
rect 127072 233232 127124 233238
rect 127072 233174 127124 233180
rect 126980 224868 127032 224874
rect 126980 224810 127032 224816
rect 128372 211041 128400 238726
rect 129568 238678 129596 239430
rect 129648 239284 129700 239290
rect 129648 239226 129700 239232
rect 129556 238672 129608 238678
rect 129556 238614 129608 238620
rect 129004 232620 129056 232626
rect 129004 232562 129056 232568
rect 128358 211032 128414 211041
rect 128358 210967 128414 210976
rect 129016 200054 129044 232562
rect 129660 202745 129688 239226
rect 129844 232937 129872 239906
rect 130396 239834 130424 241590
rect 130488 241590 130824 241618
rect 131560 241590 131896 241618
rect 132296 241590 132356 241618
rect 133032 241590 133368 241618
rect 130488 239970 130516 241590
rect 131868 240038 131896 241590
rect 131856 240032 131908 240038
rect 131856 239974 131908 239980
rect 130476 239964 130528 239970
rect 130476 239906 130528 239912
rect 130384 239828 130436 239834
rect 130384 239770 130436 239776
rect 131028 239828 131080 239834
rect 131028 239770 131080 239776
rect 129830 232928 129886 232937
rect 129830 232863 129886 232872
rect 131040 205601 131068 239770
rect 132328 217938 132356 241590
rect 133340 240038 133368 241590
rect 133432 241590 133768 241618
rect 134504 241590 135116 241618
rect 135240 241590 135576 241618
rect 135976 241590 136588 241618
rect 132408 240032 132460 240038
rect 132408 239974 132460 239980
rect 133328 240032 133380 240038
rect 133328 239974 133380 239980
rect 132316 217932 132368 217938
rect 132316 217874 132368 217880
rect 132420 209710 132448 239974
rect 133432 239970 133460 241590
rect 133788 240032 133840 240038
rect 133788 239974 133840 239980
rect 132592 239964 132644 239970
rect 132592 239906 132644 239912
rect 133420 239964 133472 239970
rect 133420 239906 133472 239912
rect 132604 233889 132632 239906
rect 132590 233880 132646 233889
rect 132590 233815 132646 233824
rect 132408 209704 132460 209710
rect 132408 209646 132460 209652
rect 133800 206990 133828 239974
rect 135088 238754 135116 241590
rect 135548 239290 135576 241590
rect 136364 240780 136416 240786
rect 136364 240722 136416 240728
rect 135536 239284 135588 239290
rect 135536 239226 135588 239232
rect 135088 238726 135208 238754
rect 135180 228721 135208 238726
rect 136376 235890 136404 240722
rect 136456 239284 136508 239290
rect 136456 239226 136508 239232
rect 136364 235884 136416 235890
rect 136364 235826 136416 235832
rect 135166 228712 135222 228721
rect 135166 228647 135222 228656
rect 136468 215257 136496 239226
rect 136454 215248 136510 215257
rect 136454 215183 136510 215192
rect 133788 206984 133840 206990
rect 133788 206926 133840 206932
rect 131026 205592 131082 205601
rect 131026 205527 131082 205536
rect 129646 202736 129702 202745
rect 129646 202671 129702 202680
rect 136560 201249 136588 241590
rect 136652 241590 136712 241618
rect 136836 241590 137448 241618
rect 138124 241590 138184 241618
rect 138584 241590 138920 241618
rect 139412 241590 139656 241618
rect 140392 241590 140728 241618
rect 141128 241590 141464 241618
rect 141864 241590 142108 241618
rect 136546 201240 136602 201249
rect 136546 201175 136602 201184
rect 129004 200048 129056 200054
rect 129004 199990 129056 199996
rect 126888 198620 126940 198626
rect 126888 198562 126940 198568
rect 122746 196616 122802 196625
rect 122746 196551 122802 196560
rect 119988 195288 120040 195294
rect 119988 195230 120040 195236
rect 113088 193860 113140 193866
rect 113088 193802 113140 193808
rect 115204 191888 115256 191894
rect 115204 191830 115256 191836
rect 107566 189680 107622 189689
rect 107566 189615 107622 189624
rect 99286 186960 99342 186969
rect 99286 186895 99342 186904
rect 113088 186448 113140 186454
rect 113088 186390 113140 186396
rect 95146 186280 95202 186289
rect 95146 186215 95202 186224
rect 103426 183696 103482 183705
rect 103426 183631 103482 183640
rect 99470 182200 99526 182209
rect 99470 182135 99526 182144
rect 98458 180976 98514 180985
rect 98458 180911 98514 180920
rect 97354 179480 97410 179489
rect 97354 179415 97410 179424
rect 97368 176905 97396 179415
rect 98472 177585 98500 180911
rect 98458 177576 98514 177585
rect 98458 177511 98514 177520
rect 97354 176896 97410 176905
rect 97354 176831 97410 176840
rect 99484 176769 99512 182135
rect 100758 180840 100814 180849
rect 100758 180775 100814 180784
rect 100772 177585 100800 180775
rect 100758 177576 100814 177585
rect 100758 177511 100814 177520
rect 103440 176769 103468 183631
rect 107568 183592 107620 183598
rect 107568 183534 107620 183540
rect 105912 180940 105964 180946
rect 105912 180882 105964 180888
rect 105924 177585 105952 180882
rect 107580 177585 107608 183534
rect 105910 177576 105966 177585
rect 105910 177511 105966 177520
rect 107566 177576 107622 177585
rect 107566 177511 107622 177520
rect 113100 177177 113128 186390
rect 114374 179616 114430 179625
rect 114374 179551 114430 179560
rect 114192 177608 114244 177614
rect 114190 177576 114192 177585
rect 114244 177576 114246 177585
rect 114190 177511 114246 177520
rect 114388 177177 114416 179551
rect 115216 177614 115244 191830
rect 136652 190466 136680 241590
rect 136836 229094 136864 241590
rect 138020 240168 138072 240174
rect 138020 240110 138072 240116
rect 138032 237386 138060 240110
rect 138124 237386 138152 241590
rect 138584 240174 138612 241590
rect 138572 240168 138624 240174
rect 138572 240110 138624 240116
rect 138020 237380 138072 237386
rect 138020 237322 138072 237328
rect 138112 237380 138164 237386
rect 138112 237322 138164 237328
rect 138032 237289 138060 237322
rect 138018 237280 138074 237289
rect 138018 237215 138074 237224
rect 138388 231124 138440 231130
rect 138388 231066 138440 231072
rect 136836 229066 137324 229094
rect 137296 226137 137324 229066
rect 137282 226128 137338 226137
rect 137282 226063 137338 226072
rect 137296 202842 137324 226063
rect 138400 223514 138428 231066
rect 138388 223508 138440 223514
rect 138388 223450 138440 223456
rect 139412 222193 139440 241590
rect 140700 231742 140728 241590
rect 141436 239426 141464 241590
rect 141424 239420 141476 239426
rect 141424 239362 141476 239368
rect 141976 239420 142028 239426
rect 141976 239362 142028 239368
rect 140688 231736 140740 231742
rect 140688 231678 140740 231684
rect 139398 222184 139454 222193
rect 139398 222119 139454 222128
rect 137284 202836 137336 202842
rect 137284 202778 137336 202784
rect 141988 202162 142016 239362
rect 141976 202156 142028 202162
rect 141976 202098 142028 202104
rect 136640 190460 136692 190466
rect 136640 190402 136692 190408
rect 125508 189100 125560 189106
rect 125508 189042 125560 189048
rect 118608 184952 118660 184958
rect 118608 184894 118660 184900
rect 115846 182336 115902 182345
rect 115846 182271 115902 182280
rect 115204 177608 115256 177614
rect 115860 177585 115888 182271
rect 118620 177585 118648 184894
rect 121920 182232 121972 182238
rect 121920 182174 121972 182180
rect 119896 179512 119948 179518
rect 119896 179454 119948 179460
rect 115204 177550 115256 177556
rect 115846 177576 115902 177585
rect 115846 177511 115902 177520
rect 118606 177576 118662 177585
rect 118606 177511 118662 177520
rect 119908 177177 119936 179454
rect 121932 177585 121960 182174
rect 123300 178152 123352 178158
rect 123300 178094 123352 178100
rect 121918 177576 121974 177585
rect 121918 177511 121974 177520
rect 113086 177168 113142 177177
rect 113086 177103 113142 177112
rect 114374 177168 114430 177177
rect 114374 177103 114430 177112
rect 119894 177168 119950 177177
rect 119894 177103 119950 177112
rect 123312 176769 123340 178094
rect 125520 177585 125548 189042
rect 133144 187740 133196 187746
rect 133144 187682 133196 187688
rect 129004 183660 129056 183666
rect 129004 183602 129056 183608
rect 126796 179444 126848 179450
rect 126796 179386 126848 179392
rect 125506 177576 125562 177585
rect 125506 177511 125562 177520
rect 126808 176769 126836 179386
rect 129016 177614 129044 183602
rect 132408 180872 132460 180878
rect 132408 180814 132460 180820
rect 129464 178016 129516 178022
rect 129464 177958 129516 177964
rect 127992 177608 128044 177614
rect 127990 177576 127992 177585
rect 129004 177608 129056 177614
rect 128044 177576 128046 177585
rect 129004 177550 129056 177556
rect 127990 177511 128046 177520
rect 129476 176769 129504 177958
rect 132420 177585 132448 180814
rect 133156 178022 133184 187682
rect 133788 186380 133840 186386
rect 133788 186322 133840 186328
rect 133144 178016 133196 178022
rect 133144 177958 133196 177964
rect 133800 177585 133828 186322
rect 142080 185609 142108 241590
rect 142172 241590 142600 241618
rect 143152 241590 143488 241618
rect 143888 241590 144224 241618
rect 142172 230450 142200 241590
rect 142986 237280 143042 237289
rect 142986 237215 143042 237224
rect 142802 236600 142858 236609
rect 142802 236535 142858 236544
rect 142160 230444 142212 230450
rect 142160 230386 142212 230392
rect 142816 226234 142844 236535
rect 143000 235793 143028 237215
rect 142986 235784 143042 235793
rect 142986 235719 143042 235728
rect 143354 235240 143410 235249
rect 143354 235175 143410 235184
rect 143368 233170 143396 235175
rect 143356 233164 143408 233170
rect 143356 233106 143408 233112
rect 142804 226228 142856 226234
rect 142804 226170 142856 226176
rect 143460 220697 143488 241590
rect 144196 239426 144224 241590
rect 144288 241590 144624 241618
rect 144932 241590 145360 241618
rect 145760 241590 146096 241618
rect 144184 239420 144236 239426
rect 144184 239362 144236 239368
rect 144288 239290 144316 241590
rect 144828 239420 144880 239426
rect 144828 239362 144880 239368
rect 143540 239284 143592 239290
rect 143540 239226 143592 239232
rect 144276 239284 144328 239290
rect 144276 239226 144328 239232
rect 143552 237153 143580 239226
rect 143538 237144 143594 237153
rect 143538 237079 143594 237088
rect 143446 220688 143502 220697
rect 143446 220623 143502 220632
rect 144840 211818 144868 239362
rect 144932 227497 144960 241590
rect 145760 239426 145788 241590
rect 146818 241369 146846 241604
rect 147568 241590 147628 241618
rect 146804 241360 146860 241369
rect 146804 241295 146860 241304
rect 147218 240272 147274 240281
rect 147218 240207 147274 240216
rect 145012 239420 145064 239426
rect 145012 239362 145064 239368
rect 145748 239420 145800 239426
rect 145748 239362 145800 239368
rect 145024 234598 145052 239362
rect 146850 236736 146906 236745
rect 146850 236671 146906 236680
rect 146208 235272 146260 235278
rect 146208 235214 146260 235220
rect 145012 234592 145064 234598
rect 145012 234534 145064 234540
rect 146220 234433 146248 235214
rect 146206 234424 146262 234433
rect 146206 234359 146262 234368
rect 146864 231849 146892 236671
rect 147232 235958 147260 240207
rect 147220 235952 147272 235958
rect 147220 235894 147272 235900
rect 146850 231840 146906 231849
rect 146850 231775 146906 231784
rect 147496 229764 147548 229770
rect 147496 229706 147548 229712
rect 144918 227488 144974 227497
rect 144918 227423 144974 227432
rect 146942 226944 146998 226953
rect 146942 226879 146998 226888
rect 146956 216345 146984 226879
rect 147508 223553 147536 229706
rect 147494 223544 147550 223553
rect 147494 223479 147550 223488
rect 146942 216336 146998 216345
rect 146942 216271 146998 216280
rect 144828 211812 144880 211818
rect 144828 211754 144880 211760
rect 146942 207088 146998 207097
rect 146942 207023 146998 207032
rect 146956 206825 146984 207023
rect 146942 206816 146998 206825
rect 146942 206751 146998 206760
rect 147600 202842 147628 241590
rect 147692 241590 148304 241618
rect 149040 241590 149376 241618
rect 149776 241590 150388 241618
rect 150512 241590 150848 241618
rect 151248 241590 151768 241618
rect 151984 241590 152044 241618
rect 147692 237017 147720 241590
rect 149348 240038 149376 241590
rect 149336 240032 149388 240038
rect 149336 239974 149388 239980
rect 150256 240032 150308 240038
rect 150256 239974 150308 239980
rect 147678 237008 147734 237017
rect 147678 236943 147734 236952
rect 150268 230382 150296 239974
rect 150256 230376 150308 230382
rect 150256 230318 150308 230324
rect 150360 219065 150388 241590
rect 150820 239970 150848 241590
rect 150808 239964 150860 239970
rect 150808 239906 150860 239912
rect 150438 235240 150494 235249
rect 150438 235175 150494 235184
rect 150452 234530 150480 235175
rect 150440 234524 150492 234530
rect 150440 234466 150492 234472
rect 150346 219056 150402 219065
rect 150346 218991 150402 219000
rect 151740 204105 151768 241590
rect 151910 240816 151966 240825
rect 151910 240751 151966 240760
rect 151924 238610 151952 240751
rect 152016 240038 152044 241590
rect 152108 241590 152720 241618
rect 153456 241590 153792 241618
rect 152004 240032 152056 240038
rect 152004 239974 152056 239980
rect 151912 238604 151964 238610
rect 151912 238546 151964 238552
rect 152108 237289 152136 241590
rect 153764 239290 153792 241590
rect 154178 241505 154206 241604
rect 154164 241496 154220 241505
rect 154164 241431 154220 241440
rect 155130 241224 155186 241233
rect 155130 241159 155186 241168
rect 154488 240780 154540 240786
rect 154488 240722 154540 240728
rect 154500 239970 154528 240722
rect 154488 239964 154540 239970
rect 154488 239906 154540 239912
rect 153752 239284 153804 239290
rect 153752 239226 153804 239232
rect 154488 239284 154540 239290
rect 154488 239226 154540 239232
rect 152094 237280 152150 237289
rect 152094 237215 152150 237224
rect 151726 204096 151782 204105
rect 151726 204031 151782 204040
rect 147588 202836 147640 202842
rect 147588 202778 147640 202784
rect 142066 185600 142122 185609
rect 142066 185535 142122 185544
rect 154500 184249 154528 239226
rect 155144 238754 155172 241159
rect 155236 240145 155264 241998
rect 156694 241632 156750 241641
rect 155664 241590 155908 241618
rect 156400 241590 156694 241618
rect 155316 241528 155368 241534
rect 155316 241470 155368 241476
rect 155222 240136 155278 240145
rect 155222 240071 155278 240080
rect 155144 238726 155264 238754
rect 155236 223514 155264 238726
rect 155328 235890 155356 241470
rect 155774 240136 155830 240145
rect 155774 240071 155830 240080
rect 155316 235884 155368 235890
rect 155316 235826 155368 235832
rect 155788 223514 155816 240071
rect 155224 223508 155276 223514
rect 155224 223450 155276 223456
rect 155776 223508 155828 223514
rect 155776 223450 155828 223456
rect 155880 200705 155908 241590
rect 156694 241567 156750 241576
rect 156800 229022 156828 271079
rect 157996 264761 158024 308382
rect 158088 291854 158116 331298
rect 158168 328636 158220 328642
rect 158168 328578 158220 328584
rect 158180 325009 158208 328578
rect 158166 325000 158222 325009
rect 158166 324935 158222 324944
rect 158732 324426 158760 352514
rect 158904 349920 158956 349926
rect 158904 349862 158956 349868
rect 158916 345014 158944 349862
rect 158916 344986 159036 345014
rect 158810 343632 158866 343641
rect 158810 343567 158866 343576
rect 158824 342310 158852 343567
rect 158904 342916 158956 342922
rect 158904 342858 158956 342864
rect 158812 342304 158864 342310
rect 158812 342246 158864 342252
rect 158916 335354 158944 342858
rect 158824 335326 158944 335354
rect 158720 324420 158772 324426
rect 158720 324362 158772 324368
rect 158720 324284 158772 324290
rect 158720 324226 158772 324232
rect 158732 323241 158760 324226
rect 158718 323232 158774 323241
rect 158718 323167 158774 323176
rect 158720 322312 158772 322318
rect 158720 322254 158772 322260
rect 158732 322153 158760 322254
rect 158718 322144 158774 322153
rect 158718 322079 158774 322088
rect 158718 317792 158774 317801
rect 158718 317727 158774 317736
rect 158732 317626 158760 317727
rect 158720 317620 158772 317626
rect 158720 317562 158772 317568
rect 158720 317416 158772 317422
rect 158720 317358 158772 317364
rect 158732 316713 158760 317358
rect 158718 316704 158774 316713
rect 158718 316639 158774 316648
rect 158718 313440 158774 313449
rect 158718 313375 158720 313384
rect 158772 313375 158774 313384
rect 158720 313346 158772 313352
rect 158718 311264 158774 311273
rect 158718 311199 158774 311208
rect 158732 310554 158760 311199
rect 158720 310548 158772 310554
rect 158720 310490 158772 310496
rect 158824 310185 158852 335326
rect 158902 328672 158958 328681
rect 158902 328607 158958 328616
rect 158916 328574 158944 328607
rect 158904 328568 158956 328574
rect 158904 328510 158956 328516
rect 159008 328386 159036 344986
rect 159468 342961 159496 449890
rect 160020 356794 160048 558894
rect 161388 549364 161440 549370
rect 161388 549306 161440 549312
rect 160008 356788 160060 356794
rect 160008 356730 160060 356736
rect 160834 356008 160890 356017
rect 160834 355943 160890 355952
rect 159454 342952 159510 342961
rect 159454 342887 159510 342896
rect 160744 334824 160796 334830
rect 160744 334766 160796 334772
rect 158916 328358 159036 328386
rect 158916 327593 158944 328358
rect 158902 327584 158958 327593
rect 158902 327519 158958 327528
rect 158916 324442 158944 327519
rect 158994 326496 159050 326505
rect 158994 326431 159050 326440
rect 159008 325718 159036 326431
rect 158996 325712 159048 325718
rect 158996 325654 159048 325660
rect 159088 325644 159140 325650
rect 159088 325586 159140 325592
rect 159100 325417 159128 325586
rect 159086 325408 159142 325417
rect 159086 325343 159142 325352
rect 158916 324414 159036 324442
rect 158902 324320 158958 324329
rect 158902 324255 158958 324264
rect 158916 322998 158944 324255
rect 158904 322992 158956 322998
rect 158904 322934 158956 322940
rect 159008 322386 159036 324414
rect 159088 324420 159140 324426
rect 159088 324362 159140 324368
rect 158996 322380 159048 322386
rect 158996 322322 159048 322328
rect 159100 317422 159128 324362
rect 159272 319524 159324 319530
rect 159272 319466 159324 319472
rect 159916 319524 159968 319530
rect 159916 319466 159968 319472
rect 159284 318889 159312 319466
rect 159362 319424 159418 319433
rect 159362 319359 159418 319368
rect 159270 318880 159326 318889
rect 159270 318815 159326 318824
rect 159088 317416 159140 317422
rect 159088 317358 159140 317364
rect 159376 316034 159404 319359
rect 159284 316006 159404 316034
rect 158810 310176 158866 310185
rect 158810 310111 158866 310120
rect 158824 309806 158852 310111
rect 158812 309800 158864 309806
rect 158812 309742 158864 309748
rect 158720 308508 158772 308514
rect 158720 308450 158772 308456
rect 158732 308009 158760 308450
rect 158718 308000 158774 308009
rect 158718 307935 158774 307944
rect 158718 306912 158774 306921
rect 158718 306847 158774 306856
rect 158732 306406 158760 306847
rect 158720 306400 158772 306406
rect 158720 306342 158772 306348
rect 158718 305824 158774 305833
rect 158718 305759 158774 305768
rect 158732 305114 158760 305759
rect 158720 305108 158772 305114
rect 158720 305050 158772 305056
rect 158812 304972 158864 304978
rect 158812 304914 158864 304920
rect 158718 304736 158774 304745
rect 158718 304671 158774 304680
rect 158732 301510 158760 304671
rect 158824 303657 158852 304914
rect 158810 303648 158866 303657
rect 158810 303583 158866 303592
rect 158720 301504 158772 301510
rect 158720 301446 158772 301452
rect 158810 301472 158866 301481
rect 158810 301407 158866 301416
rect 158824 298761 158852 301407
rect 158810 298752 158866 298761
rect 158810 298687 158866 298696
rect 158720 298104 158772 298110
rect 158720 298046 158772 298052
rect 158628 297424 158680 297430
rect 158628 297366 158680 297372
rect 158076 291848 158128 291854
rect 158076 291790 158128 291796
rect 158442 284880 158498 284889
rect 158442 284815 158498 284824
rect 157982 264752 158038 264761
rect 157982 264687 158038 264696
rect 158076 262948 158128 262954
rect 158076 262890 158128 262896
rect 157984 261520 158036 261526
rect 157984 261462 158036 261468
rect 156972 243568 157024 243574
rect 156972 243510 157024 243516
rect 156880 241596 156932 241602
rect 156880 241538 156932 241544
rect 156788 229016 156840 229022
rect 156788 228958 156840 228964
rect 156604 228404 156656 228410
rect 156604 228346 156656 228352
rect 156616 227730 156644 228346
rect 156604 227724 156656 227730
rect 156604 227666 156656 227672
rect 156604 226636 156656 226642
rect 156604 226578 156656 226584
rect 156616 219366 156644 226578
rect 156892 226234 156920 241538
rect 156984 237386 157012 243510
rect 157338 240816 157394 240825
rect 157338 240751 157394 240760
rect 157352 240038 157380 240751
rect 157340 240032 157392 240038
rect 157340 239974 157392 239980
rect 157996 238610 158024 261462
rect 157984 238604 158036 238610
rect 157984 238546 158036 238552
rect 156972 237380 157024 237386
rect 156972 237322 157024 237328
rect 157340 237176 157392 237182
rect 157340 237118 157392 237124
rect 157352 233170 157380 237118
rect 158088 237017 158116 262890
rect 158456 261497 158484 284815
rect 158536 269816 158588 269822
rect 158536 269758 158588 269764
rect 158442 261488 158498 261497
rect 158442 261423 158498 261432
rect 158166 243536 158222 243545
rect 158166 243471 158222 243480
rect 158074 237008 158130 237017
rect 158074 236943 158130 236952
rect 157432 235272 157484 235278
rect 157432 235214 157484 235220
rect 157340 233164 157392 233170
rect 157340 233106 157392 233112
rect 157444 230382 157472 235214
rect 157432 230376 157484 230382
rect 157432 230318 157484 230324
rect 158180 229090 158208 243471
rect 158548 240786 158576 269758
rect 158640 245857 158668 297366
rect 158732 297129 158760 298046
rect 158718 297120 158774 297129
rect 158718 297055 158774 297064
rect 158718 296032 158774 296041
rect 158718 295967 158774 295976
rect 158732 295390 158760 295967
rect 158720 295384 158772 295390
rect 158720 295326 158772 295332
rect 158718 293856 158774 293865
rect 158718 293791 158774 293800
rect 158732 292670 158760 293791
rect 158720 292664 158772 292670
rect 158720 292606 158772 292612
rect 158718 291952 158774 291961
rect 158718 291887 158774 291896
rect 158732 291242 158760 291887
rect 158720 291236 158772 291242
rect 158720 291178 158772 291184
rect 158718 290864 158774 290873
rect 158718 290799 158774 290808
rect 158732 289882 158760 290799
rect 158720 289876 158772 289882
rect 158720 289818 158772 289824
rect 158810 289776 158866 289785
rect 158810 289711 158866 289720
rect 158824 288454 158852 289711
rect 158812 288448 158864 288454
rect 158812 288390 158864 288396
rect 158718 287600 158774 287609
rect 158718 287535 158774 287544
rect 158732 287162 158760 287535
rect 158720 287156 158772 287162
rect 158720 287098 158772 287104
rect 158720 287020 158772 287026
rect 158720 286962 158772 286968
rect 158732 286521 158760 286962
rect 158718 286512 158774 286521
rect 158718 286447 158774 286456
rect 158720 286340 158772 286346
rect 158720 286282 158772 286288
rect 158732 285433 158760 286282
rect 158718 285424 158774 285433
rect 158718 285359 158774 285368
rect 158718 284336 158774 284345
rect 158718 284271 158774 284280
rect 158812 284300 158864 284306
rect 158732 283626 158760 284271
rect 158812 284242 158864 284248
rect 158720 283620 158772 283626
rect 158720 283562 158772 283568
rect 158824 283257 158852 284242
rect 158810 283248 158866 283257
rect 158810 283183 158866 283192
rect 158720 282872 158772 282878
rect 158720 282814 158772 282820
rect 158732 282169 158760 282814
rect 158718 282160 158774 282169
rect 158718 282095 158774 282104
rect 158810 281072 158866 281081
rect 158810 281007 158866 281016
rect 158720 280152 158772 280158
rect 158720 280094 158772 280100
rect 158732 279993 158760 280094
rect 158718 279984 158774 279993
rect 158718 279919 158774 279928
rect 158718 278896 158774 278905
rect 158718 278831 158774 278840
rect 158732 278798 158760 278831
rect 158720 278792 158772 278798
rect 158720 278734 158772 278740
rect 158824 278050 158852 281007
rect 158812 278044 158864 278050
rect 158812 277986 158864 277992
rect 158720 277364 158772 277370
rect 158720 277306 158772 277312
rect 158732 276729 158760 277306
rect 158718 276720 158774 276729
rect 158718 276655 158774 276664
rect 158810 275632 158866 275641
rect 158810 275567 158866 275576
rect 158824 274718 158852 275567
rect 158812 274712 158864 274718
rect 158812 274654 158864 274660
rect 158720 274644 158772 274650
rect 158720 274586 158772 274592
rect 158732 274553 158760 274586
rect 158718 274544 158774 274553
rect 158718 274479 158774 274488
rect 158718 273456 158774 273465
rect 158718 273391 158774 273400
rect 158732 271182 158760 273391
rect 158720 271176 158772 271182
rect 158720 271118 158772 271124
rect 158718 269104 158774 269113
rect 158718 269039 158774 269048
rect 158732 269006 158760 269039
rect 158720 269000 158772 269006
rect 158720 268942 158772 268948
rect 158718 268016 158774 268025
rect 158718 267951 158720 267960
rect 158772 267951 158774 267960
rect 158720 267922 158772 267928
rect 158718 263664 158774 263673
rect 158718 263599 158720 263608
rect 158772 263599 158774 263608
rect 158720 263570 158772 263576
rect 158720 258732 158772 258738
rect 158720 258674 158772 258680
rect 158732 258233 158760 258674
rect 158718 258224 158774 258233
rect 158718 258159 158774 258168
rect 158810 256320 158866 256329
rect 158810 256255 158866 256264
rect 158824 255338 158852 256255
rect 158812 255332 158864 255338
rect 158812 255274 158864 255280
rect 158720 255264 158772 255270
rect 158718 255232 158720 255241
rect 158772 255232 158774 255241
rect 158718 255167 158774 255176
rect 158718 253056 158774 253065
rect 158718 252991 158774 253000
rect 158732 252618 158760 252991
rect 158720 252612 158772 252618
rect 158720 252554 158772 252560
rect 158810 249792 158866 249801
rect 158810 249727 158866 249736
rect 158718 248704 158774 248713
rect 158718 248639 158774 248648
rect 158732 248470 158760 248639
rect 158824 248538 158852 249727
rect 158812 248532 158864 248538
rect 158812 248474 158864 248480
rect 158720 248464 158772 248470
rect 158720 248406 158772 248412
rect 158626 245848 158682 245857
rect 158626 245783 158682 245792
rect 158812 245676 158864 245682
rect 158812 245618 158864 245624
rect 158718 244352 158774 244361
rect 158718 244287 158720 244296
rect 158772 244287 158774 244296
rect 158720 244258 158772 244264
rect 158718 243264 158774 243273
rect 158718 243199 158774 243208
rect 158732 242962 158760 243199
rect 158720 242956 158772 242962
rect 158720 242898 158772 242904
rect 158824 241233 158852 245618
rect 158810 241224 158866 241233
rect 158810 241159 158866 241168
rect 158536 240780 158588 240786
rect 158536 240722 158588 240728
rect 159284 236065 159312 316006
rect 159928 311137 159956 319466
rect 159914 311128 159970 311137
rect 159914 311063 159970 311072
rect 159454 300384 159510 300393
rect 159454 300319 159510 300328
rect 159362 293040 159418 293049
rect 159362 292975 159418 292984
rect 159376 282305 159404 292975
rect 159468 292505 159496 300319
rect 159640 300144 159692 300150
rect 159640 300086 159692 300092
rect 159652 298790 159680 300086
rect 159640 298784 159692 298790
rect 159640 298726 159692 298732
rect 159652 298217 159680 298726
rect 159638 298208 159694 298217
rect 159638 298143 159694 298152
rect 159454 292496 159510 292505
rect 159454 292431 159510 292440
rect 159362 282296 159418 282305
rect 159362 282231 159418 282240
rect 159362 277808 159418 277817
rect 159362 277743 159418 277752
rect 159376 275330 159404 277743
rect 159364 275324 159416 275330
rect 159364 275266 159416 275272
rect 159362 271280 159418 271289
rect 159362 271215 159418 271224
rect 159376 262886 159404 271215
rect 159454 265840 159510 265849
rect 159454 265775 159510 265784
rect 159364 262880 159416 262886
rect 159364 262822 159416 262828
rect 159362 261488 159418 261497
rect 159362 261423 159418 261432
rect 159270 236056 159326 236065
rect 159270 235991 159326 236000
rect 158626 233880 158682 233889
rect 158626 233815 158682 233824
rect 158168 229084 158220 229090
rect 158168 229026 158220 229032
rect 156880 226228 156932 226234
rect 156880 226170 156932 226176
rect 156604 219360 156656 219366
rect 156604 219302 156656 219308
rect 155866 200696 155922 200705
rect 155866 200631 155922 200640
rect 158640 199481 158668 233815
rect 159376 221921 159404 261423
rect 159468 257378 159496 265775
rect 159914 259584 159970 259593
rect 159914 259519 159970 259528
rect 159456 257372 159508 257378
rect 159456 257314 159508 257320
rect 159546 236056 159602 236065
rect 159546 235991 159602 236000
rect 159362 221912 159418 221921
rect 159362 221847 159418 221856
rect 159376 214606 159404 221847
rect 159560 221513 159588 235991
rect 159546 221504 159602 221513
rect 159546 221439 159602 221448
rect 159364 214600 159416 214606
rect 159364 214542 159416 214548
rect 158626 199472 158682 199481
rect 158626 199407 158682 199416
rect 154486 184240 154542 184249
rect 154486 184175 154542 184184
rect 159928 182889 159956 259519
rect 160100 256760 160152 256766
rect 160100 256702 160152 256708
rect 160006 254144 160062 254153
rect 160112 254130 160140 256702
rect 160062 254102 160140 254130
rect 160006 254079 160062 254088
rect 160756 250510 160784 334766
rect 160848 316713 160876 355943
rect 161296 352572 161348 352578
rect 161296 352514 161348 352520
rect 160926 337512 160982 337521
rect 160926 337447 160982 337456
rect 160940 328409 160968 337447
rect 160926 328400 160982 328409
rect 160926 328335 160982 328344
rect 160834 316704 160890 316713
rect 160834 316639 160890 316648
rect 160834 311944 160890 311953
rect 160834 311879 160836 311888
rect 160888 311879 160890 311888
rect 160836 311850 160888 311856
rect 160836 294636 160888 294642
rect 160836 294578 160888 294584
rect 160848 262585 160876 294578
rect 160834 262576 160890 262585
rect 160834 262511 160890 262520
rect 160836 253224 160888 253230
rect 160836 253166 160888 253172
rect 160744 250504 160796 250510
rect 160744 250446 160796 250452
rect 160742 247208 160798 247217
rect 160742 247143 160798 247152
rect 160756 220697 160784 247143
rect 160848 237289 160876 253166
rect 161202 251152 161258 251161
rect 161202 251087 161258 251096
rect 160834 237280 160890 237289
rect 160834 237215 160890 237224
rect 160742 220688 160798 220697
rect 160742 220623 160798 220632
rect 161216 209817 161244 251087
rect 161308 244905 161336 352514
rect 161400 337385 161428 549306
rect 164148 533384 164200 533390
rect 164148 533326 164200 533332
rect 164160 532778 164188 533326
rect 162860 532772 162912 532778
rect 162860 532714 162912 532720
rect 164148 532772 164200 532778
rect 164148 532714 164200 532720
rect 162124 518968 162176 518974
rect 162124 518910 162176 518916
rect 161386 337376 161442 337385
rect 161386 337311 161442 337320
rect 161388 311840 161440 311846
rect 161388 311782 161440 311788
rect 161400 247217 161428 311782
rect 162136 269385 162164 518910
rect 162768 370524 162820 370530
rect 162768 370466 162820 370472
rect 162214 355328 162270 355337
rect 162214 355263 162270 355272
rect 162228 332042 162256 355263
rect 162308 339516 162360 339522
rect 162308 339458 162360 339464
rect 162216 332036 162268 332042
rect 162216 331978 162268 331984
rect 162216 329860 162268 329866
rect 162216 329802 162268 329808
rect 162228 294710 162256 329802
rect 162320 327078 162348 339458
rect 162308 327072 162360 327078
rect 162308 327014 162360 327020
rect 162216 294704 162268 294710
rect 162216 294646 162268 294652
rect 162674 285696 162730 285705
rect 162674 285631 162730 285640
rect 162122 269376 162178 269385
rect 162122 269311 162178 269320
rect 162124 267980 162176 267986
rect 162124 267922 162176 267928
rect 162136 247518 162164 267922
rect 162216 265668 162268 265674
rect 162216 265610 162268 265616
rect 162124 247512 162176 247518
rect 162124 247454 162176 247460
rect 161386 247208 161442 247217
rect 161386 247143 161442 247152
rect 161294 244896 161350 244905
rect 161294 244831 161350 244840
rect 162228 237182 162256 265610
rect 162398 251832 162454 251841
rect 162398 251767 162454 251776
rect 162308 245744 162360 245750
rect 162308 245686 162360 245692
rect 162216 237176 162268 237182
rect 162216 237118 162268 237124
rect 162124 236020 162176 236026
rect 162124 235962 162176 235968
rect 161202 209808 161258 209817
rect 161202 209743 161258 209752
rect 162136 202745 162164 235962
rect 162320 226642 162348 245686
rect 162412 235793 162440 251767
rect 162398 235784 162454 235793
rect 162398 235719 162454 235728
rect 162308 226636 162360 226642
rect 162308 226578 162360 226584
rect 162688 209774 162716 285631
rect 162780 263702 162808 370466
rect 162872 311846 162900 532714
rect 165528 467900 165580 467906
rect 165528 467842 165580 467848
rect 164884 447840 164936 447846
rect 164884 447782 164936 447788
rect 164148 411324 164200 411330
rect 164148 411266 164200 411272
rect 162952 344548 163004 344554
rect 162952 344490 163004 344496
rect 162964 322318 162992 344490
rect 163504 335368 163556 335374
rect 163504 335310 163556 335316
rect 162952 322312 163004 322318
rect 162952 322254 163004 322260
rect 163516 319462 163544 335310
rect 163504 319456 163556 319462
rect 163504 319398 163556 319404
rect 163596 317620 163648 317626
rect 163596 317562 163648 317568
rect 163504 313404 163556 313410
rect 163504 313346 163556 313352
rect 162860 311840 162912 311846
rect 162860 311782 162912 311788
rect 162768 263696 162820 263702
rect 162768 263638 162820 263644
rect 163516 260166 163544 313346
rect 163608 297401 163636 317562
rect 164160 313993 164188 411266
rect 164240 356720 164292 356726
rect 164240 356662 164292 356668
rect 164700 356720 164752 356726
rect 164700 356662 164752 356668
rect 164146 313984 164202 313993
rect 164146 313919 164202 313928
rect 163594 297392 163650 297401
rect 163594 297327 163650 297336
rect 164252 294642 164280 356662
rect 164712 356153 164740 356662
rect 164698 356144 164754 356153
rect 164698 356079 164754 356088
rect 164896 309777 164924 447782
rect 164976 332036 165028 332042
rect 164976 331978 165028 331984
rect 164882 309768 164938 309777
rect 164882 309703 164938 309712
rect 164884 295996 164936 296002
rect 164884 295938 164936 295944
rect 164240 294636 164292 294642
rect 164240 294578 164292 294584
rect 163594 279440 163650 279449
rect 163594 279375 163650 279384
rect 163504 260160 163556 260166
rect 163504 260102 163556 260108
rect 163504 233912 163556 233918
rect 163504 233854 163556 233860
rect 162688 209746 162808 209774
rect 162122 202736 162178 202745
rect 162122 202671 162178 202680
rect 162780 195974 162808 209746
rect 163516 197334 163544 233854
rect 163608 230217 163636 279375
rect 164146 266384 164202 266393
rect 164146 266319 164202 266328
rect 164054 261488 164110 261497
rect 164054 261423 164110 261432
rect 164068 234705 164096 261423
rect 164160 237289 164188 266319
rect 164240 263696 164292 263702
rect 164240 263638 164292 263644
rect 164146 237280 164202 237289
rect 164146 237215 164202 237224
rect 164160 236026 164188 237215
rect 164148 236020 164200 236026
rect 164148 235962 164200 235968
rect 164054 234696 164110 234705
rect 164054 234631 164110 234640
rect 164252 232937 164280 263638
rect 164896 253230 164924 295938
rect 164884 253224 164936 253230
rect 164884 253166 164936 253172
rect 164988 251161 165016 331978
rect 165540 305046 165568 467842
rect 165620 382968 165672 382974
rect 165620 382910 165672 382916
rect 165632 308514 165660 382910
rect 166828 366382 166856 564402
rect 166908 542496 166960 542502
rect 166908 542438 166960 542444
rect 166816 366376 166868 366382
rect 166816 366318 166868 366324
rect 166354 364984 166410 364993
rect 166354 364919 166410 364928
rect 166264 311908 166316 311914
rect 166264 311850 166316 311856
rect 165620 308508 165672 308514
rect 165620 308450 165672 308456
rect 165068 305040 165120 305046
rect 165068 304982 165120 304988
rect 165528 305040 165580 305046
rect 165528 304982 165580 304988
rect 165080 286346 165108 304982
rect 165632 302938 165660 308450
rect 165620 302932 165672 302938
rect 165620 302874 165672 302880
rect 165158 287736 165214 287745
rect 165158 287671 165214 287680
rect 165068 286340 165120 286346
rect 165068 286282 165120 286288
rect 165068 278792 165120 278798
rect 165068 278734 165120 278740
rect 164974 251152 165030 251161
rect 164974 251087 165030 251096
rect 165080 244934 165108 278734
rect 165172 277370 165200 287671
rect 165160 277364 165212 277370
rect 165160 277306 165212 277312
rect 165160 252544 165212 252550
rect 165160 252486 165212 252492
rect 165068 244928 165120 244934
rect 165068 244870 165120 244876
rect 164976 242956 165028 242962
rect 164976 242898 165028 242904
rect 164884 240780 164936 240786
rect 164884 240722 164936 240728
rect 164238 232928 164294 232937
rect 164238 232863 164294 232872
rect 163594 230208 163650 230217
rect 163594 230143 163650 230152
rect 163504 197328 163556 197334
rect 163504 197270 163556 197276
rect 162768 195968 162820 195974
rect 162768 195910 162820 195916
rect 162780 195362 162808 195910
rect 162768 195356 162820 195362
rect 162768 195298 162820 195304
rect 164896 188426 164924 240722
rect 164988 215286 165016 242898
rect 165172 240825 165200 252486
rect 165158 240816 165214 240825
rect 165158 240751 165214 240760
rect 164976 215280 165028 215286
rect 164976 215222 165028 215228
rect 166276 202201 166304 311850
rect 166368 295225 166396 364919
rect 166446 332752 166502 332761
rect 166446 332687 166502 332696
rect 166460 312662 166488 332687
rect 166448 312656 166500 312662
rect 166448 312598 166500 312604
rect 166354 295216 166410 295225
rect 166354 295151 166410 295160
rect 166448 290488 166500 290494
rect 166448 290430 166500 290436
rect 166356 286340 166408 286346
rect 166356 286282 166408 286288
rect 166368 245750 166396 286282
rect 166460 262954 166488 290430
rect 166920 273057 166948 542438
rect 175924 538960 175976 538966
rect 175924 538902 175976 538908
rect 173162 536888 173218 536897
rect 173162 536823 173218 536832
rect 169114 535664 169170 535673
rect 169114 535599 169170 535608
rect 169024 506524 169076 506530
rect 169024 506466 169076 506472
rect 168288 448588 168340 448594
rect 168288 448530 168340 448536
rect 167000 403640 167052 403646
rect 167000 403582 167052 403588
rect 166906 273048 166962 273057
rect 166906 272983 166962 272992
rect 166920 272513 166948 272983
rect 166906 272504 166962 272513
rect 166906 272439 166962 272448
rect 166908 269884 166960 269890
rect 166908 269826 166960 269832
rect 166448 262948 166500 262954
rect 166448 262890 166500 262896
rect 166540 262540 166592 262546
rect 166540 262482 166592 262488
rect 166552 252550 166580 262482
rect 166540 252544 166592 252550
rect 166540 252486 166592 252492
rect 166356 245744 166408 245750
rect 166356 245686 166408 245692
rect 166446 245712 166502 245721
rect 166446 245647 166502 245656
rect 166460 228410 166488 245647
rect 166814 240136 166870 240145
rect 166814 240071 166870 240080
rect 166448 228404 166500 228410
rect 166448 228346 166500 228352
rect 166828 223417 166856 240071
rect 166920 235278 166948 269826
rect 167012 255270 167040 403582
rect 167092 385688 167144 385694
rect 167092 385630 167144 385636
rect 167104 325650 167132 385630
rect 168194 355328 168250 355337
rect 168194 355263 168250 355272
rect 167092 325644 167144 325650
rect 167092 325586 167144 325592
rect 167104 324358 167132 325586
rect 167092 324352 167144 324358
rect 167092 324294 167144 324300
rect 167644 306400 167696 306406
rect 167644 306342 167696 306348
rect 167656 279478 167684 306342
rect 168208 304978 168236 355263
rect 168196 304972 168248 304978
rect 168196 304914 168248 304920
rect 168208 304298 168236 304914
rect 168196 304292 168248 304298
rect 168196 304234 168248 304240
rect 167644 279472 167696 279478
rect 167644 279414 167696 279420
rect 167644 274712 167696 274718
rect 167644 274654 167696 274660
rect 167000 255264 167052 255270
rect 167000 255206 167052 255212
rect 167012 254590 167040 255206
rect 167000 254584 167052 254590
rect 167000 254526 167052 254532
rect 166908 235272 166960 235278
rect 166908 235214 166960 235220
rect 166998 234696 167054 234705
rect 166998 234631 167054 234640
rect 166814 223408 166870 223417
rect 166814 223343 166870 223352
rect 166828 219434 166856 223343
rect 166368 219406 166856 219434
rect 166262 202192 166318 202201
rect 166262 202127 166318 202136
rect 166368 201249 166396 219406
rect 166354 201240 166410 201249
rect 166354 201175 166410 201184
rect 167012 191146 167040 234631
rect 167656 229770 167684 274654
rect 168300 272542 168328 448530
rect 168380 443692 168432 443698
rect 168380 443634 168432 443640
rect 168392 443018 168420 443634
rect 168380 443012 168432 443018
rect 168380 442954 168432 442960
rect 168392 329769 168420 442954
rect 169036 334665 169064 506466
rect 169128 431934 169156 535599
rect 171048 465112 171100 465118
rect 171048 465054 171100 465060
rect 169116 431928 169168 431934
rect 169116 431870 169168 431876
rect 169668 396092 169720 396098
rect 169668 396034 169720 396040
rect 169114 368384 169170 368393
rect 169114 368319 169170 368328
rect 169022 334656 169078 334665
rect 169022 334591 169078 334600
rect 168378 329760 168434 329769
rect 168378 329695 168434 329704
rect 169036 301481 169064 334591
rect 169128 319530 169156 368319
rect 169680 357649 169708 396034
rect 171060 385694 171088 465054
rect 173176 429146 173204 536823
rect 175188 534812 175240 534818
rect 175188 534754 175240 534760
rect 173900 460964 173952 460970
rect 173900 460906 173952 460912
rect 173164 429140 173216 429146
rect 173164 429082 173216 429088
rect 171140 396772 171192 396778
rect 171140 396714 171192 396720
rect 171048 385688 171100 385694
rect 169758 385656 169814 385665
rect 171048 385630 171100 385636
rect 169758 385591 169814 385600
rect 169298 357640 169354 357649
rect 169298 357575 169354 357584
rect 169666 357640 169722 357649
rect 169666 357575 169722 357584
rect 169208 349852 169260 349858
rect 169208 349794 169260 349800
rect 169116 319524 169168 319530
rect 169116 319466 169168 319472
rect 169220 317422 169248 349794
rect 169312 349761 169340 357575
rect 169298 349752 169354 349761
rect 169298 349687 169354 349696
rect 169300 320884 169352 320890
rect 169300 320826 169352 320832
rect 169208 317416 169260 317422
rect 169208 317358 169260 317364
rect 169116 306400 169168 306406
rect 169116 306342 169168 306348
rect 169022 301472 169078 301481
rect 169022 301407 169078 301416
rect 169022 300248 169078 300257
rect 169022 300183 169078 300192
rect 168288 272536 168340 272542
rect 168288 272478 168340 272484
rect 168654 268424 168710 268433
rect 168654 268359 168710 268368
rect 167828 264240 167880 264246
rect 167828 264182 167880 264188
rect 167840 247625 167868 264182
rect 168668 262546 168696 268359
rect 168656 262540 168708 262546
rect 168656 262482 168708 262488
rect 168288 251184 168340 251190
rect 168288 251126 168340 251132
rect 167826 247616 167882 247625
rect 167826 247551 167882 247560
rect 167736 247104 167788 247110
rect 167736 247046 167788 247052
rect 167748 231742 167776 247046
rect 168300 243574 168328 251126
rect 168380 247512 168432 247518
rect 168380 247454 168432 247460
rect 168288 243568 168340 243574
rect 168288 243510 168340 243516
rect 167826 241768 167882 241777
rect 167826 241703 167882 241712
rect 167840 232801 167868 241703
rect 168392 240825 168420 247454
rect 168378 240816 168434 240825
rect 168378 240751 168434 240760
rect 167826 232792 167882 232801
rect 167826 232727 167882 232736
rect 167736 231736 167788 231742
rect 167736 231678 167788 231684
rect 167644 229764 167696 229770
rect 167644 229706 167696 229712
rect 168288 202768 168340 202774
rect 168288 202710 168340 202716
rect 168300 202162 168328 202710
rect 168288 202156 168340 202162
rect 168288 202098 168340 202104
rect 167000 191140 167052 191146
rect 167000 191082 167052 191088
rect 167012 190454 167040 191082
rect 166920 190426 167040 190454
rect 164884 188420 164936 188426
rect 164884 188362 164936 188368
rect 164976 187740 165028 187746
rect 164976 187682 165028 187688
rect 159914 182880 159970 182889
rect 159914 182815 159970 182824
rect 134800 182300 134852 182306
rect 134800 182242 134852 182248
rect 162860 182300 162912 182306
rect 162860 182242 162912 182248
rect 132406 177576 132462 177585
rect 132406 177511 132462 177520
rect 133786 177576 133842 177585
rect 133786 177511 133842 177520
rect 134812 177177 134840 182242
rect 148232 178084 148284 178090
rect 148232 178026 148284 178032
rect 134798 177168 134854 177177
rect 134798 177103 134854 177112
rect 148244 176769 148272 178026
rect 158996 176792 159048 176798
rect 99470 176760 99526 176769
rect 99470 176695 99526 176704
rect 103426 176760 103482 176769
rect 103426 176695 103482 176704
rect 123298 176760 123354 176769
rect 123298 176695 123354 176704
rect 126794 176760 126850 176769
rect 129462 176760 129518 176769
rect 126794 176695 126850 176704
rect 128176 176724 128228 176730
rect 129462 176695 129518 176704
rect 148230 176760 148286 176769
rect 148230 176695 148286 176704
rect 158994 176760 158996 176769
rect 159048 176760 159050 176769
rect 158994 176695 159050 176704
rect 128176 176666 128228 176672
rect 128188 176497 128216 176666
rect 135720 176656 135772 176662
rect 135720 176598 135772 176604
rect 128174 176488 128230 176497
rect 128174 176423 128230 176432
rect 130752 175976 130804 175982
rect 130752 175918 130804 175924
rect 130764 175681 130792 175918
rect 135732 175681 135760 176598
rect 130750 175672 130806 175681
rect 130750 175607 130806 175616
rect 135718 175672 135774 175681
rect 135718 175607 135774 175616
rect 162872 175098 162900 182242
rect 164882 178392 164938 178401
rect 164882 178327 164938 178336
rect 162860 175092 162912 175098
rect 162860 175034 162912 175040
rect 164896 162858 164924 178327
rect 164988 172514 165016 187682
rect 166920 184385 166948 190426
rect 166906 184376 166962 184385
rect 166906 184311 166962 184320
rect 167828 183660 167880 183666
rect 167828 183602 167880 183608
rect 166356 183592 166408 183598
rect 166356 183534 166408 183540
rect 166262 179480 166318 179489
rect 166262 179415 166318 179424
rect 165528 175976 165580 175982
rect 165528 175918 165580 175924
rect 165540 173874 165568 175918
rect 165528 173868 165580 173874
rect 165528 173810 165580 173816
rect 164976 172508 165028 172514
rect 164976 172450 165028 172456
rect 164884 162852 164936 162858
rect 164884 162794 164936 162800
rect 166276 155922 166304 179415
rect 166368 161430 166396 183534
rect 167642 182200 167698 182209
rect 167642 182135 167698 182144
rect 166446 179616 166502 179625
rect 166446 179551 166502 179560
rect 166460 165578 166488 179551
rect 166538 175536 166594 175545
rect 166538 175471 166594 175480
rect 166552 168366 166580 175471
rect 166540 168360 166592 168366
rect 166540 168302 166592 168308
rect 166448 165572 166500 165578
rect 166448 165514 166500 165520
rect 166356 161424 166408 161430
rect 166356 161366 166408 161372
rect 167656 157350 167684 182135
rect 167736 179512 167788 179518
rect 167736 179454 167788 179460
rect 167748 167006 167776 179454
rect 167840 171086 167868 183602
rect 168300 175273 168328 202098
rect 169036 200802 169064 300183
rect 169128 287026 169156 306342
rect 169116 287020 169168 287026
rect 169116 286962 169168 286968
rect 169116 284980 169168 284986
rect 169116 284922 169168 284928
rect 169128 202774 169156 284922
rect 169220 269074 169248 317358
rect 169312 311166 169340 320826
rect 169300 311160 169352 311166
rect 169300 311102 169352 311108
rect 169298 303784 169354 303793
rect 169298 303719 169354 303728
rect 169312 280158 169340 303719
rect 169300 280152 169352 280158
rect 169300 280094 169352 280100
rect 169300 274712 169352 274718
rect 169300 274654 169352 274660
rect 169208 269068 169260 269074
rect 169208 269010 169260 269016
rect 169208 262948 169260 262954
rect 169208 262890 169260 262896
rect 169220 202881 169248 262890
rect 169312 251190 169340 274654
rect 169300 251184 169352 251190
rect 169300 251126 169352 251132
rect 169772 248402 169800 385591
rect 169852 381540 169904 381546
rect 169852 381482 169904 381488
rect 169864 368393 169892 381482
rect 169850 368384 169906 368393
rect 169850 368319 169906 368328
rect 170404 357468 170456 357474
rect 170404 357410 170456 357416
rect 170416 337414 170444 357410
rect 170404 337408 170456 337414
rect 170404 337350 170456 337356
rect 169852 336796 169904 336802
rect 169852 336738 169904 336744
rect 169864 329186 169892 336738
rect 169852 329180 169904 329186
rect 169852 329122 169904 329128
rect 170404 328500 170456 328506
rect 170404 328442 170456 328448
rect 169852 327140 169904 327146
rect 169852 327082 169904 327088
rect 169864 325689 169892 327082
rect 169850 325680 169906 325689
rect 169850 325615 169906 325624
rect 170416 324970 170444 328442
rect 170496 327072 170548 327078
rect 170496 327014 170548 327020
rect 170404 324964 170456 324970
rect 170404 324906 170456 324912
rect 170508 311234 170536 327014
rect 170496 311228 170548 311234
rect 170496 311170 170548 311176
rect 170404 310548 170456 310554
rect 170404 310490 170456 310496
rect 169852 295384 169904 295390
rect 169852 295326 169904 295332
rect 169864 289814 169892 295326
rect 169852 289808 169904 289814
rect 169852 289750 169904 289756
rect 169850 269240 169906 269249
rect 169850 269175 169906 269184
rect 169760 248396 169812 248402
rect 169760 248338 169812 248344
rect 169772 247110 169800 248338
rect 169760 247104 169812 247110
rect 169760 247046 169812 247052
rect 169864 222873 169892 269175
rect 169850 222864 169906 222873
rect 169850 222799 169906 222808
rect 170416 219366 170444 310490
rect 171152 297430 171180 396714
rect 171784 388476 171836 388482
rect 171784 388418 171836 388424
rect 171140 297424 171192 297430
rect 171140 297366 171192 297372
rect 170496 287088 170548 287094
rect 170496 287030 170548 287036
rect 170508 269006 170536 287030
rect 170496 269000 170548 269006
rect 170496 268942 170548 268948
rect 170496 267708 170548 267714
rect 170496 267650 170548 267656
rect 170508 267617 170536 267650
rect 170494 267608 170550 267617
rect 170494 267543 170550 267552
rect 171796 226137 171824 388418
rect 173164 380928 173216 380934
rect 173164 380870 173216 380876
rect 172610 349752 172666 349761
rect 172610 349687 172666 349696
rect 172520 328568 172572 328574
rect 172520 328510 172572 328516
rect 171876 324352 171928 324358
rect 171876 324294 171928 324300
rect 171888 273873 171916 324294
rect 172532 295361 172560 328510
rect 172624 327185 172652 349687
rect 173176 334626 173204 380870
rect 173912 361593 173940 460906
rect 173898 361584 173954 361593
rect 173898 361519 173954 361528
rect 173912 360330 173940 361519
rect 175096 361480 175148 361486
rect 175096 361422 175148 361428
rect 173348 360324 173400 360330
rect 173348 360266 173400 360272
rect 173900 360324 173952 360330
rect 173900 360266 173952 360272
rect 173164 334620 173216 334626
rect 173164 334562 173216 334568
rect 172704 334008 172756 334014
rect 172704 333950 172756 333956
rect 172716 329118 172744 333950
rect 173254 330168 173310 330177
rect 173254 330103 173310 330112
rect 172704 329112 172756 329118
rect 172704 329054 172756 329060
rect 172610 327176 172666 327185
rect 172610 327111 172666 327120
rect 173162 311128 173218 311137
rect 173162 311063 173218 311072
rect 172518 295352 172574 295361
rect 172518 295287 172574 295296
rect 171968 287156 172020 287162
rect 171968 287098 172020 287104
rect 171874 273864 171930 273873
rect 171874 273799 171930 273808
rect 171980 243642 172008 287098
rect 172060 275324 172112 275330
rect 172060 275266 172112 275272
rect 171968 243636 172020 243642
rect 171968 243578 172020 243584
rect 172072 235793 172100 275266
rect 173176 256698 173204 311063
rect 173268 283257 173296 330103
rect 173360 319433 173388 360266
rect 175002 356824 175058 356833
rect 175002 356759 175058 356768
rect 174544 336864 174596 336870
rect 174544 336806 174596 336812
rect 174556 329798 174584 336806
rect 174544 329792 174596 329798
rect 174544 329734 174596 329740
rect 174544 329180 174596 329186
rect 174544 329122 174596 329128
rect 174556 319530 174584 329122
rect 174544 319524 174596 319530
rect 174544 319466 174596 319472
rect 173346 319424 173402 319433
rect 173346 319359 173402 319368
rect 175016 316033 175044 356759
rect 175002 316024 175058 316033
rect 175002 315959 175058 315968
rect 175016 315353 175044 315959
rect 175002 315344 175058 315353
rect 175002 315279 175058 315288
rect 174636 309800 174688 309806
rect 174636 309742 174688 309748
rect 174544 298784 174596 298790
rect 174544 298726 174596 298732
rect 174556 289105 174584 298726
rect 174542 289096 174598 289105
rect 174542 289031 174598 289040
rect 173254 283248 173310 283257
rect 173254 283183 173310 283192
rect 173256 280832 173308 280838
rect 173256 280774 173308 280780
rect 173164 256692 173216 256698
rect 173164 256634 173216 256640
rect 173162 249792 173218 249801
rect 173162 249727 173218 249736
rect 173176 246265 173204 249727
rect 173162 246256 173218 246265
rect 173162 246191 173218 246200
rect 172058 235784 172114 235793
rect 172058 235719 172114 235728
rect 171876 235272 171928 235278
rect 171876 235214 171928 235220
rect 171782 226128 171838 226137
rect 171782 226063 171838 226072
rect 170404 219360 170456 219366
rect 170404 219302 170456 219308
rect 169206 202872 169262 202881
rect 169206 202807 169262 202816
rect 169116 202768 169168 202774
rect 169116 202710 169168 202716
rect 169390 202328 169446 202337
rect 169390 202263 169446 202272
rect 169024 200796 169076 200802
rect 169024 200738 169076 200744
rect 169404 186318 169432 202263
rect 169392 186312 169444 186318
rect 169392 186254 169444 186260
rect 170404 180940 170456 180946
rect 170404 180882 170456 180888
rect 169116 178152 169168 178158
rect 169116 178094 169168 178100
rect 169022 176896 169078 176905
rect 169022 176831 169078 176840
rect 168286 175264 168342 175273
rect 168286 175199 168342 175208
rect 167918 171592 167974 171601
rect 167918 171527 167974 171536
rect 167932 171154 167960 171527
rect 167920 171148 167972 171154
rect 167920 171090 167972 171096
rect 167828 171080 167880 171086
rect 167828 171022 167880 171028
rect 167736 167000 167788 167006
rect 167736 166942 167788 166948
rect 169036 158710 169064 176831
rect 169128 169726 169156 178094
rect 169116 169720 169168 169726
rect 169116 169662 169168 169668
rect 170416 160070 170444 180882
rect 171782 178256 171838 178265
rect 171782 178191 171838 178200
rect 170494 175400 170550 175409
rect 170494 175335 170550 175344
rect 170508 161362 170536 175335
rect 171796 166938 171824 178191
rect 171888 175953 171916 235214
rect 173176 203590 173204 246191
rect 173268 237153 173296 280774
rect 174542 276720 174598 276729
rect 174542 276655 174598 276664
rect 173716 255400 173768 255406
rect 173716 255342 173768 255348
rect 173728 248414 173756 255342
rect 173808 255332 173860 255338
rect 173808 255274 173860 255280
rect 173820 251870 173848 255274
rect 173808 251864 173860 251870
rect 173808 251806 173860 251812
rect 173728 248386 173848 248414
rect 173254 237144 173310 237153
rect 173254 237079 173310 237088
rect 173820 233073 173848 248386
rect 173806 233064 173862 233073
rect 173806 232999 173862 233008
rect 173820 232665 173848 232999
rect 173806 232656 173862 232665
rect 173806 232591 173862 232600
rect 173164 203584 173216 203590
rect 173164 203526 173216 203532
rect 173256 182232 173308 182238
rect 173256 182174 173308 182180
rect 173164 176792 173216 176798
rect 173164 176734 173216 176740
rect 171874 175944 171930 175953
rect 171874 175879 171930 175888
rect 171784 166932 171836 166938
rect 171784 166874 171836 166880
rect 170496 161356 170548 161362
rect 170496 161298 170548 161304
rect 170404 160064 170456 160070
rect 170404 160006 170456 160012
rect 169024 158704 169076 158710
rect 169024 158646 169076 158652
rect 167644 157344 167696 157350
rect 167644 157286 167696 157292
rect 166264 155916 166316 155922
rect 166264 155858 166316 155864
rect 169116 150476 169168 150482
rect 169116 150418 169168 150424
rect 166264 146328 166316 146334
rect 166264 146270 166316 146276
rect 67638 128072 67694 128081
rect 67638 128007 67694 128016
rect 67652 82657 67680 128007
rect 164884 104168 164936 104174
rect 164884 104110 164936 104116
rect 67730 100736 67786 100745
rect 67730 100671 67786 100680
rect 67744 87650 67772 100671
rect 107750 94752 107806 94761
rect 107750 94687 107806 94696
rect 117134 94752 117190 94761
rect 117134 94687 117190 94696
rect 107764 93906 107792 94687
rect 117148 93974 117176 94687
rect 117136 93968 117188 93974
rect 117136 93910 117188 93916
rect 107752 93900 107804 93906
rect 107752 93842 107804 93848
rect 95054 93528 95110 93537
rect 95054 93463 95110 93472
rect 115846 93528 115902 93537
rect 115846 93463 115902 93472
rect 95068 93158 95096 93463
rect 103334 93256 103390 93265
rect 103334 93191 103390 93200
rect 110326 93256 110382 93265
rect 115860 93226 115888 93463
rect 110326 93191 110382 93200
rect 115848 93220 115900 93226
rect 90364 93152 90416 93158
rect 90364 93094 90416 93100
rect 95056 93152 95108 93158
rect 95056 93094 95108 93100
rect 86776 92540 86828 92546
rect 86776 92482 86828 92488
rect 86788 92449 86816 92482
rect 86774 92440 86830 92449
rect 86774 92375 86830 92384
rect 89074 92440 89130 92449
rect 89074 92375 89130 92384
rect 86130 92304 86186 92313
rect 86130 92239 86186 92248
rect 75734 91216 75790 91225
rect 75734 91151 75790 91160
rect 85486 91216 85542 91225
rect 85486 91151 85542 91160
rect 67732 87644 67784 87650
rect 67732 87586 67784 87592
rect 67638 82648 67694 82657
rect 67638 82583 67694 82592
rect 67546 68232 67602 68241
rect 67546 68167 67602 68176
rect 70306 62792 70362 62801
rect 70306 62727 70362 62736
rect 68926 44840 68982 44849
rect 68926 44775 68982 44784
rect 65524 18624 65576 18630
rect 65524 18566 65576 18572
rect 65536 3874 65564 18566
rect 67548 10396 67600 10402
rect 67548 10338 67600 10344
rect 65524 3868 65576 3874
rect 65524 3810 65576 3816
rect 67560 3534 67588 10338
rect 68940 3534 68968 44775
rect 70216 3596 70268 3602
rect 70216 3538 70268 3544
rect 66720 3528 66772 3534
rect 66720 3470 66772 3476
rect 67548 3528 67600 3534
rect 67548 3470 67600 3476
rect 67916 3528 67968 3534
rect 67916 3470 67968 3476
rect 68928 3528 68980 3534
rect 68928 3470 68980 3476
rect 69112 3528 69164 3534
rect 69112 3470 69164 3476
rect 64328 3460 64380 3466
rect 64328 3402 64380 3408
rect 64788 3460 64840 3466
rect 64788 3402 64840 3408
rect 64340 480 64368 3402
rect 65524 2100 65576 2106
rect 65524 2042 65576 2048
rect 65536 480 65564 2042
rect 66732 480 66760 3470
rect 67928 480 67956 3470
rect 69124 480 69152 3470
rect 70228 1850 70256 3538
rect 70320 3534 70348 62727
rect 75748 55214 75776 91151
rect 85500 82822 85528 91151
rect 86144 90409 86172 92239
rect 88984 91792 89036 91798
rect 88984 91734 89036 91740
rect 88062 91216 88118 91225
rect 88062 91151 88118 91160
rect 86130 90400 86186 90409
rect 86130 90335 86186 90344
rect 88076 86873 88104 91151
rect 88062 86864 88118 86873
rect 88062 86799 88118 86808
rect 85488 82816 85540 82822
rect 85488 82758 85540 82764
rect 75826 67008 75882 67017
rect 75826 66943 75882 66952
rect 75736 55208 75788 55214
rect 75736 55150 75788 55156
rect 71044 37936 71096 37942
rect 71044 37878 71096 37884
rect 71056 3670 71084 37878
rect 74448 31068 74500 31074
rect 74448 31010 74500 31016
rect 73068 25560 73120 25566
rect 73068 25502 73120 25508
rect 71504 7676 71556 7682
rect 71504 7618 71556 7624
rect 71044 3664 71096 3670
rect 71044 3606 71096 3612
rect 70308 3528 70360 3534
rect 70308 3470 70360 3476
rect 70228 1822 70348 1850
rect 70320 480 70348 1822
rect 71516 480 71544 7618
rect 73080 3534 73108 25502
rect 74460 3534 74488 31010
rect 72608 3528 72660 3534
rect 72608 3470 72660 3476
rect 73068 3528 73120 3534
rect 73068 3470 73120 3476
rect 73804 3528 73856 3534
rect 73804 3470 73856 3476
rect 74448 3528 74500 3534
rect 74448 3470 74500 3476
rect 72620 480 72648 3470
rect 73816 480 73844 3470
rect 75840 3262 75868 66943
rect 78586 65648 78642 65657
rect 78586 65583 78642 65592
rect 77208 40792 77260 40798
rect 77208 40734 77260 40740
rect 77220 3534 77248 40734
rect 76196 3528 76248 3534
rect 76196 3470 76248 3476
rect 77208 3528 77260 3534
rect 77208 3470 77260 3476
rect 75000 3256 75052 3262
rect 75000 3198 75052 3204
rect 75828 3256 75880 3262
rect 75828 3198 75880 3204
rect 75012 480 75040 3198
rect 76208 480 76236 3470
rect 77392 3392 77444 3398
rect 77392 3334 77444 3340
rect 77404 480 77432 3334
rect 78600 480 78628 65583
rect 86868 64184 86920 64190
rect 86868 64126 86920 64132
rect 79966 61568 80022 61577
rect 79966 61503 80022 61512
rect 79980 6914 80008 61503
rect 84108 53100 84160 53106
rect 84108 53042 84160 53048
rect 82726 26888 82782 26897
rect 82726 26823 82782 26832
rect 81348 11824 81400 11830
rect 81348 11766 81400 11772
rect 79704 6886 80008 6914
rect 79704 480 79732 6886
rect 81360 3534 81388 11766
rect 80888 3528 80940 3534
rect 80888 3470 80940 3476
rect 81348 3528 81400 3534
rect 81348 3470 81400 3476
rect 80900 480 80928 3470
rect 82740 3058 82768 26823
rect 84120 3466 84148 53042
rect 86776 44872 86828 44878
rect 86776 44814 86828 44820
rect 85488 28348 85540 28354
rect 85488 28290 85540 28296
rect 85500 3534 85528 28290
rect 86788 16574 86816 44814
rect 86696 16546 86816 16574
rect 85672 3596 85724 3602
rect 85672 3538 85724 3544
rect 84476 3528 84528 3534
rect 84476 3470 84528 3476
rect 85488 3528 85540 3534
rect 85488 3470 85540 3476
rect 83280 3460 83332 3466
rect 83280 3402 83332 3408
rect 84108 3460 84160 3466
rect 84108 3402 84160 3408
rect 82084 3052 82136 3058
rect 82084 2994 82136 3000
rect 82728 3052 82780 3058
rect 82728 2994 82780 3000
rect 82096 480 82124 2994
rect 83292 480 83320 3402
rect 84488 480 84516 3470
rect 85684 480 85712 3538
rect 86696 3482 86724 16546
rect 86880 6914 86908 64126
rect 88996 53174 89024 91734
rect 89088 91118 89116 92375
rect 89076 91112 89128 91118
rect 89076 91054 89128 91060
rect 89626 62928 89682 62937
rect 89626 62863 89682 62872
rect 88984 53168 89036 53174
rect 88984 53110 89036 53116
rect 87604 43512 87656 43518
rect 87604 43454 87656 43460
rect 86788 6886 86908 6914
rect 86788 3602 86816 6886
rect 87616 3670 87644 43454
rect 88248 22772 88300 22778
rect 88248 22714 88300 22720
rect 88260 6914 88288 22714
rect 87984 6886 88288 6914
rect 87604 3664 87656 3670
rect 87604 3606 87656 3612
rect 86776 3596 86828 3602
rect 86776 3538 86828 3544
rect 86696 3454 86908 3482
rect 86880 480 86908 3454
rect 87984 480 88012 6886
rect 89640 3534 89668 62863
rect 90376 47666 90404 93094
rect 102046 92440 102102 92449
rect 102046 92375 102102 92384
rect 97814 91352 97870 91361
rect 97814 91287 97870 91296
rect 99286 91352 99342 91361
rect 99286 91287 99342 91296
rect 101862 91352 101918 91361
rect 101862 91287 101918 91296
rect 91006 91216 91062 91225
rect 91006 91151 91062 91160
rect 93766 91216 93822 91225
rect 93766 91151 93822 91160
rect 94686 91216 94742 91225
rect 94686 91151 94742 91160
rect 96526 91216 96582 91225
rect 96526 91151 96582 91160
rect 91020 56574 91048 91151
rect 93780 84182 93808 91151
rect 94700 85513 94728 91151
rect 94686 85504 94742 85513
rect 94686 85439 94742 85448
rect 93768 84176 93820 84182
rect 96540 84153 96568 91151
rect 93768 84118 93820 84124
rect 96526 84144 96582 84153
rect 96526 84079 96582 84088
rect 97828 82793 97856 91287
rect 97906 91216 97962 91225
rect 97906 91151 97962 91160
rect 99194 91216 99250 91225
rect 99194 91151 99250 91160
rect 97814 82784 97870 82793
rect 97814 82719 97870 82728
rect 95146 79656 95202 79665
rect 95146 79591 95202 79600
rect 93766 76664 93822 76673
rect 93766 76599 93822 76608
rect 91008 56568 91060 56574
rect 91008 56510 91060 56516
rect 90364 47660 90416 47666
rect 90364 47602 90416 47608
rect 91008 42084 91060 42090
rect 91008 42026 91060 42032
rect 91020 3534 91048 42026
rect 92388 25628 92440 25634
rect 92388 25570 92440 25576
rect 92400 3534 92428 25570
rect 93780 3534 93808 76599
rect 95056 3596 95108 3602
rect 95056 3538 95108 3544
rect 89168 3528 89220 3534
rect 89168 3470 89220 3476
rect 89628 3528 89680 3534
rect 89628 3470 89680 3476
rect 90364 3528 90416 3534
rect 90364 3470 90416 3476
rect 91008 3528 91060 3534
rect 91008 3470 91060 3476
rect 91560 3528 91612 3534
rect 91560 3470 91612 3476
rect 92388 3528 92440 3534
rect 92388 3470 92440 3476
rect 92756 3528 92808 3534
rect 92756 3470 92808 3476
rect 93768 3528 93820 3534
rect 93768 3470 93820 3476
rect 93952 3528 94004 3534
rect 93952 3470 94004 3476
rect 89180 480 89208 3470
rect 90376 480 90404 3470
rect 91572 480 91600 3470
rect 92768 480 92796 3470
rect 93964 480 93992 3470
rect 95068 1850 95096 3538
rect 95160 3534 95188 79591
rect 97920 63510 97948 91151
rect 99208 81394 99236 91151
rect 99196 81388 99248 81394
rect 99196 81330 99248 81336
rect 97908 63504 97960 63510
rect 97908 63446 97960 63452
rect 97908 60036 97960 60042
rect 97908 59978 97960 59984
rect 96252 15972 96304 15978
rect 96252 15914 96304 15920
rect 95148 3528 95200 3534
rect 95148 3470 95200 3476
rect 95068 1822 95188 1850
rect 95160 480 95188 1822
rect 96264 480 96292 15914
rect 97920 3534 97948 59978
rect 99300 59362 99328 91287
rect 100574 91216 100630 91225
rect 100574 91151 100630 91160
rect 100588 87553 100616 91151
rect 100574 87544 100630 87553
rect 100574 87479 100630 87488
rect 101876 66230 101904 91287
rect 101954 91216 102010 91225
rect 102060 91186 102088 92375
rect 101954 91151 102010 91160
rect 102048 91180 102100 91186
rect 101968 71738 101996 91151
rect 102048 91122 102100 91128
rect 103348 89010 103376 93191
rect 106922 91760 106978 91769
rect 106922 91695 106978 91704
rect 106646 91624 106702 91633
rect 106646 91559 106702 91568
rect 103426 91216 103482 91225
rect 103426 91151 103482 91160
rect 104254 91216 104310 91225
rect 104254 91151 104310 91160
rect 104806 91216 104862 91225
rect 104806 91151 104862 91160
rect 105542 91216 105598 91225
rect 105542 91151 105598 91160
rect 106094 91216 106150 91225
rect 106094 91151 106150 91160
rect 103336 89004 103388 89010
rect 103336 88946 103388 88952
rect 101956 71732 102008 71738
rect 101956 71674 102008 71680
rect 101864 66224 101916 66230
rect 101864 66166 101916 66172
rect 99288 59356 99340 59362
rect 99288 59298 99340 59304
rect 102048 58676 102100 58682
rect 102048 58618 102100 58624
rect 98644 46300 98696 46306
rect 98644 46242 98696 46248
rect 98656 18698 98684 46242
rect 98644 18692 98696 18698
rect 98644 18634 98696 18640
rect 99288 18692 99340 18698
rect 99288 18634 99340 18640
rect 99300 3534 99328 18634
rect 100668 13184 100720 13190
rect 100668 13126 100720 13132
rect 100680 3534 100708 13126
rect 102060 3534 102088 58618
rect 103440 52426 103468 91151
rect 104268 85542 104296 91151
rect 104256 85536 104308 85542
rect 104256 85478 104308 85484
rect 104820 78577 104848 91151
rect 105556 87961 105584 91151
rect 105542 87952 105598 87961
rect 105542 87887 105598 87896
rect 105544 87644 105596 87650
rect 105544 87586 105596 87592
rect 104806 78568 104862 78577
rect 104806 78503 104862 78512
rect 104806 73944 104862 73953
rect 104806 73879 104862 73888
rect 103428 52420 103480 52426
rect 103428 52362 103480 52368
rect 103428 39432 103480 39438
rect 103428 39374 103480 39380
rect 103440 6914 103468 39374
rect 104820 6914 104848 73879
rect 105556 67590 105584 87586
rect 106108 74526 106136 91151
rect 106660 89593 106688 91559
rect 106646 89584 106702 89593
rect 106646 89519 106702 89528
rect 106186 82104 106242 82113
rect 106186 82039 106242 82048
rect 106096 74520 106148 74526
rect 106096 74462 106148 74468
rect 105544 67584 105596 67590
rect 105544 67526 105596 67532
rect 103348 6886 103468 6914
rect 104544 6886 104848 6914
rect 102232 6248 102284 6254
rect 102232 6190 102284 6196
rect 97448 3528 97500 3534
rect 97448 3470 97500 3476
rect 97908 3528 97960 3534
rect 97908 3470 97960 3476
rect 98644 3528 98696 3534
rect 98644 3470 98696 3476
rect 99288 3528 99340 3534
rect 99288 3470 99340 3476
rect 99840 3528 99892 3534
rect 99840 3470 99892 3476
rect 100668 3528 100720 3534
rect 100668 3470 100720 3476
rect 101036 3528 101088 3534
rect 101036 3470 101088 3476
rect 102048 3528 102100 3534
rect 102048 3470 102100 3476
rect 97460 480 97488 3470
rect 98656 480 98684 3470
rect 99852 480 99880 3470
rect 101048 480 101076 3470
rect 102244 480 102272 6190
rect 103348 480 103376 6886
rect 104544 480 104572 6886
rect 106200 3466 106228 82039
rect 106936 57934 106964 91695
rect 110234 91352 110290 91361
rect 110234 91287 110290 91296
rect 108946 91216 109002 91225
rect 108946 91151 109002 91160
rect 110142 91216 110198 91225
rect 110142 91151 110198 91160
rect 108960 84017 108988 91151
rect 108946 84008 109002 84017
rect 108946 83943 109002 83952
rect 108946 76528 109002 76537
rect 108946 76463 109002 76472
rect 106924 57928 106976 57934
rect 106924 57870 106976 57876
rect 106924 8968 106976 8974
rect 106924 8910 106976 8916
rect 105728 3460 105780 3466
rect 105728 3402 105780 3408
rect 106188 3460 106240 3466
rect 106188 3402 106240 3408
rect 105740 480 105768 3402
rect 106936 480 106964 8910
rect 108960 3466 108988 76463
rect 110156 64870 110184 91151
rect 110248 68950 110276 91287
rect 110340 90982 110368 93191
rect 115848 93162 115900 93168
rect 162214 92576 162270 92585
rect 115296 92540 115348 92546
rect 162214 92511 162270 92520
rect 115296 92482 115348 92488
rect 112350 92440 112406 92449
rect 112350 92375 112406 92384
rect 111246 91352 111302 91361
rect 111246 91287 111302 91296
rect 110328 90976 110380 90982
rect 110328 90918 110380 90924
rect 111064 90364 111116 90370
rect 111064 90306 111116 90312
rect 111076 78441 111104 90306
rect 111260 86970 111288 91287
rect 111706 91216 111762 91225
rect 111706 91151 111762 91160
rect 111248 86964 111300 86970
rect 111248 86906 111300 86912
rect 111156 86284 111208 86290
rect 111156 86226 111208 86232
rect 111062 78432 111118 78441
rect 111062 78367 111118 78376
rect 111168 75818 111196 86226
rect 111156 75812 111208 75818
rect 111156 75754 111208 75760
rect 111720 73166 111748 91151
rect 112364 91050 112392 92375
rect 114374 91352 114430 91361
rect 114374 91287 114430 91296
rect 112994 91216 113050 91225
rect 112994 91151 113050 91160
rect 112352 91044 112404 91050
rect 112352 90986 112404 90992
rect 111708 73160 111760 73166
rect 111708 73102 111760 73108
rect 113008 70310 113036 91151
rect 114388 88262 114416 91287
rect 114466 91216 114522 91225
rect 114466 91151 114522 91160
rect 115204 91180 115256 91186
rect 114376 88256 114428 88262
rect 114376 88198 114428 88204
rect 112996 70304 113048 70310
rect 112996 70246 113048 70252
rect 110236 68944 110288 68950
rect 110236 68886 110288 68892
rect 110144 64864 110196 64870
rect 110144 64806 110196 64812
rect 111708 57248 111760 57254
rect 111708 57190 111760 57196
rect 111614 53136 111670 53145
rect 111614 53071 111670 53080
rect 110328 32496 110380 32502
rect 110328 32438 110380 32444
rect 110340 3466 110368 32438
rect 111628 16574 111656 53071
rect 111536 16546 111656 16574
rect 108120 3460 108172 3466
rect 108120 3402 108172 3408
rect 108948 3460 109000 3466
rect 108948 3402 109000 3408
rect 109316 3460 109368 3466
rect 109316 3402 109368 3408
rect 110328 3460 110380 3466
rect 110328 3402 110380 3408
rect 108132 480 108160 3402
rect 109328 480 109356 3402
rect 111536 3058 111564 16546
rect 111720 6914 111748 57190
rect 112444 53168 112496 53174
rect 112444 53110 112496 53116
rect 112456 11665 112484 53110
rect 114480 51066 114508 91151
rect 115204 91122 115256 91128
rect 115216 69018 115244 91122
rect 115308 75886 115336 92482
rect 136088 92472 136140 92478
rect 132406 92440 132462 92449
rect 132406 92375 132462 92384
rect 134706 92440 134762 92449
rect 134706 92375 134762 92384
rect 136086 92440 136088 92449
rect 136140 92440 136142 92449
rect 136086 92375 136142 92384
rect 119710 91760 119766 91769
rect 119710 91695 119766 91704
rect 121734 91760 121790 91769
rect 121734 91695 121790 91704
rect 123758 91760 123814 91769
rect 123758 91695 123814 91704
rect 115846 91216 115902 91225
rect 115846 91151 115902 91160
rect 117226 91216 117282 91225
rect 117226 91151 117282 91160
rect 118054 91216 118110 91225
rect 118054 91151 118110 91160
rect 118606 91216 118662 91225
rect 118606 91151 118662 91160
rect 115860 80034 115888 91151
rect 115848 80028 115900 80034
rect 115848 79970 115900 79976
rect 117240 77178 117268 91151
rect 118068 85377 118096 91151
rect 118054 85368 118110 85377
rect 118054 85303 118110 85312
rect 117228 77172 117280 77178
rect 117228 77114 117280 77120
rect 115296 75880 115348 75886
rect 115296 75822 115348 75828
rect 115204 69012 115256 69018
rect 115204 68954 115256 68960
rect 115848 55888 115900 55894
rect 115848 55830 115900 55836
rect 114468 51060 114520 51066
rect 114468 51002 114520 51008
rect 114468 20052 114520 20058
rect 114468 19994 114520 20000
rect 112442 11656 112498 11665
rect 112442 11591 112498 11600
rect 111628 6886 111748 6914
rect 110512 3052 110564 3058
rect 110512 2994 110564 3000
rect 111524 3052 111576 3058
rect 111524 2994 111576 3000
rect 110524 480 110552 2994
rect 111628 480 111656 6886
rect 114480 3466 114508 19994
rect 115860 3466 115888 55830
rect 118620 53786 118648 91151
rect 119724 89690 119752 91695
rect 119894 91216 119950 91225
rect 119894 91151 119950 91160
rect 120446 91216 120502 91225
rect 120446 91151 120502 91160
rect 120814 91216 120870 91225
rect 120814 91151 120870 91160
rect 119712 89684 119764 89690
rect 119712 89626 119764 89632
rect 119908 62014 119936 91151
rect 120080 89004 120132 89010
rect 120080 88946 120132 88952
rect 120092 86737 120120 88946
rect 120078 86728 120134 86737
rect 120078 86663 120134 86672
rect 120460 86601 120488 91151
rect 120828 88330 120856 91151
rect 121748 89622 121776 91695
rect 122104 91112 122156 91118
rect 122104 91054 122156 91060
rect 121736 89616 121788 89622
rect 121736 89558 121788 89564
rect 120816 88324 120868 88330
rect 120816 88266 120868 88272
rect 120446 86592 120502 86601
rect 120446 86527 120502 86536
rect 120724 84856 120776 84862
rect 120724 84798 120776 84804
rect 119986 80880 120042 80889
rect 119986 80815 120042 80824
rect 119896 62008 119948 62014
rect 119896 61950 119948 61956
rect 118608 53780 118660 53786
rect 118608 53722 118660 53728
rect 116584 35284 116636 35290
rect 116584 35226 116636 35232
rect 116400 4072 116452 4078
rect 116400 4014 116452 4020
rect 114008 3460 114060 3466
rect 114008 3402 114060 3408
rect 114468 3460 114520 3466
rect 114468 3402 114520 3408
rect 115204 3460 115256 3466
rect 115204 3402 115256 3408
rect 115848 3460 115900 3466
rect 115848 3402 115900 3408
rect 112812 2168 112864 2174
rect 112812 2110 112864 2116
rect 112824 480 112852 2110
rect 114020 480 114048 3402
rect 115216 480 115244 3402
rect 116412 480 116440 4014
rect 116596 3398 116624 35226
rect 119896 17264 119948 17270
rect 119896 17206 119948 17212
rect 119908 16574 119936 17206
rect 119816 16546 119936 16574
rect 118608 14544 118660 14550
rect 118608 14486 118660 14492
rect 118620 3466 118648 14486
rect 119816 3466 119844 16546
rect 120000 6914 120028 80815
rect 120736 70378 120764 84798
rect 120724 70372 120776 70378
rect 120724 70314 120776 70320
rect 122116 63442 122144 91054
rect 123772 89729 123800 91695
rect 124034 91488 124090 91497
rect 124034 91423 124090 91432
rect 126794 91488 126850 91497
rect 126794 91423 126850 91432
rect 123942 91216 123998 91225
rect 123942 91151 123998 91160
rect 123758 89720 123814 89729
rect 123758 89655 123814 89664
rect 123482 89040 123538 89049
rect 123482 88975 123538 88984
rect 122746 74080 122802 74089
rect 122746 74015 122802 74024
rect 122104 63436 122156 63442
rect 122104 63378 122156 63384
rect 121368 51740 121420 51746
rect 121368 51682 121420 51688
rect 121380 6914 121408 51682
rect 119908 6886 120028 6914
rect 121104 6886 121408 6914
rect 117596 3460 117648 3466
rect 117596 3402 117648 3408
rect 118608 3460 118660 3466
rect 118608 3402 118660 3408
rect 118792 3460 118844 3466
rect 118792 3402 118844 3408
rect 119804 3460 119856 3466
rect 119804 3402 119856 3408
rect 116584 3392 116636 3398
rect 116584 3334 116636 3340
rect 117608 480 117636 3402
rect 118804 480 118832 3402
rect 119908 480 119936 6886
rect 121104 480 121132 6886
rect 122760 3466 122788 74015
rect 123496 73098 123524 88975
rect 123484 73092 123536 73098
rect 123484 73034 123536 73040
rect 123484 54528 123536 54534
rect 123484 54470 123536 54476
rect 123496 4078 123524 54470
rect 123956 49706 123984 91151
rect 124048 74458 124076 91423
rect 125506 91352 125562 91361
rect 125506 91287 125562 91296
rect 125414 91216 125470 91225
rect 125414 91151 125470 91160
rect 124036 74452 124088 74458
rect 124036 74394 124088 74400
rect 125428 66162 125456 91151
rect 125416 66156 125468 66162
rect 125416 66098 125468 66104
rect 125520 60722 125548 91287
rect 126702 91216 126758 91225
rect 126702 91151 126758 91160
rect 126242 84824 126298 84833
rect 126242 84759 126298 84768
rect 125508 60716 125560 60722
rect 125508 60658 125560 60664
rect 123944 49700 123996 49706
rect 123944 49642 123996 49648
rect 125508 36644 125560 36650
rect 125508 36586 125560 36592
rect 123484 4072 123536 4078
rect 123484 4014 123536 4020
rect 125520 3534 125548 36586
rect 126256 3602 126284 84759
rect 126716 84114 126744 91151
rect 126704 84108 126756 84114
rect 126704 84050 126756 84056
rect 126808 82754 126836 91423
rect 126886 91352 126942 91361
rect 126886 91287 126942 91296
rect 126796 82748 126848 82754
rect 126796 82690 126848 82696
rect 126900 81326 126928 91287
rect 128266 91216 128322 91225
rect 128266 91151 128322 91160
rect 130750 91216 130806 91225
rect 130750 91151 130806 91160
rect 126888 81320 126940 81326
rect 126888 81262 126940 81268
rect 128280 71670 128308 91151
rect 130764 88097 130792 91151
rect 132420 91118 132448 92375
rect 133786 91216 133842 91225
rect 133786 91151 133842 91160
rect 132408 91112 132460 91118
rect 132408 91054 132460 91060
rect 130750 88088 130806 88097
rect 130750 88023 130806 88032
rect 129002 87544 129058 87553
rect 129002 87479 129058 87488
rect 129016 78606 129044 87479
rect 133800 79966 133828 91151
rect 134720 91118 134748 92375
rect 160744 91792 160796 91798
rect 160744 91734 160796 91740
rect 151542 91488 151598 91497
rect 151542 91423 151598 91432
rect 134524 91112 134576 91118
rect 134524 91054 134576 91060
rect 134708 91112 134760 91118
rect 134708 91054 134760 91060
rect 133788 79960 133840 79966
rect 133788 79902 133840 79908
rect 129004 78600 129056 78606
rect 129004 78542 129056 78548
rect 128268 71664 128320 71670
rect 128268 71606 128320 71612
rect 130382 69728 130438 69737
rect 130382 69663 130438 69672
rect 126244 3596 126296 3602
rect 126244 3538 126296 3544
rect 130396 3534 130424 69663
rect 134536 62082 134564 91054
rect 151556 85474 151584 91423
rect 151726 91352 151782 91361
rect 151726 91287 151782 91296
rect 151634 91216 151690 91225
rect 151634 91151 151690 91160
rect 151544 85468 151596 85474
rect 151544 85410 151596 85416
rect 151648 78674 151676 91151
rect 151636 78668 151688 78674
rect 151636 78610 151688 78616
rect 151082 76800 151138 76809
rect 151082 76735 151138 76744
rect 134524 62076 134576 62082
rect 134524 62018 134576 62024
rect 151096 36650 151124 76735
rect 151740 67522 151768 91287
rect 152094 91216 152150 91225
rect 152094 91151 152096 91160
rect 152148 91151 152150 91160
rect 158720 91180 158772 91186
rect 152096 91122 152148 91128
rect 158720 91122 158772 91128
rect 153108 91112 153160 91118
rect 153106 91080 153108 91089
rect 153160 91080 153162 91089
rect 153106 91015 153162 91024
rect 157982 90536 158038 90545
rect 157982 90471 158038 90480
rect 157996 78606 158024 90471
rect 158732 86902 158760 91122
rect 160098 90400 160154 90409
rect 160098 90335 160154 90344
rect 160112 88233 160140 90335
rect 160098 88224 160154 88233
rect 160098 88159 160154 88168
rect 158720 86896 158772 86902
rect 158720 86838 158772 86844
rect 157984 78600 158036 78606
rect 157984 78542 158036 78548
rect 159364 77988 159416 77994
rect 159364 77930 159416 77936
rect 151728 67516 151780 67522
rect 151728 67458 151780 67464
rect 151084 36644 151136 36650
rect 151084 36586 151136 36592
rect 132498 21312 132554 21321
rect 132498 21247 132554 21256
rect 132512 16574 132540 21247
rect 142802 20088 142858 20097
rect 142802 20023 142858 20032
rect 132512 16546 133000 16574
rect 124680 3528 124732 3534
rect 124680 3470 124732 3476
rect 125508 3528 125560 3534
rect 129372 3528 129424 3534
rect 125508 3470 125560 3476
rect 125874 3496 125930 3505
rect 122288 3460 122340 3466
rect 122288 3402 122340 3408
rect 122748 3460 122800 3466
rect 122748 3402 122800 3408
rect 123484 3460 123536 3466
rect 123484 3402 123536 3408
rect 122300 480 122328 3402
rect 123496 480 123524 3402
rect 124692 480 124720 3470
rect 129372 3470 129424 3476
rect 130384 3528 130436 3534
rect 130384 3470 130436 3476
rect 125874 3431 125930 3440
rect 125888 480 125916 3431
rect 129384 480 129412 3470
rect 132972 480 133000 16546
rect 136454 11656 136510 11665
rect 136454 11591 136510 11600
rect 136468 480 136496 11591
rect 142816 2689 142844 20023
rect 159376 19990 159404 77930
rect 160756 77178 160784 91734
rect 162122 89856 162178 89865
rect 162122 89791 162178 89800
rect 162136 78577 162164 89791
rect 162228 82754 162256 92511
rect 162216 82748 162268 82754
rect 162216 82690 162268 82696
rect 164896 81326 164924 104110
rect 165528 96688 165580 96694
rect 165528 96630 165580 96636
rect 165436 95940 165488 95946
rect 165436 95882 165488 95888
rect 165448 94874 165476 95882
rect 165540 95033 165568 96630
rect 165526 95024 165582 95033
rect 165526 94959 165582 94968
rect 165448 94846 165568 94874
rect 165434 94208 165490 94217
rect 165434 94143 165490 94152
rect 165448 90545 165476 94143
rect 165540 92585 165568 94846
rect 165526 92576 165582 92585
rect 165526 92511 165582 92520
rect 165434 90536 165490 90545
rect 165434 90471 165490 90480
rect 164974 90400 165030 90409
rect 164974 90335 165030 90344
rect 164884 81320 164936 81326
rect 164884 81262 164936 81268
rect 162122 78568 162178 78577
rect 162122 78503 162178 78512
rect 160744 77172 160796 77178
rect 160744 77114 160796 77120
rect 164988 71738 165016 90335
rect 166276 79966 166304 146270
rect 167644 144220 167696 144226
rect 167644 144162 167696 144168
rect 166356 107704 166408 107710
rect 166356 107646 166408 107652
rect 166368 93158 166396 107646
rect 166448 99408 166500 99414
rect 166448 99350 166500 99356
rect 166356 93152 166408 93158
rect 166356 93094 166408 93100
rect 166460 86873 166488 99350
rect 166540 98048 166592 98054
rect 166540 97990 166592 97996
rect 166552 88233 166580 97990
rect 166538 88224 166594 88233
rect 166538 88159 166594 88168
rect 167656 88097 167684 144162
rect 167828 135924 167880 135930
rect 167828 135866 167880 135872
rect 167736 124228 167788 124234
rect 167736 124170 167788 124176
rect 167642 88088 167698 88097
rect 167642 88023 167698 88032
rect 166446 86864 166502 86873
rect 166446 86799 166502 86808
rect 166264 79960 166316 79966
rect 166264 79902 166316 79908
rect 167748 74458 167776 124170
rect 167840 113174 167868 135866
rect 167840 113146 167960 113174
rect 167828 111784 167880 111790
rect 167826 111752 167828 111761
rect 167880 111752 167882 111761
rect 167826 111687 167882 111696
rect 167932 108769 167960 113146
rect 169024 112464 169076 112470
rect 169024 112406 169076 112412
rect 168196 110424 168248 110430
rect 168196 110366 168248 110372
rect 168208 110129 168236 110366
rect 168194 110120 168250 110129
rect 168194 110055 168250 110064
rect 167918 108760 167974 108769
rect 167918 108695 167974 108704
rect 167920 107772 167972 107778
rect 167920 107714 167972 107720
rect 167828 106344 167880 106350
rect 167828 106286 167880 106292
rect 167840 93945 167868 106286
rect 167826 93936 167882 93945
rect 167826 93871 167882 93880
rect 167932 85513 167960 107714
rect 167918 85504 167974 85513
rect 167918 85439 167974 85448
rect 167736 74452 167788 74458
rect 167736 74394 167788 74400
rect 164976 71732 165028 71738
rect 164976 71674 165028 71680
rect 169036 67522 169064 112406
rect 169128 110430 169156 150418
rect 173176 149734 173204 176734
rect 173268 168298 173296 182174
rect 173256 168292 173308 168298
rect 173256 168234 173308 168240
rect 173164 149728 173216 149734
rect 173164 149670 173216 149676
rect 173256 147688 173308 147694
rect 173256 147630 173308 147636
rect 171784 136672 171836 136678
rect 171784 136614 171836 136620
rect 170404 127016 170456 127022
rect 170404 126958 170456 126964
rect 169208 120148 169260 120154
rect 169208 120090 169260 120096
rect 169116 110424 169168 110430
rect 169116 110366 169168 110372
rect 169116 104916 169168 104922
rect 169116 104858 169168 104864
rect 169128 82657 169156 104858
rect 169220 93974 169248 120090
rect 169300 100020 169352 100026
rect 169300 99962 169352 99968
rect 169208 93968 169260 93974
rect 169208 93910 169260 93916
rect 169312 85377 169340 99962
rect 169298 85368 169354 85377
rect 169298 85303 169354 85312
rect 169114 82648 169170 82657
rect 169114 82583 169170 82592
rect 169024 67516 169076 67522
rect 169024 67458 169076 67464
rect 170416 59362 170444 126958
rect 170496 122868 170548 122874
rect 170496 122810 170548 122816
rect 170508 89622 170536 122810
rect 170588 117360 170640 117366
rect 170588 117302 170640 117308
rect 170600 90982 170628 117302
rect 170680 109064 170732 109070
rect 170680 109006 170732 109012
rect 170588 90976 170640 90982
rect 170588 90918 170640 90924
rect 170496 89616 170548 89622
rect 170496 89558 170548 89564
rect 170692 84153 170720 109006
rect 171796 91798 171824 136614
rect 173164 133952 173216 133958
rect 173164 133894 173216 133900
rect 171876 114572 171928 114578
rect 171876 114514 171928 114520
rect 171784 91792 171836 91798
rect 171784 91734 171836 91740
rect 171888 89593 171916 114514
rect 172152 111852 172204 111858
rect 172152 111794 172204 111800
rect 171966 94480 172022 94489
rect 171966 94415 172022 94424
rect 171874 89584 171930 89593
rect 171874 89519 171930 89528
rect 171784 89004 171836 89010
rect 171784 88946 171836 88952
rect 170678 84144 170734 84153
rect 170678 84079 170734 84088
rect 171796 81433 171824 88946
rect 171782 81424 171838 81433
rect 171782 81359 171838 81368
rect 171980 77246 172008 94415
rect 172164 94217 172192 111794
rect 172150 94208 172206 94217
rect 172150 94143 172206 94152
rect 171968 77240 172020 77246
rect 171968 77182 172020 77188
rect 173176 73166 173204 133894
rect 173268 92478 173296 147630
rect 173440 113824 173492 113830
rect 173440 113766 173492 113772
rect 173348 98660 173400 98666
rect 173348 98602 173400 98608
rect 173256 92472 173308 92478
rect 173256 92414 173308 92420
rect 173164 73160 173216 73166
rect 173164 73102 173216 73108
rect 173360 63442 173388 98602
rect 173452 80034 173480 113766
rect 173440 80028 173492 80034
rect 173440 79970 173492 79976
rect 173348 63436 173400 63442
rect 173348 63378 173400 63384
rect 170404 59356 170456 59362
rect 170404 59298 170456 59304
rect 159364 19984 159416 19990
rect 174556 19961 174584 276655
rect 174648 247353 174676 309742
rect 175108 261594 175136 361422
rect 175200 332081 175228 534754
rect 175280 391264 175332 391270
rect 175280 391206 175332 391212
rect 175186 332072 175242 332081
rect 175186 332007 175242 332016
rect 175292 298110 175320 391206
rect 175936 372706 175964 538902
rect 177316 538121 177344 564470
rect 177946 557560 178002 557569
rect 177946 557495 178002 557504
rect 177394 538792 177450 538801
rect 177394 538727 177450 538736
rect 177302 538112 177358 538121
rect 177302 538047 177358 538056
rect 177408 529922 177436 538727
rect 177396 529916 177448 529922
rect 177396 529858 177448 529864
rect 177304 528624 177356 528630
rect 177304 528566 177356 528572
rect 176016 516180 176068 516186
rect 176016 516122 176068 516128
rect 176028 504393 176056 516122
rect 176014 504384 176070 504393
rect 176014 504319 176070 504328
rect 177316 500954 177344 528566
rect 177304 500948 177356 500954
rect 177304 500890 177356 500896
rect 176660 477556 176712 477562
rect 176660 477498 176712 477504
rect 176014 373280 176070 373289
rect 176014 373215 176070 373224
rect 175924 372700 175976 372706
rect 175924 372642 175976 372648
rect 175936 330614 175964 372642
rect 175924 330608 175976 330614
rect 175924 330550 175976 330556
rect 175924 304292 175976 304298
rect 175924 304234 175976 304240
rect 175280 298104 175332 298110
rect 175280 298046 175332 298052
rect 175740 298104 175792 298110
rect 175740 298046 175792 298052
rect 175752 297537 175780 298046
rect 175738 297528 175794 297537
rect 175738 297463 175794 297472
rect 175280 274780 175332 274786
rect 175280 274722 175332 274728
rect 175292 268433 175320 274722
rect 175278 268424 175334 268433
rect 175278 268359 175334 268368
rect 175096 261588 175148 261594
rect 175096 261530 175148 261536
rect 175188 259412 175240 259418
rect 175188 259354 175240 259360
rect 174726 250064 174782 250073
rect 174726 249999 174782 250008
rect 174634 247344 174690 247353
rect 174634 247279 174690 247288
rect 174740 195945 174768 249999
rect 175200 232529 175228 259354
rect 175186 232520 175242 232529
rect 175186 232455 175242 232464
rect 175200 231810 175228 232455
rect 175188 231804 175240 231810
rect 175188 231746 175240 231752
rect 175278 216064 175334 216073
rect 175278 215999 175334 216008
rect 175292 215966 175320 215999
rect 175280 215960 175332 215966
rect 175280 215902 175332 215908
rect 174726 195936 174782 195945
rect 174726 195871 174782 195880
rect 174636 189100 174688 189106
rect 174636 189042 174688 189048
rect 174648 169658 174676 189042
rect 174636 169652 174688 169658
rect 174636 169594 174688 169600
rect 174636 133204 174688 133210
rect 174636 133146 174688 133152
rect 174648 85474 174676 133146
rect 174728 120216 174780 120222
rect 174728 120158 174780 120164
rect 174740 93226 174768 120158
rect 174728 93220 174780 93226
rect 174728 93162 174780 93168
rect 174636 85468 174688 85474
rect 174636 85410 174688 85416
rect 175936 21321 175964 304234
rect 176028 292777 176056 373215
rect 176106 332888 176162 332897
rect 176106 332823 176162 332832
rect 176120 320958 176148 332823
rect 176108 320952 176160 320958
rect 176108 320894 176160 320900
rect 176014 292768 176070 292777
rect 176014 292703 176070 292712
rect 176028 280838 176056 292703
rect 176566 282296 176622 282305
rect 176566 282231 176622 282240
rect 176016 280832 176068 280838
rect 176016 280774 176068 280780
rect 176474 252648 176530 252657
rect 176016 252612 176068 252618
rect 176474 252583 176530 252592
rect 176016 252554 176068 252560
rect 176028 231810 176056 252554
rect 176016 231804 176068 231810
rect 176016 231746 176068 231752
rect 176488 217841 176516 252583
rect 176580 252550 176608 282231
rect 176672 255406 176700 477498
rect 177304 418192 177356 418198
rect 177304 418134 177356 418140
rect 176750 338056 176806 338065
rect 176750 337991 176806 338000
rect 176764 337385 176792 337991
rect 176750 337376 176806 337385
rect 176750 337311 176806 337320
rect 176660 255400 176712 255406
rect 176660 255342 176712 255348
rect 176568 252544 176620 252550
rect 176568 252486 176620 252492
rect 177316 249801 177344 418134
rect 177486 338328 177542 338337
rect 177486 338263 177542 338272
rect 177396 325032 177448 325038
rect 177396 324974 177448 324980
rect 177408 259418 177436 324974
rect 177500 316810 177528 338263
rect 177960 337385 177988 557495
rect 181536 556232 181588 556238
rect 181536 556174 181588 556180
rect 184386 556200 184442 556209
rect 180156 550656 180208 550662
rect 180156 550598 180208 550604
rect 180064 548004 180116 548010
rect 180064 547946 180116 547952
rect 178776 536852 178828 536858
rect 178776 536794 178828 536800
rect 178684 427848 178736 427854
rect 178684 427790 178736 427796
rect 177946 337376 178002 337385
rect 177946 337311 178002 337320
rect 178038 330032 178094 330041
rect 178038 329967 178094 329976
rect 178052 326466 178080 329967
rect 178040 326460 178092 326466
rect 178040 326402 178092 326408
rect 178038 325000 178094 325009
rect 178038 324935 178094 324944
rect 178052 320890 178080 324935
rect 178040 320884 178092 320890
rect 178040 320826 178092 320832
rect 177488 316804 177540 316810
rect 177488 316746 177540 316752
rect 178038 316704 178094 316713
rect 178038 316639 178094 316648
rect 177488 309188 177540 309194
rect 177488 309130 177540 309136
rect 177500 290494 177528 309130
rect 177488 290488 177540 290494
rect 177488 290430 177540 290436
rect 178052 274786 178080 316639
rect 178132 283620 178184 283626
rect 178132 283562 178184 283568
rect 178144 282946 178172 283562
rect 178132 282940 178184 282946
rect 178132 282882 178184 282888
rect 178040 274780 178092 274786
rect 178040 274722 178092 274728
rect 177396 259412 177448 259418
rect 177396 259354 177448 259360
rect 177396 257372 177448 257378
rect 177396 257314 177448 257320
rect 177302 249792 177358 249801
rect 177302 249727 177358 249736
rect 176568 248532 176620 248538
rect 176568 248474 176620 248480
rect 176580 243681 176608 248474
rect 177408 245041 177436 257314
rect 177948 256828 178000 256834
rect 177948 256770 178000 256776
rect 177856 245880 177908 245886
rect 177856 245822 177908 245828
rect 177868 245682 177896 245822
rect 177856 245676 177908 245682
rect 177856 245618 177908 245624
rect 177394 245032 177450 245041
rect 177394 244967 177450 244976
rect 177488 244928 177540 244934
rect 177488 244870 177540 244876
rect 176566 243672 176622 243681
rect 176566 243607 176622 243616
rect 177396 243568 177448 243574
rect 177396 243510 177448 243516
rect 177302 227760 177358 227769
rect 177302 227695 177358 227704
rect 176474 217832 176530 217841
rect 176474 217767 176530 217776
rect 177316 200122 177344 227695
rect 177304 200116 177356 200122
rect 177304 200058 177356 200064
rect 177304 195288 177356 195294
rect 177304 195230 177356 195236
rect 176016 138712 176068 138718
rect 176016 138654 176068 138660
rect 176028 86601 176056 138654
rect 176200 110492 176252 110498
rect 176200 110434 176252 110440
rect 176108 94580 176160 94586
rect 176108 94522 176160 94528
rect 176014 86592 176070 86601
rect 176014 86527 176070 86536
rect 176120 66230 176148 94522
rect 176212 94081 176240 110434
rect 176198 94072 176254 94081
rect 176198 94007 176254 94016
rect 176108 66224 176160 66230
rect 176108 66166 176160 66172
rect 175922 21312 175978 21321
rect 175922 21247 175978 21256
rect 159364 19926 159416 19932
rect 174542 19952 174598 19961
rect 174542 19887 174598 19896
rect 177316 4146 177344 195230
rect 177408 192506 177436 243510
rect 177500 216578 177528 244870
rect 177868 240786 177896 245618
rect 177856 240780 177908 240786
rect 177856 240722 177908 240728
rect 177960 228721 177988 256770
rect 178040 252544 178092 252550
rect 178040 252486 178092 252492
rect 178052 234433 178080 252486
rect 178696 245886 178724 427790
rect 178788 421598 178816 536794
rect 178868 423700 178920 423706
rect 178868 423642 178920 423648
rect 178776 421592 178828 421598
rect 178776 421534 178828 421540
rect 178774 359000 178830 359009
rect 178774 358935 178830 358944
rect 178788 324290 178816 358935
rect 178880 347993 178908 423642
rect 180076 357406 180104 547946
rect 180168 365809 180196 550598
rect 180800 487824 180852 487830
rect 180800 487766 180852 487772
rect 180248 463752 180300 463758
rect 180248 463694 180300 463700
rect 180260 372570 180288 463694
rect 180706 373280 180762 373289
rect 180706 373215 180762 373224
rect 180248 372564 180300 372570
rect 180248 372506 180300 372512
rect 180154 365800 180210 365809
rect 180154 365735 180210 365744
rect 180064 357400 180116 357406
rect 180064 357342 180116 357348
rect 180064 351960 180116 351966
rect 180064 351902 180116 351908
rect 178866 347984 178922 347993
rect 178866 347919 178922 347928
rect 178880 330449 178908 347919
rect 178866 330440 178922 330449
rect 178866 330375 178922 330384
rect 178776 324284 178828 324290
rect 178776 324226 178828 324232
rect 178866 285832 178922 285841
rect 178866 285767 178922 285776
rect 178776 268388 178828 268394
rect 178776 268330 178828 268336
rect 178684 245880 178736 245886
rect 178684 245822 178736 245828
rect 178788 241369 178816 268330
rect 178880 265674 178908 285767
rect 179328 282940 179380 282946
rect 179328 282882 179380 282888
rect 178868 265668 178920 265674
rect 178868 265610 178920 265616
rect 179340 250578 179368 282882
rect 180076 278089 180104 351902
rect 180168 327826 180196 365735
rect 180156 327820 180208 327826
rect 180156 327762 180208 327768
rect 180156 302932 180208 302938
rect 180156 302874 180208 302880
rect 180168 281518 180196 302874
rect 180260 300150 180288 372506
rect 180720 361457 180748 373215
rect 180706 361448 180762 361457
rect 180706 361383 180762 361392
rect 180340 357400 180392 357406
rect 180340 357342 180392 357348
rect 180352 356726 180380 357342
rect 180340 356720 180392 356726
rect 180340 356662 180392 356668
rect 180352 331945 180380 356662
rect 180338 331936 180394 331945
rect 180338 331871 180394 331880
rect 180340 329792 180392 329798
rect 180340 329734 180392 329740
rect 180248 300144 180300 300150
rect 180248 300086 180300 300092
rect 180352 291825 180380 329734
rect 180616 298784 180668 298790
rect 180616 298726 180668 298732
rect 180338 291816 180394 291825
rect 180338 291751 180394 291760
rect 180246 287600 180302 287609
rect 180246 287535 180302 287544
rect 180156 281512 180208 281518
rect 180156 281454 180208 281460
rect 180156 278112 180208 278118
rect 180062 278080 180118 278089
rect 180156 278054 180208 278060
rect 180062 278015 180118 278024
rect 180064 273352 180116 273358
rect 180064 273294 180116 273300
rect 179328 250572 179380 250578
rect 179328 250514 179380 250520
rect 180076 241466 180104 273294
rect 180064 241460 180116 241466
rect 180064 241402 180116 241408
rect 178774 241360 178830 241369
rect 178774 241295 178830 241304
rect 178038 234424 178094 234433
rect 178038 234359 178094 234368
rect 178052 234161 178080 234359
rect 178038 234152 178094 234161
rect 178038 234087 178094 234096
rect 178682 234152 178738 234161
rect 178682 234087 178738 234096
rect 177946 228712 178002 228721
rect 177946 228647 178002 228656
rect 177960 227769 177988 228647
rect 177946 227760 178002 227769
rect 177946 227695 178002 227704
rect 177488 216572 177540 216578
rect 177488 216514 177540 216520
rect 178696 197985 178724 234087
rect 180168 219201 180196 278054
rect 180260 269890 180288 287535
rect 180248 269884 180300 269890
rect 180248 269826 180300 269832
rect 180340 269884 180392 269890
rect 180340 269826 180392 269832
rect 180352 258074 180380 269826
rect 180260 258046 180380 258074
rect 180260 257961 180288 258046
rect 180246 257952 180302 257961
rect 180246 257887 180302 257896
rect 180260 250481 180288 257887
rect 180246 250472 180302 250481
rect 180246 250407 180302 250416
rect 180628 241641 180656 298726
rect 180812 256834 180840 487766
rect 181442 361040 181498 361049
rect 181442 360975 181498 360984
rect 180800 256828 180852 256834
rect 180800 256770 180852 256776
rect 180708 248464 180760 248470
rect 180708 248406 180760 248412
rect 180338 241632 180394 241641
rect 180338 241567 180394 241576
rect 180614 241632 180670 241641
rect 180614 241567 180670 241576
rect 180248 241460 180300 241466
rect 180248 241402 180300 241408
rect 180154 219192 180210 219201
rect 180154 219127 180210 219136
rect 180062 203552 180118 203561
rect 180062 203487 180118 203496
rect 178682 197976 178738 197985
rect 178682 197911 178738 197920
rect 177396 192500 177448 192506
rect 177396 192442 177448 192448
rect 177396 186448 177448 186454
rect 177396 186390 177448 186396
rect 177408 164218 177436 186390
rect 177396 164212 177448 164218
rect 177396 164154 177448 164160
rect 177488 142180 177540 142186
rect 177488 142122 177540 142128
rect 177396 116612 177448 116618
rect 177396 116554 177448 116560
rect 177408 74526 177436 116554
rect 177500 104174 177528 142122
rect 180076 141438 180104 203487
rect 180260 199617 180288 241402
rect 180352 238513 180380 241567
rect 180338 238504 180394 238513
rect 180338 238439 180394 238448
rect 180246 199608 180302 199617
rect 180246 199543 180302 199552
rect 180720 182918 180748 248406
rect 180708 182912 180760 182918
rect 180708 182854 180760 182860
rect 180154 182336 180210 182345
rect 180154 182271 180210 182280
rect 180168 165510 180196 182271
rect 180156 165504 180208 165510
rect 180156 165446 180208 165452
rect 181456 146946 181484 360975
rect 181548 360262 181576 556174
rect 184386 556135 184442 556144
rect 184204 547936 184256 547942
rect 184204 547878 184256 547884
rect 182822 539744 182878 539753
rect 182822 539679 182878 539688
rect 182088 487824 182140 487830
rect 182088 487766 182140 487772
rect 182100 487218 182128 487766
rect 182088 487212 182140 487218
rect 182088 487154 182140 487160
rect 181536 360256 181588 360262
rect 181536 360198 181588 360204
rect 181548 314129 181576 360198
rect 181628 325712 181680 325718
rect 181628 325654 181680 325660
rect 181640 315314 181668 325654
rect 181628 315308 181680 315314
rect 181628 315250 181680 315256
rect 181534 314120 181590 314129
rect 181534 314055 181590 314064
rect 182088 304292 182140 304298
rect 182088 304234 182140 304240
rect 181536 271176 181588 271182
rect 181536 271118 181588 271124
rect 181548 249762 181576 271118
rect 181536 249756 181588 249762
rect 181536 249698 181588 249704
rect 181718 247208 181774 247217
rect 181718 247143 181774 247152
rect 181534 244896 181590 244905
rect 181534 244831 181590 244840
rect 181444 146940 181496 146946
rect 181444 146882 181496 146888
rect 180064 141432 180116 141438
rect 180064 141374 180116 141380
rect 180064 135312 180116 135318
rect 180064 135254 180116 135260
rect 178776 129056 178828 129062
rect 178776 128998 178828 129004
rect 177580 124908 177632 124914
rect 177580 124850 177632 124856
rect 177488 104168 177540 104174
rect 177488 104110 177540 104116
rect 177488 100768 177540 100774
rect 177488 100710 177540 100716
rect 177500 82822 177528 100710
rect 177592 92177 177620 124850
rect 178684 121508 178736 121514
rect 178684 121450 178736 121456
rect 177578 92168 177634 92177
rect 177578 92103 177634 92112
rect 177488 82816 177540 82822
rect 177488 82758 177540 82764
rect 177396 74520 177448 74526
rect 177396 74462 177448 74468
rect 177394 69728 177450 69737
rect 177394 69663 177450 69672
rect 177304 4140 177356 4146
rect 177304 4082 177356 4088
rect 177408 3369 177436 69663
rect 178696 53786 178724 121450
rect 178788 62014 178816 128998
rect 178868 103556 178920 103562
rect 178868 103498 178920 103504
rect 178880 73098 178908 103498
rect 178868 73092 178920 73098
rect 178868 73034 178920 73040
rect 180076 70310 180104 135254
rect 181444 132524 181496 132530
rect 181444 132466 181496 132472
rect 180156 129804 180208 129810
rect 180156 129746 180208 129752
rect 180168 86737 180196 129746
rect 180154 86728 180210 86737
rect 180154 86663 180210 86672
rect 181456 84017 181484 132466
rect 181548 93129 181576 244831
rect 181628 243636 181680 243642
rect 181628 243578 181680 243584
rect 181640 229090 181668 243578
rect 181732 243574 181760 247143
rect 181720 243568 181772 243574
rect 181720 243510 181772 243516
rect 182100 235890 182128 304234
rect 182836 267714 182864 539679
rect 184216 354793 184244 547878
rect 184294 537024 184350 537033
rect 184294 536959 184350 536968
rect 184308 443698 184336 536959
rect 184400 518226 184428 556135
rect 187056 554872 187108 554878
rect 187056 554814 187108 554820
rect 187514 554840 187570 554849
rect 185584 545216 185636 545222
rect 185584 545158 185636 545164
rect 184388 518220 184440 518226
rect 184388 518162 184440 518168
rect 184296 443692 184348 443698
rect 184296 443634 184348 443640
rect 184388 443692 184440 443698
rect 184388 443634 184440 443640
rect 184296 383716 184348 383722
rect 184296 383658 184348 383664
rect 184308 373318 184336 383658
rect 184400 376038 184428 443634
rect 184388 376032 184440 376038
rect 184388 375974 184440 375980
rect 184296 373312 184348 373318
rect 184296 373254 184348 373260
rect 184400 369073 184428 375974
rect 184386 369064 184442 369073
rect 184386 368999 184442 369008
rect 184296 368620 184348 368626
rect 184296 368562 184348 368568
rect 184202 354784 184258 354793
rect 184202 354719 184258 354728
rect 183190 349208 183246 349217
rect 183190 349143 183246 349152
rect 183006 322280 183062 322289
rect 183006 322215 183062 322224
rect 182916 282192 182968 282198
rect 182916 282134 182968 282140
rect 182824 267708 182876 267714
rect 182824 267650 182876 267656
rect 182824 263696 182876 263702
rect 182824 263638 182876 263644
rect 182836 248470 182864 263638
rect 182824 248464 182876 248470
rect 182824 248406 182876 248412
rect 182270 245848 182326 245857
rect 182270 245783 182326 245792
rect 182284 244254 182312 245783
rect 182272 244248 182324 244254
rect 182272 244190 182324 244196
rect 182088 235884 182140 235890
rect 182088 235826 182140 235832
rect 181628 229084 181680 229090
rect 181628 229026 181680 229032
rect 182928 222154 182956 282134
rect 183020 264246 183048 322215
rect 183204 322153 183232 349143
rect 183190 322144 183246 322153
rect 183190 322079 183246 322088
rect 184216 298081 184244 354719
rect 184308 331158 184336 368562
rect 185398 365528 185454 365537
rect 185398 365463 185454 365472
rect 185412 365022 185440 365463
rect 185400 365016 185452 365022
rect 185400 364958 185452 364964
rect 185596 361865 185624 545158
rect 186962 538248 187018 538257
rect 186962 538183 187018 538192
rect 185676 455456 185728 455462
rect 185676 455398 185728 455404
rect 185688 441590 185716 455398
rect 185676 441584 185728 441590
rect 185676 441526 185728 441532
rect 185676 414044 185728 414050
rect 185676 413986 185728 413992
rect 185582 361856 185638 361865
rect 185582 361791 185638 361800
rect 184386 342408 184442 342417
rect 184386 342343 184442 342352
rect 184296 331152 184348 331158
rect 184296 331094 184348 331100
rect 184400 314022 184428 342343
rect 184480 330540 184532 330546
rect 184480 330482 184532 330488
rect 184388 314016 184440 314022
rect 184388 313958 184440 313964
rect 184492 310486 184520 330482
rect 185596 326398 185624 361791
rect 185584 326392 185636 326398
rect 185584 326334 185636 326340
rect 185584 322312 185636 322318
rect 185584 322254 185636 322260
rect 185596 312594 185624 322254
rect 185688 314265 185716 413986
rect 185768 387116 185820 387122
rect 185768 387058 185820 387064
rect 185780 377369 185808 387058
rect 185766 377360 185822 377369
rect 185766 377295 185822 377304
rect 186134 364440 186190 364449
rect 186134 364375 186190 364384
rect 186148 361554 186176 364375
rect 186136 361548 186188 361554
rect 186136 361490 186188 361496
rect 185674 314256 185730 314265
rect 185674 314191 185730 314200
rect 185584 312588 185636 312594
rect 185584 312530 185636 312536
rect 184480 310480 184532 310486
rect 184480 310422 184532 310428
rect 184294 307048 184350 307057
rect 184294 306983 184350 306992
rect 184202 298072 184258 298081
rect 184202 298007 184258 298016
rect 184308 293185 184336 306983
rect 184388 302320 184440 302326
rect 184388 302262 184440 302268
rect 184400 296002 184428 302262
rect 186042 301472 186098 301481
rect 186042 301407 186098 301416
rect 184846 298072 184902 298081
rect 184846 298007 184902 298016
rect 184860 296857 184888 298007
rect 184846 296848 184902 296857
rect 184846 296783 184902 296792
rect 184388 295996 184440 296002
rect 184388 295938 184440 295944
rect 184294 293176 184350 293185
rect 184294 293111 184350 293120
rect 183100 292596 183152 292602
rect 183100 292538 183152 292544
rect 183112 282742 183140 292538
rect 184020 289944 184072 289950
rect 184020 289886 184072 289892
rect 184032 287745 184060 289886
rect 184018 287736 184074 287745
rect 184018 287671 184074 287680
rect 184204 287156 184256 287162
rect 184204 287098 184256 287104
rect 183100 282736 183152 282742
rect 183100 282678 183152 282684
rect 183098 273864 183154 273873
rect 183098 273799 183154 273808
rect 183008 264240 183060 264246
rect 183008 264182 183060 264188
rect 183112 234433 183140 273799
rect 183560 272536 183612 272542
rect 183560 272478 183612 272484
rect 183572 260953 183600 272478
rect 183558 260944 183614 260953
rect 183558 260879 183614 260888
rect 184216 258738 184244 287098
rect 184860 273222 184888 296783
rect 185674 287328 185730 287337
rect 185674 287263 185730 287272
rect 185688 282305 185716 287263
rect 185674 282296 185730 282305
rect 185674 282231 185730 282240
rect 185582 278080 185638 278089
rect 185582 278015 185638 278024
rect 184848 273216 184900 273222
rect 184848 273158 184900 273164
rect 184480 261588 184532 261594
rect 184480 261530 184532 261536
rect 184204 258732 184256 258738
rect 184204 258674 184256 258680
rect 184216 258074 184244 258674
rect 184216 258046 184336 258074
rect 183468 249756 183520 249762
rect 183468 249698 183520 249704
rect 183480 248470 183508 249698
rect 183468 248464 183520 248470
rect 183468 248406 183520 248412
rect 183098 234424 183154 234433
rect 183098 234359 183154 234368
rect 182916 222148 182968 222154
rect 182916 222090 182968 222096
rect 183284 213920 183336 213926
rect 183282 213888 183284 213897
rect 183336 213888 183338 213897
rect 183282 213823 183338 213832
rect 182822 199472 182878 199481
rect 182822 199407 182878 199416
rect 181628 102808 181680 102814
rect 181628 102750 181680 102756
rect 181534 93120 181590 93129
rect 181534 93055 181590 93064
rect 181442 84008 181498 84017
rect 181442 83943 181498 83952
rect 181640 71670 181668 102750
rect 181628 71664 181680 71670
rect 181628 71606 181680 71612
rect 180064 70304 180116 70310
rect 180064 70246 180116 70252
rect 178776 62008 178828 62014
rect 178776 61950 178828 61956
rect 178684 53780 178736 53786
rect 178684 53722 178736 53728
rect 182836 30977 182864 199407
rect 183480 180713 183508 248406
rect 184204 229764 184256 229770
rect 184204 229706 184256 229712
rect 184216 222154 184244 229706
rect 184204 222148 184256 222154
rect 184204 222090 184256 222096
rect 184204 203584 184256 203590
rect 184204 203526 184256 203532
rect 183466 180704 183522 180713
rect 183466 180639 183522 180648
rect 182916 171148 182968 171154
rect 182916 171090 182968 171096
rect 182928 150414 182956 171090
rect 182916 150408 182968 150414
rect 182916 150350 182968 150356
rect 182916 125656 182968 125662
rect 182916 125598 182968 125604
rect 182928 84114 182956 125598
rect 182916 84108 182968 84114
rect 182916 84050 182968 84056
rect 182916 35216 182968 35222
rect 182916 35158 182968 35164
rect 182822 30968 182878 30977
rect 182822 30903 182878 30912
rect 182928 20058 182956 35158
rect 182916 20052 182968 20058
rect 182916 19994 182968 20000
rect 184216 19990 184244 203526
rect 184308 181490 184336 258046
rect 184386 250472 184442 250481
rect 184386 250407 184442 250416
rect 184296 181484 184348 181490
rect 184296 181426 184348 181432
rect 184400 180033 184428 250407
rect 184492 247042 184520 261530
rect 184848 250504 184900 250510
rect 184848 250446 184900 250452
rect 184480 247036 184532 247042
rect 184480 246978 184532 246984
rect 184860 244934 184888 250446
rect 184848 244928 184900 244934
rect 184848 244870 184900 244876
rect 184756 241596 184808 241602
rect 184756 241538 184808 241544
rect 184768 241369 184796 241538
rect 184754 241360 184810 241369
rect 184754 241295 184810 241304
rect 184756 226296 184808 226302
rect 184754 226264 184756 226273
rect 184808 226264 184810 226273
rect 184754 226199 184810 226208
rect 184768 225010 184796 226199
rect 184756 225004 184808 225010
rect 184756 224946 184808 224952
rect 184480 213920 184532 213926
rect 184480 213862 184532 213868
rect 184386 180024 184442 180033
rect 184386 179959 184442 179968
rect 184492 162178 184520 213862
rect 184860 210526 184888 244870
rect 185596 237153 185624 278015
rect 186056 277370 186084 301407
rect 186148 296177 186176 361490
rect 186976 347721 187004 538183
rect 187068 517478 187096 554814
rect 187514 554775 187570 554784
rect 187056 517472 187108 517478
rect 187056 517414 187108 517420
rect 187528 467838 187556 554775
rect 187516 467832 187568 467838
rect 187516 467774 187568 467780
rect 187056 398880 187108 398886
rect 187056 398822 187108 398828
rect 187068 397526 187096 398822
rect 187056 397520 187108 397526
rect 187056 397462 187108 397468
rect 187068 381177 187096 397462
rect 187240 386436 187292 386442
rect 187240 386378 187292 386384
rect 187054 381168 187110 381177
rect 187054 381103 187110 381112
rect 187056 376780 187108 376786
rect 187056 376722 187108 376728
rect 186962 347712 187018 347721
rect 186962 347647 187018 347656
rect 186228 328976 186280 328982
rect 186228 328918 186280 328924
rect 186134 296168 186190 296177
rect 186134 296103 186190 296112
rect 186044 277364 186096 277370
rect 186044 277306 186096 277312
rect 185676 274780 185728 274786
rect 185676 274722 185728 274728
rect 185688 248402 185716 274722
rect 186136 256760 186188 256766
rect 186136 256702 186188 256708
rect 185676 248396 185728 248402
rect 185676 248338 185728 248344
rect 185674 245032 185730 245041
rect 185674 244967 185730 244976
rect 185582 237144 185638 237153
rect 185582 237079 185638 237088
rect 185688 219201 185716 244967
rect 185674 219192 185730 219201
rect 185674 219127 185730 219136
rect 184848 210520 184900 210526
rect 184848 210462 184900 210468
rect 186148 187105 186176 256702
rect 186240 255338 186268 328918
rect 187068 264926 187096 376722
rect 187148 331288 187200 331294
rect 187148 331230 187200 331236
rect 187056 264920 187108 264926
rect 187056 264862 187108 264868
rect 186964 263628 187016 263634
rect 186964 263570 187016 263576
rect 186228 255332 186280 255338
rect 186228 255274 186280 255280
rect 186226 245848 186282 245857
rect 186226 245783 186282 245792
rect 186240 241369 186268 245783
rect 186226 241360 186282 241369
rect 186226 241295 186282 241304
rect 186134 187096 186190 187105
rect 186134 187031 186190 187040
rect 185584 184952 185636 184958
rect 185584 184894 185636 184900
rect 184570 180976 184626 180985
rect 184570 180911 184626 180920
rect 184480 162172 184532 162178
rect 184480 162114 184532 162120
rect 184584 155854 184612 180911
rect 185596 170377 185624 184894
rect 185582 170368 185638 170377
rect 185582 170303 185638 170312
rect 184572 155848 184624 155854
rect 184572 155790 184624 155796
rect 184296 145580 184348 145586
rect 184296 145522 184348 145528
rect 184308 91089 184336 145522
rect 184388 143608 184440 143614
rect 184388 143550 184440 143556
rect 184400 93673 184428 143550
rect 184480 117428 184532 117434
rect 184480 117370 184532 117376
rect 184386 93664 184442 93673
rect 184386 93599 184442 93608
rect 184294 91080 184350 91089
rect 184294 91015 184350 91024
rect 184492 86970 184520 117370
rect 185584 102196 185636 102202
rect 185584 102138 185636 102144
rect 184480 86964 184532 86970
rect 184480 86906 184532 86912
rect 184296 86284 184348 86290
rect 184296 86226 184348 86232
rect 184308 35290 184336 86226
rect 185596 75818 185624 102138
rect 185584 75812 185636 75818
rect 185584 75754 185636 75760
rect 184296 35284 184348 35290
rect 184296 35226 184348 35232
rect 184204 19984 184256 19990
rect 184204 19926 184256 19932
rect 186976 14521 187004 263570
rect 187160 251938 187188 331230
rect 187252 325038 187280 386378
rect 187620 374649 187648 589290
rect 197176 567248 197228 567254
rect 197176 567190 197228 567196
rect 195888 563168 195940 563174
rect 195888 563110 195940 563116
rect 193218 559600 193274 559609
rect 193218 559535 193274 559544
rect 193232 559065 193260 559535
rect 193218 559056 193274 559065
rect 192484 559020 192536 559026
rect 193218 558991 193274 559000
rect 192484 558962 192536 558968
rect 188344 553444 188396 553450
rect 188344 553386 188396 553392
rect 187606 374640 187662 374649
rect 187606 374575 187662 374584
rect 188356 363050 188384 553386
rect 189816 549296 189868 549302
rect 189816 549238 189868 549244
rect 188436 545148 188488 545154
rect 188436 545090 188488 545096
rect 188448 523734 188476 545090
rect 188436 523728 188488 523734
rect 188436 523670 188488 523676
rect 189724 522300 189776 522306
rect 189724 522242 189776 522248
rect 188436 495508 188488 495514
rect 188436 495450 188488 495456
rect 188344 363044 188396 363050
rect 188344 362986 188396 362992
rect 188448 354113 188476 495450
rect 188528 395344 188580 395350
rect 188528 395286 188580 395292
rect 188540 379574 188568 395286
rect 188618 381032 188674 381041
rect 188618 380967 188674 380976
rect 188528 379568 188580 379574
rect 188528 379510 188580 379516
rect 188526 357776 188582 357785
rect 188526 357711 188582 357720
rect 188434 354104 188490 354113
rect 188434 354039 188490 354048
rect 188344 331152 188396 331158
rect 188344 331094 188396 331100
rect 187240 325032 187292 325038
rect 187240 324974 187292 324980
rect 187238 291816 187294 291825
rect 187238 291751 187294 291760
rect 187252 258738 187280 291751
rect 187608 284436 187660 284442
rect 187608 284378 187660 284384
rect 187620 280922 187648 284378
rect 187620 280894 187740 280922
rect 187240 258732 187292 258738
rect 187240 258674 187292 258680
rect 187608 257100 187660 257106
rect 187608 257042 187660 257048
rect 187148 251932 187200 251938
rect 187148 251874 187200 251880
rect 187620 251841 187648 257042
rect 187606 251832 187662 251841
rect 187606 251767 187662 251776
rect 187056 250572 187108 250578
rect 187056 250514 187108 250520
rect 187068 180130 187096 250514
rect 187240 249824 187292 249830
rect 187240 249766 187292 249772
rect 187146 243672 187202 243681
rect 187146 243607 187202 243616
rect 187160 227730 187188 243607
rect 187252 233918 187280 249766
rect 187240 233912 187292 233918
rect 187240 233854 187292 233860
rect 187148 227724 187200 227730
rect 187148 227666 187200 227672
rect 187712 227662 187740 280894
rect 188356 267714 188384 331094
rect 188434 319424 188490 319433
rect 188434 319359 188490 319368
rect 188344 267708 188396 267714
rect 188344 267650 188396 267656
rect 188344 260160 188396 260166
rect 188344 260102 188396 260108
rect 187792 255332 187844 255338
rect 187792 255274 187844 255280
rect 187700 227656 187752 227662
rect 187700 227598 187752 227604
rect 187712 226370 187740 227598
rect 187700 226364 187752 226370
rect 187700 226306 187752 226312
rect 187698 216472 187754 216481
rect 187698 216407 187754 216416
rect 187712 216073 187740 216407
rect 187698 216064 187754 216073
rect 187698 215999 187754 216008
rect 187148 214668 187200 214674
rect 187148 214610 187200 214616
rect 187160 208282 187188 214610
rect 187804 209409 187832 255274
rect 188356 230382 188384 260102
rect 188448 257106 188476 319359
rect 188540 300257 188568 357711
rect 188632 331906 188660 380967
rect 188712 363044 188764 363050
rect 188712 362986 188764 362992
rect 188620 331900 188672 331906
rect 188620 331842 188672 331848
rect 188724 323649 188752 362986
rect 189736 335617 189764 522242
rect 189828 520266 189856 549238
rect 191102 547904 191158 547913
rect 191102 547839 191158 547848
rect 190366 533488 190422 533497
rect 190366 533423 190422 533432
rect 189816 520260 189868 520266
rect 189816 520202 189868 520208
rect 189908 399492 189960 399498
rect 189908 399434 189960 399440
rect 189816 379568 189868 379574
rect 189816 379510 189868 379516
rect 189722 335608 189778 335617
rect 189722 335543 189778 335552
rect 188710 323640 188766 323649
rect 188710 323575 188766 323584
rect 189078 320240 189134 320249
rect 189078 320175 189134 320184
rect 189092 318170 189120 320175
rect 189080 318164 189132 318170
rect 189080 318106 189132 318112
rect 189736 307086 189764 335543
rect 189724 307080 189776 307086
rect 189724 307022 189776 307028
rect 188526 300248 188582 300257
rect 188526 300183 188582 300192
rect 188988 297424 189040 297430
rect 188988 297366 189040 297372
rect 188526 291272 188582 291281
rect 188526 291207 188582 291216
rect 188540 286346 188568 291207
rect 188528 286340 188580 286346
rect 188528 286282 188580 286288
rect 188436 257100 188488 257106
rect 188436 257042 188488 257048
rect 188344 230376 188396 230382
rect 188344 230318 188396 230324
rect 188528 226364 188580 226370
rect 188528 226306 188580 226312
rect 188344 210452 188396 210458
rect 188344 210394 188396 210400
rect 187790 209400 187846 209409
rect 187790 209335 187846 209344
rect 187804 208457 187832 209335
rect 187790 208448 187846 208457
rect 187790 208383 187846 208392
rect 187148 208276 187200 208282
rect 187148 208218 187200 208224
rect 188356 204202 188384 210394
rect 188344 204196 188396 204202
rect 188344 204138 188396 204144
rect 188342 203552 188398 203561
rect 188342 203487 188398 203496
rect 187056 180124 187108 180130
rect 187056 180066 187108 180072
rect 187148 150544 187200 150550
rect 187148 150486 187200 150492
rect 187056 116000 187108 116006
rect 187056 115942 187108 115948
rect 187068 68950 187096 115942
rect 187160 111790 187188 150486
rect 187240 114640 187292 114646
rect 187240 114582 187292 114588
rect 187148 111784 187200 111790
rect 187148 111726 187200 111732
rect 187252 87961 187280 114582
rect 187238 87952 187294 87961
rect 187238 87887 187294 87896
rect 187056 68944 187108 68950
rect 187056 68886 187108 68892
rect 188356 20097 188384 203487
rect 188434 196752 188490 196761
rect 188434 196687 188490 196696
rect 188448 28257 188476 196687
rect 188540 193934 188568 226306
rect 189000 219434 189028 297366
rect 189080 278044 189132 278050
rect 189080 277986 189132 277992
rect 189092 276690 189120 277986
rect 189080 276684 189132 276690
rect 189080 276626 189132 276632
rect 189828 269006 189856 379510
rect 189920 376718 189948 399434
rect 189908 376712 189960 376718
rect 189908 376654 189960 376660
rect 190380 369170 190408 533423
rect 191116 514078 191144 547839
rect 191194 545456 191250 545465
rect 191194 545391 191250 545400
rect 191208 533390 191236 545391
rect 191746 541376 191802 541385
rect 191746 541311 191802 541320
rect 191196 533384 191248 533390
rect 191196 533326 191248 533332
rect 191104 514072 191156 514078
rect 191104 514014 191156 514020
rect 191104 480480 191156 480486
rect 191104 480422 191156 480428
rect 191116 388482 191144 480422
rect 191196 467832 191248 467838
rect 191196 467774 191248 467780
rect 191104 388476 191156 388482
rect 191104 388418 191156 388424
rect 191104 385688 191156 385694
rect 191104 385630 191156 385636
rect 190368 369164 190420 369170
rect 190368 369106 190420 369112
rect 190092 357536 190144 357542
rect 190092 357478 190144 357484
rect 189906 339824 189962 339833
rect 189906 339759 189962 339768
rect 189920 334694 189948 339759
rect 189908 334688 189960 334694
rect 189908 334630 189960 334636
rect 190104 331809 190132 357478
rect 190090 331800 190146 331809
rect 190090 331735 190146 331744
rect 190368 285796 190420 285802
rect 190368 285738 190420 285744
rect 190276 276684 190328 276690
rect 190276 276626 190328 276632
rect 189080 269000 189132 269006
rect 189080 268942 189132 268948
rect 189816 269000 189868 269006
rect 189816 268942 189868 268948
rect 189092 268394 189120 268942
rect 189080 268388 189132 268394
rect 189080 268330 189132 268336
rect 189080 266416 189132 266422
rect 189080 266358 189132 266364
rect 189092 260137 189120 266358
rect 189078 260128 189134 260137
rect 189078 260063 189134 260072
rect 190182 252512 190238 252521
rect 190182 252447 190238 252456
rect 189724 247716 189776 247722
rect 189724 247658 189776 247664
rect 189736 224942 189764 247658
rect 190196 238746 190224 252447
rect 190288 242894 190316 276626
rect 190276 242888 190328 242894
rect 190276 242830 190328 242836
rect 190184 238740 190236 238746
rect 190184 238682 190236 238688
rect 189724 224936 189776 224942
rect 189724 224878 189776 224884
rect 188816 219406 189028 219434
rect 188816 216073 188844 219406
rect 188802 216064 188858 216073
rect 188802 215999 188858 216008
rect 189080 212628 189132 212634
rect 189080 212570 189132 212576
rect 189092 212537 189120 212570
rect 189078 212528 189134 212537
rect 189078 212463 189134 212472
rect 188618 208448 188674 208457
rect 188618 208383 188674 208392
rect 188632 195401 188660 208383
rect 188618 195392 188674 195401
rect 188618 195327 188674 195336
rect 188528 193928 188580 193934
rect 188528 193870 188580 193876
rect 188526 180840 188582 180849
rect 188526 180775 188582 180784
rect 188540 157282 188568 180775
rect 189736 177449 189764 224878
rect 190380 212634 190408 285738
rect 191116 271862 191144 385630
rect 191208 378457 191236 467774
rect 191656 394732 191708 394738
rect 191656 394674 191708 394680
rect 191194 378448 191250 378457
rect 191194 378383 191250 378392
rect 191196 372632 191248 372638
rect 191196 372574 191248 372580
rect 191208 338745 191236 372574
rect 191668 353433 191696 394674
rect 191760 373425 191788 541311
rect 191746 373416 191802 373425
rect 191746 373351 191802 373360
rect 192496 358834 192524 558962
rect 192574 549536 192630 549545
rect 192574 549471 192630 549480
rect 192588 447846 192616 549471
rect 192576 447840 192628 447846
rect 192576 447782 192628 447788
rect 192576 433356 192628 433362
rect 192576 433298 192628 433304
rect 192484 358828 192536 358834
rect 192484 358770 192536 358776
rect 191654 353424 191710 353433
rect 191654 353359 191710 353368
rect 191668 347070 191696 353359
rect 191746 351112 191802 351121
rect 191746 351047 191802 351056
rect 191656 347064 191708 347070
rect 191656 347006 191708 347012
rect 191194 338736 191250 338745
rect 191194 338671 191250 338680
rect 191194 332072 191250 332081
rect 191194 332007 191250 332016
rect 191208 294545 191236 332007
rect 191288 295384 191340 295390
rect 191288 295326 191340 295332
rect 191194 294536 191250 294545
rect 191194 294471 191250 294480
rect 191194 284064 191250 284073
rect 191194 283999 191250 284008
rect 191208 274650 191236 283999
rect 191196 274644 191248 274650
rect 191196 274586 191248 274592
rect 191104 271856 191156 271862
rect 191104 271798 191156 271804
rect 191196 271244 191248 271250
rect 191196 271186 191248 271192
rect 191208 252521 191236 271186
rect 191300 262954 191328 295326
rect 191288 262948 191340 262954
rect 191288 262890 191340 262896
rect 191380 262200 191432 262206
rect 191380 262142 191432 262148
rect 191288 254584 191340 254590
rect 191288 254526 191340 254532
rect 191194 252512 191250 252521
rect 191194 252447 191250 252456
rect 191104 242888 191156 242894
rect 191104 242830 191156 242836
rect 190368 212628 190420 212634
rect 190368 212570 190420 212576
rect 190460 200864 190512 200870
rect 190460 200806 190512 200812
rect 190472 197169 190500 200806
rect 190458 197160 190514 197169
rect 190458 197095 190514 197104
rect 191116 184210 191144 242830
rect 191300 237017 191328 254526
rect 191286 237008 191342 237017
rect 191286 236943 191342 236952
rect 191392 195294 191420 262142
rect 191760 259418 191788 351047
rect 192496 320793 192524 358770
rect 192588 328982 192616 433298
rect 193232 400926 193260 558991
rect 195428 557592 195480 557598
rect 195428 557534 195480 557540
rect 193864 552152 193916 552158
rect 193864 552094 193916 552100
rect 193220 400920 193272 400926
rect 193220 400862 193272 400868
rect 193232 400246 193260 400862
rect 193220 400240 193272 400246
rect 193220 400182 193272 400188
rect 192668 382288 192720 382294
rect 192668 382230 192720 382236
rect 192680 365809 192708 382230
rect 192666 365800 192722 365809
rect 192666 365735 192722 365744
rect 193876 364585 193904 552094
rect 195334 548040 195390 548049
rect 195334 547975 195390 547984
rect 194140 543856 194192 543862
rect 194140 543798 194192 543804
rect 194152 538966 194180 543798
rect 195244 542428 195296 542434
rect 195244 542370 195296 542376
rect 194140 538960 194192 538966
rect 194140 538902 194192 538908
rect 195256 538898 195284 542370
rect 195244 538892 195296 538898
rect 195244 538834 195296 538840
rect 193954 538384 194010 538393
rect 193954 538319 194010 538328
rect 193968 382945 193996 538319
rect 195244 538280 195296 538286
rect 195244 538222 195296 538228
rect 194048 401668 194100 401674
rect 194048 401610 194100 401616
rect 193954 382936 194010 382945
rect 193954 382871 194010 382880
rect 193862 364576 193918 364585
rect 193862 364511 193918 364520
rect 193876 364334 193904 364511
rect 193876 364306 193996 364334
rect 192668 334620 192720 334626
rect 192668 334562 192720 334568
rect 192576 328976 192628 328982
rect 192576 328918 192628 328924
rect 192482 320784 192538 320793
rect 192482 320719 192538 320728
rect 192484 311160 192536 311166
rect 192484 311102 192536 311108
rect 191840 271856 191892 271862
rect 191840 271798 191892 271804
rect 191852 261526 191880 271798
rect 191840 261520 191892 261526
rect 191840 261462 191892 261468
rect 191748 259412 191800 259418
rect 191748 259354 191800 259360
rect 191656 251864 191708 251870
rect 191656 251806 191708 251812
rect 191668 210361 191696 251806
rect 191748 247172 191800 247178
rect 191748 247114 191800 247120
rect 191760 243545 191788 247114
rect 191746 243536 191802 243545
rect 191746 243471 191802 243480
rect 192496 240310 192524 311102
rect 192574 289912 192630 289921
rect 192574 289847 192630 289856
rect 192588 282198 192616 289847
rect 192576 282192 192628 282198
rect 192576 282134 192628 282140
rect 192680 273154 192708 334562
rect 193864 320952 193916 320958
rect 193864 320894 193916 320900
rect 192760 282124 192812 282130
rect 192760 282066 192812 282072
rect 192668 273148 192720 273154
rect 192668 273090 192720 273096
rect 192574 251152 192630 251161
rect 192574 251087 192630 251096
rect 192484 240304 192536 240310
rect 192484 240246 192536 240252
rect 191746 236056 191802 236065
rect 191746 235991 191802 236000
rect 191760 231577 191788 235991
rect 191746 231568 191802 231577
rect 191746 231503 191802 231512
rect 192484 216708 192536 216714
rect 192484 216650 192536 216656
rect 191654 210352 191710 210361
rect 191654 210287 191710 210296
rect 191380 195288 191432 195294
rect 191380 195230 191432 195236
rect 191196 193860 191248 193866
rect 191196 193802 191248 193808
rect 191104 184204 191156 184210
rect 191104 184146 191156 184152
rect 189722 177440 189778 177449
rect 189722 177375 189778 177384
rect 188528 157276 188580 157282
rect 188528 157218 188580 157224
rect 191102 142760 191158 142769
rect 191102 142695 191158 142704
rect 189724 139460 189776 139466
rect 189724 139402 189776 139408
rect 188528 123480 188580 123486
rect 188528 123422 188580 123428
rect 188540 49706 188568 123422
rect 189736 92313 189764 139402
rect 189722 92304 189778 92313
rect 189722 92239 189778 92248
rect 188528 49700 188580 49706
rect 188528 49642 188580 49648
rect 188434 28248 188490 28257
rect 188434 28183 188490 28192
rect 188342 20088 188398 20097
rect 187056 20052 187108 20058
rect 188342 20023 188398 20032
rect 187056 19994 187108 20000
rect 186962 14512 187018 14521
rect 186962 14447 187018 14456
rect 187068 3466 187096 19994
rect 191116 4865 191144 142695
rect 191208 91089 191236 193802
rect 192496 191146 192524 216650
rect 192588 200841 192616 251087
rect 192772 247178 192800 282066
rect 193220 279472 193272 279478
rect 193220 279414 193272 279420
rect 193232 278798 193260 279414
rect 193220 278792 193272 278798
rect 193220 278734 193272 278740
rect 193232 262206 193260 278734
rect 193220 262200 193272 262206
rect 193220 262142 193272 262148
rect 193128 259480 193180 259486
rect 193128 259422 193180 259428
rect 193036 252612 193088 252618
rect 193036 252554 193088 252560
rect 193048 251161 193076 252554
rect 193034 251152 193090 251161
rect 193034 251087 193090 251096
rect 192760 247172 192812 247178
rect 192760 247114 192812 247120
rect 192668 247104 192720 247110
rect 192668 247046 192720 247052
rect 192680 217938 192708 247046
rect 193140 220726 193168 259422
rect 193876 249762 193904 320894
rect 193968 305697 193996 364306
rect 193954 305688 194010 305697
rect 193954 305623 194010 305632
rect 194060 297430 194088 401610
rect 194140 400240 194192 400246
rect 194140 400182 194192 400188
rect 194152 328545 194180 400182
rect 195256 380225 195284 538222
rect 195348 520946 195376 547975
rect 195440 531282 195468 557534
rect 195428 531276 195480 531282
rect 195428 531218 195480 531224
rect 195336 520940 195388 520946
rect 195336 520882 195388 520888
rect 195796 470756 195848 470762
rect 195796 470698 195848 470704
rect 195242 380216 195298 380225
rect 195242 380151 195298 380160
rect 194598 379536 194654 379545
rect 194598 379471 194654 379480
rect 194612 375290 194640 379471
rect 195244 378208 195296 378214
rect 195244 378150 195296 378156
rect 194600 375284 194652 375290
rect 194600 375226 194652 375232
rect 195256 373969 195284 378150
rect 195702 376544 195758 376553
rect 195702 376479 195758 376488
rect 195336 374060 195388 374066
rect 195336 374002 195388 374008
rect 195242 373960 195298 373969
rect 195242 373895 195298 373904
rect 195348 371210 195376 374002
rect 195336 371204 195388 371210
rect 195336 371146 195388 371152
rect 195244 368552 195296 368558
rect 195244 368494 195296 368500
rect 195256 367849 195284 368494
rect 195242 367840 195298 367849
rect 195242 367775 195298 367784
rect 195716 351393 195744 376479
rect 195702 351384 195758 351393
rect 195702 351319 195758 351328
rect 195244 351212 195296 351218
rect 195244 351154 195296 351160
rect 195256 347177 195284 351154
rect 195242 347168 195298 347177
rect 195242 347103 195298 347112
rect 195244 341556 195296 341562
rect 195244 341498 195296 341504
rect 194138 328536 194194 328545
rect 194138 328471 194194 328480
rect 194152 325694 194180 328471
rect 194152 325666 194548 325694
rect 194140 301572 194192 301578
rect 194140 301514 194192 301520
rect 194048 297424 194100 297430
rect 194048 297366 194100 297372
rect 194048 291848 194100 291854
rect 194048 291790 194100 291796
rect 193954 282160 194010 282169
rect 193954 282095 194010 282104
rect 193864 249756 193916 249762
rect 193864 249698 193916 249704
rect 193968 241466 193996 282095
rect 194060 274582 194088 291790
rect 194152 282130 194180 301514
rect 194140 282124 194192 282130
rect 194140 282066 194192 282072
rect 194520 279313 194548 325666
rect 195256 325038 195284 341498
rect 195244 325032 195296 325038
rect 195244 324974 195296 324980
rect 195244 319524 195296 319530
rect 195244 319466 195296 319472
rect 194506 279304 194562 279313
rect 194506 279239 194562 279248
rect 194048 274576 194100 274582
rect 194048 274518 194100 274524
rect 195152 270564 195204 270570
rect 195152 270506 195204 270512
rect 195164 269822 195192 270506
rect 195152 269816 195204 269822
rect 195152 269758 195204 269764
rect 194416 258732 194468 258738
rect 194416 258674 194468 258680
rect 194048 251932 194100 251938
rect 194048 251874 194100 251880
rect 193956 241460 194008 241466
rect 193956 241402 194008 241408
rect 194060 226234 194088 251874
rect 194324 240780 194376 240786
rect 194324 240722 194376 240728
rect 194336 234297 194364 240722
rect 194322 234288 194378 234297
rect 194322 234223 194378 234232
rect 194048 226228 194100 226234
rect 194048 226170 194100 226176
rect 193128 220720 193180 220726
rect 193128 220662 193180 220668
rect 193140 220114 193168 220662
rect 193128 220108 193180 220114
rect 193128 220050 193180 220056
rect 192668 217932 192720 217938
rect 192668 217874 192720 217880
rect 192680 216714 192708 217874
rect 192668 216708 192720 216714
rect 192668 216650 192720 216656
rect 194428 202162 194456 258674
rect 194508 249756 194560 249762
rect 194508 249698 194560 249704
rect 194520 248742 194548 249698
rect 194508 248736 194560 248742
rect 194508 248678 194560 248684
rect 194416 202156 194468 202162
rect 194416 202098 194468 202104
rect 192574 200832 192630 200841
rect 192574 200767 192630 200776
rect 192668 195356 192720 195362
rect 192668 195298 192720 195304
rect 192576 191208 192628 191214
rect 192576 191150 192628 191156
rect 192484 191140 192536 191146
rect 192484 191082 192536 191088
rect 192482 183696 192538 183705
rect 192482 183631 192538 183640
rect 192496 158642 192524 183631
rect 192484 158636 192536 158642
rect 192484 158578 192536 158584
rect 192588 146946 192616 191150
rect 192680 177313 192708 195298
rect 194520 178809 194548 248678
rect 195256 238066 195284 319466
rect 195808 300937 195836 470698
rect 195900 376009 195928 563110
rect 197084 560380 197136 560386
rect 197084 560322 197136 560328
rect 196622 542600 196678 542609
rect 196622 542535 196678 542544
rect 196636 387025 196664 542535
rect 196622 387016 196678 387025
rect 196622 386951 196678 386960
rect 196624 384328 196676 384334
rect 196624 384270 196676 384276
rect 195886 376000 195942 376009
rect 195886 375935 195942 375944
rect 196636 374785 196664 384270
rect 197096 377534 197124 560322
rect 197084 377528 197136 377534
rect 197084 377470 197136 377476
rect 196808 375284 196860 375290
rect 196808 375226 196860 375232
rect 196622 374776 196678 374785
rect 196622 374711 196678 374720
rect 196624 367124 196676 367130
rect 196624 367066 196676 367072
rect 195888 355360 195940 355366
rect 195888 355302 195940 355308
rect 195900 354754 195928 355302
rect 195888 354748 195940 354754
rect 195888 354690 195940 354696
rect 195794 300928 195850 300937
rect 195794 300863 195850 300872
rect 195796 298852 195848 298858
rect 195796 298794 195848 298800
rect 195426 284336 195482 284345
rect 195426 284271 195482 284280
rect 195334 267336 195390 267345
rect 195334 267271 195390 267280
rect 195348 266422 195376 267271
rect 195336 266416 195388 266422
rect 195336 266358 195388 266364
rect 195336 264988 195388 264994
rect 195336 264930 195388 264936
rect 195348 242865 195376 264930
rect 195334 242856 195390 242865
rect 195334 242791 195390 242800
rect 195244 238060 195296 238066
rect 195244 238002 195296 238008
rect 195334 232656 195390 232665
rect 195334 232591 195390 232600
rect 195242 225720 195298 225729
rect 195242 225655 195298 225664
rect 195152 225004 195204 225010
rect 195152 224946 195204 224952
rect 195164 219434 195192 224946
rect 195256 224942 195284 225655
rect 195348 225593 195376 232591
rect 195334 225584 195390 225593
rect 195334 225519 195390 225528
rect 195244 224936 195296 224942
rect 195244 224878 195296 224884
rect 195164 219406 195284 219434
rect 195150 215928 195206 215937
rect 195150 215863 195206 215872
rect 195164 213761 195192 215863
rect 195150 213752 195206 213761
rect 195150 213687 195206 213696
rect 194506 178800 194562 178809
rect 194506 178735 194562 178744
rect 192666 177304 192722 177313
rect 192666 177239 192722 177248
rect 193954 152416 194010 152425
rect 193954 152351 194010 152360
rect 192484 146940 192536 146946
rect 192484 146882 192536 146888
rect 192576 146940 192628 146946
rect 192576 146882 192628 146888
rect 191288 104984 191340 104990
rect 191288 104926 191340 104932
rect 191194 91080 191250 91089
rect 191194 91015 191250 91024
rect 191300 56574 191328 104926
rect 191288 56568 191340 56574
rect 191288 56510 191340 56516
rect 192496 35290 192524 146882
rect 192576 134564 192628 134570
rect 192576 134506 192628 134512
rect 192588 89729 192616 134506
rect 193864 125724 193916 125730
rect 193864 125666 193916 125672
rect 192574 89720 192630 89729
rect 192574 89655 192630 89664
rect 193876 66162 193904 125666
rect 193968 119513 193996 152351
rect 193954 119504 194010 119513
rect 193954 119439 194010 119448
rect 193956 113212 194008 113218
rect 193956 113154 194008 113160
rect 193968 85542 193996 113154
rect 193956 85536 194008 85542
rect 193956 85478 194008 85484
rect 193864 66156 193916 66162
rect 193864 66098 193916 66104
rect 192484 35284 192536 35290
rect 192484 35226 192536 35232
rect 191102 4856 191158 4865
rect 191102 4791 191158 4800
rect 195256 3466 195284 219406
rect 195334 207224 195390 207233
rect 195334 207159 195390 207168
rect 195348 11665 195376 207159
rect 195440 187649 195468 284271
rect 195808 251870 195836 298794
rect 195900 282878 195928 354690
rect 195888 282872 195940 282878
rect 195888 282814 195940 282820
rect 196636 280158 196664 367066
rect 196714 356960 196770 356969
rect 196714 356895 196770 356904
rect 196728 292641 196756 356895
rect 196820 348430 196848 375226
rect 197188 365702 197216 567190
rect 197280 443714 197308 702646
rect 218992 700330 219020 703520
rect 233884 702772 233936 702778
rect 233884 702714 233936 702720
rect 218980 700324 219032 700330
rect 218980 700266 219032 700272
rect 204260 590708 204312 590714
rect 204260 590650 204312 590656
rect 198832 558204 198884 558210
rect 198832 558146 198884 558152
rect 198556 554056 198608 554062
rect 198556 553998 198608 554004
rect 198096 537532 198148 537538
rect 198096 537474 198148 537480
rect 198002 535528 198058 535537
rect 198002 535463 198058 535472
rect 197360 532704 197412 532710
rect 197360 532646 197412 532652
rect 197372 532273 197400 532646
rect 197358 532264 197414 532273
rect 197358 532199 197414 532208
rect 197360 529916 197412 529922
rect 197360 529858 197412 529864
rect 197372 529825 197400 529858
rect 197358 529816 197414 529825
rect 197358 529751 197414 529760
rect 197360 528556 197412 528562
rect 197360 528498 197412 528504
rect 197372 527377 197400 528498
rect 197358 527368 197414 527377
rect 197358 527303 197414 527312
rect 198016 525094 198044 535463
rect 198004 525088 198056 525094
rect 198004 525030 198056 525036
rect 197450 524784 197506 524793
rect 197450 524719 197506 524728
rect 197358 522336 197414 522345
rect 197464 522306 197492 524719
rect 197358 522271 197414 522280
rect 197452 522300 197504 522306
rect 197372 521694 197400 522271
rect 197452 522242 197504 522248
rect 197360 521688 197412 521694
rect 197360 521630 197412 521636
rect 197358 519888 197414 519897
rect 197358 519823 197414 519832
rect 197372 518974 197400 519823
rect 197360 518968 197412 518974
rect 197360 518910 197412 518916
rect 197358 517440 197414 517449
rect 197358 517375 197414 517384
rect 197372 516186 197400 517375
rect 197360 516180 197412 516186
rect 197360 516122 197412 516128
rect 197360 510604 197412 510610
rect 197360 510546 197412 510552
rect 197372 510241 197400 510546
rect 197358 510232 197414 510241
rect 197358 510167 197414 510176
rect 197358 507648 197414 507657
rect 197358 507583 197414 507592
rect 197372 506530 197400 507583
rect 197360 506524 197412 506530
rect 197360 506466 197412 506472
rect 197360 500948 197412 500954
rect 197360 500890 197412 500896
rect 197372 500449 197400 500890
rect 197358 500440 197414 500449
rect 197358 500375 197414 500384
rect 197358 495544 197414 495553
rect 197358 495479 197360 495488
rect 197412 495479 197414 495488
rect 197360 495450 197412 495456
rect 197358 492960 197414 492969
rect 197358 492895 197414 492904
rect 197372 492726 197400 492895
rect 197360 492720 197412 492726
rect 197360 492662 197412 492668
rect 197358 490512 197414 490521
rect 197358 490447 197414 490456
rect 197372 489938 197400 490447
rect 197360 489932 197412 489938
rect 197360 489874 197412 489880
rect 197358 488064 197414 488073
rect 197358 487999 197414 488008
rect 197372 487218 197400 487999
rect 197360 487212 197412 487218
rect 197360 487154 197412 487160
rect 198002 483168 198058 483177
rect 198002 483103 198058 483112
rect 197358 480720 197414 480729
rect 197358 480655 197414 480664
rect 197372 480486 197400 480655
rect 197360 480480 197412 480486
rect 197360 480422 197412 480428
rect 197358 478272 197414 478281
rect 197358 478207 197414 478216
rect 197372 477562 197400 478207
rect 197360 477556 197412 477562
rect 197360 477498 197412 477504
rect 197358 475824 197414 475833
rect 197358 475759 197414 475768
rect 197372 474774 197400 475759
rect 197360 474768 197412 474774
rect 197360 474710 197412 474716
rect 197360 473408 197412 473414
rect 197358 473376 197360 473385
rect 197412 473376 197414 473385
rect 197358 473311 197414 473320
rect 197634 470928 197690 470937
rect 197634 470863 197690 470872
rect 197648 470762 197676 470863
rect 197636 470756 197688 470762
rect 197636 470698 197688 470704
rect 197358 468480 197414 468489
rect 197358 468415 197414 468424
rect 197372 467906 197400 468415
rect 197360 467900 197412 467906
rect 197360 467842 197412 467848
rect 197358 466032 197414 466041
rect 197358 465967 197414 465976
rect 197372 465118 197400 465967
rect 197360 465112 197412 465118
rect 197360 465054 197412 465060
rect 197358 463312 197414 463321
rect 197358 463247 197414 463256
rect 197372 462398 197400 463247
rect 197360 462392 197412 462398
rect 197360 462334 197412 462340
rect 197358 460864 197414 460873
rect 197358 460799 197414 460808
rect 197372 460222 197400 460799
rect 197360 460216 197412 460222
rect 197360 460158 197412 460164
rect 197358 458416 197414 458425
rect 197358 458351 197414 458360
rect 197372 458250 197400 458351
rect 197360 458244 197412 458250
rect 197360 458186 197412 458192
rect 197358 448624 197414 448633
rect 197358 448559 197360 448568
rect 197412 448559 197414 448568
rect 197360 448530 197412 448536
rect 197358 446176 197414 446185
rect 197358 446111 197414 446120
rect 197372 445806 197400 446111
rect 197360 445800 197412 445806
rect 197360 445742 197412 445748
rect 197358 443728 197414 443737
rect 197280 443686 197358 443714
rect 197358 443663 197360 443672
rect 197412 443663 197414 443672
rect 197360 443634 197412 443640
rect 197360 441584 197412 441590
rect 197360 441526 197412 441532
rect 197372 441425 197400 441526
rect 197358 441416 197414 441425
rect 197358 441351 197414 441360
rect 197358 433936 197414 433945
rect 197358 433871 197414 433880
rect 197372 433362 197400 433871
rect 197360 433356 197412 433362
rect 197360 433298 197412 433304
rect 197358 429040 197414 429049
rect 197358 428975 197414 428984
rect 197372 427854 197400 428975
rect 197360 427848 197412 427854
rect 197360 427790 197412 427796
rect 197358 426592 197414 426601
rect 197358 426527 197414 426536
rect 197372 426494 197400 426527
rect 197360 426488 197412 426494
rect 197360 426430 197412 426436
rect 197358 424144 197414 424153
rect 197358 424079 197414 424088
rect 197372 423706 197400 424079
rect 197360 423700 197412 423706
rect 197360 423642 197412 423648
rect 197358 419248 197414 419257
rect 197358 419183 197414 419192
rect 197372 418198 197400 419183
rect 197360 418192 197412 418198
rect 197360 418134 197412 418140
rect 197358 414352 197414 414361
rect 197358 414287 197414 414296
rect 197372 414050 197400 414287
rect 197360 414044 197412 414050
rect 197360 413986 197412 413992
rect 197358 411904 197414 411913
rect 197358 411839 197414 411848
rect 197372 411330 197400 411839
rect 197360 411324 197412 411330
rect 197360 411266 197412 411272
rect 197360 409828 197412 409834
rect 197360 409770 197412 409776
rect 197372 409601 197400 409770
rect 197358 409592 197414 409601
rect 197358 409527 197414 409536
rect 197358 407008 197414 407017
rect 197358 406943 197414 406952
rect 197372 405754 197400 406943
rect 197360 405748 197412 405754
rect 197360 405690 197412 405696
rect 197358 402112 197414 402121
rect 197358 402047 197414 402056
rect 197372 401674 197400 402047
rect 197360 401668 197412 401674
rect 197360 401610 197412 401616
rect 197358 399664 197414 399673
rect 197358 399599 197414 399608
rect 197372 398886 197400 399599
rect 197360 398880 197412 398886
rect 197360 398822 197412 398828
rect 197358 397216 197414 397225
rect 197358 397151 197414 397160
rect 197372 396098 197400 397151
rect 197360 396092 197412 396098
rect 197360 396034 197412 396040
rect 197358 394768 197414 394777
rect 197358 394703 197360 394712
rect 197412 394703 197414 394712
rect 197360 394674 197412 394680
rect 197358 392320 197414 392329
rect 197358 392255 197414 392264
rect 197372 392018 197400 392255
rect 197360 392012 197412 392018
rect 197360 391954 197412 391960
rect 197358 387424 197414 387433
rect 197358 387359 197414 387368
rect 197372 386442 197400 387359
rect 197360 386436 197412 386442
rect 197360 386378 197412 386384
rect 197266 384976 197322 384985
rect 197266 384911 197322 384920
rect 197280 372570 197308 384911
rect 197358 380080 197414 380089
rect 197358 380015 197414 380024
rect 197372 379574 197400 380015
rect 197360 379568 197412 379574
rect 197360 379510 197412 379516
rect 197268 372564 197320 372570
rect 197268 372506 197320 372512
rect 197176 365696 197228 365702
rect 197176 365638 197228 365644
rect 196808 348424 196860 348430
rect 196808 348366 196860 348372
rect 196808 338156 196860 338162
rect 196808 338098 196860 338104
rect 196714 292632 196770 292641
rect 196714 292567 196770 292576
rect 196716 280492 196768 280498
rect 196716 280434 196768 280440
rect 196624 280152 196676 280158
rect 196624 280094 196676 280100
rect 196728 269890 196756 280434
rect 196820 278730 196848 338098
rect 198016 325689 198044 483103
rect 198108 476814 198136 537474
rect 198568 529825 198596 553998
rect 198648 551336 198700 551342
rect 198648 551278 198700 551284
rect 198554 529816 198610 529825
rect 198554 529751 198610 529760
rect 198660 500449 198688 551278
rect 198740 535628 198792 535634
rect 198740 535570 198792 535576
rect 198752 530641 198780 535570
rect 198738 530632 198794 530641
rect 198738 530567 198794 530576
rect 198646 500440 198702 500449
rect 198646 500375 198702 500384
rect 198096 476808 198148 476814
rect 198096 476750 198148 476756
rect 198844 463321 198872 558146
rect 204272 556850 204300 590650
rect 213920 568608 213972 568614
rect 213920 568550 213972 568556
rect 209044 567316 209096 567322
rect 209044 567258 209096 567264
rect 206284 563100 206336 563106
rect 206284 563042 206336 563048
rect 204260 556844 204312 556850
rect 204260 556786 204312 556792
rect 204272 541686 204300 556786
rect 206296 545465 206324 563042
rect 205638 545456 205694 545465
rect 205638 545391 205694 545400
rect 206282 545456 206338 545465
rect 206282 545391 206338 545400
rect 199476 541680 199528 541686
rect 199476 541622 199528 541628
rect 204260 541680 204312 541686
rect 204260 541622 204312 541628
rect 199384 538348 199436 538354
rect 199384 538290 199436 538296
rect 199106 505200 199162 505209
rect 199106 505135 199162 505144
rect 198830 463312 198886 463321
rect 198830 463247 198886 463256
rect 198830 458416 198886 458425
rect 198830 458351 198886 458360
rect 198646 455968 198702 455977
rect 198646 455903 198702 455912
rect 198554 453520 198610 453529
rect 198554 453455 198610 453464
rect 198462 393408 198518 393417
rect 198462 393343 198464 393352
rect 198516 393343 198518 393352
rect 198464 393314 198516 393320
rect 198462 392320 198518 392329
rect 198462 392255 198518 392264
rect 198002 325680 198058 325689
rect 198002 325615 198058 325624
rect 197176 307080 197228 307086
rect 197176 307022 197228 307028
rect 197188 299538 197216 307022
rect 197176 299532 197228 299538
rect 197176 299474 197228 299480
rect 197188 282985 197216 299474
rect 198016 296714 198044 325615
rect 198372 296744 198424 296750
rect 198016 296692 198372 296714
rect 198016 296686 198424 296692
rect 197174 282976 197230 282985
rect 197174 282911 197230 282920
rect 197268 282940 197320 282946
rect 197268 282882 197320 282888
rect 197280 280498 197308 282882
rect 198004 282872 198056 282878
rect 198004 282814 198056 282820
rect 197360 282804 197412 282810
rect 197360 282746 197412 282752
rect 197372 282441 197400 282746
rect 197358 282432 197414 282441
rect 197358 282367 197414 282376
rect 198016 281625 198044 282814
rect 198002 281616 198058 281625
rect 198002 281551 198058 281560
rect 197360 281512 197412 281518
rect 197360 281454 197412 281460
rect 197372 280809 197400 281454
rect 197358 280800 197414 280809
rect 197358 280735 197414 280744
rect 198278 280528 198334 280537
rect 197268 280492 197320 280498
rect 198278 280463 198280 280472
rect 197268 280434 197320 280440
rect 198332 280463 198334 280472
rect 198280 280434 198332 280440
rect 197358 279576 197414 279585
rect 197358 279511 197414 279520
rect 197372 278798 197400 279511
rect 197360 278792 197412 278798
rect 197360 278734 197412 278740
rect 196808 278724 196860 278730
rect 196808 278666 196860 278672
rect 197268 278724 197320 278730
rect 197268 278666 197320 278672
rect 197280 278610 197308 278666
rect 197358 278624 197414 278633
rect 197280 278582 197358 278610
rect 197084 274576 197136 274582
rect 197084 274518 197136 274524
rect 196716 269884 196768 269890
rect 196716 269826 196768 269832
rect 196624 262880 196676 262886
rect 196624 262822 196676 262828
rect 196636 256834 196664 262822
rect 196624 256828 196676 256834
rect 196624 256770 196676 256776
rect 196622 253056 196678 253065
rect 196622 252991 196678 253000
rect 195796 251864 195848 251870
rect 195796 251806 195848 251812
rect 195704 249892 195756 249898
rect 195704 249834 195756 249840
rect 195716 247722 195744 249834
rect 195704 247716 195756 247722
rect 195704 247658 195756 247664
rect 195612 244316 195664 244322
rect 195612 244258 195664 244264
rect 195520 241528 195572 241534
rect 195520 241470 195572 241476
rect 195532 200054 195560 241470
rect 195624 235958 195652 244258
rect 196636 241602 196664 252991
rect 197096 246158 197124 274518
rect 197176 256828 197228 256834
rect 197176 256770 197228 256776
rect 197084 246152 197136 246158
rect 197084 246094 197136 246100
rect 197084 243568 197136 243574
rect 197084 243510 197136 243516
rect 197096 241641 197124 243510
rect 197082 241632 197138 241641
rect 195980 241596 196032 241602
rect 195980 241538 196032 241544
rect 196624 241596 196676 241602
rect 197082 241567 197138 241576
rect 196624 241538 196676 241544
rect 195992 240174 196020 241538
rect 196992 241460 197044 241466
rect 196992 241402 197044 241408
rect 197004 240961 197032 241402
rect 196990 240952 197046 240961
rect 196990 240887 197046 240896
rect 195980 240168 196032 240174
rect 195980 240110 196032 240116
rect 195612 235952 195664 235958
rect 195612 235894 195664 235900
rect 197004 229094 197032 240887
rect 197082 240816 197138 240825
rect 197082 240751 197138 240760
rect 197096 237386 197124 240751
rect 197084 237380 197136 237386
rect 197084 237322 197136 237328
rect 197004 229066 197124 229094
rect 196624 227044 196676 227050
rect 196624 226986 196676 226992
rect 195888 221468 195940 221474
rect 195888 221410 195940 221416
rect 195900 217938 195928 221410
rect 195888 217932 195940 217938
rect 195888 217874 195940 217880
rect 195520 200048 195572 200054
rect 195520 199990 195572 199996
rect 195532 191185 195560 199990
rect 195518 191176 195574 191185
rect 195518 191111 195574 191120
rect 195426 187640 195482 187649
rect 195426 187575 195482 187584
rect 195440 183161 195468 187575
rect 195426 183152 195482 183161
rect 195426 183087 195482 183096
rect 195426 177032 195482 177041
rect 195426 176967 195482 176976
rect 195440 160721 195468 176967
rect 195426 160712 195482 160721
rect 195426 160647 195482 160656
rect 195520 131164 195572 131170
rect 195520 131106 195572 131112
rect 195532 116618 195560 131106
rect 195520 116612 195572 116618
rect 195520 116554 195572 116560
rect 195428 116068 195480 116074
rect 195428 116010 195480 116016
rect 195440 93906 195468 116010
rect 195428 93900 195480 93906
rect 195428 93842 195480 93848
rect 195334 11656 195390 11665
rect 195334 11591 195390 11600
rect 196636 3505 196664 226986
rect 197096 199481 197124 229066
rect 197188 214606 197216 256770
rect 197176 214600 197228 214606
rect 197176 214542 197228 214548
rect 197082 199472 197138 199481
rect 197082 199407 197138 199416
rect 196808 191888 196860 191894
rect 196808 191830 196860 191836
rect 196714 183016 196770 183025
rect 196714 182951 196770 182960
rect 196728 101454 196756 182951
rect 196820 164150 196848 191830
rect 197280 176594 197308 278582
rect 197358 278559 197414 278568
rect 197360 277364 197412 277370
rect 197360 277306 197412 277312
rect 197372 277273 197400 277306
rect 197358 277264 197414 277273
rect 197358 277199 197414 277208
rect 197358 276720 197414 276729
rect 197358 276655 197360 276664
rect 197412 276655 197414 276664
rect 197360 276626 197412 276632
rect 197450 275904 197506 275913
rect 197450 275839 197506 275848
rect 197358 275088 197414 275097
rect 197358 275023 197414 275032
rect 197372 274718 197400 275023
rect 197464 274786 197492 275839
rect 197452 274780 197504 274786
rect 197452 274722 197504 274728
rect 197360 274712 197412 274718
rect 197360 274654 197412 274660
rect 197360 274576 197412 274582
rect 197358 274544 197360 274553
rect 197412 274544 197414 274553
rect 197358 274479 197414 274488
rect 197358 273728 197414 273737
rect 197358 273663 197414 273672
rect 197372 273358 197400 273663
rect 197360 273352 197412 273358
rect 197360 273294 197412 273300
rect 197360 273216 197412 273222
rect 197360 273158 197412 273164
rect 197372 272921 197400 273158
rect 197452 273148 197504 273154
rect 197452 273090 197504 273096
rect 197358 272912 197414 272921
rect 197358 272847 197414 272856
rect 197464 272377 197492 273090
rect 197450 272368 197506 272377
rect 197450 272303 197506 272312
rect 197358 271552 197414 271561
rect 197358 271487 197414 271496
rect 197372 270570 197400 271487
rect 198384 271017 198412 296686
rect 198370 271008 198426 271017
rect 198370 270943 198426 270952
rect 197360 270564 197412 270570
rect 197360 270506 197412 270512
rect 197360 269068 197412 269074
rect 197360 269010 197412 269016
rect 197372 268841 197400 269010
rect 197452 269000 197504 269006
rect 197452 268942 197504 268948
rect 197358 268832 197414 268841
rect 197358 268767 197414 268776
rect 197464 268025 197492 268942
rect 197450 268016 197506 268025
rect 197450 267951 197506 267960
rect 197360 267708 197412 267714
rect 197360 267650 197412 267656
rect 197372 266665 197400 267650
rect 197358 266656 197414 266665
rect 197358 266591 197414 266600
rect 197450 265296 197506 265305
rect 197450 265231 197506 265240
rect 197464 264994 197492 265231
rect 197452 264988 197504 264994
rect 197452 264930 197504 264936
rect 197360 264920 197412 264926
rect 197360 264862 197412 264868
rect 197372 264489 197400 264862
rect 197358 264480 197414 264489
rect 197358 264415 197414 264424
rect 197360 263696 197412 263702
rect 197358 263664 197360 263673
rect 197412 263664 197414 263673
rect 197358 263599 197414 263608
rect 197360 261520 197412 261526
rect 197358 261488 197360 261497
rect 197412 261488 197414 261497
rect 197358 261423 197414 261432
rect 197358 260128 197414 260137
rect 197358 260063 197414 260072
rect 197372 259486 197400 260063
rect 197360 259480 197412 259486
rect 197360 259422 197412 259428
rect 197452 259412 197504 259418
rect 197452 259354 197504 259360
rect 197358 259312 197414 259321
rect 197358 259247 197414 259256
rect 197372 258738 197400 259247
rect 197464 258777 197492 259354
rect 197450 258768 197506 258777
rect 197360 258732 197412 258738
rect 197450 258703 197506 258712
rect 197360 258674 197412 258680
rect 197450 257952 197506 257961
rect 197450 257887 197506 257896
rect 197464 256766 197492 257887
rect 198094 257408 198150 257417
rect 198094 257343 198150 257352
rect 198108 256834 198136 257343
rect 198096 256828 198148 256834
rect 198096 256770 198148 256776
rect 197452 256760 197504 256766
rect 197452 256702 197504 256708
rect 197360 256692 197412 256698
rect 197360 256634 197412 256640
rect 197372 255785 197400 256634
rect 197450 256592 197506 256601
rect 197450 256527 197506 256536
rect 197358 255776 197414 255785
rect 197358 255711 197414 255720
rect 197464 255338 197492 256527
rect 197452 255332 197504 255338
rect 197452 255274 197504 255280
rect 197360 255264 197412 255270
rect 197358 255232 197360 255241
rect 197412 255232 197414 255241
rect 197358 255167 197414 255176
rect 197358 253600 197414 253609
rect 197358 253535 197414 253544
rect 197372 252618 197400 253535
rect 197360 252612 197412 252618
rect 197360 252554 197412 252560
rect 197360 251864 197412 251870
rect 197360 251806 197412 251812
rect 198002 251832 198058 251841
rect 197372 251705 197400 251806
rect 198002 251767 198058 251776
rect 197358 251696 197414 251705
rect 197358 251631 197414 251640
rect 197910 250880 197966 250889
rect 197910 250815 197966 250824
rect 197358 250064 197414 250073
rect 197358 249999 197414 250008
rect 197372 249830 197400 249999
rect 197924 249898 197952 250815
rect 197912 249892 197964 249898
rect 197912 249834 197964 249840
rect 197360 249824 197412 249830
rect 197360 249766 197412 249772
rect 197358 249520 197414 249529
rect 197358 249455 197414 249464
rect 197372 248470 197400 249455
rect 197452 248736 197504 248742
rect 197450 248704 197452 248713
rect 197504 248704 197506 248713
rect 197450 248639 197506 248648
rect 197360 248464 197412 248470
rect 197360 248406 197412 248412
rect 197450 247888 197506 247897
rect 197450 247823 197506 247832
rect 197464 247110 197492 247823
rect 197452 247104 197504 247110
rect 197452 247046 197504 247052
rect 197360 247036 197412 247042
rect 197360 246978 197412 246984
rect 197372 245993 197400 246978
rect 197358 245984 197414 245993
rect 197358 245919 197414 245928
rect 197358 245168 197414 245177
rect 197358 245103 197414 245112
rect 197372 244934 197400 245103
rect 197360 244928 197412 244934
rect 197360 244870 197412 244876
rect 197360 244248 197412 244254
rect 197360 244190 197412 244196
rect 197372 243001 197400 244190
rect 198016 243817 198044 251767
rect 198476 244361 198504 392255
rect 198568 262313 198596 453455
rect 198660 263129 198688 455903
rect 198740 376848 198792 376854
rect 198740 376790 198792 376796
rect 198752 376038 198780 376790
rect 198740 376032 198792 376038
rect 198740 375974 198792 375980
rect 198740 374332 198792 374338
rect 198740 374274 198792 374280
rect 198752 271250 198780 374274
rect 198844 366489 198872 458351
rect 198922 416800 198978 416809
rect 198922 416735 198978 416744
rect 198936 374678 198964 416735
rect 199014 382528 199070 382537
rect 199014 382463 199070 382472
rect 198924 374672 198976 374678
rect 198924 374614 198976 374620
rect 199028 373386 199056 382463
rect 199120 376854 199148 505135
rect 199396 384849 199424 538290
rect 199488 512650 199516 541622
rect 205652 538214 205680 545391
rect 209056 542366 209084 567258
rect 212538 553480 212594 553489
rect 212538 553415 212594 553424
rect 209044 542360 209096 542366
rect 209044 542302 209096 542308
rect 210424 542360 210476 542366
rect 210424 542302 210476 542308
rect 207020 541680 207072 541686
rect 207020 541622 207072 541628
rect 205652 538186 205772 538214
rect 205744 535908 205772 538186
rect 207032 535922 207060 541622
rect 210436 535922 210464 542302
rect 207032 535894 207414 535922
rect 210436 535894 210910 535922
rect 212552 535908 212580 553415
rect 213458 538520 213514 538529
rect 213458 538455 213514 538464
rect 213472 538257 213500 538455
rect 213458 538248 213514 538257
rect 213458 538183 213514 538192
rect 213932 535922 213960 568550
rect 230478 556200 230534 556209
rect 230478 556135 230534 556144
rect 225326 552120 225382 552129
rect 225326 552055 225382 552064
rect 226984 552084 227036 552090
rect 215392 549364 215444 549370
rect 215392 549306 215444 549312
rect 215404 535922 215432 549306
rect 218702 548040 218758 548049
rect 218702 547975 218758 547984
rect 216586 538792 216642 538801
rect 216586 538727 216642 538736
rect 213932 535894 214222 535922
rect 215404 535894 215878 535922
rect 200408 535634 200790 535650
rect 200396 535628 200790 535634
rect 200448 535622 200790 535628
rect 200396 535570 200448 535576
rect 203706 535528 203762 535537
rect 201408 535492 201460 535498
rect 203762 535486 204102 535514
rect 208688 535498 209070 535514
rect 208676 535492 209070 535498
rect 203706 535463 203762 535472
rect 201408 535434 201460 535440
rect 208728 535486 209070 535492
rect 208676 535434 208728 535440
rect 201420 535401 201448 535434
rect 216600 535401 216628 538727
rect 217138 538520 217194 538529
rect 217138 538455 217194 538464
rect 216680 538280 216732 538286
rect 216678 538248 216680 538257
rect 216732 538248 216734 538257
rect 216678 538183 216734 538192
rect 217152 535922 217180 538455
rect 218716 535922 218744 547975
rect 220820 545216 220872 545222
rect 220820 545158 220872 545164
rect 217152 535894 217534 535922
rect 218716 535894 219190 535922
rect 220832 535908 220860 545158
rect 223672 543856 223724 543862
rect 223672 543798 223724 543804
rect 222474 538384 222530 538393
rect 222474 538319 222530 538328
rect 220912 538280 220964 538286
rect 220912 538222 220964 538228
rect 220924 537538 220952 538222
rect 220912 537532 220964 537538
rect 220912 537474 220964 537480
rect 222488 535908 222516 538319
rect 223684 535922 223712 543798
rect 225340 535922 225368 552055
rect 226984 552026 227036 552032
rect 226996 535922 227024 552026
rect 229100 550656 229152 550662
rect 229100 550598 229152 550604
rect 223684 535894 224158 535922
rect 225340 535894 225814 535922
rect 226996 535894 227470 535922
rect 229112 535908 229140 550598
rect 230492 535922 230520 556135
rect 231950 549536 232006 549545
rect 231950 549471 232006 549480
rect 231964 535922 231992 549471
rect 233896 536858 233924 702714
rect 235184 702574 235212 703520
rect 267660 702914 267688 703520
rect 281540 702976 281592 702982
rect 281540 702918 281592 702924
rect 267648 702908 267700 702914
rect 267648 702850 267700 702856
rect 276020 702908 276072 702914
rect 276020 702850 276072 702856
rect 273260 702840 273312 702846
rect 273260 702782 273312 702788
rect 235172 702568 235224 702574
rect 235172 702510 235224 702516
rect 264244 702568 264296 702574
rect 264244 702510 264296 702516
rect 255964 589348 256016 589354
rect 255964 589290 256016 589296
rect 241518 559056 241574 559065
rect 241518 558991 241574 559000
rect 237378 557560 237434 557569
rect 241532 557534 241560 558991
rect 241532 557506 241928 557534
rect 237378 557495 237434 557504
rect 235262 545320 235318 545329
rect 235262 545255 235318 545264
rect 233884 536852 233936 536858
rect 233884 536794 233936 536800
rect 234068 536852 234120 536858
rect 234068 536794 234120 536800
rect 230492 535894 230782 535922
rect 231964 535894 232438 535922
rect 234080 535908 234108 536794
rect 235276 535922 235304 545255
rect 235276 535894 235750 535922
rect 237392 535908 237420 557495
rect 240230 554840 240286 554849
rect 240230 554775 240286 554784
rect 238758 541376 238814 541385
rect 238758 541311 238814 541320
rect 238772 535922 238800 541311
rect 240244 535922 240272 554775
rect 241900 535922 241928 557506
rect 251824 556232 251876 556238
rect 251824 556174 251876 556180
rect 244924 554804 244976 554810
rect 244924 554746 244976 554752
rect 243542 547904 243598 547913
rect 243542 547839 243598 547848
rect 243556 535922 243584 547839
rect 244936 542366 244964 554746
rect 245660 547188 245712 547194
rect 245660 547130 245712 547136
rect 244924 542360 244976 542366
rect 244924 542302 244976 542308
rect 238772 535894 239062 535922
rect 240244 535894 240718 535922
rect 241900 535894 242374 535922
rect 243556 535894 244030 535922
rect 245672 535908 245700 547130
rect 248510 546680 248566 546689
rect 248510 546615 248566 546624
rect 247040 542360 247092 542366
rect 247040 542302 247092 542308
rect 247052 535922 247080 542302
rect 248524 535922 248552 546615
rect 250628 539640 250680 539646
rect 250628 539582 250680 539588
rect 247052 535894 247632 535922
rect 248524 535894 248998 535922
rect 250640 535908 250668 539582
rect 251836 535922 251864 556174
rect 253938 542600 253994 542609
rect 253938 542535 253994 542544
rect 251836 535894 252310 535922
rect 253952 535908 253980 542535
rect 255976 541657 256004 589290
rect 259460 564528 259512 564534
rect 259460 564470 259512 564476
rect 259472 557534 259500 564470
rect 264256 561678 264284 702510
rect 266360 571396 266412 571402
rect 266360 571338 266412 571344
rect 263600 561672 263652 561678
rect 263600 561614 263652 561620
rect 264244 561672 264296 561678
rect 264244 561614 264296 561620
rect 263612 560318 263640 561614
rect 263600 560312 263652 560318
rect 263600 560254 263652 560260
rect 259472 557506 260144 557534
rect 255962 541648 256018 541657
rect 255962 541583 256018 541592
rect 257342 541648 257398 541657
rect 257342 541583 257398 541592
rect 255596 538348 255648 538354
rect 255596 538290 255648 538296
rect 255608 535908 255636 538290
rect 257356 535922 257384 541583
rect 258448 541000 258500 541006
rect 258448 540942 258500 540948
rect 257278 535894 257384 535922
rect 258460 535922 258488 540942
rect 260116 535922 260144 557506
rect 262218 541240 262274 541249
rect 262218 541175 262274 541184
rect 258460 535894 258934 535922
rect 260116 535894 260590 535922
rect 262232 535908 262260 541175
rect 263612 535922 263640 560254
rect 266372 557534 266400 571338
rect 273272 567730 273300 702782
rect 273260 567724 273312 567730
rect 273260 567666 273312 567672
rect 273904 567724 273956 567730
rect 273904 567666 273956 567672
rect 273272 567254 273300 567666
rect 273260 567248 273312 567254
rect 273260 567190 273312 567196
rect 271880 563168 271932 563174
rect 271880 563110 271932 563116
rect 266372 557506 266768 557534
rect 265530 538248 265586 538257
rect 265530 538183 265586 538192
rect 263612 535894 263902 535922
rect 265544 535908 265572 538183
rect 266740 535922 266768 557506
rect 270500 553444 270552 553450
rect 270500 553386 270552 553392
rect 268566 546544 268622 546553
rect 268566 546479 268622 546488
rect 268580 535922 268608 546479
rect 270512 535922 270540 553386
rect 270866 543824 270922 543833
rect 270866 543759 270922 543768
rect 270880 539510 270908 543759
rect 270868 539504 270920 539510
rect 270868 539446 270920 539452
rect 271892 535922 271920 563110
rect 273916 539578 273944 567666
rect 273904 539572 273956 539578
rect 273904 539514 273956 539520
rect 275652 539572 275704 539578
rect 275652 539514 275704 539520
rect 273996 539504 274048 539510
rect 273996 539446 274048 539452
rect 266740 535894 267214 535922
rect 268580 535894 269054 535922
rect 270512 535894 270710 535922
rect 271892 535894 272366 535922
rect 274008 535908 274036 539446
rect 275664 535908 275692 539514
rect 247604 535498 247632 535894
rect 276032 535673 276060 702850
rect 281552 557534 281580 702918
rect 283852 700330 283880 703520
rect 300136 702642 300164 703520
rect 332520 703050 332548 703520
rect 331220 703044 331272 703050
rect 331220 702986 331272 702992
rect 332508 703044 332560 703050
rect 332508 702986 332560 702992
rect 300124 702636 300176 702642
rect 300124 702578 300176 702584
rect 300768 702636 300820 702642
rect 300768 702578 300820 702584
rect 300780 700330 300808 702578
rect 283840 700324 283892 700330
rect 283840 700266 283892 700272
rect 295340 700324 295392 700330
rect 295340 700266 295392 700272
rect 300768 700324 300820 700330
rect 300768 700266 300820 700272
rect 295352 594862 295380 700266
rect 327724 698964 327776 698970
rect 327724 698906 327776 698912
rect 295340 594856 295392 594862
rect 295340 594798 295392 594804
rect 295984 594856 296036 594862
rect 295984 594798 296036 594804
rect 291200 565888 291252 565894
rect 291200 565830 291252 565836
rect 288440 560380 288492 560386
rect 288440 560322 288492 560328
rect 287060 559020 287112 559026
rect 287060 558962 287112 558968
rect 281552 557506 281856 557534
rect 278042 549400 278098 549409
rect 278042 549335 278098 549344
rect 278056 539578 278084 549335
rect 280618 539744 280674 539753
rect 280618 539679 280674 539688
rect 278044 539572 278096 539578
rect 278044 539514 278096 539520
rect 278964 539572 279016 539578
rect 278964 539514 279016 539520
rect 278976 535908 279004 539514
rect 280632 535908 280660 539679
rect 281828 535922 281856 557506
rect 285128 548004 285180 548010
rect 285128 547946 285180 547952
rect 284300 543788 284352 543794
rect 284300 543730 284352 543736
rect 284312 543017 284340 543730
rect 284298 543008 284354 543017
rect 284298 542943 284354 542952
rect 283470 542464 283526 542473
rect 283470 542399 283526 542408
rect 283484 535922 283512 542399
rect 285140 535922 285168 547946
rect 287072 535922 287100 558962
rect 288452 535922 288480 560322
rect 291212 557534 291240 565830
rect 291212 557506 291792 557534
rect 290096 545148 290148 545154
rect 290096 545090 290148 545096
rect 290108 535922 290136 545090
rect 291764 535922 291792 557506
rect 295996 549914 296024 594798
rect 298100 564460 298152 564466
rect 298100 564402 298152 564408
rect 298112 557534 298140 564402
rect 309140 558952 309192 558958
rect 309140 558894 309192 558900
rect 309152 557534 309180 558894
rect 298112 557506 298416 557534
rect 309152 557506 310008 557534
rect 296720 552152 296772 552158
rect 296720 552094 296772 552100
rect 295984 549908 296036 549914
rect 295984 549850 296036 549856
rect 295522 539744 295578 539753
rect 295522 539679 295578 539688
rect 293866 537160 293922 537169
rect 293866 537095 293922 537104
rect 281828 535894 282302 535922
rect 283484 535894 283958 535922
rect 285140 535894 285614 535922
rect 287072 535894 287270 535922
rect 288452 535894 288926 535922
rect 290108 535894 290582 535922
rect 291764 535894 292238 535922
rect 293880 535908 293908 537095
rect 295536 535908 295564 539679
rect 296732 535922 296760 552094
rect 298388 535922 298416 557506
rect 303618 550760 303674 550769
rect 303618 550695 303674 550704
rect 300030 545184 300086 545193
rect 300030 545119 300086 545128
rect 300044 535922 300072 545119
rect 302146 537160 302202 537169
rect 302146 537095 302202 537104
rect 296732 535894 297206 535922
rect 298388 535894 298862 535922
rect 300044 535894 300518 535922
rect 302160 535908 302188 537095
rect 303632 535922 303660 550695
rect 305000 549296 305052 549302
rect 305000 549238 305052 549244
rect 305012 535922 305040 549238
rect 306656 542496 306708 542502
rect 306656 542438 306708 542444
rect 306668 535922 306696 542438
rect 309980 535922 310008 557506
rect 327736 555286 327764 698906
rect 331232 558210 331260 702986
rect 348804 698970 348832 703520
rect 349804 702840 349856 702846
rect 349804 702782 349856 702788
rect 348792 698964 348844 698970
rect 348792 698906 348844 698912
rect 349816 598942 349844 702782
rect 364996 702710 365024 703520
rect 397472 702794 397500 703520
rect 397380 702778 397500 702794
rect 397368 702772 397500 702778
rect 397420 702766 397500 702772
rect 397368 702714 397420 702720
rect 364984 702704 365036 702710
rect 364984 702646 365036 702652
rect 382924 702704 382976 702710
rect 382924 702646 382976 702652
rect 363604 702636 363656 702642
rect 363604 702578 363656 702584
rect 360200 700324 360252 700330
rect 360200 700266 360252 700272
rect 349160 598936 349212 598942
rect 349160 598878 349212 598884
rect 349804 598936 349856 598942
rect 349804 598878 349856 598884
rect 349172 597582 349200 598878
rect 349160 597576 349212 597582
rect 349160 597518 349212 597524
rect 331220 558204 331272 558210
rect 331220 558146 331272 558152
rect 324320 555280 324372 555286
rect 324320 555222 324372 555228
rect 324872 555280 324924 555286
rect 324872 555222 324924 555228
rect 327724 555280 327776 555286
rect 327724 555222 327776 555228
rect 324332 554878 324360 555222
rect 324320 554872 324372 554878
rect 324320 554814 324372 554820
rect 320178 545184 320234 545193
rect 320178 545119 320234 545128
rect 311900 543788 311952 543794
rect 311900 543730 311952 543736
rect 311912 535922 311940 543730
rect 316592 541000 316644 541006
rect 316592 540942 316644 540948
rect 316604 535922 316632 540942
rect 318706 538248 318762 538257
rect 318706 538183 318762 538192
rect 303632 535894 303830 535922
rect 305012 535894 305486 535922
rect 306668 535894 307142 535922
rect 309980 535894 310454 535922
rect 311912 535894 312110 535922
rect 316604 535894 317078 535922
rect 318720 535908 318748 538183
rect 320192 535922 320220 545119
rect 321558 543960 321614 543969
rect 321558 543895 321614 543904
rect 321572 535922 321600 543895
rect 323582 541104 323638 541113
rect 323582 541039 323638 541048
rect 323596 538214 323624 541039
rect 323596 538186 323716 538214
rect 323688 537538 323716 538186
rect 323676 537532 323728 537538
rect 323676 537474 323728 537480
rect 320192 535894 320390 535922
rect 321572 535894 322046 535922
rect 323688 535908 323716 537474
rect 324884 535922 324912 555222
rect 343640 547936 343692 547942
rect 343640 547878 343692 547884
rect 339960 546508 340012 546514
rect 339960 546450 340012 546456
rect 328460 545148 328512 545154
rect 328460 545090 328512 545096
rect 328472 535922 328500 545090
rect 330024 543856 330076 543862
rect 330024 543798 330076 543804
rect 330036 535922 330064 543798
rect 338304 542496 338356 542502
rect 338304 542438 338356 542444
rect 331680 541068 331732 541074
rect 331680 541010 331732 541016
rect 331692 535922 331720 541010
rect 335450 537024 335506 537033
rect 335450 536959 335506 536968
rect 333794 536888 333850 536897
rect 333794 536823 333850 536832
rect 324884 535894 325358 535922
rect 328472 535894 328854 535922
rect 330036 535894 330510 535922
rect 331692 535894 332166 535922
rect 333808 535908 333836 536823
rect 335464 535908 335492 536959
rect 337108 536852 337160 536858
rect 337108 536794 337160 536800
rect 337120 535908 337148 536794
rect 338316 535922 338344 542438
rect 339972 535922 340000 546450
rect 342074 539608 342130 539617
rect 342074 539543 342130 539552
rect 338316 535894 338790 535922
rect 339972 535894 340446 535922
rect 342088 535908 342116 539543
rect 343652 538214 343680 547878
rect 348698 539880 348754 539889
rect 348698 539815 348754 539824
rect 347688 539640 347740 539646
rect 347688 539582 347740 539588
rect 345386 539472 345442 539481
rect 345386 539407 345442 539416
rect 343652 538186 343772 538214
rect 343744 535908 343772 538186
rect 345400 535908 345428 539407
rect 347700 538801 347728 539582
rect 347686 538792 347742 538801
rect 347686 538727 347742 538736
rect 347044 538348 347096 538354
rect 347044 538290 347096 538296
rect 347056 535908 347084 538290
rect 348712 535908 348740 539815
rect 349172 539481 349200 597518
rect 353300 569968 353352 569974
rect 353300 569910 353352 569916
rect 351920 549908 351972 549914
rect 351920 549850 351972 549856
rect 349158 539472 349214 539481
rect 349158 539407 349214 539416
rect 350354 538384 350410 538393
rect 350354 538319 350410 538328
rect 350368 535908 350396 538319
rect 351932 538214 351960 549850
rect 351932 538186 352052 538214
rect 352024 535908 352052 538186
rect 353312 535922 353340 569910
rect 358912 561740 358964 561746
rect 358912 561682 358964 561688
rect 357440 557592 357492 557598
rect 357440 557534 357492 557540
rect 356244 543788 356296 543794
rect 356244 543730 356296 543736
rect 356152 542428 356204 542434
rect 356152 542370 356204 542376
rect 355322 538248 355378 538257
rect 355322 538183 355378 538192
rect 353312 535894 353694 535922
rect 355336 535908 355364 538183
rect 313370 535800 313426 535809
rect 313426 535758 313766 535786
rect 313370 535735 313426 535744
rect 276018 535664 276074 535673
rect 276018 535599 276074 535608
rect 276938 535664 276994 535673
rect 276994 535622 277334 535650
rect 276938 535599 276994 535608
rect 308404 535560 308456 535566
rect 327448 535560 327500 535566
rect 315670 535528 315726 535537
rect 308456 535508 308798 535514
rect 308404 535502 308798 535508
rect 247592 535492 247644 535498
rect 308416 535486 308798 535502
rect 315422 535486 315670 535514
rect 327198 535508 327448 535514
rect 327198 535502 327500 535508
rect 327198 535486 327488 535502
rect 315670 535463 315726 535472
rect 247592 535434 247644 535440
rect 201406 535392 201462 535401
rect 216586 535392 216642 535401
rect 201406 535327 201462 535336
rect 202064 535350 202446 535378
rect 202064 535294 202092 535350
rect 216586 535327 216642 535336
rect 202052 535288 202104 535294
rect 202052 535230 202104 535236
rect 199842 534984 199898 534993
rect 199842 534919 199898 534928
rect 199856 534041 199884 534919
rect 199842 534032 199898 534041
rect 199842 533967 199898 533976
rect 199476 512644 199528 512650
rect 199476 512586 199528 512592
rect 356164 497162 356192 542370
rect 356256 497434 356284 543730
rect 356336 538280 356388 538286
rect 356336 538222 356388 538228
rect 356348 499574 356376 538222
rect 357452 522345 357480 557534
rect 357622 543008 357678 543017
rect 357622 542943 357678 542952
rect 357532 539708 357584 539714
rect 357532 539650 357584 539656
rect 357438 522336 357494 522345
rect 357438 522271 357494 522280
rect 357544 512689 357572 539650
rect 357636 534721 357664 542943
rect 357622 534712 357678 534721
rect 357622 534647 357678 534656
rect 358726 532128 358782 532137
rect 358726 532063 358782 532072
rect 358740 532030 358768 532063
rect 358924 532030 358952 561682
rect 359096 538348 359148 538354
rect 359096 538290 359148 538296
rect 358728 532024 358780 532030
rect 358728 531966 358780 531972
rect 358912 532024 358964 532030
rect 358912 531966 358964 531972
rect 358910 529680 358966 529689
rect 358910 529615 358966 529624
rect 358726 527232 358782 527241
rect 358726 527167 358728 527176
rect 358780 527167 358782 527176
rect 358728 527138 358780 527144
rect 358726 524784 358782 524793
rect 358726 524719 358782 524728
rect 358740 524482 358768 524719
rect 358728 524476 358780 524482
rect 358728 524418 358780 524424
rect 358726 522336 358782 522345
rect 358726 522271 358728 522280
rect 358780 522271 358782 522280
rect 358728 522242 358780 522248
rect 357900 520056 357952 520062
rect 357898 520024 357900 520033
rect 357952 520024 357954 520033
rect 357898 519959 357954 519968
rect 358726 517440 358782 517449
rect 358726 517375 358782 517384
rect 358740 516186 358768 517375
rect 358728 516180 358780 516186
rect 358728 516122 358780 516128
rect 358634 514992 358690 515001
rect 358634 514927 358690 514936
rect 358648 514826 358676 514927
rect 358636 514820 358688 514826
rect 358636 514762 358688 514768
rect 357530 512680 357586 512689
rect 357530 512615 357586 512624
rect 357622 510096 357678 510105
rect 357622 510031 357678 510040
rect 357636 505782 357664 510031
rect 357624 505776 357676 505782
rect 357624 505718 357676 505724
rect 358726 505200 358782 505209
rect 358726 505135 358728 505144
rect 358780 505135 358782 505144
rect 358728 505106 358780 505112
rect 358726 502752 358782 502761
rect 358726 502687 358782 502696
rect 358740 502382 358768 502687
rect 358728 502376 358780 502382
rect 358728 502318 358780 502324
rect 358726 500304 358782 500313
rect 358726 500239 358782 500248
rect 358740 499594 358768 500239
rect 358728 499588 358780 499594
rect 356348 499546 356652 499574
rect 356256 497406 356560 497434
rect 356164 497134 356376 497162
rect 356348 496806 356376 497134
rect 356336 496800 356388 496806
rect 356336 496742 356388 496748
rect 356242 492688 356298 492697
rect 356164 492646 356242 492674
rect 199382 384840 199438 384849
rect 199382 384775 199438 384784
rect 199842 378448 199898 378457
rect 199842 378383 199898 378392
rect 199856 377233 199884 378383
rect 204442 377632 204498 377641
rect 199842 377224 199898 377233
rect 199842 377159 199898 377168
rect 199108 376848 199160 376854
rect 199108 376790 199160 376796
rect 200040 374338 200068 377604
rect 201512 377590 201710 377618
rect 202892 377590 203366 377618
rect 201406 377224 201462 377233
rect 201406 377159 201462 377168
rect 200302 375320 200358 375329
rect 200302 375255 200358 375264
rect 200316 374785 200344 375255
rect 200302 374776 200358 374785
rect 200302 374711 200358 374720
rect 200028 374332 200080 374338
rect 200028 374274 200080 374280
rect 200118 373416 200174 373425
rect 199016 373380 199068 373386
rect 200118 373351 200174 373360
rect 199016 373322 199068 373328
rect 198830 366480 198886 366489
rect 198830 366415 198886 366424
rect 198832 365696 198884 365702
rect 198832 365638 198884 365644
rect 198844 296721 198872 365638
rect 200132 364410 200160 373351
rect 200120 364404 200172 364410
rect 200120 364346 200172 364352
rect 199382 353560 199438 353569
rect 199382 353495 199438 353504
rect 199396 353394 199424 353495
rect 199384 353388 199436 353394
rect 199384 353330 199436 353336
rect 199396 315382 199424 353330
rect 199476 316736 199528 316742
rect 199476 316678 199528 316684
rect 199384 315376 199436 315382
rect 199384 315318 199436 315324
rect 198830 296712 198886 296721
rect 198830 296647 198886 296656
rect 198844 296041 198872 296647
rect 198830 296032 198886 296041
rect 198830 295967 198886 295976
rect 198832 285728 198884 285734
rect 198832 285670 198884 285676
rect 198844 284986 198872 285670
rect 198832 284980 198884 284986
rect 198832 284922 198884 284928
rect 198830 284608 198886 284617
rect 198830 284543 198886 284552
rect 198844 278118 198872 284543
rect 199488 282946 199516 316678
rect 200118 309768 200174 309777
rect 200118 309703 200174 309712
rect 200028 291848 200080 291854
rect 200028 291790 200080 291796
rect 199476 282940 199528 282946
rect 199476 282882 199528 282888
rect 199384 280152 199436 280158
rect 199384 280094 199436 280100
rect 198832 278112 198884 278118
rect 198832 278054 198884 278060
rect 198740 271244 198792 271250
rect 198740 271186 198792 271192
rect 199396 265849 199424 280094
rect 200040 275913 200068 291790
rect 200132 285326 200160 309703
rect 200120 285320 200172 285326
rect 200120 285262 200172 285268
rect 200316 284889 200344 374711
rect 201420 356726 201448 377159
rect 201408 356720 201460 356726
rect 201408 356662 201460 356668
rect 201408 338768 201460 338774
rect 201406 338736 201408 338745
rect 201460 338736 201462 338745
rect 201406 338671 201462 338680
rect 200764 312656 200816 312662
rect 200764 312598 200816 312604
rect 200776 309777 200804 312598
rect 200762 309768 200818 309777
rect 200762 309703 200818 309712
rect 201420 298110 201448 338671
rect 201512 298790 201540 377590
rect 201592 377528 201644 377534
rect 201592 377470 201644 377476
rect 201604 347818 201632 377470
rect 202050 377360 202106 377369
rect 202234 377360 202290 377369
rect 202106 377318 202184 377346
rect 202050 377295 202106 377304
rect 202156 359582 202184 377318
rect 202234 377295 202290 377304
rect 202248 375358 202276 377295
rect 202236 375352 202288 375358
rect 202236 375294 202288 375300
rect 202892 367810 202920 377590
rect 204442 377567 204498 377576
rect 203524 375352 203576 375358
rect 203524 375294 203576 375300
rect 202880 367804 202932 367810
rect 202880 367746 202932 367752
rect 202144 359576 202196 359582
rect 202144 359518 202196 359524
rect 202144 356788 202196 356794
rect 202144 356730 202196 356736
rect 201592 347812 201644 347818
rect 201592 347754 201644 347760
rect 202156 308514 202184 356730
rect 202236 347812 202288 347818
rect 202236 347754 202288 347760
rect 202248 312633 202276 347754
rect 202880 331900 202932 331906
rect 202880 331842 202932 331848
rect 202234 312624 202290 312633
rect 202234 312559 202290 312568
rect 202236 311160 202288 311166
rect 202236 311102 202288 311108
rect 202144 308508 202196 308514
rect 202144 308450 202196 308456
rect 201500 298784 201552 298790
rect 201500 298726 201552 298732
rect 201408 298104 201460 298110
rect 201408 298046 201460 298052
rect 201682 292632 201738 292641
rect 201682 292567 201738 292576
rect 201406 288552 201462 288561
rect 201406 288487 201462 288496
rect 200394 285832 200450 285841
rect 200394 285767 200450 285776
rect 200302 284880 200358 284889
rect 200302 284815 200358 284824
rect 200408 284172 200436 285767
rect 200762 285696 200818 285705
rect 200762 285631 200818 285640
rect 200776 283914 200804 285631
rect 200948 285320 201000 285326
rect 200948 285262 201000 285268
rect 200960 284186 200988 285262
rect 200960 284158 201342 284186
rect 201420 284073 201448 288487
rect 201696 284172 201724 292567
rect 202248 291281 202276 311102
rect 202788 298104 202840 298110
rect 202788 298046 202840 298052
rect 202234 291272 202290 291281
rect 202234 291207 202290 291216
rect 202248 284172 202276 291207
rect 202800 284172 202828 298046
rect 202892 285841 202920 331842
rect 203536 301578 203564 375294
rect 204352 374672 204404 374678
rect 204352 374614 204404 374620
rect 203616 366376 203668 366382
rect 203616 366318 203668 366324
rect 203628 302841 203656 366318
rect 203614 302832 203670 302841
rect 203614 302767 203670 302776
rect 203524 301572 203576 301578
rect 203524 301514 203576 301520
rect 204364 298858 204392 374614
rect 204352 298852 204404 298858
rect 204352 298794 204404 298800
rect 204456 290465 204484 377567
rect 204902 375456 204958 375465
rect 204902 375391 204958 375400
rect 204916 330682 204944 375391
rect 205008 375358 205036 377604
rect 204996 375352 205048 375358
rect 206664 375329 206692 377604
rect 207110 376000 207166 376009
rect 207110 375935 207166 375944
rect 204996 375294 205048 375300
rect 206650 375320 206706 375329
rect 206650 375255 206706 375264
rect 206468 374332 206520 374338
rect 206468 374274 206520 374280
rect 206376 365016 206428 365022
rect 206376 364958 206428 364964
rect 206284 364404 206336 364410
rect 206284 364346 206336 364352
rect 204994 337512 205050 337521
rect 204994 337447 205050 337456
rect 204904 330676 204956 330682
rect 204904 330618 204956 330624
rect 204904 326392 204956 326398
rect 204904 326334 204956 326340
rect 204442 290456 204498 290465
rect 204442 290391 204498 290400
rect 203154 287328 203210 287337
rect 203154 287263 203210 287272
rect 202878 285832 202934 285841
rect 202878 285767 202934 285776
rect 203168 284172 203196 287263
rect 204628 285728 204680 285734
rect 204916 285705 204944 326334
rect 205008 306374 205036 337447
rect 205178 306504 205234 306513
rect 205178 306439 205234 306448
rect 205192 306374 205220 306439
rect 205008 306346 205220 306374
rect 204628 285670 204680 285676
rect 204902 285696 204958 285705
rect 204258 284472 204314 284481
rect 204258 284407 204314 284416
rect 203706 284336 203762 284345
rect 203706 284271 203762 284280
rect 203720 284172 203748 284271
rect 204272 284172 204300 284407
rect 204640 284172 204668 285670
rect 204902 285631 204958 285640
rect 205192 284172 205220 306346
rect 206296 296818 206324 364346
rect 206388 304298 206416 364958
rect 206480 364410 206508 374274
rect 207020 373380 207072 373386
rect 207020 373322 207072 373328
rect 206468 364404 206520 364410
rect 206468 364346 206520 364352
rect 206480 362273 206508 364346
rect 206466 362264 206522 362273
rect 206466 362199 206522 362208
rect 206468 358148 206520 358154
rect 206468 358090 206520 358096
rect 206480 318073 206508 358090
rect 206558 330440 206614 330449
rect 206558 330375 206614 330384
rect 206466 318064 206522 318073
rect 206466 317999 206522 318008
rect 206468 313268 206520 313274
rect 206468 313210 206520 313216
rect 206376 304292 206428 304298
rect 206376 304234 206428 304240
rect 206284 296812 206336 296818
rect 206284 296754 206336 296760
rect 206480 295361 206508 313210
rect 206572 306374 206600 330375
rect 207032 311166 207060 373322
rect 207124 343602 207152 375935
rect 208320 374338 208348 377604
rect 209792 377590 209990 377618
rect 211172 377590 211646 377618
rect 212552 377590 213302 377618
rect 214576 377590 214958 377618
rect 215956 377590 216614 377618
rect 208308 374332 208360 374338
rect 208308 374274 208360 374280
rect 209136 367804 209188 367810
rect 209136 367746 209188 367752
rect 209044 366376 209096 366382
rect 209044 366318 209096 366324
rect 207112 343596 207164 343602
rect 207112 343538 207164 343544
rect 207124 342378 207152 343538
rect 207112 342372 207164 342378
rect 207112 342314 207164 342320
rect 207664 342372 207716 342378
rect 207664 342314 207716 342320
rect 207020 311160 207072 311166
rect 207020 311102 207072 311108
rect 206572 306346 206692 306374
rect 206664 303754 206692 306346
rect 206652 303748 206704 303754
rect 206652 303690 206704 303696
rect 206466 295352 206522 295361
rect 206466 295287 206522 295296
rect 206098 286104 206154 286113
rect 206098 286039 206154 286048
rect 205546 285968 205602 285977
rect 205546 285903 205602 285912
rect 205560 284172 205588 285903
rect 206112 284172 206140 286039
rect 206664 284172 206692 303690
rect 207676 301578 207704 342314
rect 207756 338836 207808 338842
rect 207756 338778 207808 338784
rect 207664 301572 207716 301578
rect 207664 301514 207716 301520
rect 207768 299441 207796 338778
rect 208492 302252 208544 302258
rect 208492 302194 208544 302200
rect 207018 299432 207074 299441
rect 207018 299367 207074 299376
rect 207754 299432 207810 299441
rect 207754 299367 207810 299376
rect 207032 298353 207060 299367
rect 207018 298344 207074 298353
rect 207018 298279 207074 298288
rect 207032 284172 207060 298279
rect 208032 295996 208084 296002
rect 208032 295938 208084 295944
rect 207584 285734 207612 285765
rect 207572 285728 207624 285734
rect 207570 285696 207572 285705
rect 207624 285696 207626 285705
rect 207570 285631 207626 285640
rect 207584 284172 207612 285631
rect 208044 284345 208072 295938
rect 208122 289232 208178 289241
rect 208122 289167 208178 289176
rect 208030 284336 208086 284345
rect 208030 284271 208086 284280
rect 208136 284172 208164 289167
rect 208504 284172 208532 302194
rect 209056 289814 209084 366318
rect 209148 315353 209176 367746
rect 209228 364404 209280 364410
rect 209228 364346 209280 364352
rect 209240 330546 209268 364346
rect 209792 337657 209820 377590
rect 211172 361486 211200 377590
rect 211804 369164 211856 369170
rect 211804 369106 211856 369112
rect 211160 361480 211212 361486
rect 211160 361422 211212 361428
rect 211066 342952 211122 342961
rect 211066 342887 211122 342896
rect 211080 342281 211108 342887
rect 209870 342272 209926 342281
rect 209870 342207 209926 342216
rect 211066 342272 211122 342281
rect 211066 342207 211122 342216
rect 209778 337648 209834 337657
rect 209778 337583 209834 337592
rect 209320 330608 209372 330614
rect 209320 330550 209372 330556
rect 209228 330540 209280 330546
rect 209228 330482 209280 330488
rect 209228 327820 209280 327826
rect 209228 327762 209280 327768
rect 209240 317529 209268 327762
rect 209226 317520 209282 317529
rect 209226 317455 209282 317464
rect 209134 315344 209190 315353
rect 209134 315279 209190 315288
rect 209332 302258 209360 330550
rect 209410 317520 209466 317529
rect 209410 317455 209466 317464
rect 209320 302252 209372 302258
rect 209320 302194 209372 302200
rect 209044 289808 209096 289814
rect 209044 289750 209096 289756
rect 209056 284172 209084 289750
rect 209424 284172 209452 317455
rect 209884 313274 209912 342207
rect 210424 315308 210476 315314
rect 210424 315250 210476 315256
rect 210516 315308 210568 315314
rect 210516 315250 210568 315256
rect 209872 313268 209924 313274
rect 209872 313210 209924 313216
rect 209964 302320 210016 302326
rect 209964 302262 210016 302268
rect 209976 284172 210004 302262
rect 210436 287026 210464 315250
rect 210528 302326 210556 315250
rect 211816 303686 211844 369106
rect 212552 365022 212580 377590
rect 214576 374105 214604 377590
rect 214562 374096 214618 374105
rect 214562 374031 214618 374040
rect 213184 371272 213236 371278
rect 213184 371214 213236 371220
rect 212540 365016 212592 365022
rect 212540 364958 212592 364964
rect 211986 358864 212042 358873
rect 211986 358799 212042 358808
rect 211894 329080 211950 329089
rect 211894 329015 211950 329024
rect 211804 303680 211856 303686
rect 211804 303622 211856 303628
rect 210516 302320 210568 302326
rect 210516 302262 210568 302268
rect 211436 296812 211488 296818
rect 211436 296754 211488 296760
rect 211448 295390 211476 296754
rect 211068 295384 211120 295390
rect 211068 295326 211120 295332
rect 211436 295384 211488 295390
rect 211436 295326 211488 295332
rect 211080 295225 211108 295326
rect 211066 295216 211122 295225
rect 211066 295151 211122 295160
rect 210424 287020 210476 287026
rect 210424 286962 210476 286968
rect 210436 284186 210464 286962
rect 210884 285796 210936 285802
rect 210884 285738 210936 285744
rect 210436 284158 210542 284186
rect 210896 284172 210924 285738
rect 211448 284172 211476 295326
rect 211816 287473 211844 303622
rect 211908 291145 211936 329015
rect 212000 325009 212028 358799
rect 211986 325000 212042 325009
rect 211986 324935 212042 324944
rect 213196 311273 213224 371214
rect 213276 365016 213328 365022
rect 213276 364958 213328 364964
rect 213288 316169 213316 364958
rect 213274 316160 213330 316169
rect 213274 316095 213330 316104
rect 213288 316034 213316 316095
rect 213288 316006 213500 316034
rect 213182 311264 213238 311273
rect 213182 311199 213238 311208
rect 212906 296168 212962 296177
rect 212906 296103 212962 296112
rect 211894 291136 211950 291145
rect 211894 291071 211950 291080
rect 212446 291136 212502 291145
rect 212446 291071 212502 291080
rect 211802 287464 211858 287473
rect 211802 287399 211858 287408
rect 211816 284186 211844 287399
rect 212460 287054 212488 291071
rect 212368 287026 212488 287054
rect 212368 284481 212396 287026
rect 212354 284472 212410 284481
rect 212354 284407 212410 284416
rect 211816 284158 212014 284186
rect 212368 284172 212396 284407
rect 212920 284172 212948 296103
rect 213472 284172 213500 316006
rect 214576 312497 214604 374031
rect 215956 345817 215984 377590
rect 218256 376718 218284 377604
rect 219452 377590 219926 377618
rect 220832 377590 221582 377618
rect 222212 377590 223238 377618
rect 223592 377590 224894 377618
rect 226352 377590 226550 377618
rect 227732 377590 228206 377618
rect 218060 376712 218112 376718
rect 218060 376654 218112 376660
rect 218244 376712 218296 376718
rect 218244 376654 218296 376660
rect 217414 369064 217470 369073
rect 217414 368999 217470 369008
rect 215942 345808 215998 345817
rect 215942 345743 215998 345752
rect 216034 334112 216090 334121
rect 216034 334047 216090 334056
rect 215392 331900 215444 331906
rect 215392 331842 215444 331848
rect 215404 328409 215432 331842
rect 215390 328400 215446 328409
rect 215390 328335 215446 328344
rect 214562 312488 214618 312497
rect 214562 312423 214618 312432
rect 215300 299668 215352 299674
rect 215300 299610 215352 299616
rect 213828 294704 213880 294710
rect 213828 294646 213880 294652
rect 213840 284172 213868 294646
rect 214746 285832 214802 285841
rect 214746 285767 214802 285776
rect 214378 285696 214434 285705
rect 214378 285631 214434 285640
rect 214392 284172 214420 285631
rect 214760 284345 214788 285767
rect 214746 284336 214802 284345
rect 214746 284271 214802 284280
rect 214760 284172 214788 284271
rect 215312 284172 215340 299610
rect 215404 285841 215432 328335
rect 215944 326392 215996 326398
rect 215944 326334 215996 326340
rect 215956 289241 215984 326334
rect 216048 299674 216076 334047
rect 216036 299668 216088 299674
rect 216036 299610 216088 299616
rect 215942 289232 215998 289241
rect 215942 289167 215998 289176
rect 217324 288516 217376 288522
rect 217324 288458 217376 288464
rect 216772 287156 216824 287162
rect 216772 287098 216824 287104
rect 215390 285832 215446 285841
rect 215390 285767 215446 285776
rect 215850 285696 215906 285705
rect 215850 285631 215906 285640
rect 201406 284064 201462 284073
rect 215864 284050 215892 285631
rect 216784 284172 216812 287098
rect 217336 284172 217364 288458
rect 217428 287337 217456 368999
rect 218072 366382 218100 376654
rect 218150 366480 218206 366489
rect 218150 366415 218206 366424
rect 218060 366376 218112 366382
rect 218060 366318 218112 366324
rect 218164 309194 218192 366415
rect 218702 362400 218758 362409
rect 218702 362335 218758 362344
rect 218152 309188 218204 309194
rect 218152 309130 218204 309136
rect 218164 306374 218192 309130
rect 218164 306346 218284 306374
rect 217414 287328 217470 287337
rect 217414 287263 217470 287272
rect 218060 287156 218112 287162
rect 218060 287098 218112 287104
rect 218072 287026 218100 287098
rect 218060 287020 218112 287026
rect 218060 286962 218112 286968
rect 217692 284436 217744 284442
rect 217692 284378 217744 284384
rect 217704 284172 217732 284378
rect 218256 284172 218284 306346
rect 218716 302977 218744 362335
rect 218702 302968 218758 302977
rect 218702 302903 218758 302912
rect 219452 296313 219480 377590
rect 220832 365537 220860 377590
rect 222106 365800 222162 365809
rect 222106 365735 222162 365744
rect 222120 365537 222148 365735
rect 220818 365528 220874 365537
rect 220818 365463 220874 365472
rect 222106 365528 222162 365537
rect 222106 365463 222162 365472
rect 220084 353320 220136 353326
rect 220084 353262 220136 353268
rect 220096 323610 220124 353262
rect 222212 352578 222240 377590
rect 222934 370016 222990 370025
rect 222934 369951 222990 369960
rect 222200 352572 222252 352578
rect 222200 352514 222252 352520
rect 221464 346452 221516 346458
rect 221464 346394 221516 346400
rect 220084 323604 220136 323610
rect 220084 323546 220136 323552
rect 220084 315376 220136 315382
rect 220084 315318 220136 315324
rect 220096 296714 220124 315318
rect 219728 296686 220124 296714
rect 219438 296304 219494 296313
rect 219438 296239 219494 296248
rect 219728 292738 219756 296686
rect 221476 294030 221504 346394
rect 222842 337376 222898 337385
rect 222842 337311 222898 337320
rect 221554 323640 221610 323649
rect 221554 323575 221610 323584
rect 221568 298790 221596 323575
rect 221648 301572 221700 301578
rect 221648 301514 221700 301520
rect 221556 298784 221608 298790
rect 221556 298726 221608 298732
rect 221464 294024 221516 294030
rect 221186 293992 221242 294001
rect 221464 293966 221516 293972
rect 221186 293927 221242 293936
rect 219716 292732 219768 292738
rect 219716 292674 219768 292680
rect 218610 284608 218666 284617
rect 218610 284543 218666 284552
rect 218624 284172 218652 284543
rect 219728 284172 219756 292674
rect 220176 292664 220228 292670
rect 220176 292606 220228 292612
rect 220082 287192 220138 287201
rect 220082 287127 220138 287136
rect 220096 284172 220124 287127
rect 220188 285841 220216 292606
rect 220174 285832 220230 285841
rect 220174 285767 220230 285776
rect 220634 285832 220690 285841
rect 220634 285767 220690 285776
rect 220648 284172 220676 285767
rect 221200 284172 221228 293927
rect 221568 284172 221596 298726
rect 221660 294001 221688 301514
rect 222856 294001 222884 337311
rect 222948 327826 222976 369951
rect 223592 358057 223620 377590
rect 223578 358048 223634 358057
rect 223578 357983 223634 357992
rect 223026 357504 223082 357513
rect 223026 357439 223082 357448
rect 223040 334626 223068 357439
rect 224408 336048 224460 336054
rect 224408 335990 224460 335996
rect 223028 334620 223080 334626
rect 223028 334562 223080 334568
rect 224224 330676 224276 330682
rect 224224 330618 224276 330624
rect 222936 327820 222988 327826
rect 222936 327762 222988 327768
rect 222936 311228 222988 311234
rect 222936 311170 222988 311176
rect 221646 293992 221702 294001
rect 221646 293927 221702 293936
rect 222842 293992 222898 294001
rect 222842 293927 222898 293936
rect 222856 285802 222884 293927
rect 222948 285977 222976 311170
rect 223026 297528 223082 297537
rect 223026 297463 223082 297472
rect 223040 295225 223068 297463
rect 223026 295216 223082 295225
rect 223026 295151 223082 295160
rect 222934 285968 222990 285977
rect 222934 285903 222990 285912
rect 222108 285796 222160 285802
rect 222108 285738 222160 285744
rect 222844 285796 222896 285802
rect 222844 285738 222896 285744
rect 222120 284172 222148 285738
rect 222948 284186 222976 285903
rect 222502 284158 222976 284186
rect 223040 284172 223068 295151
rect 224236 294710 224264 330618
rect 224314 320784 224370 320793
rect 224314 320719 224370 320728
rect 224224 294704 224276 294710
rect 224224 294646 224276 294652
rect 223948 294024 224000 294030
rect 223948 293966 224000 293972
rect 223580 289876 223632 289882
rect 223580 289818 223632 289824
rect 223592 286142 223620 289818
rect 223670 287328 223726 287337
rect 223670 287263 223726 287272
rect 223684 287094 223712 287263
rect 223672 287088 223724 287094
rect 223672 287030 223724 287036
rect 223580 286136 223632 286142
rect 223580 286078 223632 286084
rect 223684 284186 223712 287030
rect 223606 284158 223712 284186
rect 223960 284172 223988 293966
rect 224328 290057 224356 320719
rect 224420 311914 224448 335990
rect 225972 312588 226024 312594
rect 225972 312530 226024 312536
rect 224408 311908 224460 311914
rect 224408 311850 224460 311856
rect 224868 311908 224920 311914
rect 224868 311850 224920 311856
rect 224880 291122 224908 311850
rect 225142 303784 225198 303793
rect 225142 303719 225198 303728
rect 224880 291094 225000 291122
rect 224314 290048 224370 290057
rect 224314 289983 224370 289992
rect 224500 286136 224552 286142
rect 224500 286078 224552 286084
rect 216034 284064 216090 284073
rect 215864 284036 216034 284050
rect 215878 284022 216034 284036
rect 201406 283999 201462 284008
rect 216034 283999 216090 284008
rect 201130 283928 201186 283937
rect 200776 283900 201130 283914
rect 200790 283886 201130 283900
rect 201130 283863 201186 283872
rect 215942 283928 215998 283937
rect 219346 283928 219402 283937
rect 215998 283886 216246 283914
rect 219190 283886 219346 283914
rect 215942 283863 215998 283872
rect 224512 283914 224540 286078
rect 224972 284186 225000 291094
rect 225156 285705 225184 303719
rect 225420 285796 225472 285802
rect 225420 285738 225472 285744
rect 225142 285696 225198 285705
rect 225142 285631 225198 285640
rect 224972 284158 225078 284186
rect 225432 284172 225460 285738
rect 225984 284172 226012 312530
rect 226352 296002 226380 377590
rect 226984 374060 227036 374066
rect 226984 374002 227036 374008
rect 226430 311128 226486 311137
rect 226430 311063 226486 311072
rect 226444 310486 226472 311063
rect 226432 310480 226484 310486
rect 226432 310422 226484 310428
rect 226340 295996 226392 296002
rect 226340 295938 226392 295944
rect 226444 285802 226472 310422
rect 226996 307057 227024 374002
rect 227076 342304 227128 342310
rect 227076 342246 227128 342252
rect 227088 312594 227116 342246
rect 227166 312624 227222 312633
rect 227076 312588 227128 312594
rect 227166 312559 227222 312568
rect 227076 312530 227128 312536
rect 226982 307048 227038 307057
rect 226982 306983 227038 306992
rect 226890 290048 226946 290057
rect 226890 289983 226946 289992
rect 226522 289776 226578 289785
rect 226522 289711 226578 289720
rect 226536 288697 226564 289711
rect 226522 288688 226578 288697
rect 226522 288623 226578 288632
rect 226432 285796 226484 285802
rect 226432 285738 226484 285744
rect 226536 284172 226564 288623
rect 226904 284172 226932 289983
rect 227180 289785 227208 312559
rect 227732 305833 227760 377590
rect 229848 374066 229876 377604
rect 230492 377590 231518 377618
rect 231872 377590 233174 377618
rect 234632 377590 234830 377618
rect 229836 374060 229888 374066
rect 229836 374002 229888 374008
rect 229742 363216 229798 363225
rect 229742 363151 229798 363160
rect 228364 359576 228416 359582
rect 228364 359518 228416 359524
rect 228376 305833 228404 359518
rect 229756 340270 229784 363151
rect 230492 355366 230520 377590
rect 231872 366858 231900 377590
rect 233884 375284 233936 375290
rect 233884 375226 233936 375232
rect 231860 366852 231912 366858
rect 231860 366794 231912 366800
rect 232596 366852 232648 366858
rect 232596 366794 232648 366800
rect 232608 365770 232636 366794
rect 232596 365764 232648 365770
rect 232596 365706 232648 365712
rect 230480 355360 230532 355366
rect 230480 355302 230532 355308
rect 232502 351928 232558 351937
rect 232502 351863 232558 351872
rect 231124 348424 231176 348430
rect 231124 348366 231176 348372
rect 229744 340264 229796 340270
rect 229744 340206 229796 340212
rect 229742 335472 229798 335481
rect 229742 335407 229798 335416
rect 229192 332648 229244 332654
rect 229192 332590 229244 332596
rect 228456 313948 228508 313954
rect 228456 313890 228508 313896
rect 227718 305824 227774 305833
rect 227718 305759 227774 305768
rect 228362 305824 228418 305833
rect 228362 305759 228418 305768
rect 227444 294704 227496 294710
rect 227444 294646 227496 294652
rect 227166 289776 227222 289785
rect 227166 289711 227222 289720
rect 227456 284172 227484 294646
rect 227902 292496 227958 292505
rect 227902 292431 227958 292440
rect 227916 292097 227944 292431
rect 228468 292097 228496 313890
rect 228638 305688 228694 305697
rect 228638 305623 228694 305632
rect 227902 292088 227958 292097
rect 227902 292023 227958 292032
rect 228454 292088 228510 292097
rect 228454 292023 228510 292032
rect 227916 284186 227944 292023
rect 228652 291281 228680 305623
rect 228638 291272 228694 291281
rect 228638 291207 228694 291216
rect 228914 291272 228970 291281
rect 228914 291207 228970 291216
rect 227916 284158 228390 284186
rect 228928 284172 228956 291207
rect 224682 283928 224738 283937
rect 224512 283900 224682 283914
rect 224526 283886 224682 283900
rect 219346 283863 219402 283872
rect 227994 283928 228050 283937
rect 227838 283886 227994 283914
rect 224682 283863 224738 283872
rect 229204 283914 229232 332590
rect 229756 306374 229784 335407
rect 231136 319530 231164 348366
rect 231216 329112 231268 329118
rect 231216 329054 231268 329060
rect 231124 319524 231176 319530
rect 231124 319466 231176 319472
rect 230386 311264 230442 311273
rect 230386 311199 230442 311208
rect 229756 306346 229876 306374
rect 229848 302326 229876 306346
rect 229836 302320 229888 302326
rect 229836 302262 229888 302268
rect 229848 284172 229876 302262
rect 230400 284172 230428 311199
rect 231124 308508 231176 308514
rect 231124 308450 231176 308456
rect 230754 287600 230810 287609
rect 230754 287535 230810 287544
rect 230768 284172 230796 287535
rect 231136 285870 231164 308450
rect 231228 307766 231256 329054
rect 232516 308514 232544 351863
rect 232608 331974 232636 365706
rect 233148 350532 233200 350538
rect 233148 350474 233200 350480
rect 233160 349178 233188 350474
rect 233148 349172 233200 349178
rect 233148 349114 233200 349120
rect 232596 331968 232648 331974
rect 232596 331910 232648 331916
rect 232504 308508 232556 308514
rect 232504 308450 232556 308456
rect 231216 307760 231268 307766
rect 231216 307702 231268 307708
rect 232228 307760 232280 307766
rect 232228 307702 232280 307708
rect 232240 307154 232268 307702
rect 232228 307148 232280 307154
rect 232228 307090 232280 307096
rect 231216 305108 231268 305114
rect 231216 305050 231268 305056
rect 231228 288386 231256 305050
rect 231308 299532 231360 299538
rect 231308 299474 231360 299480
rect 231320 296002 231348 299474
rect 231308 295996 231360 296002
rect 231308 295938 231360 295944
rect 231308 288448 231360 288454
rect 231308 288390 231360 288396
rect 231216 288380 231268 288386
rect 231216 288322 231268 288328
rect 231124 285864 231176 285870
rect 231124 285806 231176 285812
rect 229466 283928 229522 283937
rect 229204 283886 229466 283914
rect 227994 283863 228050 283872
rect 229466 283863 229522 283872
rect 231030 283928 231086 283937
rect 231320 283914 231348 288390
rect 231676 285864 231728 285870
rect 231676 285806 231728 285812
rect 231688 284172 231716 285806
rect 232240 284172 232268 307090
rect 233160 300830 233188 349114
rect 233896 319433 233924 375226
rect 234632 371210 234660 377590
rect 236472 375290 236500 377604
rect 238128 375358 238156 377604
rect 236644 375352 236696 375358
rect 236644 375294 236696 375300
rect 238116 375352 238168 375358
rect 239784 375329 239812 377604
rect 240152 377590 241454 377618
rect 243110 377590 243584 377618
rect 238116 375294 238168 375300
rect 239770 375320 239826 375329
rect 236460 375284 236512 375290
rect 236460 375226 236512 375232
rect 234620 371204 234672 371210
rect 234620 371146 234672 371152
rect 234632 369918 234660 371146
rect 234620 369912 234672 369918
rect 234620 369854 234672 369860
rect 235264 369912 235316 369918
rect 235264 369854 235316 369860
rect 235276 352646 235304 369854
rect 235540 358080 235592 358086
rect 235540 358022 235592 358028
rect 235264 352640 235316 352646
rect 235264 352582 235316 352588
rect 235552 344350 235580 358022
rect 235540 344344 235592 344350
rect 235540 344286 235592 344292
rect 233974 322144 234030 322153
rect 233974 322079 234030 322088
rect 233882 319424 233938 319433
rect 233882 319359 233938 319368
rect 233884 318096 233936 318102
rect 233884 318038 233936 318044
rect 233896 305998 233924 318038
rect 233884 305992 233936 305998
rect 233884 305934 233936 305940
rect 233148 300824 233200 300830
rect 233148 300766 233200 300772
rect 233700 300824 233752 300830
rect 233700 300766 233752 300772
rect 233712 299538 233740 300766
rect 233700 299532 233752 299538
rect 233700 299474 233752 299480
rect 232778 289912 232834 289921
rect 232778 289847 232834 289856
rect 232792 284172 232820 289847
rect 233146 287736 233202 287745
rect 233146 287671 233202 287680
rect 233160 284172 233188 287671
rect 233712 284172 233740 299474
rect 233988 285705 234016 322079
rect 234252 305992 234304 305998
rect 234252 305934 234304 305940
rect 234264 305114 234292 305934
rect 234252 305108 234304 305114
rect 234252 305050 234304 305056
rect 233974 285696 234030 285705
rect 233974 285631 234030 285640
rect 234264 284172 234292 305050
rect 234618 302968 234674 302977
rect 234618 302903 234674 302912
rect 234632 284172 234660 302903
rect 235170 288416 235226 288425
rect 235170 288351 235226 288360
rect 235184 287337 235212 288351
rect 235170 287328 235226 287337
rect 235170 287263 235226 287272
rect 235184 284172 235212 287263
rect 235552 284172 235580 344286
rect 236656 338745 236684 375294
rect 239770 375255 239826 375264
rect 238022 357640 238078 357649
rect 238022 357575 238078 357584
rect 236642 338736 236698 338745
rect 236642 338671 236698 338680
rect 236736 327752 236788 327758
rect 236736 327694 236788 327700
rect 235908 325032 235960 325038
rect 235908 324974 235960 324980
rect 235920 288425 235948 324974
rect 236644 324964 236696 324970
rect 236644 324906 236696 324912
rect 235906 288416 235962 288425
rect 235906 288351 235962 288360
rect 236656 287201 236684 324906
rect 236748 318782 236776 327694
rect 238036 322153 238064 357575
rect 240152 350538 240180 377590
rect 242164 376032 242216 376038
rect 242164 375974 242216 375980
rect 240874 359408 240930 359417
rect 240874 359343 240930 359352
rect 240232 356720 240284 356726
rect 240232 356662 240284 356668
rect 240244 352238 240272 356662
rect 240784 352572 240836 352578
rect 240784 352514 240836 352520
rect 240796 352238 240824 352514
rect 240232 352232 240284 352238
rect 240232 352174 240284 352180
rect 240784 352232 240836 352238
rect 240784 352174 240836 352180
rect 240140 350532 240192 350538
rect 240140 350474 240192 350480
rect 239402 329896 239458 329905
rect 239402 329831 239458 329840
rect 238022 322144 238078 322153
rect 238022 322079 238078 322088
rect 237380 320884 237432 320890
rect 237380 320826 237432 320832
rect 237392 320210 237420 320826
rect 237380 320204 237432 320210
rect 237380 320146 237432 320152
rect 238024 320204 238076 320210
rect 238024 320146 238076 320152
rect 236736 318776 236788 318782
rect 236736 318718 236788 318724
rect 237288 318776 237340 318782
rect 237288 318718 237340 318724
rect 237300 317490 237328 318718
rect 237288 317484 237340 317490
rect 237288 317426 237340 317432
rect 237012 288380 237064 288386
rect 237012 288322 237064 288328
rect 236642 287192 236698 287201
rect 236642 287127 236698 287136
rect 236092 285796 236144 285802
rect 236092 285738 236144 285744
rect 236104 284172 236132 285738
rect 236642 285696 236698 285705
rect 236642 285631 236698 285640
rect 236656 284172 236684 285631
rect 231086 283900 231348 283914
rect 236734 283928 236790 283937
rect 231086 283886 231334 283900
rect 231030 283863 231086 283872
rect 237024 283914 237052 288322
rect 237300 285802 237328 317426
rect 238036 287054 238064 320146
rect 238116 314016 238168 314022
rect 238116 313958 238168 313964
rect 238128 287706 238156 313958
rect 239416 288454 239444 329831
rect 239494 326360 239550 326369
rect 239494 326295 239550 326304
rect 239508 309194 239536 326295
rect 240796 315314 240824 352174
rect 240888 351257 240916 359343
rect 240874 351248 240930 351257
rect 240874 351183 240930 351192
rect 240876 333260 240928 333266
rect 240876 333202 240928 333208
rect 240784 315308 240836 315314
rect 240784 315250 240836 315256
rect 239496 309188 239548 309194
rect 239496 309130 239548 309136
rect 239508 306374 239536 309130
rect 240888 308446 240916 333202
rect 240876 308440 240928 308446
rect 240876 308382 240928 308388
rect 239508 306346 239628 306374
rect 239404 288448 239456 288454
rect 239404 288390 239456 288396
rect 238116 287700 238168 287706
rect 238116 287642 238168 287648
rect 237944 287026 238064 287054
rect 237288 285796 237340 285802
rect 237288 285738 237340 285744
rect 237944 284186 237972 287026
rect 238114 285968 238170 285977
rect 238114 285903 238170 285912
rect 237590 284158 237972 284186
rect 238128 284172 238156 285903
rect 239416 284186 239444 288390
rect 239062 284158 239444 284186
rect 239600 284172 239628 306346
rect 240138 305824 240194 305833
rect 240138 305759 240194 305768
rect 239954 285696 240010 285705
rect 239954 285631 240010 285640
rect 239968 284172 239996 285631
rect 240152 285326 240180 305759
rect 240888 296714 240916 308382
rect 241428 298784 241480 298790
rect 241428 298726 241480 298732
rect 241440 298353 241468 298726
rect 241426 298344 241482 298353
rect 241426 298279 241482 298288
rect 240796 296686 240916 296714
rect 240508 290488 240560 290494
rect 240508 290430 240560 290436
rect 240140 285320 240192 285326
rect 240140 285262 240192 285268
rect 240520 284172 240548 290430
rect 240796 285190 240824 296686
rect 241980 294024 242032 294030
rect 241980 293966 242032 293972
rect 240874 288416 240930 288425
rect 240874 288351 240930 288360
rect 240888 287201 240916 288351
rect 240874 287192 240930 287201
rect 240874 287127 240930 287136
rect 240784 285184 240836 285190
rect 240784 285126 240836 285132
rect 240888 284172 240916 287127
rect 241060 285320 241112 285326
rect 241060 285262 241112 285268
rect 241072 284186 241100 285262
rect 241072 284158 241454 284186
rect 241992 284172 242020 293966
rect 242176 287054 242204 375974
rect 243556 371929 243584 377590
rect 244292 377590 244766 377618
rect 243542 371920 243598 371929
rect 243542 371855 243598 371864
rect 242256 367804 242308 367810
rect 242256 367746 242308 367752
rect 242268 345098 242296 367746
rect 242256 345092 242308 345098
rect 242256 345034 242308 345040
rect 242268 294030 242296 345034
rect 243556 323649 243584 371855
rect 244292 356046 244320 377590
rect 246408 374678 246436 377604
rect 248064 376553 248092 377604
rect 248432 377590 249734 377618
rect 247038 376544 247094 376553
rect 247038 376479 247094 376488
rect 248050 376544 248106 376553
rect 248050 376479 248106 376488
rect 246396 374672 246448 374678
rect 246396 374614 246448 374620
rect 247052 368393 247080 376479
rect 247038 368384 247094 368393
rect 247038 368319 247094 368328
rect 244280 356040 244332 356046
rect 244280 355982 244332 355988
rect 244924 356040 244976 356046
rect 244924 355982 244976 355988
rect 243636 334688 243688 334694
rect 243636 334630 243688 334636
rect 243542 323640 243598 323649
rect 243542 323575 243598 323584
rect 243648 298178 243676 334630
rect 244280 331968 244332 331974
rect 244280 331910 244332 331916
rect 243728 322992 243780 322998
rect 243728 322934 243780 322940
rect 243740 298790 243768 322934
rect 243910 313984 243966 313993
rect 243910 313919 243966 313928
rect 243728 298784 243780 298790
rect 243728 298726 243780 298732
rect 243636 298172 243688 298178
rect 243636 298114 243688 298120
rect 243648 296714 243676 298114
rect 243464 296686 243676 296714
rect 242256 294024 242308 294030
rect 242256 293966 242308 293972
rect 242900 287700 242952 287706
rect 242900 287642 242952 287648
rect 242176 287026 242388 287054
rect 242360 284617 242388 287026
rect 242912 285977 242940 287642
rect 242898 285968 242954 285977
rect 242898 285903 242954 285912
rect 243176 285320 243228 285326
rect 243176 285262 243228 285268
rect 242346 284608 242402 284617
rect 242346 284543 242402 284552
rect 242360 284172 242388 284543
rect 243188 284186 243216 285262
rect 242926 284158 243216 284186
rect 243464 284172 243492 296686
rect 243820 285184 243872 285190
rect 243820 285126 243872 285132
rect 243832 284172 243860 285126
rect 236790 283900 237052 283914
rect 238206 283928 238262 283937
rect 236790 283886 237038 283900
rect 236734 283863 236790 283872
rect 238262 283886 238510 283914
rect 238206 283863 238262 283872
rect 243924 277394 243952 313919
rect 244094 300248 244150 300257
rect 244094 300183 244150 300192
rect 244108 285326 244136 300183
rect 244186 286104 244242 286113
rect 244186 286039 244242 286048
rect 244096 285320 244148 285326
rect 244096 285262 244148 285268
rect 244200 283529 244228 286039
rect 244186 283520 244242 283529
rect 244186 283455 244242 283464
rect 244292 278089 244320 331910
rect 244936 311846 244964 355982
rect 248432 334665 248460 377590
rect 251376 375329 251404 377604
rect 252572 377590 253046 377618
rect 253952 377590 254702 377618
rect 255976 377590 256358 377618
rect 256804 377590 258014 377618
rect 259472 377590 259854 377618
rect 251362 375320 251418 375329
rect 251362 375255 251418 375264
rect 250444 374060 250496 374066
rect 250444 374002 250496 374008
rect 250456 353977 250484 374002
rect 251824 373312 251876 373318
rect 251824 373254 251876 373260
rect 250442 353968 250498 353977
rect 250442 353903 250498 353912
rect 249800 352640 249852 352646
rect 249800 352582 249852 352588
rect 248602 338192 248658 338201
rect 248602 338127 248658 338136
rect 248418 334656 248474 334665
rect 248418 334591 248474 334600
rect 247038 332616 247094 332625
rect 247038 332551 247094 332560
rect 245016 326460 245068 326466
rect 245016 326402 245068 326408
rect 244924 311840 244976 311846
rect 244924 311782 244976 311788
rect 244556 301504 244608 301510
rect 244556 301446 244608 301452
rect 244464 284368 244516 284374
rect 244464 284310 244516 284316
rect 244278 278080 244334 278089
rect 244278 278015 244334 278024
rect 243924 277366 244136 277394
rect 244108 276078 244136 277366
rect 244096 276072 244148 276078
rect 244096 276014 244148 276020
rect 200026 275904 200082 275913
rect 200026 275839 200082 275848
rect 199474 270192 199530 270201
rect 199474 270127 199530 270136
rect 199382 265840 199438 265849
rect 199382 265775 199438 265784
rect 198646 263120 198702 263129
rect 198646 263055 198702 263064
rect 198554 262304 198610 262313
rect 198554 262239 198610 262248
rect 198462 244352 198518 244361
rect 198462 244287 198518 244296
rect 198002 243808 198058 243817
rect 198002 243743 198058 243752
rect 197450 243536 197506 243545
rect 197450 243471 197506 243480
rect 197358 242992 197414 243001
rect 197358 242927 197414 242936
rect 197464 240038 197492 243471
rect 197818 242176 197874 242185
rect 197818 242111 197874 242120
rect 197832 241534 197860 242111
rect 197820 241528 197872 241534
rect 197820 241470 197872 241476
rect 197452 240032 197504 240038
rect 197452 239974 197504 239980
rect 198476 211993 198504 244287
rect 198568 230353 198596 262239
rect 199384 246152 199436 246158
rect 199384 246094 199436 246100
rect 198554 230344 198610 230353
rect 198554 230279 198610 230288
rect 198648 213920 198700 213926
rect 198648 213862 198700 213868
rect 198660 213246 198688 213862
rect 198648 213240 198700 213246
rect 198648 213182 198700 213188
rect 198462 211984 198518 211993
rect 198462 211919 198518 211928
rect 198002 196616 198058 196625
rect 198002 196551 198058 196560
rect 197268 176588 197320 176594
rect 197268 176530 197320 176536
rect 196808 164144 196860 164150
rect 196808 164086 196860 164092
rect 196808 110560 196860 110566
rect 196808 110502 196860 110508
rect 196716 101448 196768 101454
rect 196716 101390 196768 101396
rect 196714 100056 196770 100065
rect 196714 99991 196770 100000
rect 196728 70378 196756 99991
rect 196820 81394 196848 110502
rect 196808 81388 196860 81394
rect 196808 81330 196860 81336
rect 196716 70372 196768 70378
rect 196716 70314 196768 70320
rect 198016 4049 198044 196551
rect 198660 186998 198688 213182
rect 198648 186992 198700 186998
rect 198648 186934 198700 186940
rect 199396 182850 199424 246094
rect 199488 213926 199516 270127
rect 244370 255232 244426 255241
rect 244370 255167 244426 255176
rect 244278 250880 244334 250889
rect 244278 250815 244334 250824
rect 199842 246256 199898 246265
rect 199842 246191 199898 246200
rect 199856 238754 199884 246191
rect 244002 244896 244058 244905
rect 244002 244831 244058 244840
rect 199934 241768 199990 241777
rect 199934 241703 199990 241712
rect 199948 240145 199976 241703
rect 200026 241360 200082 241369
rect 200082 241318 200160 241346
rect 200026 241295 200082 241304
rect 200132 240378 200160 241318
rect 200120 240372 200172 240378
rect 200120 240314 200172 240320
rect 199934 240136 199990 240145
rect 199934 240071 199990 240080
rect 199856 238726 199976 238754
rect 200224 238746 200252 240244
rect 200304 240168 200356 240174
rect 200592 240145 200620 240244
rect 201040 240168 201092 240174
rect 200304 240110 200356 240116
rect 200578 240136 200634 240145
rect 199948 232665 199976 238726
rect 200212 238740 200264 238746
rect 200212 238682 200264 238688
rect 200224 237454 200252 238682
rect 200212 237448 200264 237454
rect 200212 237390 200264 237396
rect 200316 234530 200344 240110
rect 201144 240122 201172 240244
rect 201092 240116 201172 240122
rect 201040 240110 201172 240116
rect 201052 240094 201172 240110
rect 200578 240071 200634 240080
rect 200304 234524 200356 234530
rect 200304 234466 200356 234472
rect 199934 232656 199990 232665
rect 199934 232591 199990 232600
rect 200592 231742 200620 240071
rect 201144 238754 201172 240094
rect 201512 240038 201540 240244
rect 202064 240122 202092 240244
rect 202144 240168 202196 240174
rect 202064 240116 202144 240122
rect 202616 240145 202644 240244
rect 202788 240168 202840 240174
rect 202064 240110 202196 240116
rect 202602 240136 202658 240145
rect 202064 240094 202184 240110
rect 202602 240071 202658 240080
rect 202786 240136 202788 240145
rect 202840 240136 202842 240145
rect 202786 240071 202842 240080
rect 201500 240032 201552 240038
rect 201500 239974 201552 239980
rect 201512 239698 201540 239974
rect 201500 239692 201552 239698
rect 201500 239634 201552 239640
rect 202420 239692 202472 239698
rect 202420 239634 202472 239640
rect 201144 238726 201448 238754
rect 200764 237448 200816 237454
rect 200764 237390 200816 237396
rect 200580 231736 200632 231742
rect 200580 231678 200632 231684
rect 199476 213920 199528 213926
rect 199476 213862 199528 213868
rect 200776 192681 200804 237390
rect 201420 196722 201448 238726
rect 202328 238060 202380 238066
rect 202328 238002 202380 238008
rect 202340 237726 202368 238002
rect 202328 237720 202380 237726
rect 202328 237662 202380 237668
rect 201500 237448 201552 237454
rect 201500 237390 201552 237396
rect 201512 222057 201540 237390
rect 202144 231736 202196 231742
rect 202144 231678 202196 231684
rect 201498 222048 201554 222057
rect 201498 221983 201554 221992
rect 201408 196716 201460 196722
rect 201408 196658 201460 196664
rect 200856 195288 200908 195294
rect 200856 195230 200908 195236
rect 200762 192672 200818 192681
rect 200762 192607 200818 192616
rect 199384 182844 199436 182850
rect 199384 182786 199436 182792
rect 200868 178702 200896 195230
rect 202156 191214 202184 231678
rect 202234 222048 202290 222057
rect 202234 221983 202290 221992
rect 202144 191208 202196 191214
rect 202144 191150 202196 191156
rect 202248 186318 202276 221983
rect 202340 199442 202368 237662
rect 202432 221474 202460 239634
rect 202616 237454 202644 240071
rect 202604 237448 202656 237454
rect 202604 237390 202656 237396
rect 202984 234297 203012 240244
rect 203536 238754 203564 240244
rect 203536 238726 203656 238754
rect 203628 235890 203656 238726
rect 204088 237726 204116 240244
rect 204258 238504 204314 238513
rect 204258 238439 204314 238448
rect 204076 237720 204128 237726
rect 204076 237662 204128 237668
rect 204272 237425 204300 238439
rect 204258 237416 204314 237425
rect 204258 237351 204314 237360
rect 203616 235884 203668 235890
rect 203616 235826 203668 235832
rect 202970 234288 203026 234297
rect 202970 234223 203026 234232
rect 203522 230344 203578 230353
rect 203522 230279 203578 230288
rect 202420 221468 202472 221474
rect 202420 221410 202472 221416
rect 202328 199436 202380 199442
rect 202328 199378 202380 199384
rect 202236 186312 202288 186318
rect 202236 186254 202288 186260
rect 200856 178696 200908 178702
rect 200856 178638 200908 178644
rect 203536 178022 203564 230279
rect 203628 209137 203656 235826
rect 204166 234288 204222 234297
rect 204166 234223 204222 234232
rect 204180 230994 204208 234223
rect 204168 230988 204220 230994
rect 204168 230930 204220 230936
rect 203614 209128 203670 209137
rect 203614 209063 203670 209072
rect 204272 196654 204300 237351
rect 204456 235657 204484 240244
rect 204442 235648 204498 235657
rect 204442 235583 204498 235592
rect 205008 222873 205036 240244
rect 205376 237425 205404 240244
rect 205546 239592 205602 239601
rect 205546 239527 205602 239536
rect 205560 238746 205588 239527
rect 205928 238754 205956 240244
rect 205548 238740 205600 238746
rect 205548 238682 205600 238688
rect 205836 238726 205956 238754
rect 205836 238649 205864 238726
rect 205822 238640 205878 238649
rect 205822 238575 205878 238584
rect 205362 237416 205418 237425
rect 205362 237351 205418 237360
rect 204994 222864 205050 222873
rect 204994 222799 205050 222808
rect 204902 217424 204958 217433
rect 204902 217359 204958 217368
rect 204260 196648 204312 196654
rect 204260 196590 204312 196596
rect 204272 196058 204300 196590
rect 204180 196030 204300 196058
rect 204180 181529 204208 196030
rect 204166 181520 204222 181529
rect 204166 181455 204222 181464
rect 203616 178084 203668 178090
rect 203616 178026 203668 178032
rect 203524 178016 203576 178022
rect 203524 177958 203576 177964
rect 198188 153264 198240 153270
rect 198188 153206 198240 153212
rect 198096 136740 198148 136746
rect 198096 136682 198148 136688
rect 198108 51066 198136 136682
rect 198200 78674 198228 153206
rect 203628 149297 203656 178026
rect 203614 149288 203670 149297
rect 203614 149223 203670 149232
rect 201408 144968 201460 144974
rect 201408 144910 201460 144916
rect 201420 144226 201448 144910
rect 201408 144220 201460 144226
rect 201408 144162 201460 144168
rect 200764 141432 200816 141438
rect 200764 141374 200816 141380
rect 199476 121576 199528 121582
rect 199476 121518 199528 121524
rect 199384 109132 199436 109138
rect 199384 109074 199436 109080
rect 198188 78668 198240 78674
rect 198188 78610 198240 78616
rect 199396 63510 199424 109074
rect 199488 89690 199516 121518
rect 199476 89684 199528 89690
rect 199476 89626 199528 89632
rect 199384 63504 199436 63510
rect 199384 63446 199436 63452
rect 198096 51060 198148 51066
rect 198096 51002 198148 51008
rect 200776 43489 200804 141374
rect 203524 140820 203576 140826
rect 203524 140762 203576 140768
rect 202144 138032 202196 138038
rect 202144 137974 202196 137980
rect 202156 100026 202184 137974
rect 202234 113384 202290 113393
rect 202234 113319 202290 113328
rect 202144 100020 202196 100026
rect 202144 99962 202196 99968
rect 200854 98424 200910 98433
rect 200854 98359 200910 98368
rect 200868 75886 200896 98359
rect 202144 91792 202196 91798
rect 202144 91734 202196 91740
rect 200856 75880 200908 75886
rect 200856 75822 200908 75828
rect 200762 43480 200818 43489
rect 200762 43415 200818 43424
rect 202156 6254 202184 91734
rect 202248 52426 202276 113319
rect 202328 106412 202380 106418
rect 202328 106354 202380 106360
rect 202340 84182 202368 106354
rect 202328 84176 202380 84182
rect 202328 84118 202380 84124
rect 203536 60722 203564 140762
rect 203616 127084 203668 127090
rect 203616 127026 203668 127032
rect 203628 82793 203656 127026
rect 204916 97986 204944 217359
rect 205836 207097 205864 238575
rect 206284 230376 206336 230382
rect 206284 230318 206336 230324
rect 205822 207088 205878 207097
rect 205822 207023 205878 207032
rect 206296 195294 206324 230318
rect 206376 209774 206428 209778
rect 206480 209774 206508 240244
rect 206848 230382 206876 240244
rect 207296 240168 207348 240174
rect 207400 240122 207428 240244
rect 207952 240145 207980 240244
rect 207348 240116 207428 240122
rect 207296 240110 207428 240116
rect 207308 240094 207428 240110
rect 207018 237280 207074 237289
rect 207018 237215 207074 237224
rect 207032 236774 207060 237215
rect 207020 236768 207072 236774
rect 207020 236710 207072 236716
rect 207400 235142 207428 240094
rect 207938 240136 207994 240145
rect 207938 240071 207994 240080
rect 208214 240136 208270 240145
rect 208214 240071 208270 240080
rect 207662 239592 207718 239601
rect 207662 239527 207718 239536
rect 207676 237386 207704 239527
rect 207664 237380 207716 237386
rect 207664 237322 207716 237328
rect 207388 235136 207440 235142
rect 207388 235078 207440 235084
rect 206836 230376 206888 230382
rect 206836 230318 206888 230324
rect 208228 212566 208256 240071
rect 208320 240009 208348 240244
rect 208306 240000 208362 240009
rect 208306 239935 208362 239944
rect 207756 212560 207808 212566
rect 207756 212502 207808 212508
rect 208216 212560 208268 212566
rect 208216 212502 208268 212508
rect 207662 211984 207718 211993
rect 207662 211919 207718 211928
rect 206376 209772 206508 209774
rect 206428 209746 206508 209772
rect 206376 209714 206428 209720
rect 206284 195288 206336 195294
rect 206284 195230 206336 195236
rect 206388 188601 206416 209714
rect 206466 207088 206522 207097
rect 206466 207023 206522 207032
rect 206480 196654 206508 207023
rect 206468 196648 206520 196654
rect 206468 196590 206520 196596
rect 207676 194002 207704 211919
rect 207768 209681 207796 212502
rect 208320 211993 208348 239935
rect 208398 237280 208454 237289
rect 208398 237215 208454 237224
rect 208412 235929 208440 237215
rect 208398 235920 208454 235929
rect 208398 235855 208454 235864
rect 208872 235793 208900 240244
rect 209240 237289 209268 240244
rect 209226 237280 209282 237289
rect 209226 237215 209282 237224
rect 208858 235784 208914 235793
rect 208858 235719 208914 235728
rect 209044 235136 209096 235142
rect 209044 235078 209096 235084
rect 208490 232656 208546 232665
rect 208490 232591 208546 232600
rect 208400 232552 208452 232558
rect 208400 232494 208452 232500
rect 208412 231577 208440 232494
rect 208398 231568 208454 231577
rect 208398 231503 208454 231512
rect 208504 229770 208532 232591
rect 208492 229764 208544 229770
rect 208492 229706 208544 229712
rect 208306 211984 208362 211993
rect 208306 211919 208362 211928
rect 207754 209672 207810 209681
rect 207754 209607 207810 209616
rect 209056 200802 209084 235078
rect 209792 234569 209820 240244
rect 210344 237153 210372 240244
rect 210712 240145 210740 240244
rect 210698 240136 210754 240145
rect 210698 240071 210754 240080
rect 210712 238754 210740 240071
rect 211264 238754 211292 240244
rect 210712 238726 211108 238754
rect 211264 238726 211384 238754
rect 210330 237144 210386 237153
rect 210330 237079 210386 237088
rect 209778 234560 209834 234569
rect 209778 234495 209834 234504
rect 210974 234560 211030 234569
rect 210974 234495 211030 234504
rect 210988 231169 211016 234495
rect 210974 231160 211030 231169
rect 210974 231095 211030 231104
rect 210424 230988 210476 230994
rect 210424 230930 210476 230936
rect 209778 219464 209834 219473
rect 209778 219399 209834 219408
rect 209792 213625 209820 219399
rect 209778 213616 209834 213625
rect 209778 213551 209834 213560
rect 209688 212492 209740 212498
rect 209688 212434 209740 212440
rect 209700 211313 209728 212434
rect 209686 211304 209742 211313
rect 209686 211239 209742 211248
rect 209700 211206 209728 211239
rect 209688 211200 209740 211206
rect 209688 211142 209740 211148
rect 209044 200796 209096 200802
rect 209044 200738 209096 200744
rect 207664 193996 207716 194002
rect 207664 193938 207716 193944
rect 206374 188592 206430 188601
rect 206374 188527 206430 188536
rect 210436 181393 210464 230930
rect 211080 219473 211108 238726
rect 211356 220794 211384 238726
rect 211816 234666 211844 240244
rect 211894 234696 211950 234705
rect 211804 234660 211856 234666
rect 211894 234631 211950 234640
rect 211804 234602 211856 234608
rect 211344 220788 211396 220794
rect 211344 220730 211396 220736
rect 211066 219464 211122 219473
rect 211066 219399 211122 219408
rect 211356 215937 211384 220730
rect 211908 219434 211936 234631
rect 212184 228721 212212 240244
rect 212736 235929 212764 240244
rect 212722 235920 212778 235929
rect 212722 235855 212778 235864
rect 212736 234705 212764 235855
rect 212722 234696 212778 234705
rect 212540 234660 212592 234666
rect 212722 234631 212778 234640
rect 212540 234602 212592 234608
rect 212170 228712 212226 228721
rect 212170 228647 212226 228656
rect 212184 228313 212212 228647
rect 212170 228304 212226 228313
rect 212170 228239 212226 228248
rect 211816 219406 211936 219434
rect 211342 215928 211398 215937
rect 211342 215863 211398 215872
rect 211816 193225 211844 219406
rect 212552 217938 212580 234602
rect 213104 229094 213132 240244
rect 213656 238649 213684 240244
rect 213920 240168 213972 240174
rect 213918 240136 213920 240145
rect 214208 240145 214236 240244
rect 213972 240136 213974 240145
rect 213918 240071 213974 240080
rect 214194 240136 214250 240145
rect 214194 240071 214250 240080
rect 213826 239456 213882 239465
rect 213826 239391 213882 239400
rect 213642 238640 213698 238649
rect 213642 238575 213698 238584
rect 213656 229094 213684 238575
rect 213840 238105 213868 239391
rect 214208 238241 214236 240071
rect 214576 238814 214604 240244
rect 214564 238808 214616 238814
rect 214564 238750 214616 238756
rect 214194 238232 214250 238241
rect 214194 238167 214250 238176
rect 213826 238096 213882 238105
rect 213826 238031 213882 238040
rect 214208 229094 214236 238167
rect 215128 229094 215156 240244
rect 215680 238270 215708 240244
rect 215668 238264 215720 238270
rect 215668 238206 215720 238212
rect 216048 234569 216076 240244
rect 216496 238264 216548 238270
rect 216496 238206 216548 238212
rect 215298 234560 215354 234569
rect 215298 234495 215354 234504
rect 216034 234560 216090 234569
rect 216034 234495 216090 234504
rect 215312 231713 215340 234495
rect 215298 231704 215354 231713
rect 215298 231639 215354 231648
rect 213104 229066 213316 229094
rect 213656 229066 213868 229094
rect 214208 229066 214604 229094
rect 215128 229066 215248 229094
rect 212540 217932 212592 217938
rect 212540 217874 212592 217880
rect 212552 216714 212580 217874
rect 212540 216708 212592 216714
rect 212540 216650 212592 216656
rect 213184 216708 213236 216714
rect 213184 216650 213236 216656
rect 211802 193216 211858 193225
rect 211802 193151 211858 193160
rect 210516 186380 210568 186386
rect 210516 186322 210568 186328
rect 210422 181384 210478 181393
rect 210422 181319 210478 181328
rect 206284 179444 206336 179450
rect 206284 179386 206336 179392
rect 206296 171018 206324 179386
rect 207754 178120 207810 178129
rect 207754 178055 207810 178064
rect 207020 176724 207072 176730
rect 207020 176666 207072 176672
rect 207032 172446 207060 176666
rect 207020 172440 207072 172446
rect 207020 172382 207072 172388
rect 206284 171012 206336 171018
rect 206284 170954 206336 170960
rect 207768 162790 207796 178055
rect 210528 175234 210556 186322
rect 213196 185638 213224 216650
rect 213288 215121 213316 229066
rect 213274 215112 213330 215121
rect 213274 215047 213330 215056
rect 213288 201385 213316 215047
rect 213274 201376 213330 201385
rect 213274 201311 213330 201320
rect 213184 185632 213236 185638
rect 213184 185574 213236 185580
rect 213840 178673 213868 229066
rect 214576 207777 214604 229066
rect 215116 223508 215168 223514
rect 215116 223450 215168 223456
rect 215128 222329 215156 223450
rect 215114 222320 215170 222329
rect 215114 222255 215170 222264
rect 215220 219502 215248 229066
rect 215208 219496 215260 219502
rect 215208 219438 215260 219444
rect 215220 219366 215248 219438
rect 215208 219360 215260 219366
rect 215208 219302 215260 219308
rect 215206 214568 215262 214577
rect 215206 214503 215262 214512
rect 214656 211200 214708 211206
rect 214656 211142 214708 211148
rect 214562 207768 214618 207777
rect 214562 207703 214618 207712
rect 214668 192574 214696 211142
rect 215220 199510 215248 214503
rect 216508 209846 216536 238206
rect 216600 235793 216628 240244
rect 216586 235784 216642 235793
rect 216586 235719 216642 235728
rect 216496 209840 216548 209846
rect 216496 209782 216548 209788
rect 216508 208350 216536 209782
rect 216680 208412 216732 208418
rect 216680 208354 216732 208360
rect 216496 208344 216548 208350
rect 216496 208286 216548 208292
rect 216692 205562 216720 208354
rect 216680 205556 216732 205562
rect 216680 205498 216732 205504
rect 217152 204270 217180 240244
rect 217520 240145 217548 240244
rect 217506 240136 217562 240145
rect 217506 240071 217562 240080
rect 217966 240136 218022 240145
rect 217966 240071 218022 240080
rect 217980 208418 218008 240071
rect 218072 238754 218100 240244
rect 218440 240145 218468 240244
rect 218426 240136 218482 240145
rect 218426 240071 218482 240080
rect 218702 240136 218758 240145
rect 218992 240106 219020 240244
rect 218702 240071 218758 240080
rect 218980 240100 219032 240106
rect 218072 238726 218284 238754
rect 217968 208412 218020 208418
rect 217968 208354 218020 208360
rect 218256 204338 218284 238726
rect 218716 223553 218744 240071
rect 218980 240042 219032 240048
rect 218992 231742 219020 240042
rect 219544 238513 219572 240244
rect 219912 240106 219940 240244
rect 219900 240100 219952 240106
rect 219900 240042 219952 240048
rect 219912 238754 219940 240042
rect 219912 238726 220124 238754
rect 219912 238678 219940 238726
rect 219900 238672 219952 238678
rect 219900 238614 219952 238620
rect 219530 238504 219586 238513
rect 219530 238439 219586 238448
rect 218980 231736 219032 231742
rect 218980 231678 219032 231684
rect 218702 223544 218758 223553
rect 218702 223479 218758 223488
rect 218060 204332 218112 204338
rect 218060 204274 218112 204280
rect 218244 204332 218296 204338
rect 218244 204274 218296 204280
rect 217140 204264 217192 204270
rect 218072 204241 218100 204274
rect 217140 204206 217192 204212
rect 218058 204232 218114 204241
rect 217152 200114 217180 204206
rect 218058 204167 218114 204176
rect 217152 200086 217364 200114
rect 215208 199504 215260 199510
rect 215208 199446 215260 199452
rect 214656 192568 214708 192574
rect 214656 192510 214708 192516
rect 217336 189786 217364 200086
rect 217416 193928 217468 193934
rect 217416 193870 217468 193876
rect 217324 189780 217376 189786
rect 217324 189722 217376 189728
rect 217428 184521 217456 193870
rect 217414 184512 217470 184521
rect 217414 184447 217470 184456
rect 220096 183025 220124 238726
rect 220464 216578 220492 240244
rect 221016 238377 221044 240244
rect 221384 240145 221412 240244
rect 221832 240168 221884 240174
rect 221370 240136 221426 240145
rect 221936 240122 221964 240244
rect 221884 240116 221964 240122
rect 221832 240110 221964 240116
rect 221844 240094 221964 240110
rect 221370 240071 221426 240080
rect 221464 238808 221516 238814
rect 221464 238750 221516 238756
rect 221002 238368 221058 238377
rect 221002 238303 221058 238312
rect 221016 226302 221044 238303
rect 221476 234297 221504 238750
rect 222304 238746 222332 240244
rect 222292 238740 222344 238746
rect 222292 238682 222344 238688
rect 221462 234288 221518 234297
rect 221462 234223 221518 234232
rect 221004 226296 221056 226302
rect 221004 226238 221056 226244
rect 222856 226234 222884 240244
rect 223408 238754 223436 240244
rect 223304 238740 223356 238746
rect 223408 238726 223528 238754
rect 223304 238682 223356 238688
rect 223316 233073 223344 238682
rect 223500 238649 223528 238726
rect 223486 238640 223542 238649
rect 223486 238575 223542 238584
rect 223396 237448 223448 237454
rect 223396 237390 223448 237396
rect 223302 233064 223358 233073
rect 223302 232999 223358 233008
rect 223316 229094 223344 232999
rect 223408 232558 223436 237390
rect 223396 232552 223448 232558
rect 223396 232494 223448 232500
rect 223316 229066 223436 229094
rect 222844 226228 222896 226234
rect 222844 226170 222896 226176
rect 220176 216572 220228 216578
rect 220176 216514 220228 216520
rect 220452 216572 220504 216578
rect 220452 216514 220504 216520
rect 220082 183016 220138 183025
rect 220082 182951 220138 182960
rect 214932 180872 214984 180878
rect 214932 180814 214984 180820
rect 213826 178664 213882 178673
rect 213826 178599 213882 178608
rect 213920 176656 213972 176662
rect 213920 176598 213972 176604
rect 213932 175681 213960 176598
rect 213918 175672 213974 175681
rect 213918 175607 213974 175616
rect 214562 175264 214618 175273
rect 210516 175228 210568 175234
rect 210516 175170 210568 175176
rect 214012 175228 214064 175234
rect 214562 175199 214564 175208
rect 214012 175170 214064 175176
rect 214616 175199 214618 175208
rect 214564 175170 214616 175176
rect 213920 175092 213972 175098
rect 213920 175034 213972 175040
rect 213932 175001 213960 175034
rect 213918 174992 213974 175001
rect 213918 174927 213974 174936
rect 214024 174321 214052 175170
rect 214010 174312 214066 174321
rect 214010 174247 214066 174256
rect 213920 173868 213972 173874
rect 213920 173810 213972 173816
rect 213932 172961 213960 173810
rect 214944 173641 214972 180814
rect 220188 178770 220216 216514
rect 220266 210352 220322 210361
rect 220266 210287 220322 210296
rect 220280 193866 220308 210287
rect 220268 193860 220320 193866
rect 220268 193802 220320 193808
rect 220726 192536 220782 192545
rect 220726 192471 220782 192480
rect 220268 188352 220320 188358
rect 220268 188294 220320 188300
rect 220280 180198 220308 188294
rect 220740 185881 220768 192471
rect 220726 185872 220782 185881
rect 220726 185807 220782 185816
rect 222856 181665 222884 226170
rect 223408 192545 223436 229066
rect 223394 192536 223450 192545
rect 223394 192471 223450 192480
rect 223500 186726 223528 238575
rect 223776 229090 223804 240244
rect 224328 232626 224356 240244
rect 224880 238814 224908 240244
rect 225248 240122 225276 240244
rect 225328 240168 225380 240174
rect 225248 240116 225328 240122
rect 225248 240110 225380 240116
rect 225248 240094 225368 240110
rect 224868 238808 224920 238814
rect 224868 238750 224920 238756
rect 225800 238754 225828 240244
rect 224316 232620 224368 232626
rect 224316 232562 224368 232568
rect 223764 229084 223816 229090
rect 223764 229026 223816 229032
rect 223776 227798 223804 229026
rect 223764 227792 223816 227798
rect 223764 227734 223816 227740
rect 224328 219434 224356 232562
rect 224236 219406 224356 219434
rect 224236 216646 224264 219406
rect 224224 216640 224276 216646
rect 224224 216582 224276 216588
rect 223488 186720 223540 186726
rect 223488 186662 223540 186668
rect 222842 181656 222898 181665
rect 222842 181591 222898 181600
rect 220268 180192 220320 180198
rect 220268 180134 220320 180140
rect 220176 178764 220228 178770
rect 220176 178706 220228 178712
rect 224880 176905 224908 238750
rect 225616 238726 225828 238754
rect 225616 206922 225644 238726
rect 225800 238678 225828 238726
rect 225788 238672 225840 238678
rect 225788 238614 225840 238620
rect 226168 232529 226196 240244
rect 226720 238377 226748 240244
rect 226706 238368 226762 238377
rect 226706 238303 226762 238312
rect 226720 238105 226748 238303
rect 226706 238096 226762 238105
rect 226706 238031 226762 238040
rect 226154 232520 226210 232529
rect 226154 232455 226210 232464
rect 226168 219434 226196 232455
rect 226984 227792 227036 227798
rect 226984 227734 227036 227740
rect 225708 219406 226196 219434
rect 225604 206916 225656 206922
rect 225604 206858 225656 206864
rect 225708 203590 225736 219406
rect 225696 203584 225748 203590
rect 225696 203526 225748 203532
rect 226248 180872 226300 180878
rect 226248 180814 226300 180820
rect 226260 180713 226288 180814
rect 226246 180704 226302 180713
rect 226246 180639 226302 180648
rect 226432 180124 226484 180130
rect 226432 180066 226484 180072
rect 226340 178016 226392 178022
rect 226340 177958 226392 177964
rect 224866 176896 224922 176905
rect 224866 176831 224922 176840
rect 226352 176769 226380 177958
rect 226338 176760 226394 176769
rect 226338 176695 226394 176704
rect 226444 175982 226472 180066
rect 226996 178945 227024 227734
rect 227272 224874 227300 240244
rect 227640 226001 227668 240244
rect 227720 235272 227772 235278
rect 227720 235214 227772 235220
rect 227732 233238 227760 235214
rect 228192 234433 228220 240244
rect 228362 235648 228418 235657
rect 228362 235583 228418 235592
rect 228178 234424 228234 234433
rect 228178 234359 228234 234368
rect 227720 233232 227772 233238
rect 227720 233174 227772 233180
rect 227626 225992 227682 226001
rect 227626 225927 227682 225936
rect 227260 224868 227312 224874
rect 227260 224810 227312 224816
rect 227272 220794 227300 224810
rect 228376 221921 228404 235583
rect 228744 235278 228772 240244
rect 228732 235272 228784 235278
rect 228732 235214 228784 235220
rect 229112 227798 229140 240244
rect 229664 237454 229692 240244
rect 229652 237448 229704 237454
rect 229652 237390 229704 237396
rect 230216 235657 230244 240244
rect 230584 240145 230612 240244
rect 230570 240136 230626 240145
rect 230570 240071 230626 240080
rect 230754 240136 230810 240145
rect 230754 240071 230810 240080
rect 230202 235648 230258 235657
rect 230202 235583 230258 235592
rect 229100 227792 229152 227798
rect 229100 227734 229152 227740
rect 228362 221912 228418 221921
rect 228362 221847 228418 221856
rect 227260 220788 227312 220794
rect 227260 220730 227312 220736
rect 227076 220108 227128 220114
rect 227076 220050 227128 220056
rect 227088 184278 227116 220050
rect 227718 219600 227774 219609
rect 227718 219535 227774 219544
rect 227732 219434 227760 219535
rect 228364 219496 228416 219502
rect 228364 219438 228416 219444
rect 227720 219428 227772 219434
rect 227720 219370 227772 219376
rect 227720 193996 227772 194002
rect 227720 193938 227772 193944
rect 227732 191282 227760 193938
rect 227720 191276 227772 191282
rect 227720 191218 227772 191224
rect 227168 186720 227220 186726
rect 227168 186662 227220 186668
rect 227076 184272 227128 184278
rect 227076 184214 227128 184220
rect 227180 179450 227208 186662
rect 227168 179444 227220 179450
rect 227168 179386 227220 179392
rect 226982 178936 227038 178945
rect 226982 178871 227038 178880
rect 227718 178664 227774 178673
rect 227718 178599 227774 178608
rect 227732 177449 227760 178599
rect 226522 177440 226578 177449
rect 226522 177375 226578 177384
rect 227718 177440 227774 177449
rect 227718 177375 227774 177384
rect 226432 175976 226484 175982
rect 226432 175918 226484 175924
rect 226536 175846 226564 177375
rect 228376 177342 228404 219438
rect 229376 204332 229428 204338
rect 229376 204274 229428 204280
rect 228456 191140 228508 191146
rect 228456 191082 228508 191088
rect 228364 177336 228416 177342
rect 228364 177278 228416 177284
rect 228468 175846 228496 191082
rect 229006 181248 229062 181257
rect 229006 181183 229062 181192
rect 226524 175840 226576 175846
rect 226524 175782 226576 175788
rect 228456 175840 228508 175846
rect 228456 175782 228508 175788
rect 229020 175030 229048 181183
rect 229284 179444 229336 179450
rect 229284 179386 229336 179392
rect 229190 178936 229246 178945
rect 229190 178871 229246 178880
rect 229100 176724 229152 176730
rect 229100 176666 229152 176672
rect 229008 175024 229060 175030
rect 229008 174966 229060 174972
rect 229112 173777 229140 176666
rect 229098 173768 229154 173777
rect 229098 173703 229154 173712
rect 214930 173632 214986 173641
rect 214930 173567 214986 173576
rect 213918 172952 213974 172961
rect 213918 172887 213974 172896
rect 213920 172508 213972 172514
rect 213920 172450 213972 172456
rect 213932 172281 213960 172450
rect 214012 172440 214064 172446
rect 214012 172382 214064 172388
rect 213918 172272 213974 172281
rect 213918 172207 213974 172216
rect 214024 171601 214052 172382
rect 229204 171850 229232 178871
rect 229112 171822 229232 171850
rect 214010 171592 214066 171601
rect 214010 171527 214066 171536
rect 213920 171080 213972 171086
rect 213918 171048 213920 171057
rect 213972 171048 213974 171057
rect 213918 170983 213974 170992
rect 214012 171012 214064 171018
rect 214012 170954 214064 170960
rect 214024 170377 214052 170954
rect 214010 170368 214066 170377
rect 214010 170303 214066 170312
rect 214102 170232 214158 170241
rect 214102 170167 214158 170176
rect 214012 169720 214064 169726
rect 213918 169688 213974 169697
rect 214012 169662 214064 169668
rect 213918 169623 213920 169632
rect 213972 169623 213974 169632
rect 213920 169594 213972 169600
rect 214024 169017 214052 169662
rect 214010 169008 214066 169017
rect 214010 168943 214066 168952
rect 214012 168360 214064 168366
rect 213918 168328 213974 168337
rect 214012 168302 214064 168308
rect 213918 168263 213920 168272
rect 213972 168263 213974 168272
rect 213920 168234 213972 168240
rect 214024 167657 214052 168302
rect 214010 167648 214066 167657
rect 214010 167583 214066 167592
rect 213920 167000 213972 167006
rect 213918 166968 213920 166977
rect 213972 166968 213974 166977
rect 213918 166903 213974 166912
rect 214012 166932 214064 166938
rect 214012 166874 214064 166880
rect 214024 165753 214052 166874
rect 214116 166433 214144 170167
rect 214102 166424 214158 166433
rect 214102 166359 214158 166368
rect 214010 165744 214066 165753
rect 214010 165679 214066 165688
rect 214012 165572 214064 165578
rect 214012 165514 214064 165520
rect 213920 165504 213972 165510
rect 213920 165446 213972 165452
rect 213932 165073 213960 165446
rect 213918 165064 213974 165073
rect 213918 164999 213974 165008
rect 214024 164393 214052 165514
rect 214010 164384 214066 164393
rect 214010 164319 214066 164328
rect 214012 164212 214064 164218
rect 214012 164154 214064 164160
rect 213920 164144 213972 164150
rect 213920 164086 213972 164092
rect 213932 163713 213960 164086
rect 213918 163704 213974 163713
rect 213918 163639 213974 163648
rect 214024 163033 214052 164154
rect 214010 163024 214066 163033
rect 214010 162959 214066 162968
rect 213920 162852 213972 162858
rect 213920 162794 213972 162800
rect 207756 162784 207808 162790
rect 207756 162726 207808 162732
rect 213932 162353 213960 162794
rect 214012 162784 214064 162790
rect 214012 162726 214064 162732
rect 213918 162344 213974 162353
rect 213918 162279 213974 162288
rect 207664 162172 207716 162178
rect 207664 162114 207716 162120
rect 206376 153332 206428 153338
rect 206376 153274 206428 153280
rect 204996 146940 205048 146946
rect 204996 146882 205048 146888
rect 206284 146940 206336 146946
rect 206284 146882 206336 146888
rect 204904 97980 204956 97986
rect 204904 97922 204956 97928
rect 205008 86193 205036 146882
rect 205180 118720 205232 118726
rect 205180 118662 205232 118668
rect 205088 100020 205140 100026
rect 205088 99962 205140 99968
rect 204994 86184 205050 86193
rect 204994 86119 205050 86128
rect 204996 84856 205048 84862
rect 204996 84798 205048 84804
rect 203614 82784 203670 82793
rect 203614 82719 203670 82728
rect 204904 82136 204956 82142
rect 204904 82078 204956 82084
rect 203524 60716 203576 60722
rect 203524 60658 203576 60664
rect 202236 52420 202288 52426
rect 202236 52362 202288 52368
rect 204916 11830 204944 82078
rect 205008 17270 205036 84798
rect 205100 69018 205128 99962
rect 205192 88262 205220 118662
rect 205180 88256 205232 88262
rect 205180 88198 205232 88204
rect 206296 86902 206324 146882
rect 206388 133210 206416 153274
rect 206376 133204 206428 133210
rect 206376 133146 206428 133152
rect 206376 95260 206428 95266
rect 206376 95202 206428 95208
rect 206284 86896 206336 86902
rect 206284 86838 206336 86844
rect 206284 84924 206336 84930
rect 206284 84866 206336 84872
rect 205088 69012 205140 69018
rect 205088 68954 205140 68960
rect 206296 36582 206324 84866
rect 206388 55214 206416 95202
rect 207676 83502 207704 162114
rect 214024 161809 214052 162726
rect 214010 161800 214066 161809
rect 214010 161735 214066 161744
rect 214012 161424 214064 161430
rect 214012 161366 214064 161372
rect 213920 161356 213972 161362
rect 213920 161298 213972 161304
rect 213932 161129 213960 161298
rect 213918 161120 213974 161129
rect 213918 161055 213974 161064
rect 214024 160449 214052 161366
rect 214102 160712 214158 160721
rect 214102 160647 214158 160656
rect 214010 160440 214066 160449
rect 214010 160375 214066 160384
rect 213920 160064 213972 160070
rect 213920 160006 213972 160012
rect 213932 159769 213960 160006
rect 213918 159760 213974 159769
rect 213918 159695 213974 159704
rect 214116 159089 214144 160647
rect 214102 159080 214158 159089
rect 214102 159015 214158 159024
rect 214012 158704 214064 158710
rect 214012 158646 214064 158652
rect 213920 158636 213972 158642
rect 213920 158578 213972 158584
rect 213932 158409 213960 158578
rect 213918 158400 213974 158409
rect 213918 158335 213974 158344
rect 214024 157729 214052 158646
rect 214010 157720 214066 157729
rect 214010 157655 214066 157664
rect 214012 157344 214064 157350
rect 214012 157286 214064 157292
rect 213920 157276 213972 157282
rect 213920 157218 213972 157224
rect 213932 157185 213960 157218
rect 213918 157176 213974 157185
rect 213918 157111 213974 157120
rect 214024 156505 214052 157286
rect 214010 156496 214066 156505
rect 214010 156431 214066 156440
rect 214012 155916 214064 155922
rect 214012 155858 214064 155864
rect 213920 155848 213972 155854
rect 213918 155816 213920 155825
rect 213972 155816 213974 155825
rect 213918 155751 213974 155760
rect 214024 155145 214052 155858
rect 214010 155136 214066 155145
rect 214010 155071 214066 155080
rect 214010 154456 214066 154465
rect 214010 154391 214066 154400
rect 213918 153776 213974 153785
rect 213918 153711 213974 153720
rect 213932 153338 213960 153711
rect 213920 153332 213972 153338
rect 213920 153274 213972 153280
rect 214024 153270 214052 154391
rect 214012 153264 214064 153270
rect 214012 153206 214064 153212
rect 214010 153096 214066 153105
rect 214010 153031 214066 153040
rect 214024 152250 214052 153031
rect 214562 152552 214618 152561
rect 214562 152487 214618 152496
rect 211804 152244 211856 152250
rect 211804 152186 211856 152192
rect 214012 152244 214064 152250
rect 214012 152186 214064 152192
rect 209044 143676 209096 143682
rect 209044 143618 209096 143624
rect 207756 128376 207808 128382
rect 207756 128318 207808 128324
rect 207664 83496 207716 83502
rect 207664 83438 207716 83444
rect 207768 57934 207796 128318
rect 209056 102814 209084 143618
rect 209136 132592 209188 132598
rect 209136 132534 209188 132540
rect 209044 102808 209096 102814
rect 209044 102750 209096 102756
rect 209044 94512 209096 94518
rect 209044 94454 209096 94460
rect 207756 57928 207808 57934
rect 207756 57870 207808 57876
rect 206376 55208 206428 55214
rect 206376 55150 206428 55156
rect 206284 36576 206336 36582
rect 206284 36518 206336 36524
rect 206376 36576 206428 36582
rect 206376 36518 206428 36524
rect 206388 18698 206416 36518
rect 209056 20058 209084 94454
rect 209148 91633 209176 132534
rect 210516 131232 210568 131238
rect 210516 131174 210568 131180
rect 210528 119377 210556 131174
rect 210514 119368 210570 119377
rect 210514 119303 210570 119312
rect 210424 118788 210476 118794
rect 210424 118730 210476 118736
rect 209226 105224 209282 105233
rect 209226 105159 209282 105168
rect 209134 91624 209190 91633
rect 209134 91559 209190 91568
rect 209240 89010 209268 105159
rect 210436 91050 210464 118730
rect 211816 112470 211844 152186
rect 213182 151872 213238 151881
rect 213182 151807 213238 151816
rect 213196 135930 213224 151807
rect 214010 151192 214066 151201
rect 214010 151127 214066 151136
rect 213920 150544 213972 150550
rect 213918 150512 213920 150521
rect 213972 150512 213974 150521
rect 214024 150482 214052 151127
rect 213918 150447 213974 150456
rect 214012 150476 214064 150482
rect 214012 150418 214064 150424
rect 214104 150408 214156 150414
rect 214104 150350 214156 150356
rect 213920 149728 213972 149734
rect 213920 149670 213972 149676
rect 213932 148481 213960 149670
rect 214116 149161 214144 150350
rect 214102 149152 214158 149161
rect 214102 149087 214158 149096
rect 213918 148472 213974 148481
rect 213918 148407 213974 148416
rect 213918 147928 213974 147937
rect 213918 147863 213974 147872
rect 213932 147694 213960 147863
rect 213920 147688 213972 147694
rect 213920 147630 213972 147636
rect 214010 147248 214066 147257
rect 214010 147183 214066 147192
rect 213918 146568 213974 146577
rect 213918 146503 213974 146512
rect 213932 146334 213960 146503
rect 213920 146328 213972 146334
rect 213920 146270 213972 146276
rect 214024 145586 214052 147183
rect 214576 146946 214604 152487
rect 214564 146940 214616 146946
rect 214564 146882 214616 146888
rect 229112 146849 229140 171822
rect 229296 166994 229324 179386
rect 229388 177041 229416 204274
rect 230768 190454 230796 240071
rect 231136 223582 231164 240244
rect 231504 238754 231532 240244
rect 231952 240168 232004 240174
rect 231950 240136 231952 240145
rect 232004 240136 232006 240145
rect 231950 240071 232006 240080
rect 231228 238726 231532 238754
rect 231228 237153 231256 238726
rect 231214 237144 231270 237153
rect 231214 237079 231270 237088
rect 231228 228993 231256 237079
rect 232056 229094 232084 240244
rect 232608 238513 232636 240244
rect 232594 238504 232650 238513
rect 232594 238439 232650 238448
rect 232976 234433 233004 240244
rect 233148 240168 233200 240174
rect 233148 240110 233200 240116
rect 233160 238678 233188 240110
rect 233148 238672 233200 238678
rect 233148 238614 233200 238620
rect 232962 234424 233018 234433
rect 232962 234359 233018 234368
rect 231872 229066 232084 229094
rect 231214 228984 231270 228993
rect 231214 228919 231270 228928
rect 231124 223576 231176 223582
rect 231124 223518 231176 223524
rect 231872 222193 231900 229066
rect 232976 228857 233004 234359
rect 232962 228848 233018 228857
rect 232962 228783 233018 228792
rect 231952 227792 232004 227798
rect 231952 227734 232004 227740
rect 231858 222184 231914 222193
rect 231858 222119 231914 222128
rect 231122 219600 231178 219609
rect 231122 219535 231178 219544
rect 230768 190426 230980 190454
rect 230202 186280 230258 186289
rect 230202 186215 230258 186224
rect 230216 185706 230244 186215
rect 230204 185700 230256 185706
rect 230204 185642 230256 185648
rect 230662 184512 230718 184521
rect 230662 184447 230718 184456
rect 230572 184204 230624 184210
rect 230572 184146 230624 184152
rect 229468 182912 229520 182918
rect 229468 182854 229520 182860
rect 229374 177032 229430 177041
rect 229374 176967 229430 176976
rect 229374 175808 229430 175817
rect 229374 175743 229430 175752
rect 229388 175166 229416 175743
rect 229376 175160 229428 175166
rect 229376 175102 229428 175108
rect 229204 166966 229324 166994
rect 229204 155825 229232 166966
rect 229480 166161 229508 182854
rect 230388 172576 230440 172582
rect 230388 172518 230440 172524
rect 229466 166152 229522 166161
rect 229466 166087 229522 166096
rect 230020 164212 230072 164218
rect 230020 164154 230072 164160
rect 229190 155816 229246 155825
rect 229190 155751 229246 155760
rect 229742 147928 229798 147937
rect 229742 147863 229798 147872
rect 229098 146840 229154 146849
rect 229098 146775 229154 146784
rect 215942 145888 215998 145897
rect 215942 145823 215998 145832
rect 214012 145580 214064 145586
rect 214012 145522 214064 145528
rect 213918 145208 213974 145217
rect 213918 145143 213974 145152
rect 213932 144974 213960 145143
rect 213920 144968 213972 144974
rect 213920 144910 213972 144916
rect 214010 144528 214066 144537
rect 214010 144463 214066 144472
rect 213918 143848 213974 143857
rect 213918 143783 213974 143792
rect 213932 143682 213960 143783
rect 213920 143676 213972 143682
rect 213920 143618 213972 143624
rect 214024 143614 214052 144463
rect 214012 143608 214064 143614
rect 214012 143550 214064 143556
rect 213918 143304 213974 143313
rect 213918 143239 213974 143248
rect 213932 142186 213960 143239
rect 213920 142180 213972 142186
rect 213920 142122 213972 142128
rect 213918 141944 213974 141953
rect 213918 141879 213974 141888
rect 213932 140826 213960 141879
rect 214102 141264 214158 141273
rect 214102 141199 214158 141208
rect 213920 140820 213972 140826
rect 213920 140762 213972 140768
rect 213918 140584 213974 140593
rect 213918 140519 213974 140528
rect 213932 139466 213960 140519
rect 214010 139904 214066 139913
rect 214010 139839 214066 139848
rect 213920 139460 213972 139466
rect 213920 139402 213972 139408
rect 214024 138718 214052 139839
rect 214012 138712 214064 138718
rect 213918 138680 213974 138689
rect 214012 138654 214064 138660
rect 213918 138615 213974 138624
rect 213932 138038 213960 138615
rect 213920 138032 213972 138038
rect 213920 137974 213972 137980
rect 214010 138000 214066 138009
rect 214010 137935 214066 137944
rect 213920 136740 213972 136746
rect 213920 136682 213972 136688
rect 213366 136640 213422 136649
rect 213366 136575 213422 136584
rect 213184 135924 213236 135930
rect 213184 135866 213236 135872
rect 213274 133920 213330 133929
rect 213274 133855 213330 133864
rect 213182 119504 213238 119513
rect 213182 119439 213238 119448
rect 211804 112464 211856 112470
rect 211804 112406 211856 112412
rect 211896 111920 211948 111926
rect 211896 111862 211948 111868
rect 211804 93152 211856 93158
rect 211804 93094 211856 93100
rect 210424 91044 210476 91050
rect 210424 90986 210476 90992
rect 210422 89040 210478 89049
rect 209228 89004 209280 89010
rect 210422 88975 210478 88984
rect 209228 88946 209280 88952
rect 209136 87712 209188 87718
rect 209136 87654 209188 87660
rect 209148 54534 209176 87654
rect 209136 54528 209188 54534
rect 209136 54470 209188 54476
rect 210436 43518 210464 88975
rect 210424 43512 210476 43518
rect 210424 43454 210476 43460
rect 209044 20052 209096 20058
rect 209044 19994 209096 20000
rect 206376 18692 206428 18698
rect 206376 18634 206428 18640
rect 204996 17264 205048 17270
rect 204996 17206 205048 17212
rect 204904 11824 204956 11830
rect 204904 11766 204956 11772
rect 211816 8974 211844 93094
rect 211908 90409 211936 111862
rect 212448 102264 212500 102270
rect 212448 102206 212500 102212
rect 212460 94489 212488 102206
rect 212446 94480 212502 94489
rect 212446 94415 212502 94424
rect 211894 90400 211950 90409
rect 211894 90335 211950 90344
rect 213196 22681 213224 119439
rect 213288 64870 213316 133855
rect 213380 93809 213408 136575
rect 213932 135969 213960 136682
rect 214024 136678 214052 137935
rect 214012 136672 214064 136678
rect 214012 136614 214064 136620
rect 213918 135960 213974 135969
rect 213918 135895 213974 135904
rect 213920 135312 213972 135318
rect 213918 135280 213920 135289
rect 213972 135280 213974 135289
rect 213918 135215 213974 135224
rect 213918 134600 213974 134609
rect 214116 134570 214144 141199
rect 214838 139224 214894 139233
rect 214838 139159 214894 139168
rect 214746 137320 214802 137329
rect 214746 137255 214802 137264
rect 213918 134535 213974 134544
rect 214104 134564 214156 134570
rect 213932 133958 213960 134535
rect 214104 134506 214156 134512
rect 213920 133952 213972 133958
rect 213920 133894 213972 133900
rect 214010 133376 214066 133385
rect 214010 133311 214066 133320
rect 213918 132696 213974 132705
rect 213918 132631 213974 132640
rect 213932 132598 213960 132631
rect 213920 132592 213972 132598
rect 213920 132534 213972 132540
rect 214024 132530 214052 133311
rect 214012 132524 214064 132530
rect 214012 132466 214064 132472
rect 213918 132016 213974 132025
rect 213918 131951 213974 131960
rect 213932 131170 213960 131951
rect 214010 131336 214066 131345
rect 214010 131271 214066 131280
rect 214024 131238 214052 131271
rect 214012 131232 214064 131238
rect 214012 131174 214064 131180
rect 213920 131164 213972 131170
rect 213920 131106 213972 131112
rect 213918 130656 213974 130665
rect 213918 130591 213974 130600
rect 213932 129810 213960 130591
rect 214654 129976 214710 129985
rect 214654 129911 214710 129920
rect 213920 129804 213972 129810
rect 213920 129746 213972 129752
rect 214562 129296 214618 129305
rect 214562 129231 214618 129240
rect 213918 128752 213974 128761
rect 213918 128687 213974 128696
rect 213932 128382 213960 128687
rect 213920 128376 213972 128382
rect 213920 128318 213972 128324
rect 214010 128072 214066 128081
rect 214010 128007 214066 128016
rect 213918 127392 213974 127401
rect 213918 127327 213974 127336
rect 213932 127090 213960 127327
rect 213920 127084 213972 127090
rect 213920 127026 213972 127032
rect 214024 127022 214052 128007
rect 214012 127016 214064 127022
rect 214012 126958 214064 126964
rect 214010 126712 214066 126721
rect 214010 126647 214066 126656
rect 213918 126032 213974 126041
rect 213918 125967 213974 125976
rect 213932 125730 213960 125967
rect 213920 125724 213972 125730
rect 213920 125666 213972 125672
rect 214024 125662 214052 126647
rect 214012 125656 214064 125662
rect 214012 125598 214064 125604
rect 214010 125352 214066 125361
rect 214010 125287 214066 125296
rect 213918 124672 213974 124681
rect 213918 124607 213974 124616
rect 213932 124234 213960 124607
rect 213920 124228 213972 124234
rect 213920 124170 213972 124176
rect 213918 124128 213974 124137
rect 213918 124063 213974 124072
rect 213932 122874 213960 124063
rect 214024 123486 214052 125287
rect 214012 123480 214064 123486
rect 214012 123422 214064 123428
rect 213920 122868 213972 122874
rect 213920 122810 213972 122816
rect 214010 122768 214066 122777
rect 214010 122703 214066 122712
rect 213918 122088 213974 122097
rect 213918 122023 213974 122032
rect 213932 121514 213960 122023
rect 214024 121582 214052 122703
rect 214012 121576 214064 121582
rect 214012 121518 214064 121524
rect 213920 121508 213972 121514
rect 213920 121450 213972 121456
rect 214010 121408 214066 121417
rect 214010 121343 214066 121352
rect 213918 120728 213974 120737
rect 213918 120663 213974 120672
rect 213932 120222 213960 120663
rect 213920 120216 213972 120222
rect 213920 120158 213972 120164
rect 214024 120154 214052 121343
rect 214012 120148 214064 120154
rect 214012 120090 214064 120096
rect 214102 120048 214158 120057
rect 214102 119983 214158 119992
rect 213918 119504 213974 119513
rect 213918 119439 213974 119448
rect 213932 118726 213960 119439
rect 214010 118824 214066 118833
rect 214010 118759 214012 118768
rect 214064 118759 214066 118768
rect 214012 118730 214064 118736
rect 213920 118720 213972 118726
rect 213920 118662 213972 118668
rect 214010 118144 214066 118153
rect 214010 118079 214066 118088
rect 213918 117464 213974 117473
rect 214024 117434 214052 118079
rect 213918 117399 213974 117408
rect 214012 117428 214064 117434
rect 213932 117366 213960 117399
rect 214012 117370 214064 117376
rect 213920 117360 213972 117366
rect 213920 117302 213972 117308
rect 214010 116784 214066 116793
rect 214010 116719 214066 116728
rect 213918 116104 213974 116113
rect 213918 116039 213920 116048
rect 213972 116039 213974 116048
rect 213920 116010 213972 116016
rect 214024 116006 214052 116719
rect 214012 116000 214064 116006
rect 214012 115942 214064 115948
rect 214010 115424 214066 115433
rect 214010 115359 214066 115368
rect 213918 114880 213974 114889
rect 213918 114815 213974 114824
rect 213932 114646 213960 114815
rect 213920 114640 213972 114646
rect 213920 114582 213972 114588
rect 214024 114578 214052 115359
rect 214012 114572 214064 114578
rect 214012 114514 214064 114520
rect 213918 114200 213974 114209
rect 213918 114135 213974 114144
rect 213932 113218 213960 114135
rect 214116 113830 214144 119983
rect 214104 113824 214156 113830
rect 214104 113766 214156 113772
rect 213920 113212 213972 113218
rect 213920 113154 213972 113160
rect 214010 112840 214066 112849
rect 214010 112775 214066 112784
rect 213918 112160 213974 112169
rect 213918 112095 213974 112104
rect 213932 111858 213960 112095
rect 214024 111926 214052 112775
rect 214012 111920 214064 111926
rect 214012 111862 214064 111868
rect 213920 111852 213972 111858
rect 213920 111794 213972 111800
rect 214010 111480 214066 111489
rect 214010 111415 214066 111424
rect 213918 110800 213974 110809
rect 213918 110735 213974 110744
rect 213932 110566 213960 110735
rect 213920 110560 213972 110566
rect 213920 110502 213972 110508
rect 214024 110498 214052 111415
rect 214012 110492 214064 110498
rect 214012 110434 214064 110440
rect 214010 110256 214066 110265
rect 214010 110191 214066 110200
rect 213918 109576 213974 109585
rect 213918 109511 213974 109520
rect 213932 109070 213960 109511
rect 214024 109138 214052 110191
rect 214012 109132 214064 109138
rect 214012 109074 214064 109080
rect 213920 109064 213972 109070
rect 213920 109006 213972 109012
rect 214010 108896 214066 108905
rect 214010 108831 214066 108840
rect 213918 108216 213974 108225
rect 213918 108151 213974 108160
rect 213932 107778 213960 108151
rect 213920 107772 213972 107778
rect 213920 107714 213972 107720
rect 214024 107710 214052 108831
rect 214012 107704 214064 107710
rect 214012 107646 214064 107652
rect 214010 107536 214066 107545
rect 214010 107471 214066 107480
rect 213918 106856 213974 106865
rect 213918 106791 213974 106800
rect 213932 106350 213960 106791
rect 214024 106418 214052 107471
rect 214012 106412 214064 106418
rect 214012 106354 214064 106360
rect 213920 106344 213972 106350
rect 213920 106286 213972 106292
rect 214010 106176 214066 106185
rect 214010 106111 214066 106120
rect 214024 104990 214052 106111
rect 214012 104984 214064 104990
rect 213918 104952 213974 104961
rect 214012 104926 214064 104932
rect 213918 104887 213920 104896
rect 213972 104887 213974 104896
rect 213920 104858 213972 104864
rect 213918 104272 213974 104281
rect 213918 104207 213974 104216
rect 213932 103562 213960 104207
rect 213920 103556 213972 103562
rect 213920 103498 213972 103504
rect 213918 102912 213974 102921
rect 213918 102847 213974 102856
rect 213932 102202 213960 102847
rect 214012 102264 214064 102270
rect 214010 102232 214012 102241
rect 214064 102232 214066 102241
rect 213920 102196 213972 102202
rect 214010 102167 214066 102176
rect 213920 102138 213972 102144
rect 214010 101552 214066 101561
rect 214010 101487 214066 101496
rect 213918 101008 213974 101017
rect 213918 100943 213974 100952
rect 213932 100774 213960 100943
rect 213920 100768 213972 100774
rect 213920 100710 213972 100716
rect 214024 100065 214052 101487
rect 214102 100328 214158 100337
rect 214102 100263 214158 100272
rect 214010 100056 214066 100065
rect 214010 99991 214066 100000
rect 213918 99648 213974 99657
rect 213918 99583 213974 99592
rect 213932 99414 213960 99583
rect 213920 99408 213972 99414
rect 213920 99350 213972 99356
rect 214116 98666 214144 100263
rect 214104 98660 214156 98666
rect 214104 98602 214156 98608
rect 213918 98288 213974 98297
rect 213918 98223 213974 98232
rect 213932 98054 213960 98223
rect 213920 98048 213972 98054
rect 213920 97990 213972 97996
rect 213918 97608 213974 97617
rect 213918 97543 213974 97552
rect 213932 96694 213960 97543
rect 213920 96688 213972 96694
rect 213920 96630 213972 96636
rect 213918 96384 213974 96393
rect 213918 96319 213974 96328
rect 213932 95266 213960 96319
rect 213920 95260 213972 95266
rect 213920 95202 213972 95208
rect 214576 94586 214604 129231
rect 214668 113174 214696 129911
rect 214760 124914 214788 137255
rect 214852 129062 214880 139159
rect 214840 129056 214892 129062
rect 214840 128998 214892 129004
rect 214748 124908 214800 124914
rect 214748 124850 214800 124856
rect 214668 113146 214880 113174
rect 214852 100026 214880 113146
rect 214840 100020 214892 100026
rect 214840 99962 214892 99968
rect 214654 96928 214710 96937
rect 214654 96863 214710 96872
rect 214564 94580 214616 94586
rect 214564 94522 214616 94528
rect 213366 93800 213422 93809
rect 213366 93735 213422 93744
rect 214564 89004 214616 89010
rect 214564 88946 214616 88952
rect 213276 64864 213328 64870
rect 213276 64806 213328 64812
rect 213182 22672 213238 22681
rect 213182 22607 213238 22616
rect 211804 8968 211856 8974
rect 211804 8910 211856 8916
rect 202144 6248 202196 6254
rect 202144 6190 202196 6196
rect 214576 4894 214604 88946
rect 214668 67590 214696 96863
rect 214656 67584 214708 67590
rect 214656 67526 214708 67532
rect 215956 62082 215984 145823
rect 216034 142624 216090 142633
rect 216034 142559 216090 142568
rect 216048 95946 216076 142559
rect 229756 139233 229784 147863
rect 229928 147688 229980 147694
rect 229928 147630 229980 147636
rect 229834 145616 229890 145625
rect 229834 145551 229890 145560
rect 229742 139224 229798 139233
rect 229742 139159 229798 139168
rect 229742 135824 229798 135833
rect 229742 135759 229798 135768
rect 216126 123448 216182 123457
rect 216126 123383 216182 123392
rect 216036 95940 216088 95946
rect 216036 95882 216088 95888
rect 216036 93220 216088 93226
rect 216036 93162 216088 93168
rect 215944 62076 215996 62082
rect 215944 62018 215996 62024
rect 216048 22846 216076 93162
rect 216140 88330 216168 123383
rect 217232 101448 217284 101454
rect 217232 101390 217284 101396
rect 216128 88324 216180 88330
rect 216128 88266 216180 88272
rect 217244 87553 217272 101390
rect 229100 97980 229152 97986
rect 229100 97922 229152 97928
rect 229112 97889 229140 97922
rect 229098 97880 229154 97889
rect 229098 97815 229154 97824
rect 229192 97368 229244 97374
rect 229192 97310 229244 97316
rect 229204 97209 229232 97310
rect 229190 97200 229246 97209
rect 229190 97135 229246 97144
rect 219348 96076 219400 96082
rect 219348 96018 219400 96024
rect 219360 93945 219388 96018
rect 228362 95840 228418 95849
rect 228362 95775 228418 95784
rect 225696 95260 225748 95266
rect 225696 95202 225748 95208
rect 225602 94480 225658 94489
rect 225602 94415 225658 94424
rect 219346 93936 219402 93945
rect 219346 93871 219402 93880
rect 224224 93900 224276 93906
rect 224224 93842 224276 93848
rect 222934 93256 222990 93265
rect 222934 93191 222990 93200
rect 217324 91860 217376 91866
rect 217324 91802 217376 91808
rect 217230 87544 217286 87553
rect 217230 87479 217286 87488
rect 217336 53106 217364 91802
rect 222844 90432 222896 90438
rect 222844 90374 222896 90380
rect 220084 90364 220136 90370
rect 220084 90306 220136 90312
rect 218704 89072 218756 89078
rect 218704 89014 218756 89020
rect 217324 53100 217376 53106
rect 217324 53042 217376 53048
rect 216036 22840 216088 22846
rect 216036 22782 216088 22788
rect 214564 4888 214616 4894
rect 214564 4830 214616 4836
rect 198002 4040 198058 4049
rect 198002 3975 198058 3984
rect 196622 3496 196678 3505
rect 187056 3460 187108 3466
rect 187056 3402 187108 3408
rect 195244 3460 195296 3466
rect 196622 3431 196678 3440
rect 195244 3402 195296 3408
rect 177394 3360 177450 3369
rect 177394 3295 177450 3304
rect 140042 2680 140098 2689
rect 140042 2615 140098 2624
rect 142802 2680 142858 2689
rect 142802 2615 142858 2624
rect 140056 480 140084 2615
rect 218716 2174 218744 89014
rect 220096 31142 220124 90306
rect 220176 35284 220228 35290
rect 220176 35226 220228 35232
rect 220084 31136 220136 31142
rect 220084 31078 220136 31084
rect 220188 2174 220216 35226
rect 222856 15978 222884 90374
rect 222948 64161 222976 93191
rect 222934 64152 222990 64161
rect 222934 64087 222990 64096
rect 224236 36582 224264 93842
rect 224224 36576 224276 36582
rect 224224 36518 224276 36524
rect 225616 21486 225644 94415
rect 225708 79393 225736 95202
rect 226982 93936 227038 93945
rect 226982 93871 227038 93880
rect 225694 79384 225750 79393
rect 225694 79319 225750 79328
rect 225604 21480 225656 21486
rect 225604 21422 225656 21428
rect 222844 15972 222896 15978
rect 222844 15914 222896 15920
rect 226996 7682 227024 93871
rect 227076 87644 227128 87650
rect 227076 87586 227128 87592
rect 227088 14482 227116 87586
rect 228376 37942 228404 95775
rect 229756 76673 229784 135759
rect 229848 106185 229876 145551
rect 229940 137873 229968 147630
rect 230032 146305 230060 164154
rect 230400 162858 230428 172518
rect 230584 169969 230612 184146
rect 230676 175681 230704 184447
rect 230662 175672 230718 175681
rect 230662 175607 230718 175616
rect 230664 175228 230716 175234
rect 230664 175170 230716 175176
rect 230570 169960 230626 169969
rect 230570 169895 230626 169904
rect 230572 169516 230624 169522
rect 230572 169458 230624 169464
rect 230584 169017 230612 169458
rect 230570 169008 230626 169017
rect 230570 168943 230626 168952
rect 230676 164218 230704 175170
rect 230756 173188 230808 173194
rect 230756 173130 230808 173136
rect 230768 172417 230796 173130
rect 230754 172408 230810 172417
rect 230754 172343 230810 172352
rect 230952 166994 230980 190426
rect 231136 185745 231164 219535
rect 231872 219434 231900 222119
rect 231860 219428 231912 219434
rect 231860 219370 231912 219376
rect 231964 211041 231992 227734
rect 233240 223576 233292 223582
rect 233238 223544 233240 223553
rect 233292 223544 233294 223553
rect 233238 223479 233294 223488
rect 233332 214600 233384 214606
rect 233332 214542 233384 214548
rect 232136 212628 232188 212634
rect 232136 212570 232188 212576
rect 231950 211032 232006 211041
rect 231950 210967 232006 210976
rect 231122 185736 231178 185745
rect 231122 185671 231178 185680
rect 231952 178696 232004 178702
rect 231952 178638 232004 178644
rect 231964 176654 231992 178638
rect 231964 176626 232084 176654
rect 231306 176080 231362 176089
rect 231306 176015 231362 176024
rect 231320 175273 231348 176015
rect 231860 175840 231912 175846
rect 231860 175782 231912 175788
rect 231306 175264 231362 175273
rect 231306 175199 231362 175208
rect 231400 172508 231452 172514
rect 231400 172450 231452 172456
rect 231308 172440 231360 172446
rect 231308 172382 231360 172388
rect 231320 171465 231348 172382
rect 231412 171873 231440 172450
rect 231398 171864 231454 171873
rect 231398 171799 231454 171808
rect 231306 171456 231362 171465
rect 231306 171391 231362 171400
rect 231872 170513 231900 175782
rect 231952 175024 232004 175030
rect 231952 174966 232004 174972
rect 231858 170504 231914 170513
rect 231858 170439 231914 170448
rect 231216 169788 231268 169794
rect 231216 169730 231268 169736
rect 231124 169448 231176 169454
rect 231124 169390 231176 169396
rect 231136 168609 231164 169390
rect 231122 168600 231178 168609
rect 231122 168535 231178 168544
rect 230768 166966 230980 166994
rect 230664 164212 230716 164218
rect 230664 164154 230716 164160
rect 230388 162852 230440 162858
rect 230388 162794 230440 162800
rect 230386 156632 230442 156641
rect 230386 156567 230442 156576
rect 230400 148073 230428 156567
rect 230570 153096 230626 153105
rect 230570 153031 230626 153040
rect 230584 151609 230612 153031
rect 230570 151600 230626 151609
rect 230570 151535 230626 151544
rect 230386 148064 230442 148073
rect 230386 147999 230442 148008
rect 230018 146296 230074 146305
rect 230018 146231 230074 146240
rect 230768 139777 230796 166966
rect 231032 164212 231084 164218
rect 231032 164154 231084 164160
rect 231044 163849 231072 164154
rect 231030 163840 231086 163849
rect 231030 163775 231086 163784
rect 230848 162852 230900 162858
rect 230848 162794 230900 162800
rect 230940 162852 230992 162858
rect 230940 162794 230992 162800
rect 230860 157729 230888 162794
rect 230952 161945 230980 162794
rect 231124 162172 231176 162178
rect 231124 162114 231176 162120
rect 230938 161936 230994 161945
rect 230938 161871 230994 161880
rect 230846 157720 230902 157729
rect 230846 157655 230902 157664
rect 231136 142154 231164 162114
rect 231228 160585 231256 169730
rect 231400 168088 231452 168094
rect 231398 168056 231400 168065
rect 231452 168056 231454 168065
rect 231398 167991 231454 168000
rect 231400 167136 231452 167142
rect 231398 167104 231400 167113
rect 231452 167104 231454 167113
rect 231398 167039 231454 167048
rect 231768 166728 231820 166734
rect 231766 166696 231768 166705
rect 231820 166696 231822 166705
rect 231766 166631 231822 166640
rect 231492 165232 231544 165238
rect 231490 165200 231492 165209
rect 231544 165200 231546 165209
rect 231490 165135 231546 165144
rect 231676 164144 231728 164150
rect 231676 164086 231728 164092
rect 231688 162897 231716 164086
rect 231674 162888 231730 162897
rect 231674 162823 231730 162832
rect 231964 161474 231992 174966
rect 232056 164801 232084 176626
rect 232042 164792 232098 164801
rect 232042 164727 232098 164736
rect 231872 161446 231992 161474
rect 231676 160744 231728 160750
rect 231676 160686 231728 160692
rect 231214 160576 231270 160585
rect 231214 160511 231270 160520
rect 231400 159996 231452 160002
rect 231400 159938 231452 159944
rect 231412 159089 231440 159938
rect 231398 159080 231454 159089
rect 231398 159015 231454 159024
rect 231688 158681 231716 160686
rect 231768 160064 231820 160070
rect 231766 160032 231768 160041
rect 231820 160032 231822 160041
rect 231766 159967 231822 159976
rect 231674 158672 231730 158681
rect 231216 158636 231268 158642
rect 231674 158607 231730 158616
rect 231216 158578 231268 158584
rect 231228 158137 231256 158578
rect 231214 158128 231270 158137
rect 231214 158063 231270 158072
rect 231582 158128 231638 158137
rect 231582 158063 231638 158072
rect 231492 155848 231544 155854
rect 231492 155790 231544 155796
rect 231504 155281 231532 155790
rect 231490 155272 231546 155281
rect 231490 155207 231546 155216
rect 231492 154556 231544 154562
rect 231492 154498 231544 154504
rect 231504 153377 231532 154498
rect 231490 153368 231546 153377
rect 231490 153303 231546 153312
rect 231492 152992 231544 152998
rect 231490 152960 231492 152969
rect 231544 152960 231546 152969
rect 231490 152895 231546 152904
rect 231596 152017 231624 158063
rect 231674 157992 231730 158001
rect 231674 157927 231730 157936
rect 231688 157185 231716 157927
rect 231768 157276 231820 157282
rect 231768 157218 231820 157224
rect 231674 157176 231730 157185
rect 231674 157111 231730 157120
rect 231780 156777 231808 157218
rect 231766 156768 231822 156777
rect 231766 156703 231822 156712
rect 231766 156224 231822 156233
rect 231872 156210 231900 161446
rect 231822 156182 231900 156210
rect 231766 156159 231822 156168
rect 231676 155236 231728 155242
rect 231676 155178 231728 155184
rect 231688 154329 231716 155178
rect 231768 154488 231820 154494
rect 231768 154430 231820 154436
rect 231674 154320 231730 154329
rect 231674 154255 231730 154264
rect 231780 153921 231808 154430
rect 231766 153912 231822 153921
rect 231766 153847 231822 153856
rect 231582 152008 231638 152017
rect 231582 151943 231638 151952
rect 231492 151768 231544 151774
rect 231492 151710 231544 151716
rect 231504 151065 231532 151710
rect 231490 151056 231546 151065
rect 231490 150991 231546 151000
rect 231766 151056 231822 151065
rect 231766 150991 231822 151000
rect 231676 150952 231728 150958
rect 231676 150894 231728 150900
rect 231688 150657 231716 150894
rect 231674 150648 231730 150657
rect 231674 150583 231730 150592
rect 231492 148844 231544 148850
rect 231492 148786 231544 148792
rect 231504 148753 231532 148786
rect 231490 148744 231546 148753
rect 231490 148679 231546 148688
rect 231582 148336 231638 148345
rect 231582 148271 231638 148280
rect 231216 144900 231268 144906
rect 231216 144842 231268 144848
rect 231044 142126 231164 142154
rect 230754 139768 230810 139777
rect 230754 139703 230810 139712
rect 229926 137864 229982 137873
rect 229926 137799 229982 137808
rect 230572 136604 230624 136610
rect 230572 136546 230624 136552
rect 230584 135969 230612 136546
rect 230570 135960 230626 135969
rect 230570 135895 230626 135904
rect 230756 134564 230808 134570
rect 230756 134506 230808 134512
rect 229926 132832 229982 132841
rect 229926 132767 229982 132776
rect 229834 106176 229890 106185
rect 229834 106111 229890 106120
rect 229940 93945 229968 132767
rect 230572 131096 230624 131102
rect 230572 131038 230624 131044
rect 230584 129849 230612 131038
rect 230570 129840 230626 129849
rect 230570 129775 230626 129784
rect 230572 127696 230624 127702
rect 230572 127638 230624 127644
rect 230584 126449 230612 127638
rect 230768 127401 230796 134506
rect 231044 134473 231072 142126
rect 231122 142080 231178 142089
rect 231122 142015 231178 142024
rect 231136 141370 231164 142015
rect 231124 141364 231176 141370
rect 231124 141306 231176 141312
rect 231030 134464 231086 134473
rect 231030 134399 231086 134408
rect 230848 133884 230900 133890
rect 230848 133826 230900 133832
rect 230860 133521 230888 133826
rect 230846 133512 230902 133521
rect 230846 133447 230902 133456
rect 231124 131776 231176 131782
rect 231124 131718 231176 131724
rect 230940 129056 230992 129062
rect 230940 128998 230992 129004
rect 230754 127392 230810 127401
rect 230754 127327 230810 127336
rect 230848 126880 230900 126886
rect 230848 126822 230900 126828
rect 230570 126440 230626 126449
rect 230570 126375 230626 126384
rect 230860 126041 230888 126822
rect 230846 126032 230902 126041
rect 230846 125967 230902 125976
rect 230018 123312 230074 123321
rect 230018 123247 230074 123256
rect 229926 93936 229982 93945
rect 230032 93906 230060 123247
rect 230952 123185 230980 128998
rect 231136 128353 231164 131718
rect 231228 130257 231256 144842
rect 231596 144401 231624 148271
rect 231780 148209 231808 150991
rect 231766 148200 231822 148209
rect 231766 148135 231822 148144
rect 232148 147694 232176 212570
rect 232596 196716 232648 196722
rect 232596 196658 232648 196664
rect 232504 191208 232556 191214
rect 232504 191150 232556 191156
rect 232228 180192 232280 180198
rect 232228 180134 232280 180140
rect 232240 175234 232268 180134
rect 232516 178702 232544 191150
rect 232608 185774 232636 196658
rect 232596 185768 232648 185774
rect 232596 185710 232648 185716
rect 233056 185700 233108 185706
rect 233056 185642 233108 185648
rect 233068 185065 233096 185642
rect 233054 185056 233110 185065
rect 233054 184991 233110 185000
rect 233240 178764 233292 178770
rect 233240 178706 233292 178712
rect 232504 178696 232556 178702
rect 232504 178638 232556 178644
rect 232228 175228 232280 175234
rect 232228 175170 232280 175176
rect 232240 174729 232268 175170
rect 232226 174720 232282 174729
rect 232226 174655 232282 174664
rect 233252 169522 233280 178706
rect 233344 172582 233372 214542
rect 233528 194585 233556 240244
rect 234080 230450 234108 240244
rect 234448 238754 234476 240244
rect 234448 238726 234568 238754
rect 234068 230444 234120 230450
rect 234068 230386 234120 230392
rect 234080 228410 234108 230386
rect 234068 228404 234120 228410
rect 234068 228346 234120 228352
rect 234540 224210 234568 238726
rect 235000 224777 235028 240244
rect 235368 233238 235396 240244
rect 235920 238649 235948 240244
rect 236472 240145 236500 240244
rect 236458 240136 236514 240145
rect 236458 240071 236514 240080
rect 235906 238640 235962 238649
rect 235906 238575 235962 238584
rect 235356 233232 235408 233238
rect 235356 233174 235408 233180
rect 236840 227497 236868 240244
rect 237392 238814 237420 240244
rect 237944 240145 237972 240244
rect 237930 240136 237986 240145
rect 237930 240071 237986 240080
rect 237380 238808 237432 238814
rect 237380 238750 237432 238756
rect 237392 234598 237420 238750
rect 237944 234614 237972 240071
rect 237380 234592 237432 234598
rect 237944 234586 238064 234614
rect 237380 234534 237432 234540
rect 236826 227488 236882 227497
rect 236826 227423 236882 227432
rect 236840 226953 236868 227423
rect 236826 226944 236882 226953
rect 236826 226879 236882 226888
rect 234986 224768 235042 224777
rect 234986 224703 235042 224712
rect 234540 224182 234660 224210
rect 234632 204202 234660 224182
rect 237378 212528 237434 212537
rect 237378 212463 237434 212472
rect 237392 211818 237420 212463
rect 237380 211812 237432 211818
rect 237380 211754 237432 211760
rect 234620 204196 234672 204202
rect 234620 204138 234672 204144
rect 233514 194576 233570 194585
rect 233514 194511 233570 194520
rect 233884 192568 233936 192574
rect 233884 192510 233936 192516
rect 233896 180130 233924 192510
rect 233884 180124 233936 180130
rect 233884 180066 233936 180072
rect 233424 177336 233476 177342
rect 233424 177278 233476 177284
rect 233332 172576 233384 172582
rect 233332 172518 233384 172524
rect 233240 169516 233292 169522
rect 233240 169458 233292 169464
rect 232594 164928 232650 164937
rect 232594 164863 232650 164872
rect 232502 159080 232558 159089
rect 232502 159015 232558 159024
rect 232136 147688 232188 147694
rect 232136 147630 232188 147636
rect 231766 147112 231822 147121
rect 231766 147047 231822 147056
rect 231676 146260 231728 146266
rect 231676 146202 231728 146208
rect 231688 144945 231716 146202
rect 231674 144936 231730 144945
rect 231674 144871 231730 144880
rect 231582 144392 231638 144401
rect 231582 144327 231638 144336
rect 231676 143472 231728 143478
rect 231780 143449 231808 147047
rect 231676 143414 231728 143420
rect 231766 143440 231822 143449
rect 231688 143041 231716 143414
rect 231766 143375 231822 143384
rect 231674 143032 231730 143041
rect 231674 142967 231730 142976
rect 231308 142928 231360 142934
rect 231308 142870 231360 142876
rect 231320 131617 231348 142870
rect 231768 140752 231820 140758
rect 231766 140720 231768 140729
rect 231820 140720 231822 140729
rect 231766 140655 231822 140664
rect 231676 140072 231728 140078
rect 231676 140014 231728 140020
rect 231492 138916 231544 138922
rect 231492 138858 231544 138864
rect 231504 138281 231532 138858
rect 231490 138272 231546 138281
rect 231490 138207 231546 138216
rect 231584 137964 231636 137970
rect 231584 137906 231636 137912
rect 231596 136921 231624 137906
rect 231582 136912 231638 136921
rect 231582 136847 231638 136856
rect 231492 135924 231544 135930
rect 231492 135866 231544 135872
rect 231504 135425 231532 135866
rect 231490 135416 231546 135425
rect 231490 135351 231546 135360
rect 231584 135244 231636 135250
rect 231584 135186 231636 135192
rect 231596 134065 231624 135186
rect 231582 134056 231638 134065
rect 231582 133991 231638 134000
rect 231688 132569 231716 140014
rect 231768 133816 231820 133822
rect 231768 133758 231820 133764
rect 231780 133113 231808 133758
rect 231766 133104 231822 133113
rect 231766 133039 231822 133048
rect 231674 132560 231730 132569
rect 231674 132495 231730 132504
rect 231676 132456 231728 132462
rect 231676 132398 231728 132404
rect 231306 131608 231362 131617
rect 231306 131543 231362 131552
rect 231688 131209 231716 132398
rect 231674 131200 231730 131209
rect 231674 131135 231730 131144
rect 231214 130248 231270 130257
rect 231214 130183 231270 130192
rect 231676 129940 231728 129946
rect 231676 129882 231728 129888
rect 231688 128897 231716 129882
rect 231768 129736 231820 129742
rect 231768 129678 231820 129684
rect 231780 129305 231808 129678
rect 231766 129296 231822 129305
rect 231766 129231 231822 129240
rect 231674 128888 231730 128897
rect 231674 128823 231730 128832
rect 231122 128344 231178 128353
rect 231122 128279 231178 128288
rect 231768 127968 231820 127974
rect 231766 127936 231768 127945
rect 231820 127936 231822 127945
rect 231766 127871 231822 127880
rect 231122 127800 231178 127809
rect 231122 127735 231178 127744
rect 230938 123176 230994 123185
rect 230938 123111 230994 123120
rect 230756 122120 230808 122126
rect 230756 122062 230808 122068
rect 230572 121236 230624 121242
rect 230572 121178 230624 121184
rect 230584 120329 230612 121178
rect 230768 120737 230796 122062
rect 231136 121689 231164 127735
rect 231306 127664 231362 127673
rect 231306 127599 231362 127608
rect 231122 121680 231178 121689
rect 231122 121615 231178 121624
rect 230754 120728 230810 120737
rect 230754 120663 230810 120672
rect 230570 120320 230626 120329
rect 230570 120255 230626 120264
rect 231214 119232 231270 119241
rect 231214 119167 231270 119176
rect 230940 117292 230992 117298
rect 230940 117234 230992 117240
rect 230756 116748 230808 116754
rect 230756 116690 230808 116696
rect 230768 116113 230796 116690
rect 230952 116521 230980 117234
rect 230938 116512 230994 116521
rect 230938 116447 230994 116456
rect 231122 116512 231178 116521
rect 231122 116447 231178 116456
rect 230754 116104 230810 116113
rect 230754 116039 230810 116048
rect 231032 115864 231084 115870
rect 231032 115806 231084 115812
rect 231044 114617 231072 115806
rect 231030 114608 231086 114617
rect 231030 114543 231086 114552
rect 230572 114504 230624 114510
rect 230572 114446 230624 114452
rect 230584 113257 230612 114446
rect 230570 113248 230626 113257
rect 230570 113183 230626 113192
rect 230940 111104 230992 111110
rect 230940 111046 230992 111052
rect 230572 110900 230624 110906
rect 230572 110842 230624 110848
rect 230584 110809 230612 110842
rect 230570 110800 230626 110809
rect 230570 110735 230626 110744
rect 230756 110016 230808 110022
rect 230756 109958 230808 109964
rect 230768 109857 230796 109958
rect 230754 109848 230810 109857
rect 230754 109783 230810 109792
rect 230756 105596 230808 105602
rect 230756 105538 230808 105544
rect 230572 104168 230624 104174
rect 230572 104110 230624 104116
rect 230584 101425 230612 104110
rect 230664 102060 230716 102066
rect 230664 102002 230716 102008
rect 230676 101833 230704 102002
rect 230662 101824 230718 101833
rect 230662 101759 230718 101768
rect 230570 101416 230626 101425
rect 230570 101351 230626 101360
rect 230664 100700 230716 100706
rect 230664 100642 230716 100648
rect 230676 100473 230704 100642
rect 230662 100464 230718 100473
rect 230662 100399 230718 100408
rect 230768 97617 230796 105538
rect 230952 105233 230980 111046
rect 230938 105224 230994 105233
rect 230938 105159 230994 105168
rect 230940 104848 230992 104854
rect 230940 104790 230992 104796
rect 230952 104281 230980 104790
rect 230938 104272 230994 104281
rect 230938 104207 230994 104216
rect 231136 98977 231164 116447
rect 231228 115161 231256 119167
rect 231320 117201 231348 127599
rect 231766 126984 231822 126993
rect 231766 126919 231768 126928
rect 231820 126919 231822 126928
rect 231768 126890 231820 126896
rect 231492 125588 231544 125594
rect 231492 125530 231544 125536
rect 231504 124545 231532 125530
rect 231768 125520 231820 125526
rect 231768 125462 231820 125468
rect 231780 125089 231808 125462
rect 231766 125080 231822 125089
rect 231766 125015 231822 125024
rect 231490 124536 231546 124545
rect 231490 124471 231546 124480
rect 231768 124160 231820 124166
rect 231766 124128 231768 124137
rect 231820 124128 231822 124137
rect 231676 124092 231728 124098
rect 231766 124063 231822 124072
rect 231676 124034 231728 124040
rect 231688 123593 231716 124034
rect 231674 123584 231730 123593
rect 231674 123519 231730 123528
rect 231768 122800 231820 122806
rect 231768 122742 231820 122748
rect 231780 122233 231808 122742
rect 231766 122224 231822 122233
rect 231766 122159 231822 122168
rect 231584 120760 231636 120766
rect 231584 120702 231636 120708
rect 231492 120080 231544 120086
rect 231492 120022 231544 120028
rect 231504 118969 231532 120022
rect 231490 118960 231546 118969
rect 231490 118895 231546 118904
rect 231492 118720 231544 118726
rect 231492 118662 231544 118668
rect 231400 118652 231452 118658
rect 231400 118594 231452 118600
rect 231412 118017 231440 118594
rect 231398 118008 231454 118017
rect 231398 117943 231454 117952
rect 231306 117192 231362 117201
rect 231306 117127 231362 117136
rect 231504 117042 231532 118662
rect 231320 117014 231532 117042
rect 231214 115152 231270 115161
rect 231214 115087 231270 115096
rect 231320 103737 231348 117014
rect 231596 116906 231624 120702
rect 231766 120048 231822 120057
rect 231766 119983 231822 119992
rect 231780 119377 231808 119983
rect 231766 119368 231822 119377
rect 231766 119303 231822 119312
rect 231768 118584 231820 118590
rect 231768 118526 231820 118532
rect 231780 117473 231808 118526
rect 232516 118425 232544 159015
rect 232608 125497 232636 164863
rect 233436 164393 233464 177278
rect 233516 175976 233568 175982
rect 233516 175918 233568 175924
rect 233422 164384 233478 164393
rect 233422 164319 233478 164328
rect 233528 162858 233556 175918
rect 234632 169794 234660 204138
rect 236828 200864 236880 200870
rect 236828 200806 236880 200812
rect 236090 191176 236146 191185
rect 236090 191111 236146 191120
rect 234710 181656 234766 181665
rect 234710 181591 234766 181600
rect 234620 169788 234672 169794
rect 234620 169730 234672 169736
rect 233884 168564 233936 168570
rect 233884 168506 233936 168512
rect 233516 162852 233568 162858
rect 233516 162794 233568 162800
rect 232688 149728 232740 149734
rect 232688 149670 232740 149676
rect 232700 136610 232728 149670
rect 233896 148850 233924 168506
rect 234068 166116 234120 166122
rect 234068 166058 234120 166064
rect 234080 155854 234108 166058
rect 234160 160132 234212 160138
rect 234160 160074 234212 160080
rect 234068 155848 234120 155854
rect 234068 155790 234120 155796
rect 233974 155000 234030 155009
rect 233974 154935 234030 154944
rect 233884 148844 233936 148850
rect 233884 148786 233936 148792
rect 232872 148368 232924 148374
rect 232872 148310 232924 148316
rect 232688 136604 232740 136610
rect 232688 136546 232740 136552
rect 232594 125488 232650 125497
rect 232594 125423 232650 125432
rect 232778 124672 232834 124681
rect 232778 124607 232834 124616
rect 232502 118416 232558 118425
rect 232502 118351 232558 118360
rect 231766 117464 231822 117473
rect 231766 117399 231822 117408
rect 231412 116878 231624 116906
rect 231412 111353 231440 116878
rect 231768 115932 231820 115938
rect 231768 115874 231820 115880
rect 231780 115569 231808 115874
rect 231766 115560 231822 115569
rect 231766 115495 231822 115504
rect 231584 114368 231636 114374
rect 231584 114310 231636 114316
rect 231596 113665 231624 114310
rect 231582 113656 231638 113665
rect 231582 113591 231638 113600
rect 232686 113520 232742 113529
rect 232686 113455 232742 113464
rect 231768 113144 231820 113150
rect 231768 113086 231820 113092
rect 231676 113076 231728 113082
rect 231676 113018 231728 113024
rect 231688 112305 231716 113018
rect 231780 112713 231808 113086
rect 231766 112704 231822 112713
rect 231766 112639 231822 112648
rect 232502 112432 232558 112441
rect 232502 112367 232558 112376
rect 231674 112296 231730 112305
rect 231674 112231 231730 112240
rect 231398 111344 231454 111353
rect 231398 111279 231454 111288
rect 231768 110424 231820 110430
rect 231768 110366 231820 110372
rect 231780 109449 231808 110366
rect 231766 109440 231822 109449
rect 231766 109375 231822 109384
rect 231768 108996 231820 109002
rect 231768 108938 231820 108944
rect 231492 108928 231544 108934
rect 231492 108870 231544 108876
rect 231504 107953 231532 108870
rect 231780 108497 231808 108938
rect 231766 108488 231822 108497
rect 231766 108423 231822 108432
rect 231490 107944 231546 107953
rect 231490 107879 231546 107888
rect 231768 107636 231820 107642
rect 231768 107578 231820 107584
rect 231492 107568 231544 107574
rect 231492 107510 231544 107516
rect 231504 106593 231532 107510
rect 231780 107137 231808 107578
rect 231766 107128 231822 107137
rect 231766 107063 231822 107072
rect 231490 106584 231546 106593
rect 231490 106519 231546 106528
rect 231768 106072 231820 106078
rect 231768 106014 231820 106020
rect 231780 105641 231808 106014
rect 231766 105632 231822 105641
rect 231766 105567 231822 105576
rect 231306 103728 231362 103737
rect 231306 103663 231362 103672
rect 231768 103488 231820 103494
rect 231768 103430 231820 103436
rect 231492 103420 231544 103426
rect 231492 103362 231544 103368
rect 231504 102377 231532 103362
rect 231780 102785 231808 103430
rect 231766 102776 231822 102785
rect 231766 102711 231822 102720
rect 231490 102368 231546 102377
rect 231490 102303 231546 102312
rect 231676 102128 231728 102134
rect 231676 102070 231728 102076
rect 231306 101552 231362 101561
rect 231306 101487 231362 101496
rect 231122 98968 231178 98977
rect 231122 98903 231178 98912
rect 231216 98048 231268 98054
rect 231216 97990 231268 97996
rect 230754 97608 230810 97617
rect 230754 97543 230810 97552
rect 231122 97064 231178 97073
rect 231122 96999 231178 97008
rect 230570 96656 230626 96665
rect 230570 96591 230626 96600
rect 230478 96248 230534 96257
rect 230478 96183 230534 96192
rect 230492 95334 230520 96183
rect 230480 95328 230532 95334
rect 230480 95270 230532 95276
rect 229926 93871 229982 93880
rect 230020 93900 230072 93906
rect 230020 93842 230072 93848
rect 230584 90953 230612 96591
rect 230570 90944 230626 90953
rect 230570 90879 230626 90888
rect 229742 76664 229798 76673
rect 229742 76599 229798 76608
rect 228364 37936 228416 37942
rect 228364 37878 228416 37884
rect 231136 28286 231164 96999
rect 231228 84930 231256 97990
rect 231320 91798 231348 101487
rect 231688 100881 231716 102070
rect 231674 100872 231730 100881
rect 231674 100807 231730 100816
rect 231674 100736 231730 100745
rect 231674 100671 231730 100680
rect 231688 99929 231716 100671
rect 231768 100632 231820 100638
rect 231768 100574 231820 100580
rect 231674 99920 231730 99929
rect 231674 99855 231730 99864
rect 231780 99521 231808 100574
rect 231766 99512 231822 99521
rect 231766 99447 231822 99456
rect 231308 91792 231360 91798
rect 231308 91734 231360 91740
rect 231216 84924 231268 84930
rect 231216 84866 231268 84872
rect 231124 28280 231176 28286
rect 231124 28222 231176 28228
rect 227076 14476 227128 14482
rect 227076 14418 227128 14424
rect 226984 7676 227036 7682
rect 226984 7618 227036 7624
rect 232516 4826 232544 112367
rect 232596 95328 232648 95334
rect 232596 95270 232648 95276
rect 232504 4820 232556 4826
rect 232504 4762 232556 4768
rect 232608 4214 232636 95270
rect 232700 54505 232728 113455
rect 232792 87718 232820 124607
rect 232884 110906 232912 148310
rect 233884 141364 233936 141370
rect 233884 141306 233936 141312
rect 233896 140729 233924 141306
rect 233882 140720 233938 140729
rect 233882 140655 233938 140664
rect 233884 138032 233936 138038
rect 233884 137974 233936 137980
rect 232872 110900 232924 110906
rect 232872 110842 232924 110848
rect 232780 87712 232832 87718
rect 232780 87654 232832 87660
rect 232686 54496 232742 54505
rect 232686 54431 232742 54440
rect 233896 14550 233924 137974
rect 233988 114374 234016 154935
rect 234066 145480 234122 145489
rect 234066 145415 234122 145424
rect 233976 114368 234028 114374
rect 233976 114310 234028 114316
rect 233974 105360 234030 105369
rect 233974 105295 234030 105304
rect 233884 14544 233936 14550
rect 233884 14486 233936 14492
rect 232596 4208 232648 4214
rect 232596 4150 232648 4156
rect 218704 2168 218756 2174
rect 218704 2110 218756 2116
rect 220176 2168 220228 2174
rect 220176 2110 220228 2116
rect 233988 2106 234016 105295
rect 234080 103329 234108 145415
rect 234172 121242 234200 160074
rect 234250 153776 234306 153785
rect 234250 153711 234306 153720
rect 234264 143478 234292 153711
rect 234724 150958 234752 181591
rect 234802 180296 234858 180305
rect 234802 180231 234858 180240
rect 234816 169454 234844 180231
rect 235998 180160 236054 180169
rect 235998 180095 236054 180104
rect 235446 175128 235502 175137
rect 235446 175063 235502 175072
rect 234896 169788 234948 169794
rect 234896 169730 234948 169736
rect 234804 169448 234856 169454
rect 234804 169390 234856 169396
rect 234908 166734 234936 169730
rect 234896 166728 234948 166734
rect 234896 166670 234948 166676
rect 235354 166424 235410 166433
rect 235354 166359 235410 166368
rect 235264 165640 235316 165646
rect 235264 165582 235316 165588
rect 234712 150952 234764 150958
rect 234712 150894 234764 150900
rect 234252 143472 234304 143478
rect 234252 143414 234304 143420
rect 235276 126886 235304 165582
rect 235368 138922 235396 166359
rect 235460 165238 235488 175063
rect 235448 165232 235500 165238
rect 235448 165174 235500 165180
rect 236012 158642 236040 180095
rect 236104 175273 236132 191111
rect 236182 175808 236238 175817
rect 236182 175743 236238 175752
rect 236090 175264 236146 175273
rect 236090 175199 236146 175208
rect 236196 167113 236224 175743
rect 236644 173936 236696 173942
rect 236644 173878 236696 173884
rect 236182 167104 236238 167113
rect 236182 167039 236238 167048
rect 236000 158636 236052 158642
rect 236000 158578 236052 158584
rect 235540 155984 235592 155990
rect 235540 155926 235592 155932
rect 235448 150476 235500 150482
rect 235448 150418 235500 150424
rect 235356 138916 235408 138922
rect 235356 138858 235408 138864
rect 235356 135312 235408 135318
rect 235356 135254 235408 135260
rect 235264 126880 235316 126886
rect 235264 126822 235316 126828
rect 234160 121236 234212 121242
rect 234160 121178 234212 121184
rect 234158 117872 234214 117881
rect 234158 117807 234214 117816
rect 234066 103320 234122 103329
rect 234066 103255 234122 103264
rect 234172 93226 234200 117807
rect 235262 115968 235318 115977
rect 235262 115903 235318 115912
rect 234160 93220 234212 93226
rect 234160 93162 234212 93168
rect 235276 58585 235304 115903
rect 235368 90438 235396 135254
rect 235460 110022 235488 150418
rect 235552 116754 235580 155926
rect 236656 135930 236684 173878
rect 236840 167142 236868 200806
rect 236828 167136 236880 167142
rect 236828 167078 236880 167084
rect 236736 167068 236788 167074
rect 236736 167010 236788 167016
rect 236644 135924 236696 135930
rect 236644 135866 236696 135872
rect 236642 128752 236698 128761
rect 236642 128687 236698 128696
rect 235540 116748 235592 116754
rect 235540 116690 235592 116696
rect 235448 110016 235500 110022
rect 235448 109958 235500 109964
rect 235540 109064 235592 109070
rect 235540 109006 235592 109012
rect 235356 90432 235408 90438
rect 235356 90374 235408 90380
rect 235552 73953 235580 109006
rect 235538 73944 235594 73953
rect 235538 73879 235594 73888
rect 235262 58576 235318 58585
rect 235262 58511 235318 58520
rect 236656 36553 236684 128687
rect 236748 127974 236776 167010
rect 237392 152998 237420 211754
rect 237472 181484 237524 181490
rect 237472 181426 237524 181432
rect 237484 168094 237512 181426
rect 238036 169794 238064 234586
rect 238312 223514 238340 240244
rect 238864 234614 238892 240244
rect 239232 240009 239260 240244
rect 239218 240000 239274 240009
rect 239218 239935 239274 239944
rect 239404 237244 239456 237250
rect 239404 237186 239456 237192
rect 239220 236700 239272 236706
rect 239220 236642 239272 236648
rect 239232 235657 239260 236642
rect 239416 235929 239444 237186
rect 239402 235920 239458 235929
rect 239402 235855 239458 235864
rect 239218 235648 239274 235657
rect 239218 235583 239274 235592
rect 238864 234586 238984 234614
rect 238300 223508 238352 223514
rect 238300 223450 238352 223456
rect 238116 200796 238168 200802
rect 238116 200738 238168 200744
rect 238128 191146 238156 200738
rect 238760 199436 238812 199442
rect 238760 199378 238812 199384
rect 238116 191140 238168 191146
rect 238116 191082 238168 191088
rect 238024 169788 238076 169794
rect 238024 169730 238076 169736
rect 238300 169788 238352 169794
rect 238300 169730 238352 169736
rect 238024 168428 238076 168434
rect 238024 168370 238076 168376
rect 237472 168088 237524 168094
rect 237472 168030 237524 168036
rect 237380 152992 237432 152998
rect 237380 152934 237432 152940
rect 236920 152516 236972 152522
rect 236920 152458 236972 152464
rect 236828 144220 236880 144226
rect 236828 144162 236880 144168
rect 236736 127968 236788 127974
rect 236736 127910 236788 127916
rect 236736 116000 236788 116006
rect 236736 115942 236788 115948
rect 236748 59945 236776 115942
rect 236840 104854 236868 144162
rect 236932 117298 236960 152458
rect 238036 129946 238064 168370
rect 238116 154624 238168 154630
rect 238116 154566 238168 154572
rect 238024 129940 238076 129946
rect 238024 129882 238076 129888
rect 238022 117464 238078 117473
rect 238022 117399 238078 117408
rect 236920 117292 236972 117298
rect 236920 117234 236972 117240
rect 236828 104848 236880 104854
rect 236828 104790 236880 104796
rect 236734 59936 236790 59945
rect 236734 59871 236790 59880
rect 236642 36544 236698 36553
rect 236642 36479 236698 36488
rect 238036 11762 238064 117399
rect 238128 115870 238156 154566
rect 238208 147688 238260 147694
rect 238208 147630 238260 147636
rect 238116 115864 238168 115870
rect 238116 115806 238168 115812
rect 238220 106078 238248 147630
rect 238312 144906 238340 169730
rect 238772 168570 238800 199378
rect 238956 198694 238984 234586
rect 239784 230489 239812 240244
rect 240336 238678 240364 240244
rect 240324 238672 240376 238678
rect 240324 238614 240376 238620
rect 240704 236774 240732 240244
rect 241256 239465 241284 240244
rect 241242 239456 241298 239465
rect 241242 239391 241298 239400
rect 240784 238672 240836 238678
rect 240784 238614 240836 238620
rect 240692 236768 240744 236774
rect 240692 236710 240744 236716
rect 240704 235929 240732 236710
rect 240690 235920 240746 235929
rect 240690 235855 240746 235864
rect 239770 230480 239826 230489
rect 239770 230415 239826 230424
rect 240138 213888 240194 213897
rect 240138 213823 240194 213832
rect 238944 198688 238996 198694
rect 238944 198630 238996 198636
rect 238852 189780 238904 189786
rect 238852 189722 238904 189728
rect 238760 168564 238812 168570
rect 238760 168506 238812 168512
rect 238864 165753 238892 189722
rect 238944 185632 238996 185638
rect 238944 185574 238996 185580
rect 238956 166122 238984 185574
rect 239588 175296 239640 175302
rect 239588 175238 239640 175244
rect 238944 166116 238996 166122
rect 238944 166058 238996 166064
rect 238850 165744 238906 165753
rect 238850 165679 238906 165688
rect 238300 144900 238352 144906
rect 238300 144842 238352 144848
rect 238392 142860 238444 142866
rect 238392 142802 238444 142808
rect 238300 120148 238352 120154
rect 238300 120090 238352 120096
rect 238208 106072 238260 106078
rect 238208 106014 238260 106020
rect 238114 105496 238170 105505
rect 238114 105431 238170 105440
rect 238128 21418 238156 105431
rect 238206 104000 238262 104009
rect 238206 103935 238262 103944
rect 238220 39370 238248 103935
rect 238312 82142 238340 120090
rect 238404 118726 238432 142802
rect 239402 137184 239458 137193
rect 239402 137119 239458 137128
rect 238392 118720 238444 118726
rect 238392 118662 238444 118668
rect 238300 82136 238352 82142
rect 238300 82078 238352 82084
rect 239416 39438 239444 137119
rect 239496 133952 239548 133958
rect 239496 133894 239548 133900
rect 239508 67017 239536 133894
rect 239600 116521 239628 175238
rect 240152 172446 240180 213823
rect 240796 204105 240824 238614
rect 241256 235958 241284 239391
rect 241808 237386 241836 240244
rect 241796 237380 241848 237386
rect 241796 237322 241848 237328
rect 242176 237318 242204 240244
rect 242256 237380 242308 237386
rect 242256 237322 242308 237328
rect 242164 237312 242216 237318
rect 242164 237254 242216 237260
rect 241244 235952 241296 235958
rect 241244 235894 241296 235900
rect 240876 235612 240928 235618
rect 240876 235554 240928 235560
rect 240888 213897 240916 235554
rect 241426 215928 241482 215937
rect 241426 215863 241482 215872
rect 240874 213888 240930 213897
rect 240874 213823 240930 213832
rect 240782 204096 240838 204105
rect 240782 204031 240838 204040
rect 241440 198014 241468 215863
rect 241428 198008 241480 198014
rect 241428 197950 241480 197956
rect 241612 188420 241664 188426
rect 241612 188362 241664 188368
rect 240230 186960 240286 186969
rect 240230 186895 240286 186904
rect 240244 175273 240272 186895
rect 240322 183152 240378 183161
rect 240322 183087 240378 183096
rect 240230 175264 240286 175273
rect 240230 175199 240286 175208
rect 240140 172440 240192 172446
rect 240140 172382 240192 172388
rect 239772 167136 239824 167142
rect 239772 167078 239824 167084
rect 239678 166288 239734 166297
rect 239678 166223 239734 166232
rect 239692 129742 239720 166223
rect 239784 134570 239812 167078
rect 240336 163441 240364 183087
rect 241520 180124 241572 180130
rect 241520 180066 241572 180072
rect 240414 177440 240470 177449
rect 240414 177375 240470 177384
rect 240322 163432 240378 163441
rect 240322 163367 240378 163376
rect 240428 155242 240456 177375
rect 240966 170368 241022 170377
rect 240966 170303 241022 170312
rect 240784 164280 240836 164286
rect 240784 164222 240836 164228
rect 240416 155236 240468 155242
rect 240416 155178 240468 155184
rect 239772 134564 239824 134570
rect 239772 134506 239824 134512
rect 239680 129736 239732 129742
rect 239680 129678 239732 129684
rect 240796 125526 240824 164222
rect 240980 160002 241008 170303
rect 240968 159996 241020 160002
rect 240968 159938 241020 159944
rect 240876 158772 240928 158778
rect 240876 158714 240928 158720
rect 240784 125520 240836 125526
rect 240784 125462 240836 125468
rect 239678 124808 239734 124817
rect 239678 124743 239734 124752
rect 239586 116512 239642 116521
rect 239586 116447 239642 116456
rect 239692 89078 239720 124743
rect 240782 122088 240838 122097
rect 240782 122023 240838 122032
rect 239680 89072 239732 89078
rect 239680 89014 239732 89020
rect 239494 67008 239550 67017
rect 239494 66943 239550 66952
rect 239404 39432 239456 39438
rect 239404 39374 239456 39380
rect 238208 39364 238260 39370
rect 238208 39306 238260 39312
rect 240796 25634 240824 122023
rect 240888 120086 240916 158714
rect 240968 157412 241020 157418
rect 240968 157354 241020 157360
rect 240876 120080 240928 120086
rect 240876 120022 240928 120028
rect 240980 118590 241008 157354
rect 241532 140185 241560 180066
rect 241624 154494 241652 188362
rect 241612 154488 241664 154494
rect 241612 154430 241664 154436
rect 242176 143993 242204 237254
rect 242268 180169 242296 237322
rect 242728 237017 242756 240244
rect 242714 237008 242770 237017
rect 242714 236943 242770 236952
rect 243280 235618 243308 240244
rect 243542 238504 243598 238513
rect 243648 238490 243676 240244
rect 243598 238462 243676 238490
rect 243542 238439 243598 238448
rect 243268 235612 243320 235618
rect 243268 235554 243320 235560
rect 243556 227730 243584 238439
rect 244016 234614 244044 244831
rect 243924 234586 244044 234614
rect 243544 227724 243596 227730
rect 243544 227666 243596 227672
rect 242348 199504 242400 199510
rect 242348 199446 242400 199452
rect 242254 180160 242310 180169
rect 242254 180095 242310 180104
rect 242360 173913 242388 199446
rect 243924 190466 243952 234586
rect 244292 218006 244320 250815
rect 244384 222154 244412 255167
rect 244476 253881 244504 284310
rect 244568 271017 244596 301446
rect 244648 289944 244700 289950
rect 244648 289886 244700 289892
rect 244554 271008 244610 271017
rect 244554 270943 244610 270952
rect 244462 253872 244518 253881
rect 244462 253807 244518 253816
rect 244660 253065 244688 289886
rect 245028 289882 245056 326402
rect 246120 318164 246172 318170
rect 246120 318106 246172 318112
rect 246026 297392 246082 297401
rect 246026 297327 246082 297336
rect 245016 289876 245068 289882
rect 245016 289818 245068 289824
rect 245936 289876 245988 289882
rect 245936 289818 245988 289824
rect 245842 289096 245898 289105
rect 245842 289031 245898 289040
rect 245856 287054 245884 289031
rect 245764 287026 245884 287054
rect 245660 283960 245712 283966
rect 245660 283902 245712 283908
rect 245672 281081 245700 283902
rect 245764 282962 245792 287026
rect 245948 283966 245976 289818
rect 245936 283960 245988 283966
rect 245936 283902 245988 283908
rect 245936 283824 245988 283830
rect 245934 283792 245936 283801
rect 245988 283792 245990 283801
rect 245934 283727 245990 283736
rect 245764 282934 245884 282962
rect 245752 282804 245804 282810
rect 245752 282746 245804 282752
rect 245764 281625 245792 282746
rect 245750 281616 245806 281625
rect 245750 281551 245806 281560
rect 245658 281072 245714 281081
rect 245658 281007 245714 281016
rect 245660 280832 245712 280838
rect 245660 280774 245712 280780
rect 245672 280265 245700 280774
rect 245658 280256 245714 280265
rect 245658 280191 245714 280200
rect 245658 280120 245714 280129
rect 245658 280055 245714 280064
rect 245476 253904 245528 253910
rect 245474 253872 245476 253881
rect 245528 253872 245530 253881
rect 245474 253807 245530 253816
rect 244646 253056 244702 253065
rect 244646 252991 244702 253000
rect 245474 253056 245530 253065
rect 245474 252991 245530 253000
rect 245488 252618 245516 252991
rect 245476 252612 245528 252618
rect 245476 252554 245528 252560
rect 244556 247716 244608 247722
rect 244556 247658 244608 247664
rect 244462 247344 244518 247353
rect 244462 247279 244518 247288
rect 244476 233209 244504 247279
rect 244568 240038 244596 247658
rect 245672 246537 245700 280055
rect 245752 279540 245804 279546
rect 245752 279482 245804 279488
rect 245764 278905 245792 279482
rect 245750 278896 245806 278905
rect 245750 278831 245806 278840
rect 245752 278724 245804 278730
rect 245752 278666 245804 278672
rect 245764 277545 245792 278666
rect 245750 277536 245806 277545
rect 245750 277471 245806 277480
rect 245752 276072 245804 276078
rect 245752 276014 245804 276020
rect 245764 270586 245792 276014
rect 245856 275913 245884 282934
rect 245934 282432 245990 282441
rect 245934 282367 245990 282376
rect 245948 281586 245976 282367
rect 245936 281580 245988 281586
rect 245936 281522 245988 281528
rect 245936 279472 245988 279478
rect 245934 279440 245936 279449
rect 245988 279440 245990 279449
rect 245934 279375 245990 279384
rect 246040 277394 246068 297327
rect 245948 277366 246068 277394
rect 245842 275904 245898 275913
rect 245842 275839 245898 275848
rect 245948 274553 245976 277366
rect 246132 276729 246160 318106
rect 246946 283248 247002 283257
rect 247052 283234 247080 332551
rect 247132 319456 247184 319462
rect 247132 319398 247184 319404
rect 247002 283206 247080 283234
rect 246946 283183 247002 283192
rect 246118 276720 246174 276729
rect 246118 276655 246120 276664
rect 246172 276655 246174 276664
rect 246120 276626 246172 276632
rect 246132 276595 246160 276626
rect 245934 274544 245990 274553
rect 245934 274479 245990 274488
rect 245948 273970 245976 274479
rect 245936 273964 245988 273970
rect 245936 273906 245988 273912
rect 245934 273728 245990 273737
rect 245934 273663 245990 273672
rect 245844 273216 245896 273222
rect 245844 273158 245896 273164
rect 245856 272377 245884 273158
rect 245842 272368 245898 272377
rect 245842 272303 245898 272312
rect 245948 271182 245976 273663
rect 246946 273184 247002 273193
rect 246946 273119 247002 273128
rect 245936 271176 245988 271182
rect 245936 271118 245988 271124
rect 245764 270558 245884 270586
rect 245752 270496 245804 270502
rect 245752 270438 245804 270444
rect 245764 270201 245792 270438
rect 245750 270192 245806 270201
rect 245750 270127 245806 270136
rect 245856 269822 245884 270558
rect 245844 269816 245896 269822
rect 245844 269758 245896 269764
rect 245856 269657 245884 269758
rect 245842 269648 245898 269657
rect 245842 269583 245898 269592
rect 246764 268388 246816 268394
rect 246764 268330 246816 268336
rect 246210 268016 246266 268025
rect 246210 267951 246266 267960
rect 245934 267472 245990 267481
rect 245934 267407 245990 267416
rect 245948 266393 245976 267407
rect 245934 266384 245990 266393
rect 245934 266319 245990 266328
rect 246224 266257 246252 267951
rect 246210 266248 246266 266257
rect 246210 266183 246266 266192
rect 245934 265840 245990 265849
rect 245934 265775 245990 265784
rect 245948 265674 245976 265775
rect 245936 265668 245988 265674
rect 245936 265610 245988 265616
rect 246776 265305 246804 268330
rect 246960 267578 246988 273119
rect 246948 267572 247000 267578
rect 246948 267514 247000 267520
rect 246762 265296 246818 265305
rect 246762 265231 246818 265240
rect 245844 264920 245896 264926
rect 245844 264862 245896 264868
rect 245856 263945 245884 264862
rect 245842 263936 245898 263945
rect 245842 263871 245898 263880
rect 245750 263120 245806 263129
rect 245750 263055 245806 263064
rect 245764 258074 245792 263055
rect 245934 262304 245990 262313
rect 245934 262239 245936 262248
rect 245988 262239 245990 262248
rect 245936 262210 245988 262216
rect 246396 261520 246448 261526
rect 246396 261462 246448 261468
rect 246408 260953 246436 261462
rect 246394 260944 246450 260953
rect 246394 260879 246450 260888
rect 245844 260840 245896 260846
rect 245844 260782 245896 260788
rect 245856 260137 245884 260782
rect 245842 260128 245898 260137
rect 245842 260063 245898 260072
rect 245934 259584 245990 259593
rect 245934 259519 245990 259528
rect 245948 259486 245976 259519
rect 245936 259480 245988 259486
rect 245936 259422 245988 259428
rect 245844 259412 245896 259418
rect 245844 259354 245896 259360
rect 245856 258233 245884 259354
rect 245936 259344 245988 259350
rect 245936 259286 245988 259292
rect 245948 258777 245976 259286
rect 245934 258768 245990 258777
rect 245934 258703 245990 258712
rect 245842 258224 245898 258233
rect 245842 258159 245898 258168
rect 245764 258046 245884 258074
rect 245750 250336 245806 250345
rect 245750 250271 245806 250280
rect 245764 249830 245792 250271
rect 245752 249824 245804 249830
rect 245752 249766 245804 249772
rect 245658 246528 245714 246537
rect 245658 246463 245714 246472
rect 245672 245721 245700 246463
rect 245750 245984 245806 245993
rect 245750 245919 245806 245928
rect 245658 245712 245714 245721
rect 245764 245682 245792 245919
rect 245658 245647 245714 245656
rect 245752 245676 245804 245682
rect 245752 245618 245804 245624
rect 245750 244624 245806 244633
rect 245750 244559 245806 244568
rect 245658 240816 245714 240825
rect 245658 240751 245714 240760
rect 245672 240242 245700 240751
rect 245660 240236 245712 240242
rect 245660 240178 245712 240184
rect 244556 240032 244608 240038
rect 244556 239974 244608 239980
rect 244462 233200 244518 233209
rect 244462 233135 244518 233144
rect 244372 222148 244424 222154
rect 244372 222090 244424 222096
rect 244280 218000 244332 218006
rect 244280 217942 244332 217948
rect 244186 192672 244242 192681
rect 244186 192607 244242 192616
rect 243912 190460 243964 190466
rect 243912 190402 243964 190408
rect 243924 189145 243952 190402
rect 243910 189136 243966 189145
rect 243910 189071 243966 189080
rect 242992 186992 243044 186998
rect 242992 186934 243044 186940
rect 242900 185768 242952 185774
rect 242900 185710 242952 185716
rect 242346 173904 242402 173913
rect 242346 173839 242402 173848
rect 242254 162888 242310 162897
rect 242254 162823 242310 162832
rect 242162 143984 242218 143993
rect 242162 143919 242218 143928
rect 241518 140176 241574 140185
rect 241518 140111 241574 140120
rect 242162 136912 242218 136921
rect 242162 136847 242218 136856
rect 241060 127628 241112 127634
rect 241060 127570 241112 127576
rect 240968 118584 241020 118590
rect 240968 118526 241020 118532
rect 240876 102196 240928 102202
rect 240876 102138 240928 102144
rect 240888 77897 240916 102138
rect 241072 94489 241100 127570
rect 241152 119400 241204 119406
rect 241152 119342 241204 119348
rect 241164 103426 241192 119342
rect 241152 103420 241204 103426
rect 241152 103362 241204 103368
rect 241058 94480 241114 94489
rect 241058 94415 241114 94424
rect 240874 77888 240930 77897
rect 240874 77823 240930 77832
rect 240784 25628 240836 25634
rect 240784 25570 240836 25576
rect 238116 21412 238168 21418
rect 238116 21354 238168 21360
rect 242176 13190 242204 136847
rect 242268 122806 242296 162823
rect 242912 154562 242940 185710
rect 243004 160750 243032 186934
rect 244200 184210 244228 192607
rect 244188 184204 244240 184210
rect 244188 184146 244240 184152
rect 243544 168496 243596 168502
rect 243544 168438 243596 168444
rect 242992 160744 243044 160750
rect 242992 160686 243044 160692
rect 242900 154556 242952 154562
rect 242900 154498 242952 154504
rect 242346 143984 242402 143993
rect 242346 143919 242402 143928
rect 242256 122800 242308 122806
rect 242256 122742 242308 122748
rect 242256 114572 242308 114578
rect 242256 114514 242308 114520
rect 242164 13184 242216 13190
rect 242164 13126 242216 13132
rect 242268 13122 242296 114514
rect 242360 102066 242388 143919
rect 242438 142760 242494 142769
rect 242438 142695 242494 142704
rect 242452 104689 242480 142695
rect 243556 131102 243584 168438
rect 243912 161492 243964 161498
rect 243912 161434 243964 161440
rect 243728 153264 243780 153270
rect 243728 153206 243780 153212
rect 243636 135380 243688 135386
rect 243636 135322 243688 135328
rect 243544 131096 243596 131102
rect 243544 131038 243596 131044
rect 243542 116104 243598 116113
rect 243542 116039 243598 116048
rect 242438 104680 242494 104689
rect 242438 104615 242494 104624
rect 242348 102060 242400 102066
rect 242348 102002 242400 102008
rect 242348 98116 242400 98122
rect 242348 98058 242400 98064
rect 242360 69737 242388 98058
rect 242346 69728 242402 69737
rect 242346 69663 242402 69672
rect 242256 13116 242308 13122
rect 242256 13058 242308 13064
rect 238024 11756 238076 11762
rect 238024 11698 238076 11704
rect 243556 10334 243584 116039
rect 243648 62937 243676 135322
rect 243740 113082 243768 153206
rect 243820 128376 243872 128382
rect 243820 128318 243872 128324
rect 243728 113076 243780 113082
rect 243728 113018 243780 113024
rect 243832 93158 243860 128318
rect 243924 127809 243952 161434
rect 244292 157282 244320 217942
rect 244384 164150 244412 222090
rect 244464 210520 244516 210526
rect 244464 210462 244516 210468
rect 244476 166433 244504 210462
rect 245764 208282 245792 244559
rect 245856 227050 245884 258046
rect 246026 257408 246082 257417
rect 246026 257343 246082 257352
rect 246040 256766 246068 257343
rect 246028 256760 246080 256766
rect 246028 256702 246080 256708
rect 245936 256692 245988 256698
rect 245936 256634 245988 256640
rect 245948 256601 245976 256634
rect 245934 256592 245990 256601
rect 245934 256527 245990 256536
rect 245936 255264 245988 255270
rect 245936 255206 245988 255212
rect 245948 254425 245976 255206
rect 246948 254584 247000 254590
rect 246948 254526 247000 254532
rect 245934 254416 245990 254425
rect 245934 254351 245990 254360
rect 245936 252544 245988 252550
rect 245936 252486 245988 252492
rect 245948 251705 245976 252486
rect 245934 251696 245990 251705
rect 245934 251631 245990 251640
rect 245936 249552 245988 249558
rect 245934 249520 245936 249529
rect 245988 249520 245990 249529
rect 245934 249455 245990 249464
rect 245934 248704 245990 248713
rect 245934 248639 245936 248648
rect 245988 248639 245990 248648
rect 245936 248610 245988 248616
rect 246960 248169 246988 254526
rect 246946 248160 247002 248169
rect 246946 248095 247002 248104
rect 246960 247790 246988 248095
rect 246948 247784 247000 247790
rect 246948 247726 247000 247732
rect 246118 245712 246174 245721
rect 246118 245647 246174 245656
rect 245934 240272 245990 240281
rect 245934 240207 245990 240216
rect 245948 227633 245976 240207
rect 246132 238754 246160 245647
rect 246394 242448 246450 242457
rect 246394 242383 246450 242392
rect 246408 241534 246436 242383
rect 246396 241528 246448 241534
rect 246302 241496 246358 241505
rect 246396 241470 246448 241476
rect 246302 241431 246358 241440
rect 246040 238726 246160 238754
rect 245934 227624 245990 227633
rect 245934 227559 245990 227568
rect 245844 227044 245896 227050
rect 245844 226986 245896 226992
rect 245936 209840 245988 209846
rect 245936 209782 245988 209788
rect 245752 208276 245804 208282
rect 245752 208218 245804 208224
rect 245660 202156 245712 202162
rect 245660 202098 245712 202104
rect 244556 184272 244608 184278
rect 244556 184214 244608 184220
rect 244462 166424 244518 166433
rect 244462 166359 244518 166368
rect 244372 164144 244424 164150
rect 244372 164086 244424 164092
rect 244280 157276 244332 157282
rect 244280 157218 244332 157224
rect 244568 146985 244596 184214
rect 245108 165708 245160 165714
rect 245108 165650 245160 165656
rect 245016 162920 245068 162926
rect 245016 162862 245068 162868
rect 244924 149116 244976 149122
rect 244924 149058 244976 149064
rect 244554 146976 244610 146985
rect 244554 146911 244610 146920
rect 243910 127800 243966 127809
rect 243910 127735 243966 127744
rect 244936 108934 244964 149058
rect 245028 124098 245056 162862
rect 245120 127702 245148 165650
rect 245198 146976 245254 146985
rect 245198 146911 245254 146920
rect 245108 127696 245160 127702
rect 245108 127638 245160 127644
rect 245016 124092 245068 124098
rect 245016 124034 245068 124040
rect 245016 110492 245068 110498
rect 245016 110434 245068 110440
rect 244924 108928 244976 108934
rect 244924 108870 244976 108876
rect 243820 93152 243872 93158
rect 243820 93094 243872 93100
rect 244922 91896 244978 91905
rect 244922 91831 244978 91840
rect 243634 62928 243690 62937
rect 243634 62863 243690 62872
rect 244280 60104 244332 60110
rect 244280 60046 244332 60052
rect 244292 16574 244320 60046
rect 244292 16546 244872 16574
rect 243544 10328 243596 10334
rect 243544 10270 243596 10276
rect 242898 9072 242954 9081
rect 242898 9007 242954 9016
rect 239310 5672 239366 5681
rect 239310 5607 239366 5616
rect 235816 4208 235868 4214
rect 235816 4150 235868 4156
rect 233976 2100 234028 2106
rect 233976 2042 234028 2048
rect 235828 480 235856 4150
rect 239324 480 239352 5607
rect 241704 5568 241756 5574
rect 241704 5510 241756 5516
rect 240508 2168 240560 2174
rect 240508 2110 240560 2116
rect 240520 480 240548 2110
rect 241716 480 241744 5510
rect 242912 480 242940 9007
rect 244094 7576 244150 7585
rect 244094 7511 244150 7520
rect 244108 480 244136 7511
rect 244844 3482 244872 16546
rect 244936 5681 244964 91831
rect 245028 55894 245056 110434
rect 245106 109440 245162 109449
rect 245106 109375 245162 109384
rect 245120 60042 245148 109375
rect 245212 108905 245240 146911
rect 245672 136377 245700 202098
rect 245764 200870 245792 208218
rect 245752 200864 245804 200870
rect 245752 200806 245804 200812
rect 245844 195288 245896 195294
rect 245844 195230 245896 195236
rect 245856 146266 245884 195230
rect 245948 151774 245976 209782
rect 246040 197169 246068 238726
rect 246316 237250 246344 241431
rect 246304 237244 246356 237250
rect 246304 237186 246356 237192
rect 246026 197160 246082 197169
rect 246026 197095 246082 197104
rect 246672 170400 246724 170406
rect 246672 170342 246724 170348
rect 245936 151768 245988 151774
rect 245936 151710 245988 151716
rect 246302 150512 246358 150521
rect 246302 150447 246358 150456
rect 245844 146260 245896 146266
rect 245844 146202 245896 146208
rect 245658 136368 245714 136377
rect 245658 136303 245714 136312
rect 245198 108896 245254 108905
rect 245198 108831 245254 108840
rect 245200 105664 245252 105670
rect 245200 105606 245252 105612
rect 245212 91866 245240 105606
rect 245200 91860 245252 91866
rect 245200 91802 245252 91808
rect 245108 60036 245160 60042
rect 245108 59978 245160 59984
rect 245016 55888 245068 55894
rect 245016 55830 245068 55836
rect 244922 5672 244978 5681
rect 244922 5607 244978 5616
rect 246316 5574 246344 150447
rect 246580 144968 246632 144974
rect 246580 144910 246632 144916
rect 246394 139496 246450 139505
rect 246394 139431 246450 139440
rect 246408 51746 246436 139431
rect 246592 103494 246620 144910
rect 246684 140729 246712 170342
rect 247052 153785 247080 283206
rect 247144 273193 247172 319398
rect 248420 311840 248472 311846
rect 248420 311782 248472 311788
rect 247316 291236 247368 291242
rect 247316 291178 247368 291184
rect 247130 273184 247186 273193
rect 247130 273119 247186 273128
rect 247222 271552 247278 271561
rect 247222 271487 247278 271496
rect 247130 264480 247186 264489
rect 247130 264415 247186 264424
rect 247144 202842 247172 264415
rect 247236 235657 247264 271487
rect 247328 261526 247356 291178
rect 248432 283830 248460 311782
rect 248512 288516 248564 288522
rect 248512 288458 248564 288464
rect 248420 283824 248472 283830
rect 248420 283766 248472 283772
rect 248420 267572 248472 267578
rect 248420 267514 248472 267520
rect 247316 261520 247368 261526
rect 247316 261462 247368 261468
rect 247316 241528 247368 241534
rect 247316 241470 247368 241476
rect 247222 235648 247278 235657
rect 247222 235583 247278 235592
rect 247328 231810 247356 241470
rect 247316 231804 247368 231810
rect 247316 231746 247368 231752
rect 247132 202836 247184 202842
rect 247132 202778 247184 202784
rect 247144 200114 247172 202778
rect 247144 200086 247264 200114
rect 247132 192500 247184 192506
rect 247132 192442 247184 192448
rect 247038 153776 247094 153785
rect 247038 153711 247094 153720
rect 247144 140758 247172 192442
rect 247236 173194 247264 200086
rect 247224 173188 247276 173194
rect 247224 173130 247276 173136
rect 247684 171148 247736 171154
rect 247684 171090 247736 171096
rect 247132 140752 247184 140758
rect 246670 140720 246726 140729
rect 247132 140694 247184 140700
rect 246670 140655 246726 140664
rect 247696 140078 247724 171090
rect 248432 160070 248460 267514
rect 248524 209710 248552 288458
rect 248616 265674 248644 338127
rect 249064 337408 249116 337414
rect 249064 337350 249116 337356
rect 249076 269074 249104 337350
rect 249064 269068 249116 269074
rect 249064 269010 249116 269016
rect 248604 265668 248656 265674
rect 248604 265610 248656 265616
rect 248602 249928 248658 249937
rect 248602 249863 248658 249872
rect 248616 249830 248644 249863
rect 248604 249824 248656 249830
rect 248604 249766 248656 249772
rect 249812 249558 249840 352582
rect 250074 328672 250130 328681
rect 250074 328607 250130 328616
rect 249982 296032 250038 296041
rect 249982 295967 250038 295976
rect 249892 281580 249944 281586
rect 249892 281522 249944 281528
rect 249800 249552 249852 249558
rect 249800 249494 249852 249500
rect 249064 243364 249116 243370
rect 249064 243306 249116 243312
rect 248604 240236 248656 240242
rect 248604 240178 248656 240184
rect 248616 209774 248644 240178
rect 249076 237386 249104 243306
rect 249064 237380 249116 237386
rect 249064 237322 249116 237328
rect 249904 229094 249932 281522
rect 249996 279546 250024 295967
rect 250088 280838 250116 328607
rect 251364 323604 251416 323610
rect 251364 323546 251416 323552
rect 251180 298784 251232 298790
rect 251180 298726 251232 298732
rect 250076 280832 250128 280838
rect 250076 280774 250128 280780
rect 249984 279540 250036 279546
rect 249984 279482 250036 279488
rect 249982 278760 250038 278769
rect 249982 278695 249984 278704
rect 250036 278695 250038 278704
rect 249984 278666 250036 278672
rect 251192 273222 251220 298726
rect 251180 273216 251232 273222
rect 251180 273158 251232 273164
rect 250076 269068 250128 269074
rect 250076 269010 250128 269016
rect 249984 248668 250036 248674
rect 249984 248610 250036 248616
rect 249812 229066 249932 229094
rect 249812 224942 249840 229066
rect 249800 224936 249852 224942
rect 249800 224878 249852 224884
rect 248616 209746 248736 209774
rect 248512 209704 248564 209710
rect 248512 209646 248564 209652
rect 248524 160993 248552 209646
rect 248708 206990 248736 209746
rect 248696 206984 248748 206990
rect 248696 206926 248748 206932
rect 248604 182844 248656 182850
rect 248604 182786 248656 182792
rect 248510 160984 248566 160993
rect 248510 160919 248566 160928
rect 248420 160064 248472 160070
rect 248420 160006 248472 160012
rect 247868 156052 247920 156058
rect 247868 155994 247920 156000
rect 247776 150544 247828 150550
rect 247776 150486 247828 150492
rect 247684 140072 247736 140078
rect 247684 140014 247736 140020
rect 247684 136672 247736 136678
rect 247684 136614 247736 136620
rect 247696 128382 247724 136614
rect 247684 128376 247736 128382
rect 247684 128318 247736 128324
rect 247684 127016 247736 127022
rect 247684 126958 247736 126964
rect 246580 103488 246632 103494
rect 246580 103430 246632 103436
rect 246486 102232 246542 102241
rect 246486 102167 246542 102176
rect 246396 51740 246448 51746
rect 246396 51682 246448 51688
rect 246500 49026 246528 102167
rect 246488 49020 246540 49026
rect 246488 48962 246540 48968
rect 247696 24206 247724 126958
rect 247788 110430 247816 150486
rect 247880 119241 247908 155994
rect 248616 147801 248644 182786
rect 248708 176089 248736 206926
rect 248694 176080 248750 176089
rect 248694 176015 248750 176024
rect 249248 172576 249300 172582
rect 249248 172518 249300 172524
rect 249064 153332 249116 153338
rect 249064 153274 249116 153280
rect 248602 147792 248658 147801
rect 248602 147727 248658 147736
rect 247866 119232 247922 119241
rect 247866 119167 247922 119176
rect 247960 118720 248012 118726
rect 247960 118662 248012 118668
rect 247868 111852 247920 111858
rect 247868 111794 247920 111800
rect 247776 110424 247828 110430
rect 247776 110366 247828 110372
rect 247880 74089 247908 111794
rect 247972 89049 248000 118662
rect 249076 111761 249104 153274
rect 249154 135960 249210 135969
rect 249154 135895 249210 135904
rect 249062 111752 249118 111761
rect 249062 111687 249118 111696
rect 249062 99784 249118 99793
rect 249062 99719 249118 99728
rect 247958 89040 248014 89049
rect 247958 88975 248014 88984
rect 247866 74080 247922 74089
rect 247866 74015 247922 74024
rect 248418 71224 248474 71233
rect 248418 71159 248474 71168
rect 247684 24200 247736 24206
rect 247684 24142 247736 24148
rect 246304 5568 246356 5574
rect 246304 5510 246356 5516
rect 247590 3496 247646 3505
rect 244844 3454 245240 3482
rect 245212 480 245240 3454
rect 246396 3460 246448 3466
rect 247590 3431 247646 3440
rect 246396 3402 246448 3408
rect 246408 480 246436 3402
rect 247604 480 247632 3431
rect 248432 490 248460 71159
rect 249076 6186 249104 99719
rect 249168 64190 249196 135895
rect 249260 133822 249288 172518
rect 249812 170377 249840 224878
rect 249996 219434 250024 248610
rect 250088 243370 250116 269010
rect 251272 265668 251324 265674
rect 251272 265610 251324 265616
rect 251180 261520 251232 261526
rect 251180 261462 251232 261468
rect 250444 244316 250496 244322
rect 250444 244258 250496 244264
rect 250076 243364 250128 243370
rect 250076 243306 250128 243312
rect 250456 238678 250484 244258
rect 250444 238672 250496 238678
rect 250444 238614 250496 238620
rect 249904 219406 250024 219434
rect 249904 215286 249932 219406
rect 249892 215280 249944 215286
rect 249892 215222 249944 215228
rect 249904 215121 249932 215222
rect 249890 215112 249946 215121
rect 249890 215047 249946 215056
rect 250718 171592 250774 171601
rect 250718 171527 250774 171536
rect 249798 170368 249854 170377
rect 249798 170303 249854 170312
rect 250442 160440 250498 160449
rect 250442 160375 250498 160384
rect 249340 157480 249392 157486
rect 249340 157422 249392 157428
rect 249248 133816 249300 133822
rect 249248 133758 249300 133764
rect 249352 127673 249380 157422
rect 249432 133204 249484 133210
rect 249432 133146 249484 133152
rect 249338 127664 249394 127673
rect 249338 127599 249394 127608
rect 249338 110664 249394 110673
rect 249338 110599 249394 110608
rect 249248 106344 249300 106350
rect 249248 106286 249300 106292
rect 249156 64184 249208 64190
rect 249156 64126 249208 64132
rect 249260 61577 249288 106286
rect 249352 76537 249380 110599
rect 249444 107574 249472 133146
rect 250456 129033 250484 160375
rect 250536 154692 250588 154698
rect 250536 154634 250588 154640
rect 250442 129024 250498 129033
rect 250442 128959 250498 128968
rect 250548 114510 250576 154634
rect 250626 148472 250682 148481
rect 250626 148407 250682 148416
rect 250536 114504 250588 114510
rect 250536 114446 250588 114452
rect 250444 113212 250496 113218
rect 250444 113154 250496 113160
rect 249432 107568 249484 107574
rect 249432 107510 249484 107516
rect 249338 76528 249394 76537
rect 249338 76463 249394 76472
rect 249246 61568 249302 61577
rect 249246 61503 249302 61512
rect 250456 29714 250484 113154
rect 250534 107944 250590 107953
rect 250534 107879 250590 107888
rect 250548 44878 250576 107879
rect 250640 107545 250668 148407
rect 250732 141545 250760 171527
rect 251192 148345 251220 261462
rect 251284 158137 251312 265610
rect 251376 252550 251404 323546
rect 251836 322250 251864 373254
rect 252572 359009 252600 377590
rect 253204 374672 253256 374678
rect 253204 374614 253256 374620
rect 252558 359000 252614 359009
rect 252558 358935 252614 358944
rect 252560 332716 252612 332722
rect 252560 332658 252612 332664
rect 251824 322244 251876 322250
rect 251824 322186 251876 322192
rect 251824 314696 251876 314702
rect 251824 314638 251876 314644
rect 251836 268841 251864 314638
rect 252468 273216 252520 273222
rect 252468 273158 252520 273164
rect 252480 272542 252508 273158
rect 252468 272536 252520 272542
rect 252468 272478 252520 272484
rect 251822 268832 251878 268841
rect 251822 268767 251878 268776
rect 251364 252544 251416 252550
rect 251364 252486 251416 252492
rect 252468 252544 252520 252550
rect 252468 252486 252520 252492
rect 252480 251870 252508 252486
rect 252468 251864 252520 251870
rect 252468 251806 252520 251812
rect 251364 247784 251416 247790
rect 251364 247726 251416 247732
rect 251376 217977 251404 247726
rect 252572 237318 252600 332658
rect 252744 306400 252796 306406
rect 252744 306342 252796 306348
rect 252652 262268 252704 262274
rect 252652 262210 252704 262216
rect 252560 237312 252612 237318
rect 252560 237254 252612 237260
rect 251362 217968 251418 217977
rect 251362 217903 251418 217912
rect 252664 200114 252692 262210
rect 252756 259350 252784 306342
rect 253216 297430 253244 374614
rect 253294 359000 253350 359009
rect 253294 358935 253350 358944
rect 253308 329118 253336 358935
rect 253952 358154 253980 377590
rect 255976 374066 256004 377590
rect 256698 375320 256754 375329
rect 256698 375255 256754 375264
rect 255964 374060 256016 374066
rect 255964 374002 256016 374008
rect 253940 358148 253992 358154
rect 253940 358090 253992 358096
rect 255320 351212 255372 351218
rect 255320 351154 255372 351160
rect 255332 350606 255360 351154
rect 255320 350600 255372 350606
rect 255320 350542 255372 350548
rect 255332 345014 255360 350542
rect 255332 344986 255544 345014
rect 254032 340944 254084 340950
rect 254032 340886 254084 340892
rect 253296 329112 253348 329118
rect 253296 329054 253348 329060
rect 253940 312588 253992 312594
rect 253940 312530 253992 312536
rect 253204 297424 253256 297430
rect 253204 297366 253256 297372
rect 253204 294636 253256 294642
rect 253204 294578 253256 294584
rect 253216 263566 253244 294578
rect 253204 263560 253256 263566
rect 253204 263502 253256 263508
rect 253216 260846 253244 263502
rect 253204 260840 253256 260846
rect 253204 260782 253256 260788
rect 252744 259344 252796 259350
rect 252744 259286 252796 259292
rect 253020 259344 253072 259350
rect 253020 259286 253072 259292
rect 253032 258738 253060 259286
rect 253020 258732 253072 258738
rect 253020 258674 253072 258680
rect 253952 233238 253980 312530
rect 254044 270502 254072 340886
rect 254584 292596 254636 292602
rect 254584 292538 254636 292544
rect 254596 282878 254624 292538
rect 255318 290048 255374 290057
rect 255318 289983 255374 289992
rect 254584 282872 254636 282878
rect 254584 282814 254636 282820
rect 255136 282872 255188 282878
rect 255136 282814 255188 282820
rect 254032 270496 254084 270502
rect 254032 270438 254084 270444
rect 254400 269068 254452 269074
rect 254400 269010 254452 269016
rect 254412 268394 254440 269010
rect 254400 268388 254452 268394
rect 254400 268330 254452 268336
rect 254030 261216 254086 261225
rect 254030 261151 254086 261160
rect 253940 233232 253992 233238
rect 253940 233174 253992 233180
rect 253952 232558 253980 233174
rect 253940 232552 253992 232558
rect 253940 232494 253992 232500
rect 254044 209774 254072 261151
rect 254124 259412 254176 259418
rect 254124 259354 254176 259360
rect 254136 258806 254164 259354
rect 255148 258806 255176 282814
rect 254124 258800 254176 258806
rect 254124 258742 254176 258748
rect 255136 258800 255188 258806
rect 255136 258742 255188 258748
rect 253952 209746 254072 209774
rect 253952 205630 253980 209746
rect 253940 205624 253992 205630
rect 253940 205566 253992 205572
rect 252572 200086 252692 200114
rect 252572 198626 252600 200086
rect 252560 198620 252612 198626
rect 252560 198562 252612 198568
rect 251364 180872 251416 180878
rect 251364 180814 251416 180820
rect 251270 158128 251326 158137
rect 251270 158063 251326 158072
rect 251178 148336 251234 148345
rect 251178 148271 251234 148280
rect 250718 141536 250774 141545
rect 250718 141471 250774 141480
rect 250812 141432 250864 141438
rect 250812 141374 250864 141380
rect 250720 122868 250772 122874
rect 250720 122810 250772 122816
rect 250626 107536 250682 107545
rect 250626 107471 250682 107480
rect 250628 104236 250680 104242
rect 250628 104178 250680 104184
rect 250640 76809 250668 104178
rect 250732 101561 250760 122810
rect 250824 113150 250852 141374
rect 251376 137970 251404 180814
rect 252572 172514 252600 198562
rect 253204 191276 253256 191282
rect 253204 191218 253256 191224
rect 253216 180130 253244 191218
rect 253204 180124 253256 180130
rect 253204 180066 253256 180072
rect 252560 172508 252612 172514
rect 252560 172450 252612 172456
rect 253478 168464 253534 168473
rect 253478 168399 253534 168408
rect 253388 164348 253440 164354
rect 253388 164290 253440 164296
rect 253202 161528 253258 161537
rect 253202 161463 253258 161472
rect 251914 156496 251970 156505
rect 251914 156431 251970 156440
rect 251364 137964 251416 137970
rect 251364 137906 251416 137912
rect 251822 120184 251878 120193
rect 251822 120119 251878 120128
rect 250812 113144 250864 113150
rect 250812 113086 250864 113092
rect 250718 101552 250774 101561
rect 250718 101487 250774 101496
rect 250626 76800 250682 76809
rect 250626 76735 250682 76744
rect 250536 44872 250588 44878
rect 250536 44814 250588 44820
rect 250536 32428 250588 32434
rect 250536 32370 250588 32376
rect 250444 29708 250496 29714
rect 250444 29650 250496 29656
rect 250548 9654 250576 32370
rect 251836 31074 251864 120119
rect 251928 115938 251956 156431
rect 252008 151836 252060 151842
rect 252008 151778 252060 151784
rect 252020 120766 252048 151778
rect 252100 143608 252152 143614
rect 252100 143550 252152 143556
rect 252008 120760 252060 120766
rect 252008 120702 252060 120708
rect 252008 117360 252060 117366
rect 252008 117302 252060 117308
rect 251916 115932 251968 115938
rect 251916 115874 251968 115880
rect 251914 99648 251970 99657
rect 251914 99583 251970 99592
rect 251928 47598 251956 99583
rect 252020 69601 252048 117302
rect 252112 104174 252140 143550
rect 253216 122126 253244 161463
rect 253294 131608 253350 131617
rect 253294 131543 253350 131552
rect 253204 122120 253256 122126
rect 253204 122062 253256 122068
rect 253202 112160 253258 112169
rect 253202 112095 253258 112104
rect 252100 104168 252152 104174
rect 252100 104110 252152 104116
rect 252006 69592 252062 69601
rect 252006 69527 252062 69536
rect 251916 47592 251968 47598
rect 251916 47534 251968 47540
rect 253216 43450 253244 112095
rect 253308 72593 253336 131543
rect 253400 125594 253428 164290
rect 253492 131782 253520 168399
rect 253952 162489 253980 205566
rect 254676 171216 254728 171222
rect 254676 171158 254728 171164
rect 253938 162480 253994 162489
rect 253938 162415 253994 162424
rect 254584 158840 254636 158846
rect 254584 158782 254636 158788
rect 253480 131776 253532 131782
rect 253480 131718 253532 131724
rect 253388 125588 253440 125594
rect 253388 125530 253440 125536
rect 253480 124908 253532 124914
rect 253480 124850 253532 124856
rect 253386 100872 253442 100881
rect 253386 100807 253442 100816
rect 253400 87650 253428 100807
rect 253492 100638 253520 124850
rect 254596 118658 254624 158782
rect 254688 142934 254716 171158
rect 254858 167648 254914 167657
rect 254858 167583 254914 167592
rect 254676 142928 254728 142934
rect 254676 142870 254728 142876
rect 254766 142896 254822 142905
rect 254766 142831 254822 142840
rect 254676 129804 254728 129810
rect 254676 129746 254728 129752
rect 254584 118652 254636 118658
rect 254584 118594 254636 118600
rect 254584 116068 254636 116074
rect 254584 116010 254636 116016
rect 253480 100632 253532 100638
rect 253480 100574 253532 100580
rect 253388 87644 253440 87650
rect 253388 87586 253440 87592
rect 253294 72584 253350 72593
rect 253294 72519 253350 72528
rect 254596 46238 254624 116010
rect 254688 73817 254716 129746
rect 254780 100706 254808 142831
rect 254872 131073 254900 167583
rect 254858 131064 254914 131073
rect 254858 130999 254914 131008
rect 254768 100700 254820 100706
rect 254768 100642 254820 100648
rect 254766 98696 254822 98705
rect 254766 98631 254822 98640
rect 254780 77994 254808 98631
rect 255332 96529 255360 289983
rect 255412 287156 255464 287162
rect 255412 287098 255464 287104
rect 255424 164218 255452 287098
rect 255516 234297 255544 344986
rect 255594 280120 255650 280129
rect 255594 280055 255650 280064
rect 255608 279478 255636 280055
rect 255596 279472 255648 279478
rect 255596 279414 255648 279420
rect 255608 278798 255636 279414
rect 255596 278792 255648 278798
rect 255596 278734 255648 278740
rect 255502 234288 255558 234297
rect 255502 234223 255558 234232
rect 255976 187678 256004 374002
rect 256712 203561 256740 375255
rect 256804 325694 256832 377590
rect 258722 376680 258778 376689
rect 258722 376615 258778 376624
rect 258736 374678 258764 376615
rect 258724 374672 258776 374678
rect 258724 374614 258776 374620
rect 258078 331256 258134 331265
rect 258078 331191 258134 331200
rect 256804 325666 256924 325694
rect 256896 300121 256924 325666
rect 256882 300112 256938 300121
rect 256882 300047 256938 300056
rect 256792 299600 256844 299606
rect 256792 299542 256844 299548
rect 256698 203552 256754 203561
rect 256698 203487 256754 203496
rect 255964 187672 256016 187678
rect 255964 187614 256016 187620
rect 256804 170406 256832 299542
rect 256896 269142 256924 300047
rect 256976 271176 257028 271182
rect 256976 271118 257028 271124
rect 256884 269136 256936 269142
rect 256884 269078 256936 269084
rect 256988 175234 257016 271118
rect 258092 238746 258120 331191
rect 258172 322380 258224 322386
rect 258172 322322 258224 322328
rect 258184 255270 258212 322322
rect 258264 316804 258316 316810
rect 258264 316746 258316 316752
rect 258276 266529 258304 316746
rect 258736 297537 258764 374614
rect 259472 366353 259500 377590
rect 261496 375358 261524 377604
rect 262232 377590 263166 377618
rect 263612 377590 264822 377618
rect 266372 377590 266478 377618
rect 267752 377590 268134 377618
rect 269132 377590 269790 377618
rect 270512 377590 271446 377618
rect 260104 375352 260156 375358
rect 260104 375294 260156 375300
rect 261484 375352 261536 375358
rect 261484 375294 261536 375300
rect 259458 366344 259514 366353
rect 259458 366279 259514 366288
rect 259734 366344 259790 366353
rect 259734 366279 259790 366288
rect 259552 362228 259604 362234
rect 259552 362170 259604 362176
rect 258722 297528 258778 297537
rect 258722 297463 258778 297472
rect 259460 297424 259512 297430
rect 259460 297366 259512 297372
rect 258724 285796 258776 285802
rect 258724 285738 258776 285744
rect 258736 268433 258764 285738
rect 258722 268424 258778 268433
rect 258722 268359 258778 268368
rect 258262 266520 258318 266529
rect 258262 266455 258318 266464
rect 259366 266520 259422 266529
rect 259366 266455 259422 266464
rect 259380 264217 259408 266455
rect 259366 264208 259422 264217
rect 259366 264143 259422 264152
rect 258172 255264 258224 255270
rect 258172 255206 258224 255212
rect 258080 238740 258132 238746
rect 258080 238682 258132 238688
rect 259368 227792 259420 227798
rect 259368 227734 259420 227740
rect 259380 191214 259408 227734
rect 259472 215257 259500 297366
rect 259564 290494 259592 362170
rect 259644 308508 259696 308514
rect 259644 308450 259696 308456
rect 259552 290488 259604 290494
rect 259552 290430 259604 290436
rect 259550 288552 259606 288561
rect 259550 288487 259606 288496
rect 259564 256698 259592 288487
rect 259552 256692 259604 256698
rect 259552 256634 259604 256640
rect 259656 240009 259684 308450
rect 259748 287745 259776 366279
rect 260116 362234 260144 375294
rect 260104 362228 260156 362234
rect 260104 362170 260156 362176
rect 260932 322244 260984 322250
rect 260932 322186 260984 322192
rect 260840 311908 260892 311914
rect 260840 311850 260892 311856
rect 259734 287736 259790 287745
rect 259734 287671 259790 287680
rect 260102 287328 260158 287337
rect 260102 287263 260158 287272
rect 260116 269890 260144 287263
rect 260104 269884 260156 269890
rect 260104 269826 260156 269832
rect 260104 260160 260156 260166
rect 260104 260102 260156 260108
rect 259642 240000 259698 240009
rect 259642 239935 259698 239944
rect 259656 238746 259684 239935
rect 259644 238740 259696 238746
rect 259644 238682 259696 238688
rect 260116 227798 260144 260102
rect 260748 256692 260800 256698
rect 260748 256634 260800 256640
rect 260760 256018 260788 256634
rect 260748 256012 260800 256018
rect 260748 255954 260800 255960
rect 260196 247104 260248 247110
rect 260196 247046 260248 247052
rect 260208 238513 260236 247046
rect 260194 238504 260250 238513
rect 260194 238439 260250 238448
rect 260104 227792 260156 227798
rect 260104 227734 260156 227740
rect 259458 215248 259514 215257
rect 259458 215183 259514 215192
rect 260746 215248 260802 215257
rect 260746 215183 260802 215192
rect 260760 214606 260788 215183
rect 260748 214600 260800 214606
rect 260748 214542 260800 214548
rect 260196 198076 260248 198082
rect 260196 198018 260248 198024
rect 259368 191208 259420 191214
rect 259368 191150 259420 191156
rect 258080 187672 258132 187678
rect 258080 187614 258132 187620
rect 256976 175228 257028 175234
rect 256976 175170 257028 175176
rect 257342 174312 257398 174321
rect 257342 174247 257398 174256
rect 256792 170400 256844 170406
rect 256792 170342 256844 170348
rect 255412 164212 255464 164218
rect 255412 164154 255464 164160
rect 256056 146328 256108 146334
rect 256056 146270 256108 146276
rect 255964 121508 256016 121514
rect 255964 121450 256016 121456
rect 255318 96520 255374 96529
rect 255318 96455 255374 96464
rect 255870 96520 255926 96529
rect 255870 96455 255926 96464
rect 255884 95946 255912 96455
rect 255872 95940 255924 95946
rect 255872 95882 255924 95888
rect 254768 77988 254820 77994
rect 254768 77930 254820 77936
rect 254674 73808 254730 73817
rect 254674 73743 254730 73752
rect 254584 46232 254636 46238
rect 254584 46174 254636 46180
rect 253204 43444 253256 43450
rect 253204 43386 253256 43392
rect 251824 31068 251876 31074
rect 251824 31010 251876 31016
rect 251180 26920 251232 26926
rect 251180 26862 251232 26868
rect 249984 9648 250036 9654
rect 249984 9590 250036 9596
rect 250536 9648 250588 9654
rect 250536 9590 250588 9596
rect 249064 6180 249116 6186
rect 249064 6122 249116 6128
rect 248616 598 248828 626
rect 248616 490 248644 598
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248432 462 248644 490
rect 248800 480 248828 598
rect 249996 480 250024 9590
rect 251192 480 251220 26862
rect 255976 22778 256004 121450
rect 256068 111110 256096 146270
rect 257356 141409 257384 174247
rect 257618 172816 257674 172825
rect 257618 172751 257674 172760
rect 257436 160200 257488 160206
rect 257436 160142 257488 160148
rect 257342 141400 257398 141409
rect 257342 141335 257398 141344
rect 257344 132524 257396 132530
rect 257344 132466 257396 132472
rect 256056 111104 256108 111110
rect 256056 111046 256108 111052
rect 256148 107704 256200 107710
rect 256148 107646 256200 107652
rect 256054 106584 256110 106593
rect 256054 106519 256110 106528
rect 256068 40798 256096 106519
rect 256160 79665 256188 107646
rect 256146 79656 256202 79665
rect 256146 79591 256202 79600
rect 257356 68377 257384 132466
rect 257448 120057 257476 160142
rect 257526 149696 257582 149705
rect 257526 149631 257582 149640
rect 257434 120048 257490 120057
rect 257434 119983 257490 119992
rect 257436 114640 257488 114646
rect 257436 114582 257488 114588
rect 257342 68368 257398 68377
rect 257342 68303 257398 68312
rect 257448 55865 257476 114582
rect 257540 109002 257568 149631
rect 257632 133890 257660 172751
rect 257620 133884 257672 133890
rect 257620 133826 257672 133832
rect 257620 113280 257672 113286
rect 257620 113222 257672 113228
rect 257528 108996 257580 109002
rect 257528 108938 257580 108944
rect 257632 75313 257660 113222
rect 257618 75304 257674 75313
rect 257618 75239 257674 75248
rect 257434 55856 257490 55865
rect 257434 55791 257490 55800
rect 256056 40792 256108 40798
rect 256056 40734 256108 40740
rect 256054 33960 256110 33969
rect 256054 33895 256110 33904
rect 255964 22772 256016 22778
rect 255964 22714 256016 22720
rect 253202 22672 253258 22681
rect 253202 22607 253258 22616
rect 252374 3360 252430 3369
rect 252374 3295 252430 3304
rect 252388 480 252416 3295
rect 253216 2106 253244 22607
rect 253938 22128 253994 22137
rect 253938 22063 253994 22072
rect 253952 16574 253980 22063
rect 253952 16546 254256 16574
rect 253478 3496 253534 3505
rect 253478 3431 253534 3440
rect 253204 2100 253256 2106
rect 253204 2042 253256 2048
rect 253492 480 253520 3431
rect 254228 490 254256 16546
rect 256068 6914 256096 33895
rect 258092 16574 258120 187614
rect 260102 167104 260158 167113
rect 260102 167039 260158 167048
rect 258908 162988 258960 162994
rect 258908 162930 258960 162936
rect 258722 152008 258778 152017
rect 258722 151943 258778 151952
rect 258736 110401 258764 151943
rect 258816 142792 258868 142798
rect 258816 142734 258868 142740
rect 258722 110392 258778 110401
rect 258722 110327 258778 110336
rect 258828 102134 258856 142734
rect 258920 129062 258948 162930
rect 258908 129056 258960 129062
rect 258908 128998 258960 129004
rect 260116 126954 260144 167039
rect 260208 158001 260236 198018
rect 260288 174004 260340 174010
rect 260288 173946 260340 173952
rect 260300 162178 260328 173946
rect 260852 173369 260880 311850
rect 260944 282810 260972 322186
rect 262232 291825 262260 377590
rect 262494 377496 262550 377505
rect 262494 377431 262550 377440
rect 262508 375358 262536 377431
rect 262496 375352 262548 375358
rect 262496 375294 262548 375300
rect 263612 343913 263640 377590
rect 264978 348528 265034 348537
rect 264978 348463 265034 348472
rect 264992 347857 265020 348463
rect 264978 347848 265034 347857
rect 264978 347783 265034 347792
rect 263598 343904 263654 343913
rect 263598 343839 263654 343848
rect 264242 343904 264298 343913
rect 264242 343839 264298 343848
rect 263600 327820 263652 327826
rect 263600 327762 263652 327768
rect 262864 307080 262916 307086
rect 262864 307022 262916 307028
rect 262312 305040 262364 305046
rect 262312 304982 262364 304988
rect 262218 291816 262274 291825
rect 262218 291751 262274 291760
rect 260932 282804 260984 282810
rect 260932 282746 260984 282752
rect 262324 258074 262352 304982
rect 262140 258046 262352 258074
rect 262140 256766 262168 258046
rect 262128 256760 262180 256766
rect 262128 256702 262180 256708
rect 262140 188358 262168 256702
rect 262876 239465 262904 307022
rect 262956 275324 263008 275330
rect 262956 275266 263008 275272
rect 262862 239456 262918 239465
rect 262862 239391 262918 239400
rect 262876 200802 262904 239391
rect 262968 233073 262996 275266
rect 263612 235793 263640 327762
rect 264256 261526 264284 343839
rect 264336 273624 264388 273630
rect 264336 273566 264388 273572
rect 264244 261520 264296 261526
rect 264244 261462 264296 261468
rect 264348 247722 264376 273566
rect 264336 247716 264388 247722
rect 264336 247658 264388 247664
rect 263598 235784 263654 235793
rect 263598 235719 263654 235728
rect 262954 233064 263010 233073
rect 262954 232999 263010 233008
rect 262956 229152 263008 229158
rect 262956 229094 263008 229100
rect 262968 220794 262996 229094
rect 262956 220788 263008 220794
rect 262956 220730 263008 220736
rect 262864 200796 262916 200802
rect 262864 200738 262916 200744
rect 262128 188352 262180 188358
rect 262128 188294 262180 188300
rect 264992 177313 265020 347783
rect 266372 296177 266400 377590
rect 267648 370592 267700 370598
rect 267648 370534 267700 370540
rect 267002 301064 267058 301073
rect 267002 300999 267058 301008
rect 266358 296168 266414 296177
rect 266358 296103 266414 296112
rect 266266 283520 266322 283529
rect 266266 283455 266322 283464
rect 266280 278662 266308 283455
rect 266268 278656 266320 278662
rect 266268 278598 266320 278604
rect 266280 190369 266308 278598
rect 266452 245676 266504 245682
rect 266452 245618 266504 245624
rect 266360 244248 266412 244254
rect 266358 244216 266360 244225
rect 266412 244216 266414 244225
rect 266358 244151 266414 244160
rect 266464 238754 266492 245618
rect 266372 238726 266492 238754
rect 266372 219201 266400 238726
rect 266358 219192 266414 219201
rect 266358 219127 266414 219136
rect 267016 192506 267044 300999
rect 267660 244254 267688 370534
rect 267648 244248 267700 244254
rect 267648 244190 267700 244196
rect 267752 231742 267780 377590
rect 267832 319524 267884 319530
rect 267832 319466 267884 319472
rect 267844 266257 267872 319466
rect 269028 285796 269080 285802
rect 269028 285738 269080 285744
rect 269040 285705 269068 285738
rect 268382 285696 268438 285705
rect 268382 285631 268438 285640
rect 269026 285696 269082 285705
rect 269026 285631 269082 285640
rect 267830 266248 267886 266257
rect 267830 266183 267886 266192
rect 267832 244248 267884 244254
rect 267832 244190 267884 244196
rect 267740 231736 267792 231742
rect 267740 231678 267792 231684
rect 267844 195945 267872 244190
rect 268396 216345 268424 285631
rect 269132 273630 269160 377590
rect 269762 317520 269818 317529
rect 269762 317455 269818 317464
rect 269120 273624 269172 273630
rect 269120 273566 269172 273572
rect 269026 266248 269082 266257
rect 269026 266183 269082 266192
rect 269040 265577 269068 266183
rect 269026 265568 269082 265577
rect 269026 265503 269082 265512
rect 269028 256760 269080 256766
rect 269028 256702 269080 256708
rect 269040 253910 269068 256702
rect 269028 253904 269080 253910
rect 269028 253846 269080 253852
rect 269028 231736 269080 231742
rect 269028 231678 269080 231684
rect 269040 231130 269068 231678
rect 269028 231124 269080 231130
rect 269028 231066 269080 231072
rect 268474 229800 268530 229809
rect 268474 229735 268530 229744
rect 268382 216336 268438 216345
rect 268382 216271 268438 216280
rect 267830 195936 267886 195945
rect 267830 195871 267886 195880
rect 268382 195936 268438 195945
rect 268382 195871 268438 195880
rect 267004 192500 267056 192506
rect 267004 192442 267056 192448
rect 266266 190360 266322 190369
rect 266266 190295 266322 190304
rect 266280 189825 266308 190295
rect 266266 189816 266322 189825
rect 266266 189751 266322 189760
rect 268396 177342 268424 195871
rect 268488 180169 268516 229735
rect 269026 216336 269082 216345
rect 269026 216271 269082 216280
rect 269040 215937 269068 216271
rect 269026 215928 269082 215937
rect 269026 215863 269082 215872
rect 269776 185638 269804 317455
rect 269856 302252 269908 302258
rect 269856 302194 269908 302200
rect 269764 185632 269816 185638
rect 269764 185574 269816 185580
rect 269868 183161 269896 302194
rect 270408 267028 270460 267034
rect 270408 266970 270460 266976
rect 270420 266393 270448 266970
rect 270038 266384 270094 266393
rect 270038 266319 270094 266328
rect 270406 266384 270462 266393
rect 270406 266319 270462 266328
rect 270052 224913 270080 266319
rect 270512 234530 270540 377590
rect 273088 375358 273116 377604
rect 274744 375358 274772 377604
rect 276032 377590 276414 377618
rect 277688 377590 278070 377618
rect 273076 375352 273128 375358
rect 273076 375294 273128 375300
rect 273996 375352 274048 375358
rect 273996 375294 274048 375300
rect 274732 375352 274784 375358
rect 274732 375294 274784 375300
rect 273260 366376 273312 366382
rect 273260 366318 273312 366324
rect 273272 359514 273300 366318
rect 273260 359508 273312 359514
rect 273260 359450 273312 359456
rect 270592 302320 270644 302326
rect 270592 302262 270644 302268
rect 270500 234524 270552 234530
rect 270500 234466 270552 234472
rect 270038 224904 270094 224913
rect 270038 224839 270094 224848
rect 270406 224904 270462 224913
rect 270406 224839 270462 224848
rect 270420 224233 270448 224839
rect 270406 224224 270462 224233
rect 270406 224159 270462 224168
rect 269948 223644 270000 223650
rect 269948 223586 270000 223592
rect 269854 183152 269910 183161
rect 269854 183087 269910 183096
rect 268474 180160 268530 180169
rect 268474 180095 268530 180104
rect 268384 177336 268436 177342
rect 264978 177304 265034 177313
rect 268384 177278 268436 177284
rect 264978 177239 265034 177248
rect 269960 176662 269988 223586
rect 270604 198082 270632 302262
rect 272524 295996 272576 296002
rect 272524 295938 272576 295944
rect 271142 288688 271198 288697
rect 271142 288623 271198 288632
rect 270592 198076 270644 198082
rect 270592 198018 270644 198024
rect 271156 178809 271184 288623
rect 271236 234524 271288 234530
rect 271236 234466 271288 234472
rect 271248 181558 271276 234466
rect 272536 200870 272564 295938
rect 272616 282192 272668 282198
rect 272616 282134 272668 282140
rect 272628 234433 272656 282134
rect 273272 264926 273300 359450
rect 273904 358148 273956 358154
rect 273904 358090 273956 358096
rect 273260 264920 273312 264926
rect 273260 264862 273312 264868
rect 272614 234424 272670 234433
rect 272614 234359 272670 234368
rect 273916 232626 273944 358090
rect 274008 351218 274036 375294
rect 273996 351212 274048 351218
rect 273996 351154 274048 351160
rect 275284 337408 275336 337414
rect 275284 337350 275336 337356
rect 274640 305108 274692 305114
rect 274640 305050 274692 305056
rect 274652 301510 274680 305050
rect 274640 301504 274692 301510
rect 274640 301446 274692 301452
rect 275296 285802 275324 337350
rect 275284 285796 275336 285802
rect 275284 285738 275336 285744
rect 273904 232620 273956 232626
rect 273904 232562 273956 232568
rect 272524 200864 272576 200870
rect 272524 200806 272576 200812
rect 271236 181552 271288 181558
rect 271236 181494 271288 181500
rect 273916 181490 273944 232562
rect 275928 230444 275980 230450
rect 275928 230386 275980 230392
rect 275940 229770 275968 230386
rect 275928 229764 275980 229770
rect 275928 229706 275980 229712
rect 273994 200832 274050 200841
rect 273994 200767 274050 200776
rect 273904 181484 273956 181490
rect 273904 181426 273956 181432
rect 274008 180305 274036 200767
rect 275940 188426 275968 229706
rect 276032 226302 276060 377590
rect 277688 374066 277716 377590
rect 279712 375358 279740 377604
rect 281368 376689 281396 377604
rect 283038 377590 283604 377618
rect 281354 376680 281410 376689
rect 281354 376615 281410 376624
rect 278044 375352 278096 375358
rect 278044 375294 278096 375300
rect 279700 375352 279752 375358
rect 279700 375294 279752 375300
rect 276664 374060 276716 374066
rect 276664 374002 276716 374008
rect 277676 374060 277728 374066
rect 277676 374002 277728 374008
rect 276676 230450 276704 374002
rect 276754 294128 276810 294137
rect 276754 294063 276810 294072
rect 276664 230444 276716 230450
rect 276664 230386 276716 230392
rect 276020 226296 276072 226302
rect 276020 226238 276072 226244
rect 276032 225622 276060 226238
rect 276020 225616 276072 225622
rect 276020 225558 276072 225564
rect 276664 221468 276716 221474
rect 276664 221410 276716 221416
rect 275928 188420 275980 188426
rect 275928 188362 275980 188368
rect 273994 180296 274050 180305
rect 273994 180231 274050 180240
rect 276020 180124 276072 180130
rect 276020 180066 276072 180072
rect 273258 180024 273314 180033
rect 273258 179959 273314 179968
rect 271142 178800 271198 178809
rect 271142 178735 271198 178744
rect 273272 177313 273300 179959
rect 276032 178945 276060 180066
rect 276018 178936 276074 178945
rect 276018 178871 276074 178880
rect 273258 177304 273314 177313
rect 273258 177239 273314 177248
rect 269948 176656 270000 176662
rect 269948 176598 270000 176604
rect 276676 175982 276704 221410
rect 276768 177449 276796 294063
rect 278056 275330 278084 375294
rect 281368 374678 281396 376615
rect 281356 374672 281408 374678
rect 280894 374640 280950 374649
rect 281356 374614 281408 374620
rect 282184 374672 282236 374678
rect 282184 374614 282236 374620
rect 280894 374575 280950 374584
rect 279422 300928 279478 300937
rect 279422 300863 279478 300872
rect 278136 295384 278188 295390
rect 278136 295326 278188 295332
rect 278044 275324 278096 275330
rect 278044 275266 278096 275272
rect 278044 258800 278096 258806
rect 278044 258742 278096 258748
rect 277584 228404 277636 228410
rect 277584 228346 277636 228352
rect 277596 224262 277624 228346
rect 277584 224256 277636 224262
rect 277584 224198 277636 224204
rect 276848 193860 276900 193866
rect 276848 193802 276900 193808
rect 276860 179450 276888 193802
rect 276848 179444 276900 179450
rect 276848 179386 276900 179392
rect 276754 177440 276810 177449
rect 278056 177410 278084 258742
rect 278148 244934 278176 295326
rect 278136 244928 278188 244934
rect 278136 244870 278188 244876
rect 279436 222902 279464 300863
rect 280804 292732 280856 292738
rect 280804 292674 280856 292680
rect 279608 226364 279660 226370
rect 279608 226306 279660 226312
rect 279514 224224 279570 224233
rect 279514 224159 279570 224168
rect 279424 222896 279476 222902
rect 279424 222838 279476 222844
rect 278136 212560 278188 212566
rect 278136 212502 278188 212508
rect 278148 180198 278176 212502
rect 279422 211984 279478 211993
rect 279422 211919 279478 211928
rect 279330 192536 279386 192545
rect 279330 192471 279386 192480
rect 279238 183016 279294 183025
rect 279238 182951 279294 182960
rect 278136 180192 278188 180198
rect 278136 180134 278188 180140
rect 279148 179444 279200 179450
rect 279148 179386 279200 179392
rect 276754 177375 276810 177384
rect 278044 177404 278096 177410
rect 278044 177346 278096 177352
rect 276664 175976 276716 175982
rect 276664 175918 276716 175924
rect 264978 175672 265034 175681
rect 264978 175607 265034 175616
rect 264992 175302 265020 175607
rect 264980 175296 265032 175302
rect 264980 175238 265032 175244
rect 265622 175264 265678 175273
rect 265622 175199 265678 175208
rect 264978 174856 265034 174865
rect 264978 174791 265034 174800
rect 264992 173942 265020 174791
rect 265070 174040 265126 174049
rect 265070 173975 265072 173984
rect 265124 173975 265126 173984
rect 265072 173946 265124 173952
rect 264980 173936 265032 173942
rect 264980 173878 265032 173884
rect 264242 173632 264298 173641
rect 264242 173567 264298 173576
rect 260838 173360 260894 173369
rect 260838 173295 260894 173304
rect 261484 169856 261536 169862
rect 261484 169798 261536 169804
rect 260378 162752 260434 162761
rect 260378 162687 260434 162696
rect 260288 162172 260340 162178
rect 260288 162114 260340 162120
rect 260194 157992 260250 158001
rect 260194 157927 260250 157936
rect 260286 155272 260342 155281
rect 260286 155207 260342 155216
rect 260104 126948 260156 126954
rect 260104 126890 260156 126896
rect 260196 124228 260248 124234
rect 260196 124170 260248 124176
rect 260104 121576 260156 121582
rect 260104 121518 260156 121524
rect 259366 109168 259422 109177
rect 259366 109103 259422 109112
rect 258908 102264 258960 102270
rect 258908 102206 258960 102212
rect 258816 102128 258868 102134
rect 258816 102070 258868 102076
rect 258724 100836 258776 100842
rect 258724 100778 258776 100784
rect 258736 50386 258764 100778
rect 258920 65521 258948 102206
rect 259380 95198 259408 109103
rect 259368 95192 259420 95198
rect 259368 95134 259420 95140
rect 258906 65512 258962 65521
rect 258906 65447 258962 65456
rect 258724 50380 258776 50386
rect 258724 50322 258776 50328
rect 260116 28354 260144 121518
rect 260208 32502 260236 124170
rect 260300 114481 260328 155207
rect 260392 124166 260420 162687
rect 261496 132462 261524 169798
rect 262864 161696 262916 161702
rect 262864 161638 262916 161644
rect 262772 146396 262824 146402
rect 262772 146338 262824 146344
rect 262588 145036 262640 145042
rect 262588 144978 262640 144984
rect 262600 142866 262628 144978
rect 262784 144226 262812 146338
rect 262772 144220 262824 144226
rect 262772 144162 262824 144168
rect 262588 142860 262640 142866
rect 262588 142802 262640 142808
rect 262770 135960 262826 135969
rect 262770 135895 262826 135904
rect 262784 135425 262812 135895
rect 262770 135416 262826 135425
rect 262770 135351 262826 135360
rect 261484 132456 261536 132462
rect 261484 132398 261536 132404
rect 260472 131164 260524 131170
rect 260472 131106 260524 131112
rect 260380 124160 260432 124166
rect 260380 124102 260432 124108
rect 260286 114472 260342 114481
rect 260286 114407 260342 114416
rect 260484 112441 260512 131106
rect 261484 128376 261536 128382
rect 261484 128318 261536 128324
rect 260470 112432 260526 112441
rect 260470 112367 260526 112376
rect 260380 111920 260432 111926
rect 260380 111862 260432 111868
rect 260286 105768 260342 105777
rect 260286 105703 260342 105712
rect 260300 62801 260328 105703
rect 260392 94518 260420 111862
rect 260380 94512 260432 94518
rect 260380 94454 260432 94460
rect 260286 62792 260342 62801
rect 260286 62727 260342 62736
rect 261496 48929 261524 128318
rect 261576 125656 261628 125662
rect 261576 125598 261628 125604
rect 261588 80889 261616 125598
rect 262770 125080 262826 125089
rect 262770 125015 262826 125024
rect 262784 124681 262812 125015
rect 262770 124672 262826 124681
rect 262770 124607 262826 124616
rect 262876 121417 262904 161638
rect 263048 139460 263100 139466
rect 263048 139402 263100 139408
rect 262862 121408 262918 121417
rect 262862 121343 262918 121352
rect 261668 120216 261720 120222
rect 261668 120158 261720 120164
rect 261680 86290 261708 120158
rect 262862 118960 262918 118969
rect 262862 118895 262918 118904
rect 262126 107808 262182 107817
rect 262126 107743 262182 107752
rect 262140 105670 262168 107743
rect 262128 105664 262180 105670
rect 262128 105606 262180 105612
rect 261760 103964 261812 103970
rect 261760 103906 261812 103912
rect 261772 89010 261800 103906
rect 261760 89004 261812 89010
rect 261760 88946 261812 88952
rect 261668 86284 261720 86290
rect 261668 86226 261720 86232
rect 261574 80880 261630 80889
rect 261574 80815 261630 80824
rect 261482 48920 261538 48929
rect 261482 48855 261538 48864
rect 260196 32496 260248 32502
rect 260196 32438 260248 32444
rect 260104 28348 260156 28354
rect 260104 28290 260156 28296
rect 259458 28248 259514 28257
rect 259458 28183 259514 28192
rect 258092 16546 258304 16574
rect 257068 11756 257120 11762
rect 257068 11698 257120 11704
rect 255884 6886 256096 6914
rect 255884 4078 255912 6886
rect 257080 4146 257108 11698
rect 257068 4140 257120 4146
rect 257068 4082 257120 4088
rect 255872 4072 255924 4078
rect 255872 4014 255924 4020
rect 254504 598 254716 626
rect 254504 490 254532 598
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254228 462 254532 490
rect 254688 480 254716 598
rect 255884 480 255912 4014
rect 257080 480 257108 4082
rect 258276 480 258304 16546
rect 259472 480 259500 28183
rect 260838 21312 260894 21321
rect 260838 21247 260894 21256
rect 259552 17264 259604 17270
rect 259552 17206 259604 17212
rect 259564 16574 259592 17206
rect 260852 16574 260880 21247
rect 262876 18630 262904 118895
rect 262956 107772 263008 107778
rect 262956 107714 263008 107720
rect 262968 42090 262996 107714
rect 263060 104242 263088 139402
rect 264256 135250 264284 173567
rect 264978 172680 265034 172689
rect 264978 172615 265034 172624
rect 264992 172582 265020 172615
rect 264980 172576 265032 172582
rect 264980 172518 265032 172524
rect 265070 172272 265126 172281
rect 265070 172207 265126 172216
rect 264978 171456 265034 171465
rect 264978 171391 265034 171400
rect 264992 171222 265020 171391
rect 264980 171216 265032 171222
rect 264980 171158 265032 171164
rect 265084 171154 265112 172207
rect 265072 171148 265124 171154
rect 265072 171090 265124 171096
rect 265070 171048 265126 171057
rect 265070 170983 265126 170992
rect 264978 170096 265034 170105
rect 264978 170031 265034 170040
rect 264992 169794 265020 170031
rect 265084 169862 265112 170983
rect 265162 170504 265218 170513
rect 265162 170439 265218 170448
rect 265072 169856 265124 169862
rect 265072 169798 265124 169804
rect 264980 169788 265032 169794
rect 264980 169730 265032 169736
rect 264978 169688 265034 169697
rect 264978 169623 265034 169632
rect 264992 168502 265020 169623
rect 265070 168872 265126 168881
rect 265070 168807 265126 168816
rect 264980 168496 265032 168502
rect 264980 168438 265032 168444
rect 265084 168434 265112 168807
rect 265072 168428 265124 168434
rect 265072 168370 265124 168376
rect 265070 167920 265126 167929
rect 265070 167855 265126 167864
rect 264978 167512 265034 167521
rect 264978 167447 265034 167456
rect 264992 167142 265020 167447
rect 264980 167136 265032 167142
rect 264980 167078 265032 167084
rect 265084 167074 265112 167855
rect 265176 167657 265204 170439
rect 265254 169280 265310 169289
rect 265254 169215 265310 169224
rect 265162 167648 265218 167657
rect 265162 167583 265218 167592
rect 265072 167068 265124 167074
rect 265072 167010 265124 167016
rect 265070 166696 265126 166705
rect 265070 166631 265126 166640
rect 264978 166288 265034 166297
rect 264978 166223 265034 166232
rect 264992 165646 265020 166223
rect 265084 165714 265112 166631
rect 265268 166433 265296 169215
rect 265254 166424 265310 166433
rect 265254 166359 265310 166368
rect 265162 165880 265218 165889
rect 265162 165815 265218 165824
rect 265072 165708 265124 165714
rect 265072 165650 265124 165656
rect 264980 165640 265032 165646
rect 264980 165582 265032 165588
rect 265070 165336 265126 165345
rect 265070 165271 265126 165280
rect 264978 164928 265034 164937
rect 264978 164863 265034 164872
rect 264992 164354 265020 164863
rect 264980 164348 265032 164354
rect 264980 164290 265032 164296
rect 265084 164286 265112 165271
rect 265176 165073 265204 165815
rect 265162 165064 265218 165073
rect 265162 164999 265218 165008
rect 265254 164520 265310 164529
rect 265254 164455 265310 164464
rect 265072 164280 265124 164286
rect 265072 164222 265124 164228
rect 264978 164112 265034 164121
rect 264978 164047 265034 164056
rect 264992 162926 265020 164047
rect 265070 163704 265126 163713
rect 265070 163639 265126 163648
rect 265084 162994 265112 163639
rect 265162 163296 265218 163305
rect 265162 163231 265218 163240
rect 265072 162988 265124 162994
rect 265072 162930 265124 162936
rect 264980 162920 265032 162926
rect 264980 162862 265032 162868
rect 264978 162344 265034 162353
rect 264978 162279 265034 162288
rect 264992 161498 265020 162279
rect 265070 161936 265126 161945
rect 265070 161871 265126 161880
rect 265084 161702 265112 161871
rect 265072 161696 265124 161702
rect 265072 161638 265124 161644
rect 264980 161492 265032 161498
rect 264980 161434 265032 161440
rect 265070 161120 265126 161129
rect 265070 161055 265126 161064
rect 264978 160304 265034 160313
rect 264978 160239 265034 160248
rect 264992 160206 265020 160239
rect 264980 160200 265032 160206
rect 264980 160142 265032 160148
rect 265084 160138 265112 161055
rect 265072 160132 265124 160138
rect 265072 160074 265124 160080
rect 265070 159760 265126 159769
rect 265070 159695 265126 159704
rect 264978 158944 265034 158953
rect 264978 158879 265034 158888
rect 264992 158846 265020 158879
rect 264980 158840 265032 158846
rect 264980 158782 265032 158788
rect 265084 158778 265112 159695
rect 265072 158772 265124 158778
rect 265072 158714 265124 158720
rect 265070 158536 265126 158545
rect 265070 158471 265126 158480
rect 264978 158128 265034 158137
rect 264978 158063 265034 158072
rect 264992 157486 265020 158063
rect 264980 157480 265032 157486
rect 264334 157448 264390 157457
rect 264980 157422 265032 157428
rect 265084 157418 265112 158471
rect 265176 157457 265204 163231
rect 265268 162761 265296 164455
rect 265254 162752 265310 162761
rect 265254 162687 265310 162696
rect 265346 157720 265402 157729
rect 265346 157655 265402 157664
rect 265162 157448 265218 157457
rect 264334 157383 264390 157392
rect 265072 157412 265124 157418
rect 264244 135244 264296 135250
rect 264244 135186 264296 135192
rect 264348 122777 264376 157383
rect 265162 157383 265218 157392
rect 265072 157354 265124 157360
rect 265070 157176 265126 157185
rect 265070 157111 265126 157120
rect 264978 156360 265034 156369
rect 264978 156295 265034 156304
rect 264992 156058 265020 156295
rect 264980 156052 265032 156058
rect 264980 155994 265032 156000
rect 265084 155990 265112 157111
rect 265072 155984 265124 155990
rect 265072 155926 265124 155932
rect 265162 155952 265218 155961
rect 265162 155887 265218 155896
rect 264980 154692 265032 154698
rect 264980 154634 265032 154640
rect 264992 154601 265020 154634
rect 265176 154630 265204 155887
rect 265164 154624 265216 154630
rect 264978 154592 265034 154601
rect 265164 154566 265216 154572
rect 264978 154527 265034 154536
rect 265070 153776 265126 153785
rect 265070 153711 265126 153720
rect 264978 153368 265034 153377
rect 264978 153303 264980 153312
rect 265032 153303 265034 153312
rect 264980 153274 265032 153280
rect 265084 153270 265112 153711
rect 265072 153264 265124 153270
rect 265072 153206 265124 153212
rect 264978 152960 265034 152969
rect 264978 152895 265034 152904
rect 264992 151842 265020 152895
rect 265254 152552 265310 152561
rect 265360 152522 265388 157655
rect 265254 152487 265310 152496
rect 265348 152516 265400 152522
rect 264980 151836 265032 151842
rect 265268 151814 265296 152487
rect 265348 152458 265400 152464
rect 264980 151778 265032 151784
rect 265176 151786 265296 151814
rect 265070 151600 265126 151609
rect 265070 151535 265126 151544
rect 264978 151192 265034 151201
rect 264978 151127 265034 151136
rect 264992 150550 265020 151127
rect 264980 150544 265032 150550
rect 264980 150486 265032 150492
rect 265084 150482 265112 151535
rect 265072 150476 265124 150482
rect 265072 150418 265124 150424
rect 264978 149968 265034 149977
rect 264978 149903 265034 149912
rect 264992 149122 265020 149903
rect 265070 149560 265126 149569
rect 265070 149495 265126 149504
rect 264980 149116 265032 149122
rect 264980 149058 265032 149064
rect 265084 148481 265112 149495
rect 265070 148472 265126 148481
rect 265070 148407 265126 148416
rect 265176 148374 265204 151786
rect 265254 150784 265310 150793
rect 265254 150719 265310 150728
rect 265164 148368 265216 148374
rect 265164 148310 265216 148316
rect 265162 148200 265218 148209
rect 265162 148135 265218 148144
rect 264978 147792 265034 147801
rect 264978 147727 265034 147736
rect 264992 147694 265020 147727
rect 264980 147688 265032 147694
rect 264980 147630 265032 147636
rect 264978 147384 265034 147393
rect 264978 147319 265034 147328
rect 264992 146334 265020 147319
rect 265070 146432 265126 146441
rect 265070 146367 265072 146376
rect 265124 146367 265126 146376
rect 265072 146338 265124 146344
rect 264980 146328 265032 146334
rect 264980 146270 265032 146276
rect 265070 146024 265126 146033
rect 265070 145959 265126 145968
rect 264978 145208 265034 145217
rect 264978 145143 265034 145152
rect 264992 144974 265020 145143
rect 265084 145042 265112 145959
rect 265176 145625 265204 148135
rect 265268 146985 265296 150719
rect 265636 149734 265664 175199
rect 279160 171134 279188 179386
rect 279252 172258 279280 182951
rect 279344 172394 279372 192471
rect 279436 178770 279464 211919
rect 279528 183025 279556 224159
rect 279620 219434 279648 226306
rect 279608 219428 279660 219434
rect 279608 219370 279660 219376
rect 280158 184376 280214 184385
rect 280158 184311 280214 184320
rect 279514 183016 279570 183025
rect 279514 182951 279570 182960
rect 279424 178764 279476 178770
rect 279424 178706 279476 178712
rect 279344 172366 279556 172394
rect 279330 172272 279386 172281
rect 279252 172230 279330 172258
rect 279330 172207 279386 172216
rect 279160 171106 279280 171134
rect 279252 157334 279280 171106
rect 279528 161474 279556 172366
rect 280172 162625 280200 184311
rect 280252 180192 280304 180198
rect 280252 180134 280304 180140
rect 280264 168745 280292 180134
rect 280816 175098 280844 292674
rect 280908 291145 280936 374575
rect 281448 320884 281500 320890
rect 281448 320826 281500 320832
rect 281460 320210 281488 320826
rect 281448 320204 281500 320210
rect 281448 320146 281500 320152
rect 281356 319456 281408 319462
rect 281356 319398 281408 319404
rect 281368 307737 281396 319398
rect 281354 307728 281410 307737
rect 281354 307663 281410 307672
rect 281368 307154 281396 307663
rect 281356 307148 281408 307154
rect 281356 307090 281408 307096
rect 280894 291136 280950 291145
rect 280894 291071 280950 291080
rect 280986 287192 281042 287201
rect 280986 287127 281042 287136
rect 280894 284608 280950 284617
rect 280894 284543 280950 284552
rect 280908 182850 280936 284543
rect 281000 275330 281028 287127
rect 280988 275324 281040 275330
rect 280988 275266 281040 275272
rect 280896 182844 280948 182850
rect 280896 182786 280948 182792
rect 280894 182064 280950 182073
rect 280894 181999 280950 182008
rect 280804 175092 280856 175098
rect 280804 175034 280856 175040
rect 280250 168736 280306 168745
rect 280250 168671 280306 168680
rect 280158 162616 280214 162625
rect 280158 162551 280214 162560
rect 279068 157306 279280 157334
rect 279344 161446 279556 161474
rect 265714 154184 265770 154193
rect 265714 154119 265770 154128
rect 265624 149728 265676 149734
rect 265624 149670 265676 149676
rect 265254 146976 265310 146985
rect 265254 146911 265310 146920
rect 265438 146976 265494 146985
rect 265438 146911 265494 146920
rect 265162 145616 265218 145625
rect 265162 145551 265218 145560
rect 265072 145036 265124 145042
rect 265072 144978 265124 144984
rect 264980 144968 265032 144974
rect 264980 144910 265032 144916
rect 264610 144800 264666 144809
rect 264610 144735 264666 144744
rect 264426 140856 264482 140865
rect 264426 140791 264482 140800
rect 264334 122768 264390 122777
rect 264334 122703 264390 122712
rect 264242 119368 264298 119377
rect 264242 119303 264298 119312
rect 263140 104916 263192 104922
rect 263140 104858 263192 104864
rect 263048 104236 263100 104242
rect 263048 104178 263100 104184
rect 263048 100768 263100 100774
rect 263048 100710 263100 100716
rect 263060 83473 263088 100710
rect 263152 90370 263180 104858
rect 263140 90364 263192 90370
rect 263140 90306 263192 90312
rect 263046 83464 263102 83473
rect 263046 83399 263102 83408
rect 262956 42084 263008 42090
rect 262956 42026 263008 42032
rect 262864 18624 262916 18630
rect 262864 18566 262916 18572
rect 263598 17368 263654 17377
rect 263598 17303 263654 17312
rect 263612 16574 263640 17303
rect 259564 16546 260696 16574
rect 260852 16546 261800 16574
rect 263612 16546 264192 16574
rect 260668 480 260696 16546
rect 261772 480 261800 16546
rect 262956 7608 263008 7614
rect 262956 7550 263008 7556
rect 262968 480 262996 7550
rect 264164 480 264192 16546
rect 264256 10402 264284 119303
rect 264334 109984 264390 109993
rect 264334 109919 264390 109928
rect 264348 58682 264376 109919
rect 264440 105602 264468 140791
rect 264624 119406 264652 144735
rect 264978 143848 265034 143857
rect 264978 143783 265034 143792
rect 264992 143614 265020 143783
rect 264980 143608 265032 143614
rect 264980 143550 265032 143556
rect 264978 143440 265034 143449
rect 264978 143375 265034 143384
rect 264992 142798 265020 143375
rect 264980 142792 265032 142798
rect 265452 142769 265480 146911
rect 264980 142734 265032 142740
rect 265438 142760 265494 142769
rect 265438 142695 265494 142704
rect 265162 142624 265218 142633
rect 265162 142559 265218 142568
rect 265070 141264 265126 141273
rect 265070 141199 265126 141208
rect 264978 139224 265034 139233
rect 264978 139159 265034 139168
rect 264992 138038 265020 139159
rect 265084 138689 265112 141199
rect 265176 140049 265204 142559
rect 265622 142216 265678 142225
rect 265622 142151 265678 142160
rect 265162 140040 265218 140049
rect 265162 139975 265218 139984
rect 265346 140040 265402 140049
rect 265346 139975 265402 139984
rect 265360 139466 265388 139975
rect 265348 139460 265400 139466
rect 265348 139402 265400 139408
rect 265070 138680 265126 138689
rect 265070 138615 265126 138624
rect 264980 138032 265032 138038
rect 264980 137974 265032 137980
rect 264978 137864 265034 137873
rect 264978 137799 265034 137808
rect 264992 136678 265020 137799
rect 264980 136672 265032 136678
rect 264980 136614 265032 136620
rect 265070 136640 265126 136649
rect 265070 136575 265126 136584
rect 264978 135688 265034 135697
rect 264978 135623 265034 135632
rect 264992 135386 265020 135623
rect 264980 135380 265032 135386
rect 264980 135322 265032 135328
rect 265084 135318 265112 136575
rect 265072 135312 265124 135318
rect 265072 135254 265124 135260
rect 264978 134056 265034 134065
rect 264978 133991 265034 134000
rect 264992 133958 265020 133991
rect 264980 133952 265032 133958
rect 264980 133894 265032 133900
rect 264978 132696 265034 132705
rect 264978 132631 265034 132640
rect 264992 132530 265020 132631
rect 264980 132524 265032 132530
rect 264980 132466 265032 132472
rect 264978 132288 265034 132297
rect 264978 132223 265034 132232
rect 264992 131170 265020 132223
rect 264980 131164 265032 131170
rect 264980 131106 265032 131112
rect 264978 131064 265034 131073
rect 264978 130999 265034 131008
rect 264992 129810 265020 130999
rect 265070 130520 265126 130529
rect 265070 130455 265126 130464
rect 264980 129804 265032 129810
rect 264980 129746 265032 129752
rect 264978 129296 265034 129305
rect 264978 129231 265034 129240
rect 264992 127634 265020 129231
rect 264980 127628 265032 127634
rect 264980 127570 265032 127576
rect 264978 127528 265034 127537
rect 264978 127463 265034 127472
rect 264992 127022 265020 127463
rect 264980 127016 265032 127022
rect 264980 126958 265032 126964
rect 265084 126585 265112 130455
rect 265162 129704 265218 129713
rect 265162 129639 265218 129648
rect 265176 128382 265204 129639
rect 265164 128376 265216 128382
rect 265164 128318 265216 128324
rect 265070 126576 265126 126585
rect 265070 126511 265126 126520
rect 264978 125896 265034 125905
rect 264978 125831 265034 125840
rect 264992 125662 265020 125831
rect 264980 125656 265032 125662
rect 264980 125598 265032 125604
rect 265636 124914 265664 142151
rect 265728 141438 265756 154119
rect 279068 153194 279096 157306
rect 279344 155961 279372 161446
rect 280068 156664 280120 156670
rect 280068 156606 280120 156612
rect 279330 155952 279386 155961
rect 279330 155887 279386 155896
rect 279068 153166 279464 153194
rect 267094 149016 267150 149025
rect 267094 148951 267150 148960
rect 265806 148608 265862 148617
rect 265806 148543 265862 148552
rect 265716 141432 265768 141438
rect 265716 141374 265768 141380
rect 265716 138032 265768 138038
rect 265716 137974 265768 137980
rect 265624 124908 265676 124914
rect 265624 124850 265676 124856
rect 264978 124536 265034 124545
rect 264978 124471 265034 124480
rect 264992 124234 265020 124471
rect 264980 124228 265032 124234
rect 264980 124170 265032 124176
rect 264978 123720 265034 123729
rect 264978 123655 265034 123664
rect 264992 122874 265020 123655
rect 265622 122904 265678 122913
rect 264980 122868 265032 122874
rect 265622 122839 265678 122848
rect 264980 122810 265032 122816
rect 264978 121952 265034 121961
rect 264978 121887 265034 121896
rect 264992 121514 265020 121887
rect 265072 121576 265124 121582
rect 265070 121544 265072 121553
rect 265124 121544 265126 121553
rect 264980 121508 265032 121514
rect 265070 121479 265126 121488
rect 264980 121450 265032 121456
rect 264978 121136 265034 121145
rect 264978 121071 265034 121080
rect 264992 120154 265020 121071
rect 265070 120728 265126 120737
rect 265070 120663 265126 120672
rect 265084 120222 265112 120663
rect 265072 120216 265124 120222
rect 265072 120158 265124 120164
rect 264980 120148 265032 120154
rect 264980 120090 265032 120096
rect 264978 119776 265034 119785
rect 264978 119711 265034 119720
rect 264612 119400 264664 119406
rect 264612 119342 264664 119348
rect 264992 118726 265020 119711
rect 264980 118720 265032 118726
rect 264980 118662 265032 118668
rect 264978 118552 265034 118561
rect 264978 118487 265034 118496
rect 264992 117366 265020 118487
rect 264980 117360 265032 117366
rect 264980 117302 265032 117308
rect 265070 117192 265126 117201
rect 265070 117127 265126 117136
rect 264978 116784 265034 116793
rect 264978 116719 265034 116728
rect 264992 116006 265020 116719
rect 265084 116074 265112 117127
rect 265072 116068 265124 116074
rect 265072 116010 265124 116016
rect 264980 116000 265032 116006
rect 264980 115942 265032 115948
rect 265070 115152 265126 115161
rect 265070 115087 265126 115096
rect 265084 114646 265112 115087
rect 265072 114640 265124 114646
rect 264978 114608 265034 114617
rect 265072 114582 265124 114588
rect 264978 114543 264980 114552
rect 265032 114543 265034 114552
rect 264980 114514 265032 114520
rect 265070 113792 265126 113801
rect 265070 113727 265126 113736
rect 264978 113384 265034 113393
rect 264978 113319 265034 113328
rect 264992 113218 265020 113319
rect 265084 113286 265112 113727
rect 265072 113280 265124 113286
rect 265072 113222 265124 113228
rect 264980 113212 265032 113218
rect 264980 113154 265032 113160
rect 264978 112568 265034 112577
rect 264978 112503 265034 112512
rect 264992 111858 265020 112503
rect 264980 111852 265032 111858
rect 264980 111794 265032 111800
rect 264978 111616 265034 111625
rect 264978 111551 265034 111560
rect 264992 110498 265020 111551
rect 264980 110492 265032 110498
rect 264980 110434 265032 110440
rect 265070 110392 265126 110401
rect 265070 110327 265126 110336
rect 265084 109070 265112 110327
rect 265072 109064 265124 109070
rect 264978 109032 265034 109041
rect 265072 109006 265124 109012
rect 264978 108967 265034 108976
rect 264992 107710 265020 108967
rect 265346 108624 265402 108633
rect 265346 108559 265402 108568
rect 265360 107778 265388 108559
rect 265348 107772 265400 107778
rect 265348 107714 265400 107720
rect 264980 107704 265032 107710
rect 264980 107646 265032 107652
rect 264978 107400 265034 107409
rect 264978 107335 265034 107344
rect 264886 106448 264942 106457
rect 264886 106383 264942 106392
rect 264428 105596 264480 105602
rect 264428 105538 264480 105544
rect 264428 99408 264480 99414
rect 264428 99350 264480 99356
rect 264440 84862 264468 99350
rect 264900 93906 264928 106383
rect 264992 106350 265020 107335
rect 264980 106344 265032 106350
rect 264980 106286 265032 106292
rect 264978 105224 265034 105233
rect 264978 105159 265034 105168
rect 264992 104922 265020 105159
rect 264980 104916 265032 104922
rect 264980 104858 265032 104864
rect 264978 104408 265034 104417
rect 264978 104343 265034 104352
rect 264992 103970 265020 104343
rect 264980 103964 265032 103970
rect 264980 103906 265032 103912
rect 265070 103456 265126 103465
rect 265070 103391 265126 103400
rect 264978 102640 265034 102649
rect 264978 102575 265034 102584
rect 264992 102202 265020 102575
rect 265084 102270 265112 103391
rect 265072 102264 265124 102270
rect 265072 102206 265124 102212
rect 264980 102196 265032 102202
rect 264980 102138 265032 102144
rect 264978 101824 265034 101833
rect 264978 101759 265034 101768
rect 264992 100842 265020 101759
rect 265070 101280 265126 101289
rect 265070 101215 265126 101224
rect 264980 100836 265032 100842
rect 264980 100778 265032 100784
rect 265084 100774 265112 101215
rect 265072 100768 265124 100774
rect 265072 100710 265124 100716
rect 265070 99240 265126 99249
rect 265070 99175 265126 99184
rect 264978 98696 265034 98705
rect 264978 98631 265034 98640
rect 264992 98054 265020 98631
rect 265084 98122 265112 99175
rect 265072 98116 265124 98122
rect 265072 98058 265124 98064
rect 264980 98048 265032 98054
rect 264980 97990 265032 97996
rect 265070 97880 265126 97889
rect 265070 97815 265126 97824
rect 264980 97368 265032 97374
rect 264980 97310 265032 97316
rect 264992 96665 265020 97310
rect 265084 97306 265112 97815
rect 265072 97300 265124 97306
rect 265072 97242 265124 97248
rect 264978 96656 265034 96665
rect 264978 96591 265034 96600
rect 264978 96248 265034 96257
rect 264978 96183 265034 96192
rect 264992 95266 265020 96183
rect 264980 95260 265032 95266
rect 264980 95202 265032 95208
rect 264888 93900 264940 93906
rect 264888 93842 264940 93848
rect 264428 84856 264480 84862
rect 265636 84833 265664 122839
rect 265728 107642 265756 137974
rect 265820 133210 265848 148543
rect 267002 138272 267058 138281
rect 267002 138207 267058 138216
rect 265808 133204 265860 133210
rect 265808 133146 265860 133152
rect 265806 127936 265862 127945
rect 265806 127871 265862 127880
rect 265716 107636 265768 107642
rect 265716 107578 265768 107584
rect 265820 98841 265848 127871
rect 265898 126304 265954 126313
rect 265898 126239 265954 126248
rect 265912 111926 265940 126239
rect 265990 112024 266046 112033
rect 265990 111959 266046 111968
rect 265900 111920 265952 111926
rect 265900 111862 265952 111868
rect 266004 99414 266032 111959
rect 265992 99408 266044 99414
rect 265992 99350 266044 99356
rect 265806 98832 265862 98841
rect 265806 98767 265862 98776
rect 265990 98288 266046 98297
rect 265990 98223 266046 98232
rect 265714 97472 265770 97481
rect 265714 97407 265770 97416
rect 264428 84798 264480 84804
rect 265622 84824 265678 84833
rect 265622 84759 265678 84768
rect 265728 80753 265756 97407
rect 265714 80744 265770 80753
rect 265714 80679 265770 80688
rect 266004 79529 266032 98223
rect 265990 79520 266046 79529
rect 265990 79455 266046 79464
rect 264336 58676 264388 58682
rect 264336 58618 264388 58624
rect 267016 53145 267044 138207
rect 267108 138038 267136 148951
rect 279330 148336 279386 148345
rect 279330 148271 279386 148280
rect 279344 143534 279372 148271
rect 279436 144809 279464 153166
rect 280080 148345 280108 156606
rect 280066 148336 280122 148345
rect 280066 148271 280122 148280
rect 280908 145897 280936 181999
rect 281460 179450 281488 320146
rect 282196 282198 282224 374614
rect 283576 374105 283604 377590
rect 284312 377590 284694 377618
rect 285692 377590 286350 377618
rect 287072 377590 288006 377618
rect 283562 374096 283618 374105
rect 283562 374031 283618 374040
rect 283576 360913 283604 374031
rect 283562 360904 283618 360913
rect 283562 360839 283618 360848
rect 282276 303748 282328 303754
rect 282276 303690 282328 303696
rect 282288 286346 282316 303690
rect 282920 296744 282972 296750
rect 282920 296686 282972 296692
rect 282276 286340 282328 286346
rect 282276 286282 282328 286288
rect 282184 282192 282236 282198
rect 282184 282134 282236 282140
rect 282276 282192 282328 282198
rect 282276 282134 282328 282140
rect 282288 260166 282316 282134
rect 282276 260160 282328 260166
rect 282276 260102 282328 260108
rect 281630 202328 281686 202337
rect 281630 202263 281686 202272
rect 281540 200796 281592 200802
rect 281540 200738 281592 200744
rect 281448 179444 281500 179450
rect 281448 179386 281500 179392
rect 280988 175228 281040 175234
rect 280988 175170 281040 175176
rect 281000 166433 281028 175170
rect 280986 166424 281042 166433
rect 280986 166359 281042 166368
rect 280894 145888 280950 145897
rect 280894 145823 280950 145832
rect 279422 144800 279478 144809
rect 279422 144735 279478 144744
rect 279068 143506 279372 143534
rect 267096 138032 267148 138038
rect 267096 137974 267148 137980
rect 267094 134464 267150 134473
rect 267094 134399 267150 134408
rect 267108 65657 267136 134399
rect 267186 124128 267242 124137
rect 267186 124063 267242 124072
rect 267200 82113 267228 124063
rect 279068 113174 279096 143506
rect 281552 119241 281580 200738
rect 281644 163305 281672 202263
rect 281906 178936 281962 178945
rect 281906 178871 281962 178880
rect 281816 177336 281868 177342
rect 281816 177278 281868 177284
rect 281724 176656 281776 176662
rect 281724 176598 281776 176604
rect 281736 175545 281764 176598
rect 281722 175536 281778 175545
rect 281722 175471 281778 175480
rect 281630 163296 281686 163305
rect 281630 163231 281686 163240
rect 281828 161474 281856 177278
rect 281920 175234 281948 178871
rect 281908 175228 281960 175234
rect 281908 175170 281960 175176
rect 282184 175228 282236 175234
rect 282184 175170 282236 175176
rect 282196 174049 282224 175170
rect 282182 174040 282238 174049
rect 282182 173975 282238 173984
rect 282460 173868 282512 173874
rect 282460 173810 282512 173816
rect 282472 172553 282500 173810
rect 282458 172544 282514 172553
rect 282458 172479 282514 172488
rect 282276 170944 282328 170950
rect 282274 170912 282276 170921
rect 282328 170912 282330 170921
rect 282274 170847 282330 170856
rect 282828 169720 282880 169726
rect 282828 169662 282880 169668
rect 282840 169425 282868 169662
rect 282826 169416 282882 169425
rect 282826 169351 282882 169360
rect 282276 168360 282328 168366
rect 282276 168302 282328 168308
rect 282288 167929 282316 168302
rect 282274 167920 282330 167929
rect 282274 167855 282330 167864
rect 282826 165608 282882 165617
rect 282932 165594 282960 296686
rect 283012 294024 283064 294030
rect 283012 293966 283064 293972
rect 283024 182073 283052 293966
rect 283102 207768 283158 207777
rect 283102 207703 283158 207712
rect 283010 182064 283066 182073
rect 283010 181999 283066 182008
rect 283012 175976 283064 175982
rect 283012 175918 283064 175924
rect 282882 165566 282960 165594
rect 282826 165543 282882 165552
rect 281908 165368 281960 165374
rect 281908 165310 281960 165316
rect 281920 164937 281948 165310
rect 281906 164928 281962 164937
rect 281906 164863 281962 164872
rect 282826 164112 282882 164121
rect 282826 164047 282882 164056
rect 282840 163334 282868 164047
rect 282828 163328 282880 163334
rect 282828 163270 282880 163276
rect 282828 162852 282880 162858
rect 282828 162794 282880 162800
rect 282840 161809 282868 162794
rect 282826 161800 282882 161809
rect 282826 161735 282882 161744
rect 281644 161446 281856 161474
rect 281644 157334 281672 161446
rect 282828 161424 282880 161430
rect 282828 161366 282880 161372
rect 282840 161129 282868 161366
rect 282826 161120 282882 161129
rect 282826 161055 282882 161064
rect 281724 160608 281776 160614
rect 281724 160550 281776 160556
rect 281736 160313 281764 160550
rect 281722 160304 281778 160313
rect 281722 160239 281778 160248
rect 281908 160064 281960 160070
rect 281908 160006 281960 160012
rect 281920 159497 281948 160006
rect 282368 159996 282420 160002
rect 282368 159938 282420 159944
rect 281906 159488 281962 159497
rect 281906 159423 281962 159432
rect 282380 158817 282408 159938
rect 282366 158808 282422 158817
rect 282366 158743 282422 158752
rect 282826 157992 282882 158001
rect 282826 157927 282882 157936
rect 282840 157622 282868 157927
rect 282828 157616 282880 157622
rect 282828 157558 282880 157564
rect 281644 157306 281764 157334
rect 281632 155916 281684 155922
rect 281632 155858 281684 155864
rect 281644 155009 281672 155858
rect 281630 155000 281686 155009
rect 281630 154935 281686 154944
rect 281632 154488 281684 154494
rect 281632 154430 281684 154436
rect 281644 154193 281672 154430
rect 281630 154184 281686 154193
rect 281630 154119 281686 154128
rect 281632 153196 281684 153202
rect 281632 153138 281684 153144
rect 281644 152697 281672 153138
rect 281630 152688 281686 152697
rect 281630 152623 281686 152632
rect 281632 152516 281684 152522
rect 281632 152458 281684 152464
rect 281644 151201 281672 152458
rect 281736 151881 281764 157306
rect 282182 153776 282238 153785
rect 282182 153711 282238 153720
rect 281722 151872 281778 151881
rect 281722 151807 281778 151816
rect 281630 151192 281686 151201
rect 281630 151127 281686 151136
rect 281816 151088 281868 151094
rect 281816 151030 281868 151036
rect 281632 150408 281684 150414
rect 281630 150376 281632 150385
rect 281684 150376 281686 150385
rect 281630 150311 281686 150320
rect 281724 150340 281776 150346
rect 281724 150282 281776 150288
rect 281736 149705 281764 150282
rect 281722 149696 281778 149705
rect 281722 149631 281778 149640
rect 281632 149048 281684 149054
rect 281632 148990 281684 148996
rect 281644 148073 281672 148990
rect 281828 148889 281856 151030
rect 281814 148880 281870 148889
rect 281814 148815 281870 148824
rect 281630 148064 281686 148073
rect 281630 147999 281686 148008
rect 282092 142112 282144 142118
rect 282092 142054 282144 142060
rect 282104 141273 282132 142054
rect 282090 141264 282146 141273
rect 282090 141199 282146 141208
rect 282196 132161 282224 153711
rect 283024 151814 283052 175918
rect 283116 153513 283144 207703
rect 284312 198762 284340 377590
rect 285692 358154 285720 377590
rect 286324 373312 286376 373318
rect 286324 373254 286376 373260
rect 285680 358148 285732 358154
rect 285680 358090 285732 358096
rect 284942 298344 284998 298353
rect 284942 298279 284998 298288
rect 284392 203584 284444 203590
rect 284392 203526 284444 203532
rect 284300 198756 284352 198762
rect 284300 198698 284352 198704
rect 284312 198665 284340 198698
rect 284298 198656 284354 198665
rect 284298 198591 284354 198600
rect 284300 196648 284352 196654
rect 284300 196590 284352 196596
rect 283564 184204 283616 184210
rect 283564 184146 283616 184152
rect 283196 181552 283248 181558
rect 283196 181494 283248 181500
rect 283208 175982 283236 181494
rect 283576 176050 283604 184146
rect 283564 176044 283616 176050
rect 283564 175986 283616 175992
rect 283196 175976 283248 175982
rect 283196 175918 283248 175924
rect 283196 175840 283248 175846
rect 283196 175782 283248 175788
rect 283102 153504 283158 153513
rect 283102 153439 283158 153448
rect 282932 151786 283052 151814
rect 282828 147620 282880 147626
rect 282828 147562 282880 147568
rect 282840 147393 282868 147562
rect 282826 147384 282882 147393
rect 282826 147319 282882 147328
rect 282368 146260 282420 146266
rect 282368 146202 282420 146208
rect 282380 145081 282408 146202
rect 282366 145072 282422 145081
rect 282366 145007 282422 145016
rect 282828 143540 282880 143546
rect 282828 143482 282880 143488
rect 282840 142769 282868 143482
rect 282826 142760 282882 142769
rect 282826 142695 282882 142704
rect 282826 142080 282882 142089
rect 282826 142015 282828 142024
rect 282880 142015 282882 142024
rect 282828 141986 282880 141992
rect 282828 140752 282880 140758
rect 282828 140694 282880 140700
rect 282840 139777 282868 140694
rect 282826 139768 282882 139777
rect 282826 139703 282882 139712
rect 282828 139392 282880 139398
rect 282828 139334 282880 139340
rect 282840 138961 282868 139334
rect 282826 138952 282882 138961
rect 282826 138887 282882 138896
rect 282826 138272 282882 138281
rect 282932 138258 282960 151786
rect 283208 142154 283236 175782
rect 282882 138230 282960 138258
rect 283024 142126 283236 142154
rect 282826 138207 282882 138216
rect 282828 137964 282880 137970
rect 282828 137906 282880 137912
rect 282840 137465 282868 137906
rect 282826 137456 282882 137465
rect 282826 137391 282882 137400
rect 282826 136640 282882 136649
rect 282826 136575 282828 136584
rect 282880 136575 282882 136584
rect 282828 136546 282880 136552
rect 282826 136368 282882 136377
rect 283024 136354 283052 142126
rect 282882 136326 283052 136354
rect 282826 136303 282882 136312
rect 282460 135176 282512 135182
rect 282460 135118 282512 135124
rect 282472 134473 282500 135118
rect 282458 134464 282514 134473
rect 282458 134399 282514 134408
rect 282736 133884 282788 133890
rect 282736 133826 282788 133832
rect 282748 132841 282776 133826
rect 282828 133816 282880 133822
rect 282828 133758 282880 133764
rect 282840 133657 282868 133758
rect 282826 133648 282882 133657
rect 282826 133583 282882 133592
rect 282734 132832 282790 132841
rect 282734 132767 282790 132776
rect 282828 132456 282880 132462
rect 282828 132398 282880 132404
rect 282182 132152 282238 132161
rect 282182 132087 282238 132096
rect 282840 131345 282868 132398
rect 282826 131336 282882 131345
rect 282826 131271 282882 131280
rect 282828 131096 282880 131102
rect 282828 131038 282880 131044
rect 282736 131028 282788 131034
rect 282736 130970 282788 130976
rect 282748 129849 282776 130970
rect 282840 130665 282868 131038
rect 282826 130656 282882 130665
rect 282826 130591 282882 130600
rect 282734 129840 282790 129849
rect 282734 129775 282790 129784
rect 284312 129742 284340 196590
rect 281816 129736 281868 129742
rect 281816 129678 281868 129684
rect 284300 129736 284352 129742
rect 284300 129678 284352 129684
rect 281828 129033 281856 129678
rect 283564 129056 283616 129062
rect 281814 129024 281870 129033
rect 283564 128998 283616 129004
rect 281814 128959 281870 128968
rect 282826 128344 282882 128353
rect 282826 128279 282828 128288
rect 282880 128279 282882 128288
rect 282828 128250 282880 128256
rect 282736 128240 282788 128246
rect 282736 128182 282788 128188
rect 282748 127537 282776 128182
rect 282734 127528 282790 127537
rect 282734 127463 282790 127472
rect 282368 126948 282420 126954
rect 282368 126890 282420 126896
rect 282092 126268 282144 126274
rect 282092 126210 282144 126216
rect 282104 123049 282132 126210
rect 282380 126041 282408 126890
rect 282366 126032 282422 126041
rect 282366 125967 282422 125976
rect 282828 125588 282880 125594
rect 282828 125530 282880 125536
rect 282736 125520 282788 125526
rect 282736 125462 282788 125468
rect 282748 124545 282776 125462
rect 282840 125225 282868 125530
rect 282826 125216 282882 125225
rect 282826 125151 282882 125160
rect 282734 124536 282790 124545
rect 282734 124471 282790 124480
rect 282826 123720 282882 123729
rect 282826 123655 282828 123664
rect 282880 123655 282882 123664
rect 282828 123626 282880 123632
rect 282184 123480 282236 123486
rect 282184 123422 282236 123428
rect 282090 123040 282146 123049
rect 282090 122975 282146 122984
rect 282092 120964 282144 120970
rect 282092 120906 282144 120912
rect 282104 120737 282132 120906
rect 282090 120728 282146 120737
rect 282090 120663 282146 120672
rect 281538 119232 281594 119241
rect 281538 119167 281594 119176
rect 281724 113824 281776 113830
rect 281724 113766 281776 113772
rect 279068 113146 279372 113174
rect 267738 111208 267794 111217
rect 267738 111143 267794 111152
rect 267646 100464 267702 100473
rect 267646 100399 267702 100408
rect 267660 95266 267688 100399
rect 267648 95260 267700 95266
rect 267648 95202 267700 95208
rect 267186 82104 267242 82113
rect 267186 82039 267242 82048
rect 267094 65648 267150 65657
rect 267094 65583 267150 65592
rect 267752 57254 267780 111143
rect 279344 100609 279372 113146
rect 281736 109993 281764 113766
rect 282196 112305 282224 123422
rect 282828 122800 282880 122806
rect 282828 122742 282880 122748
rect 282840 122233 282868 122742
rect 282826 122224 282882 122233
rect 282826 122159 282882 122168
rect 282644 122120 282696 122126
rect 282644 122062 282696 122068
rect 282656 114617 282684 122062
rect 282828 121440 282880 121446
rect 282826 121408 282828 121417
rect 282880 121408 282882 121417
rect 282826 121343 282882 121352
rect 282828 120080 282880 120086
rect 282828 120022 282880 120028
rect 282840 119921 282868 120022
rect 282826 119912 282882 119921
rect 282826 119847 282882 119856
rect 282828 118652 282880 118658
rect 282828 118594 282880 118600
rect 282840 118425 282868 118594
rect 282826 118416 282882 118425
rect 282826 118351 282882 118360
rect 282734 118008 282790 118017
rect 282734 117943 282790 117952
rect 282828 117972 282880 117978
rect 282748 116113 282776 117943
rect 282828 117914 282880 117920
rect 282840 117609 282868 117914
rect 282826 117600 282882 117609
rect 282826 117535 282882 117544
rect 282826 116920 282882 116929
rect 282826 116855 282882 116864
rect 282840 116618 282868 116855
rect 282828 116612 282880 116618
rect 282828 116554 282880 116560
rect 282734 116104 282790 116113
rect 282734 116039 282790 116048
rect 282828 115932 282880 115938
rect 282828 115874 282880 115880
rect 282840 115433 282868 115874
rect 282826 115424 282882 115433
rect 282826 115359 282882 115368
rect 282642 114608 282698 114617
rect 282642 114543 282698 114552
rect 282828 114164 282880 114170
rect 282828 114106 282880 114112
rect 282840 113801 282868 114106
rect 282826 113792 282882 113801
rect 282826 113727 282882 113736
rect 282828 113144 282880 113150
rect 282826 113112 282828 113121
rect 282880 113112 282882 113121
rect 282826 113047 282882 113056
rect 282182 112296 282238 112305
rect 282182 112231 282238 112240
rect 282828 111784 282880 111790
rect 282828 111726 282880 111732
rect 282092 111648 282144 111654
rect 282090 111616 282092 111625
rect 282144 111616 282146 111625
rect 282090 111551 282146 111560
rect 282840 110809 282868 111726
rect 282826 110800 282882 110809
rect 282826 110735 282882 110744
rect 282644 110424 282696 110430
rect 282644 110366 282696 110372
rect 281722 109984 281778 109993
rect 281722 109919 281778 109928
rect 282656 109313 282684 110366
rect 282642 109304 282698 109313
rect 282642 109239 282698 109248
rect 281724 108996 281776 109002
rect 281724 108938 281776 108944
rect 281736 108497 281764 108938
rect 282828 108928 282880 108934
rect 282828 108870 282880 108876
rect 281722 108488 281778 108497
rect 281722 108423 281778 108432
rect 282840 107817 282868 108870
rect 282826 107808 282882 107817
rect 282826 107743 282882 107752
rect 282826 106992 282882 107001
rect 282826 106927 282828 106936
rect 282880 106927 282882 106936
rect 282828 106898 282880 106904
rect 282828 106276 282880 106282
rect 282828 106218 282880 106224
rect 282840 106185 282868 106218
rect 282826 106176 282882 106185
rect 282826 106111 282882 106120
rect 282826 105496 282882 105505
rect 282826 105431 282882 105440
rect 282840 105330 282868 105431
rect 282828 105324 282880 105330
rect 282828 105266 282880 105272
rect 282828 104848 282880 104854
rect 282828 104790 282880 104796
rect 281540 104780 281592 104786
rect 281540 104722 281592 104728
rect 281552 104009 281580 104722
rect 282840 104689 282868 104790
rect 282826 104680 282882 104689
rect 282826 104615 282882 104624
rect 281538 104000 281594 104009
rect 281538 103935 281594 103944
rect 282092 103488 282144 103494
rect 282092 103430 282144 103436
rect 282104 103193 282132 103430
rect 282090 103184 282146 103193
rect 282090 103119 282146 103128
rect 282276 102128 282328 102134
rect 282276 102070 282328 102076
rect 282288 101697 282316 102070
rect 282274 101688 282330 101697
rect 282274 101623 282330 101632
rect 281538 100872 281594 100881
rect 281538 100807 281594 100816
rect 279330 100600 279386 100609
rect 279330 100535 279386 100544
rect 279330 98152 279386 98161
rect 279330 98087 279386 98096
rect 267832 95940 267884 95946
rect 267832 95882 267884 95888
rect 267844 93838 267872 95882
rect 269212 95260 269264 95266
rect 269212 95202 269264 95208
rect 267924 93900 267976 93906
rect 267924 93842 267976 93848
rect 267832 93832 267884 93838
rect 267832 93774 267884 93780
rect 267936 84194 267964 93842
rect 269118 92576 269174 92585
rect 269118 92511 269174 92520
rect 267844 84166 267964 84194
rect 267740 57248 267792 57254
rect 267740 57190 267792 57196
rect 267002 53136 267058 53145
rect 267002 53071 267058 53080
rect 266358 37224 266414 37233
rect 266358 37159 266414 37168
rect 264978 22672 265034 22681
rect 264978 22607 265034 22616
rect 264244 10396 264296 10402
rect 264244 10338 264296 10344
rect 264992 490 265020 22607
rect 266372 16574 266400 37159
rect 267844 25566 267872 84166
rect 268382 43480 268438 43489
rect 268382 43415 268438 43424
rect 267832 25560 267884 25566
rect 267832 25502 267884 25508
rect 266372 16546 266584 16574
rect 265176 598 265388 626
rect 265176 490 265204 598
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 264992 462 265204 490
rect 265360 480 265388 598
rect 266556 480 266584 16546
rect 268290 13016 268346 13025
rect 268290 12951 268346 12960
rect 267738 4040 267794 4049
rect 267738 3975 267794 3984
rect 267752 480 267780 3975
rect 268304 490 268332 12951
rect 268396 3194 268424 43415
rect 269132 35222 269160 92511
rect 269224 51785 269252 95202
rect 270590 95024 270646 95033
rect 270590 94959 270646 94968
rect 270498 93256 270554 93265
rect 270498 93191 270554 93200
rect 269210 51776 269266 51785
rect 269210 51711 269266 51720
rect 270512 40730 270540 93191
rect 270604 46306 270632 94959
rect 274008 93838 274036 96084
rect 278778 95840 278834 95849
rect 278778 95775 278834 95784
rect 278792 95169 278820 95775
rect 279344 95198 279372 98087
rect 279332 95192 279384 95198
rect 278778 95160 278834 95169
rect 279332 95134 279384 95140
rect 278778 95095 278834 95104
rect 273996 93832 274048 93838
rect 273996 93774 274048 93780
rect 276756 93152 276808 93158
rect 276756 93094 276808 93100
rect 273258 91760 273314 91769
rect 273258 91695 273314 91704
rect 270592 46300 270644 46306
rect 270592 46242 270644 46248
rect 270500 40724 270552 40730
rect 270500 40666 270552 40672
rect 269120 35216 269172 35222
rect 269120 35158 269172 35164
rect 269118 30968 269174 30977
rect 269118 30903 269174 30912
rect 269132 16574 269160 30903
rect 269132 16546 270080 16574
rect 268474 10296 268530 10305
rect 268474 10231 268530 10240
rect 268488 4049 268516 10231
rect 268474 4040 268530 4049
rect 268474 3975 268530 3984
rect 268384 3188 268436 3194
rect 268384 3130 268436 3136
rect 268672 598 268884 626
rect 268672 490 268700 598
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268304 462 268700 490
rect 268856 480 268884 598
rect 270052 480 270080 16546
rect 270774 11656 270830 11665
rect 270774 11591 270830 11600
rect 270788 490 270816 11591
rect 272432 2100 272484 2106
rect 272432 2042 272484 2048
rect 271064 598 271276 626
rect 271064 490 271092 598
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 270788 462 271092 490
rect 271248 480 271276 598
rect 272444 480 272472 2042
rect 273272 490 273300 91695
rect 276768 91089 276796 93094
rect 276018 91080 276074 91089
rect 276018 91015 276074 91024
rect 276754 91080 276810 91089
rect 276754 91015 276810 91024
rect 274640 47660 274692 47666
rect 274640 47602 274692 47608
rect 274652 16574 274680 47602
rect 276032 17270 276060 91015
rect 281552 88233 281580 100807
rect 282000 100020 282052 100026
rect 282000 99962 282052 99968
rect 281630 99376 281686 99385
rect 281630 99311 281632 99320
rect 281684 99311 281686 99320
rect 281632 99282 281684 99288
rect 282012 97889 282040 99962
rect 283576 99346 283604 128998
rect 284404 104786 284432 203526
rect 284956 180130 284984 298279
rect 286048 271176 286100 271182
rect 286048 271118 286100 271124
rect 286060 270609 286088 271118
rect 285770 270600 285826 270609
rect 285770 270535 285826 270544
rect 286046 270600 286102 270609
rect 286046 270535 286102 270544
rect 285678 223000 285734 223009
rect 285678 222935 285734 222944
rect 285034 215928 285090 215937
rect 285034 215863 285090 215872
rect 284944 180124 284996 180130
rect 284944 180066 284996 180072
rect 284484 179444 284536 179450
rect 284484 179386 284536 179392
rect 284496 160614 284524 179386
rect 285048 176905 285076 215863
rect 285034 176896 285090 176905
rect 285034 176831 285090 176840
rect 284576 176044 284628 176050
rect 284576 175986 284628 175992
rect 284588 165374 284616 175986
rect 284576 165368 284628 165374
rect 284576 165310 284628 165316
rect 284484 160608 284536 160614
rect 284484 160550 284536 160556
rect 285692 120970 285720 222935
rect 285784 175234 285812 270535
rect 286336 238754 286364 373254
rect 287072 369889 287100 377590
rect 289648 375329 289676 377604
rect 291212 377590 291318 377618
rect 292592 377590 292974 377618
rect 293972 377590 294630 377618
rect 289634 375320 289690 375329
rect 289634 375255 289690 375264
rect 287058 369880 287114 369889
rect 287058 369815 287114 369824
rect 287702 369880 287758 369889
rect 287702 369815 287758 369824
rect 287060 311160 287112 311166
rect 287060 311102 287112 311108
rect 285876 238726 286364 238754
rect 285876 238377 285904 238726
rect 285862 238368 285918 238377
rect 285862 238303 285918 238312
rect 285772 175228 285824 175234
rect 285772 175170 285824 175176
rect 285772 175092 285824 175098
rect 285772 175034 285824 175040
rect 285784 170950 285812 175034
rect 285772 170944 285824 170950
rect 285772 170886 285824 170892
rect 285876 156670 285904 238303
rect 285956 185632 286008 185638
rect 285956 185574 286008 185580
rect 285864 156664 285916 156670
rect 285864 156606 285916 156612
rect 285968 135182 285996 185574
rect 285956 135176 286008 135182
rect 285956 135118 286008 135124
rect 285680 120964 285732 120970
rect 285680 120906 285732 120912
rect 284944 119400 284996 119406
rect 284944 119342 284996 119348
rect 284956 111654 284984 119342
rect 284944 111648 284996 111654
rect 284944 111590 284996 111596
rect 287072 106962 287100 311102
rect 287152 269816 287204 269822
rect 287152 269758 287204 269764
rect 287164 126954 287192 269758
rect 287716 229770 287744 369815
rect 289084 330608 289136 330614
rect 289084 330550 289136 330556
rect 289096 278662 289124 330550
rect 289084 278656 289136 278662
rect 289084 278598 289136 278604
rect 289820 273964 289872 273970
rect 289820 273906 289872 273912
rect 288440 272536 288492 272542
rect 288440 272478 288492 272484
rect 287704 229764 287756 229770
rect 287704 229706 287756 229712
rect 287244 225616 287296 225622
rect 287244 225558 287296 225564
rect 287152 126948 287204 126954
rect 287152 126890 287204 126896
rect 287256 114170 287284 225558
rect 287336 177404 287388 177410
rect 287336 177346 287388 177352
rect 287348 157622 287376 177346
rect 287336 157616 287388 157622
rect 287336 157558 287388 157564
rect 288452 123690 288480 272478
rect 288532 241460 288584 241466
rect 288532 241402 288584 241408
rect 288544 240174 288572 241402
rect 288532 240168 288584 240174
rect 288532 240110 288584 240116
rect 288440 123684 288492 123690
rect 288440 123626 288492 123632
rect 287244 114164 287296 114170
rect 287244 114106 287296 114112
rect 287060 106956 287112 106962
rect 287060 106898 287112 106904
rect 288544 105330 288572 240110
rect 288624 231124 288676 231130
rect 288624 231066 288676 231072
rect 288636 117978 288664 231066
rect 288716 181484 288768 181490
rect 288716 181426 288768 181432
rect 288728 163334 288756 181426
rect 288716 163328 288768 163334
rect 288716 163270 288768 163276
rect 289832 153785 289860 273906
rect 291212 241466 291240 377590
rect 292592 331906 292620 377590
rect 293972 373318 294000 377590
rect 296272 374678 296300 377604
rect 296260 374672 296312 374678
rect 296260 374614 296312 374620
rect 297928 374066 297956 377604
rect 299492 377590 299598 377618
rect 300872 377590 301254 377618
rect 302344 377590 302910 377618
rect 294604 374060 294656 374066
rect 294604 374002 294656 374008
rect 297916 374060 297968 374066
rect 297916 374002 297968 374008
rect 293960 373312 294012 373318
rect 293960 373254 294012 373260
rect 292580 331900 292632 331906
rect 292580 331842 292632 331848
rect 292580 298784 292632 298790
rect 292580 298726 292632 298732
rect 292592 298178 292620 298726
rect 292580 298172 292632 298178
rect 292580 298114 292632 298120
rect 291844 244928 291896 244934
rect 291844 244870 291896 244876
rect 291200 241460 291252 241466
rect 291200 241402 291252 241408
rect 291198 219464 291254 219473
rect 291198 219399 291254 219408
rect 289910 209128 289966 209137
rect 289910 209063 289966 209072
rect 289818 153776 289874 153785
rect 289818 153711 289874 153720
rect 289924 121446 289952 209063
rect 290004 200864 290056 200870
rect 290004 200806 290056 200812
rect 290016 143546 290044 200806
rect 290094 176760 290150 176769
rect 290094 176695 290150 176704
rect 290108 168366 290136 176695
rect 290096 168360 290148 168366
rect 290096 168302 290148 168308
rect 290004 143540 290056 143546
rect 290004 143482 290056 143488
rect 289912 121440 289964 121446
rect 289912 121382 289964 121388
rect 288624 117972 288676 117978
rect 288624 117914 288676 117920
rect 290646 117328 290702 117337
rect 290646 117263 290648 117272
rect 290700 117263 290702 117272
rect 290648 117234 290700 117240
rect 290660 116618 290688 117234
rect 290648 116612 290700 116618
rect 290648 116554 290700 116560
rect 291212 106282 291240 219399
rect 291292 214600 291344 214606
rect 291292 214542 291344 214548
rect 291200 106276 291252 106282
rect 291200 106218 291252 106224
rect 288532 105324 288584 105330
rect 288532 105266 288584 105272
rect 284392 104780 284444 104786
rect 284392 104722 284444 104728
rect 291304 103494 291332 214542
rect 291474 195392 291530 195401
rect 291474 195327 291530 195336
rect 291384 182844 291436 182850
rect 291384 182786 291436 182792
rect 291396 104854 291424 182786
rect 291488 146266 291516 195327
rect 291856 193866 291884 244870
rect 291844 193860 291896 193866
rect 291844 193802 291896 193808
rect 291476 146260 291528 146266
rect 291476 146202 291528 146208
rect 292592 125526 292620 298114
rect 294052 258732 294104 258738
rect 294052 258674 294104 258680
rect 293960 230444 294012 230450
rect 293960 230386 294012 230392
rect 293972 229158 294000 230386
rect 293960 229152 294012 229158
rect 293960 229094 294012 229100
rect 292672 192500 292724 192506
rect 292672 192442 292724 192448
rect 292684 150346 292712 192442
rect 292856 186380 292908 186386
rect 292856 186322 292908 186328
rect 292764 178696 292816 178702
rect 292764 178638 292816 178644
rect 292776 160002 292804 178638
rect 292868 169726 292896 186322
rect 292856 169720 292908 169726
rect 292856 169662 292908 169668
rect 292764 159996 292816 160002
rect 292764 159938 292816 159944
rect 292672 150340 292724 150346
rect 292672 150282 292724 150288
rect 292580 125520 292632 125526
rect 292580 125462 292632 125468
rect 293972 118658 294000 229094
rect 294064 149054 294092 258674
rect 294616 230450 294644 374002
rect 295982 355464 296038 355473
rect 295982 355399 296038 355408
rect 295996 325038 296024 355399
rect 295984 325032 296036 325038
rect 295984 324974 296036 324980
rect 298008 318096 298060 318102
rect 298008 318038 298060 318044
rect 298020 317490 298048 318038
rect 296904 317484 296956 317490
rect 296904 317426 296956 317432
rect 298008 317484 298060 317490
rect 298008 317426 298060 317432
rect 296810 296848 296866 296857
rect 296810 296783 296866 296792
rect 295340 269884 295392 269890
rect 295340 269826 295392 269832
rect 294604 230444 294656 230450
rect 294604 230386 294656 230392
rect 294604 198756 294656 198762
rect 294604 198698 294656 198704
rect 294142 181384 294198 181393
rect 294142 181319 294198 181328
rect 294156 150414 294184 181319
rect 294144 150408 294196 150414
rect 294144 150350 294196 150356
rect 294052 149048 294104 149054
rect 294052 148990 294104 148996
rect 293960 118652 294012 118658
rect 293960 118594 294012 118600
rect 291384 104848 291436 104854
rect 291384 104790 291436 104796
rect 291292 103488 291344 103494
rect 291292 103430 291344 103436
rect 283564 99340 283616 99346
rect 283564 99282 283616 99288
rect 281998 97880 282054 97889
rect 281998 97815 282054 97824
rect 282184 97300 282236 97306
rect 282184 97242 282236 97248
rect 281538 88224 281594 88233
rect 281538 88159 281594 88168
rect 277398 87544 277454 87553
rect 277398 87479 277454 87488
rect 276110 68232 276166 68241
rect 276110 68167 276166 68176
rect 276124 67561 276152 68167
rect 276110 67552 276166 67561
rect 276110 67487 276166 67496
rect 277306 67552 277362 67561
rect 277306 67487 277362 67496
rect 276020 17264 276072 17270
rect 276020 17206 276072 17212
rect 274652 16546 274864 16574
rect 273456 598 273668 626
rect 273456 490 273484 598
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273272 462 273484 490
rect 273640 480 273668 598
rect 274836 480 274864 16546
rect 277122 3496 277178 3505
rect 277122 3431 277178 3440
rect 276020 3188 276072 3194
rect 276020 3130 276072 3136
rect 276032 480 276060 3130
rect 277136 480 277164 3431
rect 277320 3369 277348 67487
rect 277412 16574 277440 87479
rect 280158 86184 280214 86193
rect 280158 86119 280214 86128
rect 278778 37904 278834 37913
rect 278778 37839 278834 37848
rect 278792 16574 278820 37839
rect 280172 16574 280200 86119
rect 280802 19952 280858 19961
rect 280802 19887 280858 19896
rect 277412 16546 278360 16574
rect 278792 16546 279096 16574
rect 280172 16546 280752 16574
rect 277306 3360 277362 3369
rect 277306 3295 277362 3304
rect 278332 480 278360 16546
rect 279068 490 279096 16546
rect 279344 598 279556 626
rect 279344 490 279372 598
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279068 462 279372 490
rect 279528 480 279556 598
rect 280724 480 280752 16546
rect 280816 3194 280844 19887
rect 281906 4856 281962 4865
rect 281906 4791 281962 4800
rect 280804 3188 280856 3194
rect 280804 3130 280856 3136
rect 281920 480 281948 4791
rect 282196 4078 282224 97242
rect 285678 93120 285734 93129
rect 285678 93055 285734 93064
rect 284944 83496 284996 83502
rect 284944 83438 284996 83444
rect 284956 6186 284984 83438
rect 285692 16574 285720 93055
rect 291844 19984 291896 19990
rect 289818 19952 289874 19961
rect 291844 19926 291896 19932
rect 289818 19887 289874 19896
rect 285692 16546 286640 16574
rect 284944 6180 284996 6186
rect 284944 6122 284996 6128
rect 282184 4072 282236 4078
rect 282184 4014 282236 4020
rect 284298 3360 284354 3369
rect 284298 3295 284354 3304
rect 285402 3360 285458 3369
rect 285402 3295 285458 3304
rect 283104 3188 283156 3194
rect 283104 3130 283156 3136
rect 283116 480 283144 3130
rect 284312 480 284340 3295
rect 285416 480 285444 3295
rect 286612 480 286640 16546
rect 287794 3496 287850 3505
rect 287794 3431 287850 3440
rect 288992 3460 289044 3466
rect 287808 480 287836 3431
rect 288992 3402 289044 3408
rect 289004 480 289032 3402
rect 289832 490 289860 19887
rect 291856 3534 291884 19926
rect 294616 16574 294644 198698
rect 295352 110430 295380 269826
rect 295984 249076 296036 249082
rect 295984 249018 296036 249024
rect 295996 235278 296024 249018
rect 295984 235272 296036 235278
rect 295984 235214 296036 235220
rect 295996 234666 296024 235214
rect 295524 234660 295576 234666
rect 295524 234602 295576 234608
rect 295984 234660 296036 234666
rect 295984 234602 296036 234608
rect 295432 222896 295484 222902
rect 295432 222838 295484 222844
rect 295444 111790 295472 222838
rect 295536 152522 295564 234602
rect 296718 205048 296774 205057
rect 296718 204983 296774 204992
rect 295616 188420 295668 188426
rect 295616 188362 295668 188368
rect 295628 154494 295656 188362
rect 295616 154488 295668 154494
rect 295616 154430 295668 154436
rect 295524 152516 295576 152522
rect 295524 152458 295576 152464
rect 295432 111784 295484 111790
rect 295432 111726 295484 111732
rect 295340 110424 295392 110430
rect 295340 110366 295392 110372
rect 294616 16546 294920 16574
rect 291844 3528 291896 3534
rect 291382 3496 291438 3505
rect 291844 3470 291896 3476
rect 292580 3528 292632 3534
rect 292580 3470 292632 3476
rect 293682 3496 293738 3505
rect 291382 3431 291438 3440
rect 290016 598 290228 626
rect 290016 490 290044 598
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 289832 462 290044 490
rect 290200 480 290228 598
rect 291396 480 291424 3431
rect 292592 480 292620 3470
rect 293682 3431 293738 3440
rect 293696 480 293724 3431
rect 294892 480 294920 16546
rect 296076 4140 296128 4146
rect 296076 4082 296128 4088
rect 296088 480 296116 4082
rect 296732 3466 296760 204983
rect 296824 102134 296852 296783
rect 296916 162858 296944 317426
rect 298742 296032 298798 296041
rect 298742 295967 298798 295976
rect 298190 291272 298246 291281
rect 298190 291207 298246 291216
rect 298098 216064 298154 216073
rect 298098 215999 298154 216008
rect 296996 178764 297048 178770
rect 296996 178706 297048 178712
rect 296904 162852 296956 162858
rect 296904 162794 296956 162800
rect 297008 153202 297036 178706
rect 296996 153196 297048 153202
rect 296996 153138 297048 153144
rect 296812 102128 296864 102134
rect 296812 102070 296864 102076
rect 297272 15904 297324 15910
rect 297272 15846 297324 15852
rect 296720 3460 296772 3466
rect 296720 3402 296772 3408
rect 297284 480 297312 15846
rect 298112 4146 298140 215999
rect 298204 122806 298232 291207
rect 298284 280832 298336 280838
rect 298284 280774 298336 280780
rect 298296 142050 298324 280774
rect 298756 235793 298784 295967
rect 299492 241505 299520 377590
rect 299570 293992 299626 294001
rect 299570 293927 299626 293936
rect 299478 241496 299534 241505
rect 299478 241431 299534 241440
rect 298742 235784 298798 235793
rect 298742 235719 298798 235728
rect 299480 188352 299532 188358
rect 299480 188294 299532 188300
rect 298376 180124 298428 180130
rect 298376 180066 298428 180072
rect 298284 142044 298336 142050
rect 298284 141986 298336 141992
rect 298192 122800 298244 122806
rect 298192 122742 298244 122748
rect 298388 120086 298416 180066
rect 299492 142118 299520 188294
rect 299480 142112 299532 142118
rect 299480 142054 299532 142060
rect 298376 120080 298428 120086
rect 298376 120022 298428 120028
rect 299584 113830 299612 293927
rect 300768 253224 300820 253230
rect 300768 253166 300820 253172
rect 300780 252618 300808 253166
rect 299664 252612 299716 252618
rect 299664 252554 299716 252560
rect 300768 252612 300820 252618
rect 300768 252554 300820 252560
rect 299676 137970 299704 252554
rect 300872 249082 300900 377590
rect 302238 342136 302294 342145
rect 302238 342071 302294 342080
rect 302252 340921 302280 342071
rect 302238 340912 302294 340921
rect 302238 340847 302294 340856
rect 300952 285728 301004 285734
rect 300952 285670 301004 285676
rect 300860 249076 300912 249082
rect 300860 249018 300912 249024
rect 300860 242208 300912 242214
rect 300860 242150 300912 242156
rect 300872 241534 300900 242150
rect 300860 241528 300912 241534
rect 300860 241470 300912 241476
rect 300122 200696 300178 200705
rect 300122 200631 300178 200640
rect 299664 137964 299716 137970
rect 299664 137906 299716 137912
rect 299572 113824 299624 113830
rect 299572 113766 299624 113772
rect 300136 13802 300164 200631
rect 300872 151094 300900 241470
rect 300860 151088 300912 151094
rect 300860 151030 300912 151036
rect 300964 133822 300992 285670
rect 302148 227112 302200 227118
rect 302148 227054 302200 227060
rect 302160 226953 302188 227054
rect 302146 226944 302202 226953
rect 302146 226879 302202 226888
rect 301136 193860 301188 193866
rect 301136 193802 301188 193808
rect 301042 187096 301098 187105
rect 301042 187031 301098 187040
rect 300952 133816 301004 133822
rect 300952 133758 301004 133764
rect 301056 115938 301084 187031
rect 301148 129062 301176 193802
rect 302160 188358 302188 226879
rect 302148 188352 302200 188358
rect 302148 188294 302200 188300
rect 301136 129056 301188 129062
rect 301136 128998 301188 129004
rect 301044 115932 301096 115938
rect 301044 115874 301096 115880
rect 302252 60110 302280 340847
rect 302344 282198 302372 377590
rect 304264 374876 304316 374882
rect 304264 374818 304316 374824
rect 304276 349081 304304 374818
rect 304552 374649 304580 377604
rect 306208 374882 306236 377604
rect 307878 377590 308444 377618
rect 307022 375320 307078 375329
rect 307022 375255 307078 375264
rect 306196 374876 306248 374882
rect 306196 374818 306248 374824
rect 304538 374640 304594 374649
rect 304538 374575 304594 374584
rect 305644 354000 305696 354006
rect 305644 353942 305696 353948
rect 304262 349072 304318 349081
rect 304262 349007 304318 349016
rect 304276 348401 304304 349007
rect 304262 348392 304318 348401
rect 304262 348327 304318 348336
rect 304264 341556 304316 341562
rect 304264 341498 304316 341504
rect 304276 310457 304304 341498
rect 303710 310448 303766 310457
rect 303710 310383 303766 310392
rect 304262 310448 304318 310457
rect 304262 310383 304318 310392
rect 303724 309777 303752 310383
rect 303710 309768 303766 309777
rect 303710 309703 303766 309712
rect 302424 301504 302476 301510
rect 302424 301446 302476 301452
rect 302332 282192 302384 282198
rect 302332 282134 302384 282140
rect 302332 227044 302384 227050
rect 302332 226986 302384 226992
rect 302344 226370 302372 226986
rect 302332 226364 302384 226370
rect 302332 226306 302384 226312
rect 302344 118017 302372 226306
rect 302436 173874 302464 301446
rect 302884 282192 302936 282198
rect 302884 282134 302936 282140
rect 302896 227118 302924 282134
rect 302884 227112 302936 227118
rect 302884 227054 302936 227060
rect 303618 211848 303674 211857
rect 303618 211783 303674 211792
rect 302514 189816 302570 189825
rect 302514 189751 302570 189760
rect 302424 173868 302476 173874
rect 302424 173810 302476 173816
rect 302528 139398 302556 189751
rect 302516 139392 302568 139398
rect 302516 139334 302568 139340
rect 302330 118008 302386 118017
rect 302330 117943 302386 117952
rect 302240 60104 302292 60110
rect 302240 60046 302292 60052
rect 303632 16574 303660 211783
rect 303724 122126 303752 309703
rect 305000 303680 305052 303686
rect 305000 303622 305052 303628
rect 303804 244928 303856 244934
rect 303804 244870 303856 244876
rect 303816 244322 303844 244870
rect 303804 244316 303856 244322
rect 303804 244258 303856 244264
rect 303816 161430 303844 244258
rect 303896 191140 303948 191146
rect 303896 191082 303948 191088
rect 303804 161424 303856 161430
rect 303804 161366 303856 161372
rect 303908 136610 303936 191082
rect 303896 136604 303948 136610
rect 303896 136546 303948 136552
rect 303712 122120 303764 122126
rect 303712 122062 303764 122068
rect 305012 119406 305040 303622
rect 305092 191208 305144 191214
rect 305092 191150 305144 191156
rect 305104 128246 305132 191150
rect 305092 128240 305144 128246
rect 305092 128182 305144 128188
rect 305000 119400 305052 119406
rect 305000 119342 305052 119348
rect 305656 93158 305684 353942
rect 305734 349072 305790 349081
rect 305734 349007 305790 349016
rect 305748 323610 305776 349007
rect 307036 342145 307064 375255
rect 308416 374066 308444 377590
rect 309152 377590 309534 377618
rect 310532 377590 311190 377618
rect 308404 374060 308456 374066
rect 308404 374002 308456 374008
rect 308416 364993 308444 374002
rect 308402 364984 308458 364993
rect 308402 364919 308458 364928
rect 309152 349858 309180 377590
rect 309876 374672 309928 374678
rect 309876 374614 309928 374620
rect 309140 349852 309192 349858
rect 309140 349794 309192 349800
rect 307022 342136 307078 342145
rect 307022 342071 307078 342080
rect 309784 340264 309836 340270
rect 309784 340206 309836 340212
rect 306380 330540 306432 330546
rect 306380 330482 306432 330488
rect 305736 323604 305788 323610
rect 305736 323546 305788 323552
rect 305734 206272 305790 206281
rect 305734 206207 305790 206216
rect 305644 93152 305696 93158
rect 305644 93094 305696 93100
rect 303632 16546 303936 16574
rect 302882 14512 302938 14521
rect 302882 14447 302938 14456
rect 300124 13796 300176 13802
rect 300124 13738 300176 13744
rect 300136 12510 300164 13738
rect 299664 12504 299716 12510
rect 299664 12446 299716 12452
rect 300124 12504 300176 12510
rect 300124 12446 300176 12452
rect 298466 4856 298522 4865
rect 298466 4791 298522 4800
rect 298100 4140 298152 4146
rect 298100 4082 298152 4088
rect 298480 480 298508 4791
rect 299676 480 299704 12446
rect 302896 6866 302924 14447
rect 302884 6860 302936 6866
rect 302884 6802 302936 6808
rect 301964 6180 302016 6186
rect 301964 6122 302016 6128
rect 300766 3496 300822 3505
rect 300766 3431 300822 3440
rect 300780 480 300808 3431
rect 301976 480 302004 6122
rect 302896 4570 302924 6802
rect 302896 4542 303200 4570
rect 303172 480 303200 4542
rect 303908 490 303936 16546
rect 305748 5574 305776 206207
rect 305736 5568 305788 5574
rect 305736 5510 305788 5516
rect 305552 3800 305604 3806
rect 305552 3742 305604 3748
rect 304184 598 304396 626
rect 304184 490 304212 598
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 303908 462 304212 490
rect 304368 480 304396 598
rect 305564 480 305592 3742
rect 306392 490 306420 330482
rect 307668 257372 307720 257378
rect 307668 257314 307720 257320
rect 307680 256766 307708 257314
rect 306564 256760 306616 256766
rect 306564 256702 306616 256708
rect 307668 256760 307720 256766
rect 307668 256702 307720 256708
rect 306472 229764 306524 229770
rect 306472 229706 306524 229712
rect 306484 3806 306512 229706
rect 306576 126274 306604 256702
rect 309048 250504 309100 250510
rect 309048 250446 309100 250452
rect 309060 249830 309088 250446
rect 307852 249824 307904 249830
rect 307852 249766 307904 249772
rect 309048 249824 309100 249830
rect 309048 249766 309100 249772
rect 307864 238754 307892 249766
rect 307772 238726 307892 238754
rect 306656 198008 306708 198014
rect 306656 197950 306708 197956
rect 306668 147626 306696 197950
rect 306656 147620 306708 147626
rect 306656 147562 306708 147568
rect 307772 131102 307800 238726
rect 309140 224256 309192 224262
rect 309140 224198 309192 224204
rect 307852 208412 307904 208418
rect 307852 208354 307904 208360
rect 307760 131096 307812 131102
rect 307760 131038 307812 131044
rect 307864 131034 307892 208354
rect 307852 131028 307904 131034
rect 307852 130970 307904 130976
rect 306564 126268 306616 126274
rect 306564 126210 306616 126216
rect 309152 108934 309180 224198
rect 309140 108928 309192 108934
rect 309140 108870 309192 108876
rect 307758 66872 307814 66881
rect 307758 66807 307814 66816
rect 307772 66230 307800 66807
rect 307760 66224 307812 66230
rect 307760 66166 307812 66172
rect 306472 3800 306524 3806
rect 306472 3742 306524 3748
rect 307772 3534 307800 66166
rect 309796 15978 309824 340206
rect 309888 237153 309916 374614
rect 309874 237144 309930 237153
rect 309874 237079 309930 237088
rect 309874 220144 309930 220153
rect 309874 220079 309930 220088
rect 309784 15972 309836 15978
rect 309784 15914 309836 15920
rect 307944 5568 307996 5574
rect 307944 5510 307996 5516
rect 307760 3528 307812 3534
rect 307760 3470 307812 3476
rect 306576 598 306788 626
rect 306576 490 306604 598
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306392 462 306604 490
rect 306760 480 306788 598
rect 307956 480 307984 5510
rect 309048 3528 309100 3534
rect 309048 3470 309100 3476
rect 309060 480 309088 3470
rect 309888 2990 309916 220079
rect 310532 97306 310560 377590
rect 312832 375329 312860 377604
rect 313292 377590 314502 377618
rect 316052 377590 316158 377618
rect 317524 377590 317998 377618
rect 312818 375320 312874 375329
rect 312818 375255 312874 375264
rect 311898 369064 311954 369073
rect 311898 368999 311954 369008
rect 311912 368529 311940 368999
rect 311898 368520 311954 368529
rect 311898 368455 311954 368464
rect 310612 256012 310664 256018
rect 310612 255954 310664 255960
rect 310624 100026 310652 255954
rect 310612 100020 310664 100026
rect 310612 99962 310664 99968
rect 310520 97300 310572 97306
rect 310520 97242 310572 97248
rect 310520 29640 310572 29646
rect 310520 29582 310572 29588
rect 310532 16574 310560 29582
rect 311912 16574 311940 368455
rect 313292 355337 313320 377590
rect 313924 374060 313976 374066
rect 313924 374002 313976 374008
rect 313278 355328 313334 355337
rect 313278 355263 313334 355272
rect 313372 290488 313424 290494
rect 313372 290430 313424 290436
rect 313384 289882 313412 290430
rect 313372 289876 313424 289882
rect 313372 289818 313424 289824
rect 311992 239420 312044 239426
rect 311992 239362 312044 239368
rect 312004 238814 312032 239362
rect 311992 238808 312044 238814
rect 311992 238750 312044 238756
rect 312004 133890 312032 238750
rect 313278 202192 313334 202201
rect 313278 202127 313334 202136
rect 311992 133884 312044 133890
rect 311992 133826 312044 133832
rect 313292 16574 313320 202127
rect 313384 140758 313412 289818
rect 313372 140752 313424 140758
rect 313372 140694 313424 140700
rect 310532 16546 311480 16574
rect 311912 16546 312216 16574
rect 313292 16546 313872 16574
rect 310244 4072 310296 4078
rect 310244 4014 310296 4020
rect 309876 2984 309928 2990
rect 309876 2926 309928 2932
rect 310256 480 310284 4014
rect 311452 480 311480 16546
rect 312188 490 312216 16546
rect 312464 598 312676 626
rect 312464 490 312492 598
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312188 462 312492 490
rect 312648 480 312676 598
rect 313844 480 313872 16546
rect 313936 15910 313964 374002
rect 314660 260160 314712 260166
rect 314660 260102 314712 260108
rect 314672 259486 314700 260102
rect 314660 259480 314712 259486
rect 314660 259422 314712 259428
rect 314672 123486 314700 259422
rect 316052 227050 316080 377590
rect 317420 329112 317472 329118
rect 317420 329054 317472 329060
rect 317328 309800 317380 309806
rect 317328 309742 317380 309748
rect 317340 309194 317368 309742
rect 316132 309188 316184 309194
rect 316132 309130 316184 309136
rect 317328 309188 317380 309194
rect 317328 309130 317380 309136
rect 316040 227044 316092 227050
rect 316040 226986 316092 226992
rect 314752 188352 314804 188358
rect 314752 188294 314804 188300
rect 314764 128314 314792 188294
rect 316038 184240 316094 184249
rect 316038 184175 316094 184184
rect 314752 128308 314804 128314
rect 314752 128250 314804 128256
rect 314660 123480 314712 123486
rect 314660 123422 314712 123428
rect 316052 16574 316080 184175
rect 316144 132462 316172 309130
rect 316774 302288 316830 302297
rect 316774 302223 316830 302232
rect 316682 191040 316738 191049
rect 316682 190975 316738 190984
rect 316132 132456 316184 132462
rect 316132 132398 316184 132404
rect 316052 16546 316264 16574
rect 313924 15904 313976 15910
rect 313924 15846 313976 15852
rect 315028 2984 315080 2990
rect 315028 2926 315080 2932
rect 315040 480 315068 2926
rect 316236 480 316264 16546
rect 316696 4146 316724 190975
rect 316788 184210 316816 302223
rect 316776 184204 316828 184210
rect 316776 184146 316828 184152
rect 316684 4140 316736 4146
rect 316684 4082 316736 4088
rect 317432 4078 317460 329054
rect 317524 237289 317552 377590
rect 319640 376961 319668 377604
rect 318798 376952 318854 376961
rect 318798 376887 318854 376896
rect 319626 376952 319682 376961
rect 319626 376887 319682 376896
rect 318812 352617 318840 376887
rect 321296 375358 321324 377604
rect 320180 375352 320232 375358
rect 320180 375294 320232 375300
rect 321284 375352 321336 375358
rect 321284 375294 321336 375300
rect 320192 361729 320220 375294
rect 322296 362296 322348 362302
rect 322296 362238 322348 362244
rect 320178 361720 320234 361729
rect 320178 361655 320234 361664
rect 318798 352608 318854 352617
rect 318798 352543 318854 352552
rect 318800 276684 318852 276690
rect 318800 276626 318852 276632
rect 317510 237280 317566 237289
rect 317510 237215 317566 237224
rect 317510 199472 317566 199481
rect 317510 199407 317566 199416
rect 317524 113150 317552 199407
rect 318812 160070 318840 276626
rect 318800 160064 318852 160070
rect 318800 160006 318852 160012
rect 317512 113144 317564 113150
rect 317512 113086 317564 113092
rect 317510 75168 317566 75177
rect 317510 75103 317566 75112
rect 317524 16574 317552 75103
rect 319444 19984 319496 19990
rect 319444 19926 319496 19932
rect 319456 16574 319484 19926
rect 320192 16574 320220 361655
rect 321560 315308 321612 315314
rect 321560 315250 321612 315256
rect 321572 314702 321600 315250
rect 321560 314696 321612 314702
rect 321560 314638 321612 314644
rect 320640 246356 320692 246362
rect 320640 246298 320692 246304
rect 320652 245682 320680 246298
rect 320272 245676 320324 245682
rect 320272 245618 320324 245624
rect 320640 245676 320692 245682
rect 320640 245618 320692 245624
rect 320284 125594 320312 245618
rect 321572 155922 321600 314638
rect 322202 308408 322258 308417
rect 322202 308343 322258 308352
rect 321560 155916 321612 155922
rect 321560 155858 321612 155864
rect 320272 125588 320324 125594
rect 320272 125530 320324 125536
rect 322216 25566 322244 308343
rect 322308 307086 322336 362238
rect 322296 307080 322348 307086
rect 322296 307022 322348 307028
rect 322952 224262 322980 377604
rect 324332 377590 324622 377618
rect 325712 377590 326278 377618
rect 324332 356833 324360 377590
rect 325712 368665 325740 377590
rect 327724 374876 327776 374882
rect 327724 374818 327776 374824
rect 325698 368656 325754 368665
rect 325698 368591 325754 368600
rect 326342 368656 326398 368665
rect 326342 368591 326398 368600
rect 325608 363656 325660 363662
rect 325608 363598 325660 363604
rect 325620 362982 325648 363598
rect 325608 362976 325660 362982
rect 325608 362918 325660 362924
rect 324318 356824 324374 356833
rect 324318 356759 324374 356768
rect 323584 261520 323636 261526
rect 323584 261462 323636 261468
rect 322940 224256 322992 224262
rect 322940 224198 322992 224204
rect 322938 193896 322994 193905
rect 322938 193831 322994 193840
rect 322204 25560 322256 25566
rect 322204 25502 322256 25508
rect 317524 16546 318104 16574
rect 319456 16546 319760 16574
rect 320192 16546 320496 16574
rect 317420 4072 317472 4078
rect 317420 4014 317472 4020
rect 317326 3360 317382 3369
rect 317326 3295 317382 3304
rect 317340 480 317368 3295
rect 318076 490 318104 16546
rect 319732 4146 319760 16546
rect 319720 4140 319772 4146
rect 319720 4082 319772 4088
rect 318352 598 318564 626
rect 318352 490 318380 598
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318076 462 318380 490
rect 318536 480 318564 598
rect 319732 480 319760 4082
rect 320468 490 320496 16546
rect 322112 15972 322164 15978
rect 322112 15914 322164 15920
rect 320744 598 320956 626
rect 320744 490 320772 598
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320468 462 320772 490
rect 320928 480 320956 598
rect 322124 480 322152 15914
rect 322952 490 322980 193831
rect 323596 3466 323624 261462
rect 324318 188320 324374 188329
rect 324318 188255 324374 188264
rect 324332 3534 324360 188255
rect 324412 24132 324464 24138
rect 324412 24074 324464 24080
rect 324320 3528 324372 3534
rect 324320 3470 324372 3476
rect 323584 3460 323636 3466
rect 323584 3402 323636 3408
rect 323136 598 323348 626
rect 323136 490 323164 598
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 322952 462 323164 490
rect 323320 480 323348 598
rect 324424 480 324452 24074
rect 325620 6186 325648 362918
rect 326356 247722 326384 368591
rect 327078 353424 327134 353433
rect 327078 353359 327134 353368
rect 326344 247716 326396 247722
rect 326344 247658 326396 247664
rect 326344 184204 326396 184210
rect 326344 184146 326396 184152
rect 326356 6905 326384 184146
rect 327092 16574 327120 353359
rect 327736 282198 327764 374818
rect 327920 374678 327948 377604
rect 328472 377590 329590 377618
rect 327908 374672 327960 374678
rect 327908 374614 327960 374620
rect 328472 363089 328500 377590
rect 331232 374882 331260 377604
rect 332612 377590 332902 377618
rect 334084 377590 334558 377618
rect 335372 377590 336214 377618
rect 336752 377590 337870 377618
rect 331220 374876 331272 374882
rect 331220 374818 331272 374824
rect 331956 366444 332008 366450
rect 331956 366386 332008 366392
rect 328458 363080 328514 363089
rect 328458 363015 328514 363024
rect 329102 363080 329158 363089
rect 329102 363015 329158 363024
rect 329116 302938 329144 363015
rect 331862 325000 331918 325009
rect 331862 324935 331918 324944
rect 329104 302932 329156 302938
rect 329104 302874 329156 302880
rect 327724 282192 327776 282198
rect 327724 282134 327776 282140
rect 329748 247784 329800 247790
rect 329748 247726 329800 247732
rect 329760 247110 329788 247726
rect 328460 247104 328512 247110
rect 328460 247046 328512 247052
rect 329748 247104 329800 247110
rect 329748 247046 329800 247052
rect 328472 109002 328500 247046
rect 328460 108996 328512 109002
rect 328460 108938 328512 108944
rect 328460 25560 328512 25566
rect 328460 25502 328512 25508
rect 328472 16574 328500 25502
rect 327092 16546 328040 16574
rect 328472 16546 328776 16574
rect 326342 6896 326398 6905
rect 326342 6831 326398 6840
rect 326802 6896 326858 6905
rect 326802 6831 326858 6840
rect 325608 6180 325660 6186
rect 325608 6122 325660 6128
rect 325608 3528 325660 3534
rect 325608 3470 325660 3476
rect 325620 480 325648 3470
rect 326816 480 326844 6831
rect 328012 480 328040 16546
rect 328748 490 328776 16546
rect 331220 14476 331272 14482
rect 331220 14418 331272 14424
rect 330390 3360 330446 3369
rect 330390 3295 330446 3304
rect 329024 598 329236 626
rect 329024 490 329052 598
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 328748 462 329052 490
rect 329208 480 329236 598
rect 330404 480 330432 3295
rect 331232 490 331260 14418
rect 331876 2106 331904 324935
rect 331968 320890 331996 366386
rect 331956 320884 332008 320890
rect 331956 320826 332008 320832
rect 332612 311137 332640 377590
rect 333978 345128 334034 345137
rect 333978 345063 334034 345072
rect 332598 311128 332654 311137
rect 332598 311063 332654 311072
rect 332598 185600 332654 185609
rect 332598 185535 332654 185544
rect 331864 2100 331916 2106
rect 331864 2042 331916 2048
rect 331416 598 331628 626
rect 332612 610 332640 185535
rect 333992 16574 334020 345063
rect 334084 239426 334112 377590
rect 334624 372632 334676 372638
rect 334624 372574 334676 372580
rect 334072 239420 334124 239426
rect 334072 239362 334124 239368
rect 334636 176662 334664 372574
rect 335372 338774 335400 377590
rect 336752 372638 336780 377590
rect 339512 375358 339540 377604
rect 340892 377590 341182 377618
rect 342272 377590 342838 377618
rect 340234 376000 340290 376009
rect 340234 375935 340290 375944
rect 339500 375352 339552 375358
rect 339500 375294 339552 375300
rect 340144 373312 340196 373318
rect 340144 373254 340196 373260
rect 336740 372632 336792 372638
rect 336740 372574 336792 372580
rect 338948 365084 339000 365090
rect 338948 365026 339000 365032
rect 338762 362264 338818 362273
rect 338762 362199 338818 362208
rect 338856 362228 338908 362234
rect 337384 340196 337436 340202
rect 337384 340138 337436 340144
rect 335360 338768 335412 338774
rect 335360 338710 335412 338716
rect 336004 323604 336056 323610
rect 336004 323546 336056 323552
rect 335358 209808 335414 209817
rect 335358 209743 335414 209752
rect 334624 176656 334676 176662
rect 334624 176598 334676 176604
rect 335372 16574 335400 209743
rect 333992 16546 334664 16574
rect 335372 16546 335952 16574
rect 332692 6180 332744 6186
rect 332692 6122 332744 6128
rect 331416 490 331444 598
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331232 462 331444 490
rect 331600 480 331628 598
rect 332600 604 332652 610
rect 332600 546 332652 552
rect 332704 480 332732 6122
rect 333888 604 333940 610
rect 333888 546 333940 552
rect 333900 480 333928 546
rect 334636 490 334664 16546
rect 335924 3346 335952 16546
rect 336016 3534 336044 323546
rect 336004 3528 336056 3534
rect 336004 3470 336056 3476
rect 335924 3318 336320 3346
rect 334912 598 335124 626
rect 334912 490 334940 598
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 334636 462 334940 490
rect 335096 480 335124 598
rect 336292 480 336320 3318
rect 337396 3194 337424 340138
rect 338776 66230 338804 362199
rect 338856 362170 338908 362176
rect 338868 185609 338896 362170
rect 338960 309806 338988 365026
rect 338948 309800 339000 309806
rect 338948 309742 339000 309748
rect 340156 250510 340184 373254
rect 340248 301510 340276 375935
rect 340892 354006 340920 377590
rect 341524 371884 341576 371890
rect 341524 371826 341576 371832
rect 340880 354000 340932 354006
rect 340880 353942 340932 353948
rect 340236 301504 340288 301510
rect 340236 301446 340288 301452
rect 341536 253230 341564 371826
rect 341524 253224 341576 253230
rect 341524 253166 341576 253172
rect 340144 250504 340196 250510
rect 340144 250446 340196 250452
rect 342272 244934 342300 377590
rect 344480 375358 344508 377604
rect 342352 375352 342404 375358
rect 342352 375294 342404 375300
rect 344468 375352 344520 375358
rect 346136 375329 346164 377604
rect 344468 375294 344520 375300
rect 346122 375320 346178 375329
rect 342364 374649 342392 375294
rect 342350 374640 342406 374649
rect 342350 374575 342406 374584
rect 342260 244928 342312 244934
rect 342260 244870 342312 244876
rect 342364 235929 342392 374575
rect 344480 373994 344508 375294
rect 346122 375255 346178 375264
rect 344296 373966 344508 373994
rect 344296 322250 344324 373966
rect 345664 369232 345716 369238
rect 345664 369174 345716 369180
rect 344284 322244 344336 322250
rect 344284 322186 344336 322192
rect 345676 318102 345704 369174
rect 347044 369164 347096 369170
rect 347044 369106 347096 369112
rect 347056 349761 347084 369106
rect 347792 362302 347820 377604
rect 349264 377590 349462 377618
rect 349158 375320 349214 375329
rect 348424 375284 348476 375290
rect 349158 375255 349214 375264
rect 348424 375226 348476 375232
rect 347780 362296 347832 362302
rect 347780 362238 347832 362244
rect 347042 349752 347098 349761
rect 347042 349687 347098 349696
rect 348436 326398 348464 375226
rect 348424 326392 348476 326398
rect 348424 326334 348476 326340
rect 345664 318096 345716 318102
rect 345664 318038 345716 318044
rect 345018 312488 345074 312497
rect 345018 312423 345074 312432
rect 342350 235920 342406 235929
rect 342350 235855 342406 235864
rect 340970 208992 341026 209001
rect 340970 208927 341026 208936
rect 338854 185600 338910 185609
rect 338854 185535 338910 185544
rect 338764 66224 338816 66230
rect 338764 66166 338816 66172
rect 338762 18592 338818 18601
rect 338762 18527 338818 18536
rect 338776 6914 338804 18527
rect 340984 11830 341012 208927
rect 342902 206408 342958 206417
rect 342902 206343 342958 206352
rect 342258 72448 342314 72457
rect 342258 72383 342314 72392
rect 340972 11824 341024 11830
rect 340972 11766 341024 11772
rect 342168 11824 342220 11830
rect 342168 11766 342220 11772
rect 338684 6886 338804 6914
rect 338684 5506 338712 6886
rect 338672 5500 338724 5506
rect 338672 5442 338724 5448
rect 337476 3528 337528 3534
rect 337476 3470 337528 3476
rect 337384 3188 337436 3194
rect 337384 3130 337436 3136
rect 337488 480 337516 3470
rect 338684 480 338712 5442
rect 339868 3188 339920 3194
rect 339868 3130 339920 3136
rect 339880 480 339908 3130
rect 340972 2100 341024 2106
rect 340972 2042 341024 2048
rect 340984 480 341012 2042
rect 342180 480 342208 11766
rect 342272 6914 342300 72383
rect 342916 16574 342944 206343
rect 342916 16546 343036 16574
rect 342272 6886 342944 6914
rect 342916 490 342944 6886
rect 343008 4049 343036 16546
rect 342994 4040 343050 4049
rect 342994 3975 343050 3984
rect 345032 2802 345060 312423
rect 345296 15904 345348 15910
rect 345296 15846 345348 15852
rect 344940 2774 345060 2802
rect 343192 598 343404 626
rect 343192 490 343220 598
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 342916 462 343220 490
rect 343376 480 343404 598
rect 344572 598 344784 626
rect 344572 480 344600 598
rect 344756 490 344784 598
rect 344940 490 344968 2774
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 344756 462 344968 490
rect 345308 490 345336 15846
rect 349172 13802 349200 375255
rect 349264 366382 349292 377590
rect 351104 374785 351132 377604
rect 352656 376100 352708 376106
rect 352656 376042 352708 376048
rect 352562 375320 352618 375329
rect 352562 375255 352618 375264
rect 351090 374776 351146 374785
rect 351090 374711 351146 374720
rect 349252 366376 349304 366382
rect 349252 366318 349304 366324
rect 349804 366376 349856 366382
rect 349804 366318 349856 366324
rect 349816 333266 349844 366318
rect 349804 333260 349856 333266
rect 349804 333202 349856 333208
rect 352576 242214 352604 375255
rect 352668 316742 352696 376042
rect 352760 375290 352788 377604
rect 353312 377590 354430 377618
rect 355324 377596 355376 377602
rect 352748 375284 352800 375290
rect 352748 375226 352800 375232
rect 353312 361593 353340 377590
rect 355324 377538 355376 377544
rect 354126 377496 354182 377505
rect 354126 377431 354182 377440
rect 353944 376032 353996 376038
rect 353944 375974 353996 375980
rect 353298 361584 353354 361593
rect 353298 361519 353354 361528
rect 352656 316736 352708 316742
rect 352656 316678 352708 316684
rect 353300 247716 353352 247722
rect 353300 247658 353352 247664
rect 352564 242208 352616 242214
rect 352564 242150 352616 242156
rect 351918 195256 351974 195265
rect 351918 195191 351974 195200
rect 349160 13796 349212 13802
rect 349160 13738 349212 13744
rect 346950 4040 347006 4049
rect 346950 3975 347006 3984
rect 345584 598 345796 626
rect 345584 490 345612 598
rect 345308 462 345612 490
rect 345768 480 345796 598
rect 346964 480 346992 3975
rect 349252 3528 349304 3534
rect 351932 3482 351960 195191
rect 349252 3470 349304 3476
rect 348056 3460 348108 3466
rect 348056 3402 348108 3408
rect 348068 480 348096 3402
rect 349264 480 349292 3470
rect 350448 3460 350500 3466
rect 350448 3402 350500 3408
rect 351656 3454 351960 3482
rect 350460 480 350488 3402
rect 351656 480 351684 3454
rect 353312 3369 353340 247658
rect 353956 246362 353984 375974
rect 354036 374060 354088 374066
rect 354036 374002 354088 374008
rect 354048 247790 354076 374002
rect 354140 367713 354168 377431
rect 354678 376408 354734 376417
rect 354678 376343 354734 376352
rect 354692 373289 354720 376343
rect 354678 373280 354734 373289
rect 354678 373215 354734 373224
rect 354126 367704 354182 367713
rect 354126 367639 354182 367648
rect 355336 319462 355364 377538
rect 356072 374066 356100 377604
rect 356060 374060 356112 374066
rect 356060 374002 356112 374008
rect 355416 373380 355468 373386
rect 355416 373322 355468 373328
rect 355428 330614 355456 373322
rect 356164 358086 356192 492646
rect 356242 492623 356298 492632
rect 356532 490090 356560 497406
rect 356624 490385 356652 499546
rect 358728 499530 358780 499536
rect 358082 497856 358138 497865
rect 358082 497791 358138 497800
rect 357164 496800 357216 496806
rect 357164 496742 357216 496748
rect 357176 495553 357204 496742
rect 357162 495544 357218 495553
rect 357162 495479 357218 495488
rect 356610 490376 356666 490385
rect 356610 490311 356666 490320
rect 356256 490062 356560 490090
rect 356256 377602 356284 490062
rect 357438 482896 357494 482905
rect 357438 482831 357494 482840
rect 356794 465760 356850 465769
rect 356794 465695 356850 465704
rect 356808 465118 356836 465695
rect 356336 465112 356388 465118
rect 356336 465054 356388 465060
rect 356796 465112 356848 465118
rect 356796 465054 356848 465060
rect 356244 377596 356296 377602
rect 356244 377538 356296 377544
rect 356348 365022 356376 465054
rect 356704 426828 356756 426834
rect 356704 426770 356756 426776
rect 356336 365016 356388 365022
rect 356336 364958 356388 364964
rect 356152 358080 356204 358086
rect 356152 358022 356204 358028
rect 355416 330608 355468 330614
rect 355416 330550 355468 330556
rect 355324 319456 355376 319462
rect 355324 319398 355376 319404
rect 356716 258738 356744 426770
rect 357452 315314 357480 482831
rect 358096 465050 358124 497791
rect 358636 494012 358688 494018
rect 358636 493954 358688 493960
rect 358648 493105 358676 493954
rect 358634 493096 358690 493105
rect 358634 493031 358690 493040
rect 358726 487792 358782 487801
rect 358726 487727 358782 487736
rect 358740 487218 358768 487727
rect 358728 487212 358780 487218
rect 358728 487154 358780 487160
rect 358726 485344 358782 485353
rect 358726 485279 358782 485288
rect 358740 484430 358768 485279
rect 358728 484424 358780 484430
rect 358728 484366 358780 484372
rect 358726 478000 358782 478009
rect 358726 477935 358782 477944
rect 358740 477562 358768 477935
rect 358728 477556 358780 477562
rect 358728 477498 358780 477504
rect 358726 475552 358782 475561
rect 358726 475487 358782 475496
rect 358740 474774 358768 475487
rect 358728 474768 358780 474774
rect 358728 474710 358780 474716
rect 358726 473104 358782 473113
rect 358726 473039 358782 473048
rect 358740 472054 358768 473039
rect 358728 472048 358780 472054
rect 358728 471990 358780 471996
rect 358726 470656 358782 470665
rect 358726 470591 358728 470600
rect 358780 470591 358782 470600
rect 358728 470562 358780 470568
rect 358726 468208 358782 468217
rect 358726 468143 358782 468152
rect 358740 467906 358768 468143
rect 358728 467900 358780 467906
rect 358728 467842 358780 467848
rect 358084 465044 358136 465050
rect 358084 464986 358136 464992
rect 358726 463312 358782 463321
rect 358726 463247 358782 463256
rect 358740 462398 358768 463247
rect 358728 462392 358780 462398
rect 358728 462334 358780 462340
rect 358450 460864 358506 460873
rect 358450 460799 358506 460808
rect 358464 459610 358492 460799
rect 358452 459604 358504 459610
rect 358452 459546 358504 459552
rect 358726 455968 358782 455977
rect 358726 455903 358782 455912
rect 358740 455462 358768 455903
rect 358728 455456 358780 455462
rect 358728 455398 358780 455404
rect 358726 453520 358782 453529
rect 358726 453455 358782 453464
rect 358740 452674 358768 453455
rect 358728 452668 358780 452674
rect 358728 452610 358780 452616
rect 358726 451072 358782 451081
rect 358726 451007 358782 451016
rect 358740 449954 358768 451007
rect 358728 449948 358780 449954
rect 358728 449890 358780 449896
rect 358726 448624 358782 448633
rect 358726 448559 358728 448568
rect 358780 448559 358782 448568
rect 358728 448530 358780 448536
rect 357530 446176 357586 446185
rect 357530 446111 357586 446120
rect 357544 426834 357572 446111
rect 358726 443728 358782 443737
rect 358726 443663 358782 443672
rect 358740 443018 358768 443663
rect 358728 443012 358780 443018
rect 358728 442954 358780 442960
rect 358726 441280 358782 441289
rect 358726 441215 358782 441224
rect 358740 440298 358768 441215
rect 358728 440292 358780 440298
rect 358728 440234 358780 440240
rect 358726 438968 358782 438977
rect 358726 438903 358728 438912
rect 358780 438903 358782 438912
rect 358728 438874 358780 438880
rect 358726 436384 358782 436393
rect 358726 436319 358782 436328
rect 358740 436150 358768 436319
rect 358728 436144 358780 436150
rect 358728 436086 358780 436092
rect 358726 433936 358782 433945
rect 358726 433871 358782 433880
rect 358740 433362 358768 433871
rect 358728 433356 358780 433362
rect 358728 433298 358780 433304
rect 358726 431488 358782 431497
rect 358726 431423 358782 431432
rect 358740 430642 358768 431423
rect 358728 430636 358780 430642
rect 358728 430578 358780 430584
rect 358726 429040 358782 429049
rect 358726 428975 358782 428984
rect 358740 427854 358768 428975
rect 358728 427848 358780 427854
rect 358728 427790 358780 427796
rect 357532 426828 357584 426834
rect 357532 426770 357584 426776
rect 357530 426592 357586 426601
rect 357530 426527 357586 426536
rect 357544 371890 357572 426527
rect 358726 424144 358782 424153
rect 358726 424079 358782 424088
rect 358740 423706 358768 424079
rect 358728 423700 358780 423706
rect 358728 423642 358780 423648
rect 358726 421696 358782 421705
rect 358726 421631 358782 421640
rect 358740 420986 358768 421631
rect 358728 420980 358780 420986
rect 358728 420922 358780 420928
rect 358726 419248 358782 419257
rect 358726 419183 358782 419192
rect 358740 418266 358768 419183
rect 358728 418260 358780 418266
rect 358728 418202 358780 418208
rect 357622 416800 357678 416809
rect 357622 416735 357678 416744
rect 357636 373318 357664 416735
rect 358726 414352 358782 414361
rect 358726 414287 358782 414296
rect 358740 414050 358768 414287
rect 358728 414044 358780 414050
rect 358728 413986 358780 413992
rect 358726 411904 358782 411913
rect 358726 411839 358782 411848
rect 358740 411330 358768 411839
rect 358728 411324 358780 411330
rect 358728 411266 358780 411272
rect 358726 409456 358782 409465
rect 358726 409391 358782 409400
rect 358740 408610 358768 409391
rect 358728 408604 358780 408610
rect 358728 408546 358780 408552
rect 358726 404288 358782 404297
rect 358726 404223 358782 404232
rect 358740 403578 358768 404223
rect 358728 403572 358780 403578
rect 358728 403514 358780 403520
rect 358726 401840 358782 401849
rect 358726 401775 358782 401784
rect 358740 401674 358768 401775
rect 358728 401668 358780 401674
rect 358728 401610 358780 401616
rect 357990 399392 358046 399401
rect 357990 399327 358046 399336
rect 358004 398886 358032 399327
rect 357992 398880 358044 398886
rect 357992 398822 358044 398828
rect 358726 396944 358782 396953
rect 358726 396879 358782 396888
rect 358740 396098 358768 396879
rect 358728 396092 358780 396098
rect 358728 396034 358780 396040
rect 357714 392048 357770 392057
rect 357714 391983 357770 391992
rect 357624 373312 357676 373318
rect 357624 373254 357676 373260
rect 357532 371884 357584 371890
rect 357532 371826 357584 371832
rect 357728 370598 357756 391983
rect 358818 382392 358874 382401
rect 358818 382327 358874 382336
rect 357898 379808 357954 379817
rect 357898 379743 357954 379752
rect 357912 379574 357940 379743
rect 357900 379568 357952 379574
rect 357900 379510 357952 379516
rect 358360 378140 358412 378146
rect 358360 378082 358412 378088
rect 358372 378049 358400 378082
rect 358358 378040 358414 378049
rect 358358 377975 358414 377984
rect 358832 376106 358860 382327
rect 358820 376100 358872 376106
rect 358820 376042 358872 376048
rect 358818 374776 358874 374785
rect 358818 374711 358874 374720
rect 358084 371884 358136 371890
rect 358084 371826 358136 371832
rect 357716 370592 357768 370598
rect 357716 370534 357768 370540
rect 357440 315308 357492 315314
rect 357440 315250 357492 315256
rect 357440 302932 357492 302938
rect 357440 302874 357492 302880
rect 356704 258732 356756 258738
rect 356704 258674 356756 258680
rect 354036 247784 354088 247790
rect 354036 247726 354088 247732
rect 353944 246356 353996 246362
rect 353944 246298 353996 246304
rect 357452 3534 357480 302874
rect 358096 291854 358124 371826
rect 358084 291848 358136 291854
rect 358084 291790 358136 291796
rect 358832 11762 358860 374711
rect 358924 290494 358952 529615
rect 359002 407008 359058 407017
rect 359002 406943 359058 406952
rect 359016 377505 359044 406943
rect 359002 377496 359058 377505
rect 359002 377431 359058 377440
rect 359108 367810 359136 538290
rect 360212 520062 360240 700266
rect 363616 543017 363644 702578
rect 374644 700324 374696 700330
rect 374644 700266 374696 700272
rect 364432 543856 364484 543862
rect 364432 543798 364484 543804
rect 363602 543008 363658 543017
rect 363602 542943 363658 542952
rect 363052 542496 363104 542502
rect 363052 542438 363104 542444
rect 360292 541068 360344 541074
rect 360292 541010 360344 541016
rect 360200 520056 360252 520062
rect 360200 519998 360252 520004
rect 360200 514820 360252 514826
rect 360200 514762 360252 514768
rect 359096 367804 359148 367810
rect 359096 367746 359148 367752
rect 358912 290488 358964 290494
rect 358912 290430 358964 290436
rect 360212 117298 360240 514762
rect 360304 366450 360332 541010
rect 361578 538384 361634 538393
rect 361578 538319 361634 538328
rect 360382 535528 360438 535537
rect 360382 535463 360438 535472
rect 360396 378146 360424 535463
rect 360476 398880 360528 398886
rect 360476 398822 360528 398828
rect 360384 378140 360436 378146
rect 360384 378082 360436 378088
rect 360292 366444 360344 366450
rect 360292 366386 360344 366392
rect 360488 348537 360516 398822
rect 361488 378004 361540 378010
rect 361488 377946 361540 377952
rect 360474 348528 360530 348537
rect 360474 348463 360530 348472
rect 361500 238746 361528 377946
rect 361592 298790 361620 538319
rect 361672 535560 361724 535566
rect 361672 535502 361724 535508
rect 361684 369238 361712 535502
rect 362960 477556 363012 477562
rect 362960 477498 363012 477504
rect 361764 438932 361816 438938
rect 361764 438874 361816 438880
rect 361672 369232 361724 369238
rect 361672 369174 361724 369180
rect 361776 347041 361804 438874
rect 361856 396092 361908 396098
rect 361856 396034 361908 396040
rect 361868 373969 361896 396034
rect 361854 373960 361910 373969
rect 361854 373895 361910 373904
rect 361762 347032 361818 347041
rect 361762 346967 361818 346976
rect 361580 298784 361632 298790
rect 361580 298726 361632 298732
rect 362972 267034 363000 477498
rect 363064 365090 363092 542438
rect 363144 467900 363196 467906
rect 363144 467842 363196 467848
rect 363052 365084 363104 365090
rect 363052 365026 363104 365032
rect 363156 363662 363184 467842
rect 364340 449948 364392 449954
rect 364340 449890 364392 449896
rect 363236 403572 363288 403578
rect 363236 403514 363288 403520
rect 363248 376038 363276 403514
rect 363236 376032 363288 376038
rect 363236 375974 363288 375980
rect 363144 363656 363196 363662
rect 363144 363598 363196 363604
rect 362960 267028 363012 267034
rect 362960 266970 363012 266976
rect 364352 260166 364380 449890
rect 364444 373386 364472 543798
rect 364524 541000 364576 541006
rect 364524 540942 364576 540948
rect 364536 378010 364564 540942
rect 374090 539608 374146 539617
rect 374090 539543 374146 539552
rect 371238 538248 371294 538257
rect 371238 538183 371294 538192
rect 367100 527196 367152 527202
rect 367100 527138 367152 527144
rect 365720 465044 365772 465050
rect 365720 464986 365772 464992
rect 364616 423700 364668 423706
rect 364616 423642 364668 423648
rect 364524 378004 364576 378010
rect 364524 377946 364576 377952
rect 364432 373380 364484 373386
rect 364432 373322 364484 373328
rect 364628 345681 364656 423642
rect 364614 345672 364670 345681
rect 364614 345607 364670 345616
rect 365732 272542 365760 464986
rect 365812 418260 365864 418266
rect 365812 418202 365864 418208
rect 365824 369170 365852 418202
rect 365904 408604 365956 408610
rect 365904 408546 365956 408552
rect 365916 371890 365944 408546
rect 365904 371884 365956 371890
rect 365904 371826 365956 371832
rect 365812 369164 365864 369170
rect 365812 369106 365864 369112
rect 365720 272536 365772 272542
rect 365720 272478 365772 272484
rect 364340 260160 364392 260166
rect 364340 260102 364392 260108
rect 361488 238740 361540 238746
rect 361488 238682 361540 238688
rect 360290 182880 360346 182889
rect 360290 182815 360346 182824
rect 360200 117292 360252 117298
rect 360200 117234 360252 117240
rect 358820 11756 358872 11762
rect 358820 11698 358872 11704
rect 357440 3528 357492 3534
rect 357440 3470 357492 3476
rect 360304 3466 360332 182815
rect 367112 5506 367140 527138
rect 367192 505776 367244 505782
rect 367192 505718 367244 505724
rect 367204 276690 367232 505718
rect 369952 502376 370004 502382
rect 369952 502318 370004 502324
rect 369860 484424 369912 484430
rect 369860 484366 369912 484372
rect 368572 472048 368624 472054
rect 368572 471990 368624 471996
rect 368388 449200 368440 449206
rect 368388 449142 368440 449148
rect 368400 448594 368428 449142
rect 367284 448588 367336 448594
rect 367284 448530 367336 448536
rect 368388 448588 368440 448594
rect 368388 448530 368440 448536
rect 367296 361554 367324 448530
rect 368480 440292 368532 440298
rect 368480 440234 368532 440240
rect 367376 414044 367428 414050
rect 367376 413986 367428 413992
rect 367388 377369 367416 413986
rect 367374 377360 367430 377369
rect 367374 377295 367430 377304
rect 367284 361548 367336 361554
rect 367284 361490 367336 361496
rect 367192 276684 367244 276690
rect 367192 276626 367244 276632
rect 368492 113150 368520 440234
rect 368584 366382 368612 471990
rect 368572 366376 368624 366382
rect 368572 366318 368624 366324
rect 368480 113144 368532 113150
rect 368480 113086 368532 113092
rect 369872 6866 369900 484366
rect 369964 273970 369992 502318
rect 370044 460216 370096 460222
rect 370044 460158 370096 460164
rect 370056 459610 370084 460158
rect 370044 459604 370096 459610
rect 370044 459546 370096 459552
rect 370056 365673 370084 459546
rect 370136 420980 370188 420986
rect 370136 420922 370188 420928
rect 370148 369073 370176 420922
rect 370134 369064 370190 369073
rect 370134 368999 370190 369008
rect 370042 365664 370098 365673
rect 370042 365599 370098 365608
rect 369952 273964 370004 273970
rect 369952 273906 370004 273912
rect 371252 184249 371280 538183
rect 371332 536852 371384 536858
rect 371332 536794 371384 536800
rect 371344 337414 371372 536794
rect 371424 499588 371476 499594
rect 371424 499530 371476 499536
rect 371332 337408 371384 337414
rect 371332 337350 371384 337356
rect 371436 336025 371464 499530
rect 372620 487212 372672 487218
rect 372620 487154 372672 487160
rect 371422 336016 371478 336025
rect 371422 335951 371478 335960
rect 372632 271182 372660 487154
rect 372712 427848 372764 427854
rect 372712 427790 372764 427796
rect 372724 341562 372752 427790
rect 374000 423700 374052 423706
rect 374000 423642 374052 423648
rect 372712 341556 372764 341562
rect 372712 341498 372764 341504
rect 372620 271176 372672 271182
rect 372620 271118 372672 271124
rect 371238 184240 371294 184249
rect 371238 184175 371294 184184
rect 374012 14482 374040 423642
rect 374104 362234 374132 539543
rect 374656 376553 374684 700266
rect 375472 545148 375524 545154
rect 375472 545090 375524 545096
rect 375380 516180 375432 516186
rect 375380 516122 375432 516128
rect 374642 376544 374698 376553
rect 374642 376479 374698 376488
rect 374092 362228 374144 362234
rect 374092 362170 374144 362176
rect 374000 14476 374052 14482
rect 374000 14418 374052 14424
rect 375392 7614 375420 516122
rect 375484 207641 375512 545090
rect 378232 524476 378284 524482
rect 378232 524418 378284 524424
rect 375564 474768 375616 474774
rect 375564 474710 375616 474716
rect 375576 351121 375604 474710
rect 376760 452668 376812 452674
rect 376760 452610 376812 452616
rect 375562 351112 375618 351121
rect 375562 351047 375618 351056
rect 375470 207632 375526 207641
rect 375470 207567 375526 207576
rect 376772 9654 376800 452610
rect 376852 430636 376904 430642
rect 376852 430578 376904 430584
rect 376864 257378 376892 430578
rect 378140 401668 378192 401674
rect 378140 401610 378192 401616
rect 376852 257372 376904 257378
rect 376852 257314 376904 257320
rect 378152 19990 378180 401610
rect 378244 280838 378272 524418
rect 380900 470620 380952 470626
rect 380900 470562 380952 470568
rect 379520 436144 379572 436150
rect 379520 436086 379572 436092
rect 378232 280832 378284 280838
rect 378232 280774 378284 280780
rect 379532 256018 379560 436086
rect 379520 256012 379572 256018
rect 379520 255954 379572 255960
rect 380912 219337 380940 470562
rect 380992 433356 381044 433362
rect 380992 433298 381044 433304
rect 381004 313954 381032 433298
rect 382280 379568 382332 379574
rect 382280 379510 382332 379516
rect 380992 313948 381044 313954
rect 380992 313890 381044 313896
rect 381542 284472 381598 284481
rect 381542 284407 381598 284416
rect 381556 259418 381584 284407
rect 381544 259412 381596 259418
rect 381544 259354 381596 259360
rect 381544 244316 381596 244322
rect 381544 244258 381596 244264
rect 381556 238746 381584 244258
rect 381544 238740 381596 238746
rect 381544 238682 381596 238688
rect 380898 219328 380954 219337
rect 380898 219263 380954 219272
rect 382292 115938 382320 379510
rect 382936 374649 382964 702646
rect 385040 505164 385092 505170
rect 385040 505106 385092 505112
rect 383660 443012 383712 443018
rect 383660 442954 383712 442960
rect 382922 374640 382978 374649
rect 382922 374575 382978 374584
rect 383672 282878 383700 442954
rect 383660 282872 383712 282878
rect 383660 282814 383712 282820
rect 382280 115932 382332 115938
rect 382280 115874 382332 115880
rect 378140 19984 378192 19990
rect 378140 19926 378192 19932
rect 376760 9648 376812 9654
rect 376760 9590 376812 9596
rect 375380 7608 375432 7614
rect 375380 7550 375432 7556
rect 385052 6905 385080 505106
rect 412652 494018 412680 703582
rect 413480 703474 413508 703582
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 413664 703474 413692 703520
rect 413480 703446 413692 703474
rect 429856 700330 429884 703520
rect 462332 702710 462360 703520
rect 478524 702914 478552 703520
rect 478512 702908 478564 702914
rect 478512 702850 478564 702856
rect 494808 702846 494836 703520
rect 494796 702840 494848 702846
rect 494796 702782 494848 702788
rect 462320 702704 462372 702710
rect 462320 702646 462372 702652
rect 527192 702506 527220 703520
rect 543476 702642 543504 703520
rect 543464 702636 543516 702642
rect 543464 702578 543516 702584
rect 559668 702574 559696 703520
rect 559656 702568 559708 702574
rect 559656 702510 559708 702516
rect 527180 702500 527232 702506
rect 527180 702442 527232 702448
rect 429844 700324 429896 700330
rect 429844 700266 429896 700272
rect 582470 697232 582526 697241
rect 582470 697167 582526 697176
rect 582378 564360 582434 564369
rect 582378 564295 582434 564304
rect 582392 556850 582420 564295
rect 582380 556844 582432 556850
rect 582380 556786 582432 556792
rect 580264 539640 580316 539646
rect 580264 539582 580316 539588
rect 580170 537840 580226 537849
rect 580170 537775 580226 537784
rect 580184 537538 580212 537775
rect 580172 537532 580224 537538
rect 580172 537474 580224 537480
rect 412640 494012 412692 494018
rect 412640 493954 412692 493960
rect 580276 484673 580304 539582
rect 582380 535492 582432 535498
rect 582380 535434 582432 535440
rect 582392 524521 582420 535434
rect 582378 524512 582434 524521
rect 582378 524447 582434 524456
rect 582380 522300 582432 522306
rect 582380 522242 582432 522248
rect 582392 511329 582420 522242
rect 582378 511320 582434 511329
rect 582378 511255 582434 511264
rect 580262 484664 580318 484673
rect 580262 484599 580318 484608
rect 582380 465112 582432 465118
rect 582380 465054 582432 465060
rect 385132 462392 385184 462398
rect 385132 462334 385184 462340
rect 385144 263566 385172 462334
rect 387800 455456 387852 455462
rect 387800 455398 387852 455404
rect 387812 370530 387840 455398
rect 582392 418305 582420 465054
rect 582484 449206 582512 697167
rect 582562 683904 582618 683913
rect 582562 683839 582618 683848
rect 582576 460222 582604 683839
rect 583206 670712 583262 670721
rect 583206 670647 583262 670656
rect 582746 644056 582802 644065
rect 582746 643991 582802 644000
rect 582654 577688 582710 577697
rect 582654 577623 582710 577632
rect 582564 460216 582616 460222
rect 582564 460158 582616 460164
rect 582472 449200 582524 449206
rect 582472 449142 582524 449148
rect 582378 418296 582434 418305
rect 582378 418231 582434 418240
rect 389180 411324 389232 411330
rect 389180 411266 389232 411272
rect 387800 370524 387852 370530
rect 387800 370466 387852 370472
rect 389192 278730 389220 411266
rect 582378 378448 582434 378457
rect 582378 378383 582434 378392
rect 582392 375358 582420 378383
rect 582668 376961 582696 577623
rect 582760 551342 582788 643991
rect 583022 630864 583078 630873
rect 583022 630799 583078 630808
rect 582930 591016 582986 591025
rect 582930 590951 582986 590960
rect 582840 563100 582892 563106
rect 582840 563042 582892 563048
rect 582748 551336 582800 551342
rect 582748 551278 582800 551284
rect 582748 532024 582800 532030
rect 582748 531966 582800 531972
rect 582760 404977 582788 531966
rect 582852 458153 582880 563042
rect 582944 496806 582972 590951
rect 583036 554062 583064 630799
rect 583114 617536 583170 617545
rect 583114 617471 583170 617480
rect 583024 554056 583076 554062
rect 583024 553998 583076 554004
rect 583128 541657 583156 617471
rect 583114 541648 583170 541657
rect 583114 541583 583170 541592
rect 582932 496800 582984 496806
rect 582932 496742 582984 496748
rect 582930 471472 582986 471481
rect 582930 471407 582986 471416
rect 582838 458144 582894 458153
rect 582838 458079 582894 458088
rect 582840 455456 582892 455462
rect 582840 455398 582892 455404
rect 582852 431633 582880 455398
rect 582838 431624 582894 431633
rect 582838 431559 582894 431568
rect 582746 404968 582802 404977
rect 582746 404903 582802 404912
rect 582654 376952 582710 376961
rect 582654 376887 582710 376896
rect 582380 375352 582432 375358
rect 582380 375294 582432 375300
rect 582944 372570 582972 471407
rect 583220 376689 583248 670647
rect 583206 376680 583262 376689
rect 583206 376615 583262 376624
rect 582932 372564 582984 372570
rect 582932 372506 582984 372512
rect 582378 365120 582434 365129
rect 582378 365055 582434 365064
rect 580172 352572 580224 352578
rect 580172 352514 580224 352520
rect 580184 351937 580212 352514
rect 580170 351928 580226 351937
rect 580170 351863 580226 351872
rect 582392 342961 582420 365055
rect 582378 342952 582434 342961
rect 582378 342887 582434 342896
rect 582380 334620 582432 334626
rect 582380 334562 582432 334568
rect 580722 298752 580778 298761
rect 580722 298687 580778 298696
rect 580736 296721 580764 298687
rect 580722 296712 580778 296721
rect 580722 296647 580778 296656
rect 389180 278724 389232 278730
rect 389180 278666 389232 278672
rect 389192 278050 389220 278666
rect 389180 278044 389232 278050
rect 389180 277986 389232 277992
rect 579802 272232 579858 272241
rect 579802 272167 579858 272176
rect 579816 271930 579844 272167
rect 574744 271924 574796 271930
rect 574744 271866 574796 271872
rect 579804 271924 579856 271930
rect 579804 271866 579856 271872
rect 385132 263560 385184 263566
rect 385132 263502 385184 263508
rect 566464 251864 566516 251870
rect 566464 251806 566516 251812
rect 566476 167006 566504 251806
rect 574756 234569 574784 271866
rect 580262 261488 580318 261497
rect 580262 261423 580318 261432
rect 580172 259412 580224 259418
rect 580172 259354 580224 259360
rect 580184 258913 580212 259354
rect 580170 258904 580226 258913
rect 580170 258839 580226 258848
rect 580170 245576 580226 245585
rect 580170 245511 580226 245520
rect 580184 244322 580212 245511
rect 580172 244316 580224 244322
rect 580172 244258 580224 244264
rect 574742 234560 574798 234569
rect 574742 234495 574798 234504
rect 574742 228304 574798 228313
rect 574742 228239 574798 228248
rect 566464 167000 566516 167006
rect 566464 166942 566516 166948
rect 385038 6896 385094 6905
rect 369860 6860 369912 6866
rect 574756 6866 574784 228239
rect 580276 179217 580304 261423
rect 580262 179208 580318 179217
rect 580262 179143 580318 179152
rect 580172 167000 580224 167006
rect 580172 166942 580224 166948
rect 580184 165889 580212 166942
rect 580170 165880 580226 165889
rect 580170 165815 580226 165824
rect 582392 16574 582420 334562
rect 582930 325272 582986 325281
rect 582930 325207 582986 325216
rect 582472 299532 582524 299538
rect 582472 299474 582524 299480
rect 582484 19825 582512 299474
rect 582654 292632 582710 292641
rect 582654 292567 582710 292576
rect 582564 288448 582616 288454
rect 582564 288390 582616 288396
rect 582576 73001 582604 288390
rect 582668 192545 582696 292567
rect 582840 286340 582892 286346
rect 582840 286282 582892 286288
rect 582748 232552 582800 232558
rect 582748 232494 582800 232500
rect 582654 192536 582710 192545
rect 582654 192471 582710 192480
rect 582562 72992 582618 73001
rect 582562 72927 582618 72936
rect 582760 46345 582788 232494
rect 582852 112849 582880 286282
rect 582944 254590 582972 325207
rect 583022 312080 583078 312089
rect 583022 312015 583078 312024
rect 583036 269074 583064 312015
rect 583574 287736 583630 287745
rect 583574 287671 583630 287680
rect 583206 284336 583262 284345
rect 583206 284271 583262 284280
rect 583116 278792 583168 278798
rect 583116 278734 583168 278740
rect 583024 269068 583076 269074
rect 583024 269010 583076 269016
rect 583022 264208 583078 264217
rect 583022 264143 583078 264152
rect 582932 254584 582984 254590
rect 582932 254526 582984 254532
rect 582930 231160 582986 231169
rect 582930 231095 582986 231104
rect 582838 112840 582894 112849
rect 582838 112775 582894 112784
rect 582944 59673 582972 231095
rect 583036 99521 583064 264143
rect 583128 126041 583156 278734
rect 583220 219065 583248 284271
rect 583392 278044 583444 278050
rect 583392 277986 583444 277992
rect 583300 275324 583352 275330
rect 583300 275266 583352 275272
rect 583206 219056 583262 219065
rect 583206 218991 583262 219000
rect 583312 139369 583340 275266
rect 583404 152697 583432 277986
rect 583482 265568 583538 265577
rect 583482 265503 583538 265512
rect 583496 232937 583524 265503
rect 583482 232928 583538 232937
rect 583482 232863 583538 232872
rect 583482 213208 583538 213217
rect 583482 213143 583538 213152
rect 583390 152688 583446 152697
rect 583390 152623 583446 152632
rect 583298 139360 583354 139369
rect 583298 139295 583354 139304
rect 583114 126032 583170 126041
rect 583114 125967 583170 125976
rect 583022 99512 583078 99521
rect 583022 99447 583078 99456
rect 582930 59664 582986 59673
rect 582930 59599 582986 59608
rect 582746 46336 582802 46345
rect 582746 46271 582802 46280
rect 583390 33144 583446 33153
rect 583390 33079 583392 33088
rect 583444 33079 583446 33088
rect 583392 33050 583444 33056
rect 582470 19816 582526 19825
rect 582470 19751 582526 19760
rect 582392 16546 583432 16574
rect 385038 6831 385094 6840
rect 574744 6860 574796 6866
rect 369860 6802 369912 6808
rect 574744 6802 574796 6808
rect 580172 6860 580224 6866
rect 580172 6802 580224 6808
rect 580184 6633 580212 6802
rect 580170 6624 580226 6633
rect 580170 6559 580226 6568
rect 367100 5500 367152 5506
rect 367100 5442 367152 5448
rect 581000 3528 581052 3534
rect 581000 3470 581052 3476
rect 360292 3460 360344 3466
rect 360292 3402 360344 3408
rect 353298 3360 353354 3369
rect 353298 3295 353354 3304
rect 581012 480 581040 3470
rect 582196 3324 582248 3330
rect 582196 3266 582248 3272
rect 582208 480 582236 3266
rect 583404 480 583432 16546
rect 583496 3534 583524 213143
rect 583588 206281 583616 287671
rect 583758 225584 583814 225593
rect 583758 225519 583814 225528
rect 583666 222864 583722 222873
rect 583666 222799 583722 222808
rect 583574 206272 583630 206281
rect 583574 206207 583630 206216
rect 583574 204912 583630 204921
rect 583574 204847 583630 204856
rect 583484 3528 583536 3534
rect 583484 3470 583536 3476
rect 583588 3330 583616 204847
rect 583680 33114 583708 222799
rect 583772 86737 583800 225519
rect 583758 86728 583814 86737
rect 583758 86663 583814 86672
rect 583668 33108 583720 33114
rect 583668 33050 583720 33056
rect 583576 3324 583628 3330
rect 583576 3266 583628 3272
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 684256 3478 684312
rect 3514 671200 3570 671256
rect 3422 658164 3478 658200
rect 3422 658144 3424 658164
rect 3424 658144 3476 658164
rect 3476 658144 3478 658164
rect 3422 632068 3424 632088
rect 3424 632068 3476 632088
rect 3476 632068 3478 632088
rect 3422 632032 3478 632068
rect 3146 619112 3202 619168
rect 3238 606056 3294 606112
rect 3422 579944 3478 580000
rect 3422 566888 3478 566944
rect 3422 553832 3478 553888
rect 3422 527856 3478 527912
rect 2778 514820 2834 514856
rect 2778 514800 2780 514820
rect 2780 514800 2832 514820
rect 2832 514800 2834 514820
rect 3330 475632 3386 475688
rect 3514 501744 3570 501800
rect 3514 462576 3570 462632
rect 3146 449520 3202 449576
rect 35806 526360 35862 526416
rect 3422 423580 3424 423600
rect 3424 423580 3476 423600
rect 3476 423580 3478 423600
rect 3422 423544 3478 423580
rect 3422 410488 3478 410544
rect 2778 397432 2834 397488
rect 4802 380976 4858 381032
rect 3514 371320 3570 371376
rect 3330 358400 3386 358456
rect 2778 345344 2834 345400
rect 3330 267144 3386 267200
rect 3146 254088 3202 254144
rect 4066 319232 4122 319288
rect 3514 306176 3570 306232
rect 3514 293120 3570 293176
rect 3514 241032 3570 241088
rect 3422 214920 3478 214976
rect 3422 201864 3478 201920
rect 3238 162832 3294 162888
rect 3146 110608 3202 110664
rect 3238 84632 3294 84688
rect 3330 58520 3386 58576
rect 2870 32408 2926 32464
rect 3514 188808 3570 188864
rect 3514 149776 3570 149832
rect 3514 136720 3570 136776
rect 3514 97552 3570 97608
rect 5446 79328 5502 79384
rect 3514 71576 3570 71632
rect 3514 45500 3516 45520
rect 3516 45500 3568 45520
rect 3568 45500 3570 45520
rect 3514 45464 3570 45500
rect 4066 35128 4122 35184
rect 3422 19352 3478 19408
rect 3974 17176 4030 17232
rect 570 8880 626 8936
rect 18 6840 74 6896
rect 15842 383696 15898 383752
rect 17222 329976 17278 330032
rect 32402 222808 32458 222864
rect 30286 83408 30342 83464
rect 15842 80688 15898 80744
rect 15106 61376 15162 61432
rect 10966 42064 11022 42120
rect 7654 3304 7710 3360
rect 19246 75248 19302 75304
rect 16486 33768 16542 33824
rect 23386 54440 23442 54496
rect 22006 51720 22062 51776
rect 31666 55800 31722 55856
rect 39854 384240 39910 384296
rect 41326 415384 41382 415440
rect 39946 238584 40002 238640
rect 46846 257896 46902 257952
rect 48134 240080 48190 240136
rect 43442 221448 43498 221504
rect 41326 77832 41382 77888
rect 38566 58520 38622 58576
rect 35806 57160 35862 57216
rect 33046 36488 33102 36544
rect 39946 48864 40002 48920
rect 48134 65456 48190 65512
rect 45466 59880 45522 59936
rect 44086 50224 44142 50280
rect 50802 213560 50858 213616
rect 50894 73752 50950 73808
rect 55034 445712 55090 445768
rect 53746 444488 53802 444544
rect 53654 415384 53710 415440
rect 52274 314880 52330 314936
rect 52182 235864 52238 235920
rect 53562 285640 53618 285696
rect 53470 268368 53526 268424
rect 52274 225936 52330 225992
rect 54942 373224 54998 373280
rect 56506 407088 56562 407144
rect 55034 368328 55090 368384
rect 53654 241440 53710 241496
rect 53562 217776 53618 217832
rect 54942 204176 54998 204232
rect 53746 71032 53802 71088
rect 57702 338680 57758 338736
rect 57610 335552 57666 335608
rect 56506 215872 56562 215928
rect 55862 71168 55918 71224
rect 57610 232736 57666 232792
rect 61842 462848 61898 462904
rect 60646 445848 60702 445904
rect 59174 374040 59230 374096
rect 57702 230152 57758 230208
rect 59266 334328 59322 334384
rect 59082 231376 59138 231432
rect 58990 224848 59046 224904
rect 57886 72528 57942 72584
rect 61934 363024 61990 363080
rect 60462 194520 60518 194576
rect 61842 220768 61898 220824
rect 61934 187584 61990 187640
rect 62854 416608 62910 416664
rect 62854 415384 62910 415440
rect 65890 573416 65946 573472
rect 66074 590688 66130 590744
rect 65890 542272 65946 542328
rect 63406 415384 63462 415440
rect 63406 389136 63462 389192
rect 63314 386960 63370 387016
rect 63314 378664 63370 378720
rect 63222 332696 63278 332752
rect 64786 391176 64842 391232
rect 65798 389000 65854 389056
rect 65614 388728 65670 388784
rect 64694 376624 64750 376680
rect 63222 230288 63278 230344
rect 63130 226888 63186 226944
rect 61382 79464 61438 79520
rect 59266 72392 59322 72448
rect 60646 69536 60702 69592
rect 58622 64096 58678 64152
rect 65890 388864 65946 388920
rect 66810 588376 66866 588432
rect 66258 586508 66260 586528
rect 66260 586508 66312 586528
rect 66312 586508 66314 586528
rect 66258 586472 66314 586508
rect 66810 585656 66866 585712
rect 66810 582936 66866 582992
rect 66442 581712 66498 581768
rect 66810 580216 66866 580272
rect 67270 577496 67326 577552
rect 67086 574776 67142 574832
rect 66810 572056 66866 572112
rect 67178 570696 67234 570752
rect 66810 569336 66866 569392
rect 66718 567976 66774 568032
rect 66810 564984 66866 565040
rect 66810 563624 66866 563680
rect 66810 562264 66866 562320
rect 66810 560904 66866 560960
rect 66810 559544 66866 559600
rect 66810 558184 66866 558240
rect 66810 555464 66866 555520
rect 66534 554104 66590 554160
rect 66442 550024 66498 550080
rect 66442 548664 66498 548720
rect 66166 547304 66222 547360
rect 66810 545148 66866 545184
rect 66810 545128 66812 545148
rect 66812 545128 66864 545148
rect 66864 545128 66866 545148
rect 66810 544584 66866 544640
rect 66810 543224 66866 543280
rect 67086 541864 67142 541920
rect 67362 576156 67418 576192
rect 67362 576136 67364 576156
rect 67364 576136 67416 576156
rect 67416 576136 67418 576156
rect 72882 595448 72938 595504
rect 70306 590688 70362 590744
rect 71134 590688 71190 590744
rect 73158 589872 73214 589928
rect 87602 595448 87658 595504
rect 78586 592048 78642 592104
rect 77666 589464 77722 589520
rect 83186 590960 83242 591016
rect 82266 590688 82322 590744
rect 81346 589328 81402 589384
rect 81714 588648 81770 588704
rect 88062 588512 88118 588568
rect 67638 584296 67694 584352
rect 67546 574776 67602 574832
rect 67454 566752 67510 566808
rect 67454 552744 67510 552800
rect 67546 539588 67548 539608
rect 67548 539588 67600 539608
rect 67600 539588 67602 539608
rect 67546 539552 67602 539588
rect 67362 538056 67418 538112
rect 67086 537376 67142 537432
rect 66902 523776 66958 523832
rect 66810 437824 66866 437880
rect 66718 435376 66774 435432
rect 66810 433064 66866 433120
rect 66810 431024 66866 431080
rect 66810 428576 66866 428632
rect 66718 426264 66774 426320
rect 66810 424088 66866 424144
rect 66258 421912 66314 421968
rect 66810 415112 66866 415168
rect 67086 523640 67142 523696
rect 66902 410624 66958 410680
rect 66258 406136 66314 406192
rect 66258 403688 66314 403744
rect 66258 401548 66260 401568
rect 66260 401548 66312 401568
rect 66312 401548 66314 401568
rect 66258 401512 66314 401548
rect 66258 399492 66314 399528
rect 66258 399472 66260 399492
rect 66260 399472 66312 399492
rect 66312 399472 66314 399492
rect 66994 396888 67050 396944
rect 66626 392536 66682 392592
rect 66074 360848 66130 360904
rect 65890 336776 65946 336832
rect 65798 322360 65854 322416
rect 65982 322360 66038 322416
rect 65890 303048 65946 303104
rect 65890 281288 65946 281344
rect 64694 231648 64750 231704
rect 64510 219136 64566 219192
rect 67454 412800 67510 412856
rect 67362 345616 67418 345672
rect 66626 328888 66682 328944
rect 67270 324536 67326 324592
rect 66810 321272 66866 321328
rect 66902 320184 66958 320240
rect 66902 319096 66958 319152
rect 66810 318008 66866 318064
rect 67362 316920 67418 316976
rect 66074 271768 66130 271824
rect 66074 260888 66130 260944
rect 65982 234504 66038 234560
rect 66258 315832 66314 315888
rect 66810 313928 66866 313984
rect 66442 312840 66498 312896
rect 66994 311752 67050 311808
rect 66810 309576 66866 309632
rect 66902 307400 66958 307456
rect 66810 305224 66866 305280
rect 66810 304136 66866 304192
rect 66810 301960 66866 302016
rect 66902 300872 66958 300928
rect 66626 298696 66682 298752
rect 66810 297608 66866 297664
rect 66718 295432 66774 295488
rect 66810 294344 66866 294400
rect 66810 293256 66866 293312
rect 66810 292168 66866 292224
rect 66810 291080 66866 291136
rect 66902 289992 66958 290048
rect 66810 288904 66866 288960
rect 66626 287816 66682 287872
rect 66350 286728 66406 286784
rect 66810 285640 66866 285696
rect 66718 284552 66774 284608
rect 66810 283464 66866 283520
rect 66810 278024 66866 278080
rect 66810 277208 66866 277264
rect 66626 275032 66682 275088
rect 66258 272856 66314 272912
rect 66810 268504 66866 268560
rect 66810 265240 66866 265296
rect 66810 264152 66866 264208
rect 66810 263064 66866 263120
rect 66442 261976 66498 262032
rect 66810 259800 66866 259856
rect 66810 256536 66866 256592
rect 67730 578856 67786 578912
rect 89718 586200 89774 586256
rect 88890 577496 88946 577552
rect 88890 560088 88946 560144
rect 68650 536560 68706 536616
rect 68650 535472 68706 535528
rect 69570 535472 69626 535528
rect 70214 447072 70270 447128
rect 67822 442176 67878 442232
rect 67638 439864 67694 439920
rect 67730 419600 67786 419656
rect 67546 394848 67602 394904
rect 67454 310664 67510 310720
rect 67086 306312 67142 306368
rect 68742 445848 68798 445904
rect 70398 446392 70454 446448
rect 72422 536696 72478 536752
rect 71778 445848 71834 445904
rect 78034 448568 78090 448624
rect 82818 462848 82874 462904
rect 83462 460128 83518 460184
rect 81438 456184 81494 456240
rect 79414 444488 79470 444544
rect 84198 447208 84254 447264
rect 86866 457408 86922 457464
rect 88154 536560 88210 536616
rect 86958 454688 87014 454744
rect 85578 445712 85634 445768
rect 83830 444488 83886 444544
rect 89626 560088 89682 560144
rect 89626 543768 89682 543824
rect 90362 589872 90418 589928
rect 89810 567296 89866 567352
rect 89074 459584 89130 459640
rect 87050 444624 87106 444680
rect 93766 589328 93822 589384
rect 91742 587560 91798 587616
rect 91374 584840 91430 584896
rect 91190 583652 91192 583672
rect 91192 583652 91244 583672
rect 91244 583652 91246 583672
rect 91190 583616 91246 583652
rect 91742 582120 91798 582176
rect 91742 580760 91798 580816
rect 91742 579400 91798 579456
rect 91098 576680 91154 576736
rect 91098 575320 91154 575376
rect 91098 572600 91154 572656
rect 91190 571376 91246 571432
rect 91098 570036 91154 570072
rect 91098 570016 91100 570036
rect 91100 570016 91152 570036
rect 91152 570016 91154 570036
rect 91098 568656 91154 568712
rect 91374 565836 91376 565856
rect 91376 565836 91428 565856
rect 91428 565836 91430 565856
rect 91374 565800 91430 565836
rect 91374 564460 91430 564496
rect 91374 564440 91376 564460
rect 91376 564440 91428 564460
rect 91428 564440 91430 564460
rect 91374 563100 91430 563136
rect 91374 563080 91376 563100
rect 91376 563080 91428 563100
rect 91428 563080 91430 563100
rect 91098 561448 91154 561504
rect 92386 558728 92442 558784
rect 91190 557368 91246 557424
rect 91742 556008 91798 556064
rect 91742 554648 91798 554704
rect 91742 553288 91798 553344
rect 91190 552084 91246 552120
rect 91190 552064 91192 552084
rect 91192 552064 91244 552084
rect 91244 552064 91246 552084
rect 91190 550704 91246 550760
rect 91466 547884 91468 547904
rect 91468 547884 91520 547904
rect 91520 547884 91522 547904
rect 91466 547848 91522 547884
rect 91190 546508 91246 546544
rect 91190 546488 91192 546508
rect 91192 546488 91244 546508
rect 91244 546488 91246 546508
rect 91190 545148 91246 545184
rect 91190 545128 91192 545148
rect 91192 545128 91244 545148
rect 91244 545128 91246 545148
rect 91190 542428 91246 542464
rect 91190 542408 91192 542428
rect 91192 542408 91244 542428
rect 91244 542408 91246 542428
rect 91190 541184 91246 541240
rect 91834 543904 91890 543960
rect 92386 539688 92442 539744
rect 90454 456048 90510 456104
rect 93674 534656 93730 534712
rect 93214 464344 93270 464400
rect 95146 549344 95202 549400
rect 94502 467064 94558 467120
rect 95146 460128 95202 460184
rect 94778 445712 94834 445768
rect 97354 469784 97410 469840
rect 97262 457408 97318 457464
rect 154118 702480 154174 702536
rect 103518 592048 103574 592104
rect 100758 590960 100814 591016
rect 100850 589464 100906 589520
rect 98734 470600 98790 470656
rect 97998 456864 98054 456920
rect 98642 456864 98698 456920
rect 96618 445712 96674 445768
rect 97630 445712 97686 445768
rect 96526 444896 96582 444952
rect 100114 474000 100170 474056
rect 100022 451832 100078 451888
rect 104162 453192 104218 453248
rect 100850 445748 100852 445768
rect 100852 445748 100904 445768
rect 100904 445748 100906 445768
rect 100850 445712 100906 445748
rect 109038 582936 109094 582992
rect 107014 479440 107070 479496
rect 108946 467744 109002 467800
rect 109038 447072 109094 447128
rect 112442 458768 112498 458824
rect 118698 585656 118754 585712
rect 117962 553424 118018 553480
rect 118606 553424 118662 553480
rect 115294 447208 115350 447264
rect 109038 444624 109094 444680
rect 111706 444624 111762 444680
rect 113178 445712 113234 445768
rect 114374 445712 114430 445768
rect 117594 445712 117650 445768
rect 118606 445712 118662 445768
rect 120722 429256 120778 429312
rect 120722 417016 120778 417072
rect 120630 414568 120686 414624
rect 77666 391040 77722 391096
rect 68650 389272 68706 389328
rect 69938 390360 69994 390416
rect 68742 389000 68798 389056
rect 71778 389000 71834 389056
rect 73066 389000 73122 389056
rect 69662 380160 69718 380216
rect 73158 388864 73214 388920
rect 73802 388864 73858 388920
rect 69846 344256 69902 344312
rect 67638 310664 67694 310720
rect 67546 299784 67602 299840
rect 67454 282376 67510 282432
rect 67178 280220 67234 280256
rect 67178 280200 67180 280220
rect 67180 280200 67232 280220
rect 67232 280200 67234 280220
rect 67178 279112 67234 279168
rect 66994 273944 67050 274000
rect 67270 255448 67326 255504
rect 66994 253272 67050 253328
rect 66902 251096 66958 251152
rect 66810 250008 66866 250064
rect 66902 247832 66958 247888
rect 66810 246744 66866 246800
rect 66350 244568 66406 244624
rect 67086 242800 67142 242856
rect 66166 224712 66222 224768
rect 67362 241712 67418 241768
rect 67546 266328 67602 266384
rect 67270 236544 67326 236600
rect 67086 204856 67142 204912
rect 64786 190304 64842 190360
rect 66166 129240 66222 129296
rect 65982 125160 66038 125216
rect 64970 122576 65026 122632
rect 64786 121488 64842 121544
rect 64970 121488 65026 121544
rect 65890 102312 65946 102368
rect 65890 94968 65946 95024
rect 66074 123528 66130 123584
rect 67454 126248 67510 126304
rect 67362 120808 67418 120864
rect 67454 88984 67510 89040
rect 66166 81368 66222 81424
rect 64786 68312 64842 68368
rect 70030 331744 70086 331800
rect 69846 329568 69902 329624
rect 72238 334056 72294 334112
rect 73066 365744 73122 365800
rect 76378 385600 76434 385656
rect 75826 382880 75882 382936
rect 73802 379480 73858 379536
rect 75182 331200 75238 331256
rect 79506 388728 79562 388784
rect 81438 389000 81494 389056
rect 79966 386960 80022 387016
rect 80886 386960 80942 387016
rect 81346 373360 81402 373416
rect 76746 353368 76802 353424
rect 75826 331200 75882 331256
rect 77114 337320 77170 337376
rect 76654 329840 76710 329896
rect 77482 329160 77538 329216
rect 92938 391040 92994 391096
rect 81438 339496 81494 339552
rect 83186 329160 83242 329216
rect 89810 390360 89866 390416
rect 91650 389000 91706 389056
rect 90454 388864 90510 388920
rect 85670 338136 85726 338192
rect 89626 371320 89682 371376
rect 87602 370504 87658 370560
rect 87142 342216 87198 342272
rect 89534 340992 89590 341048
rect 115754 390632 115810 390688
rect 94226 390360 94282 390416
rect 93030 388728 93086 388784
rect 90362 353232 90418 353288
rect 91006 351056 91062 351112
rect 91926 330112 91982 330168
rect 93122 369824 93178 369880
rect 97354 390360 97410 390416
rect 95238 389000 95294 389056
rect 96250 389000 96306 389056
rect 97262 374584 97318 374640
rect 93858 364384 93914 364440
rect 95146 364384 95202 364440
rect 96526 356088 96582 356144
rect 98826 390360 98882 390416
rect 102138 390360 102194 390416
rect 100758 390224 100814 390280
rect 99194 389000 99250 389056
rect 100758 389000 100814 389056
rect 102322 389000 102378 389056
rect 103334 389000 103390 389056
rect 97814 360032 97870 360088
rect 98826 356904 98882 356960
rect 97262 341400 97318 341456
rect 97814 332832 97870 332888
rect 101402 388728 101458 388784
rect 99286 371864 99342 371920
rect 99194 356904 99250 356960
rect 100022 369960 100078 370016
rect 100666 349696 100722 349752
rect 100574 346432 100630 346488
rect 104990 390360 105046 390416
rect 106554 390360 106610 390416
rect 103334 355272 103390 355328
rect 101402 337456 101458 337512
rect 102046 343984 102102 344040
rect 106922 388320 106978 388376
rect 106186 381520 106242 381576
rect 104990 380976 105046 381032
rect 105542 380976 105598 381032
rect 104162 340040 104218 340096
rect 104990 346296 105046 346352
rect 106186 346296 106242 346352
rect 106186 345752 106242 345808
rect 108026 390360 108082 390416
rect 109498 390360 109554 390416
rect 108394 389272 108450 389328
rect 110234 357448 110290 357504
rect 107750 351192 107806 351248
rect 108486 349152 108542 349208
rect 112902 389000 112958 389056
rect 113178 389000 113234 389056
rect 114374 389000 114430 389056
rect 111062 380976 111118 381032
rect 111706 348336 111762 348392
rect 111614 340856 111670 340912
rect 115662 379208 115718 379264
rect 115662 378256 115718 378312
rect 114558 376488 114614 376544
rect 113178 353368 113234 353424
rect 113822 353368 113878 353424
rect 113822 343576 113878 343632
rect 112350 339632 112406 339688
rect 114466 331200 114522 331256
rect 115938 390360 115994 390416
rect 117870 390360 117926 390416
rect 118790 390360 118846 390416
rect 120446 388320 120502 388376
rect 119342 383696 119398 383752
rect 116490 377440 116546 377496
rect 115754 376488 115810 376544
rect 115754 375400 115810 375456
rect 116582 367648 116638 367704
rect 115846 360984 115902 361040
rect 116674 364520 116730 364576
rect 118606 353368 118662 353424
rect 118514 339360 118570 339416
rect 117042 332560 117098 332616
rect 119986 378120 120042 378176
rect 119894 343848 119950 343904
rect 121182 415248 121238 415304
rect 121642 442176 121698 442232
rect 121550 440000 121606 440056
rect 121550 435376 121606 435432
rect 121458 392672 121514 392728
rect 120722 386960 120778 387016
rect 122746 428440 122802 428496
rect 121550 381520 121606 381576
rect 121458 357992 121514 358048
rect 121734 353912 121790 353968
rect 121550 345616 121606 345672
rect 123574 451832 123630 451888
rect 123482 425992 123538 426048
rect 123022 424088 123078 424144
rect 122930 421912 122986 421968
rect 123022 397296 123078 397352
rect 122930 394712 122986 394768
rect 122930 384240 122986 384296
rect 124126 442060 124182 442096
rect 124126 442040 124128 442060
rect 124128 442040 124180 442060
rect 124180 442040 124182 442060
rect 124126 437824 124182 437880
rect 124126 433064 124182 433120
rect 124126 431024 124182 431080
rect 124126 420860 124128 420880
rect 124128 420860 124180 420880
rect 124180 420860 124182 420880
rect 124126 420824 124182 420860
rect 123850 412800 123906 412856
rect 123574 410624 123630 410680
rect 123758 403688 123814 403744
rect 124126 408312 124182 408368
rect 124126 406172 124128 406192
rect 124128 406172 124180 406192
rect 124180 406172 124182 406192
rect 124126 406136 124182 406172
rect 124126 401512 124182 401568
rect 124126 399492 124182 399528
rect 124310 447208 124366 447264
rect 124862 444760 124918 444816
rect 125506 443808 125562 443864
rect 124126 399472 124128 399492
rect 124128 399472 124180 399492
rect 124180 399472 124182 399492
rect 124126 397296 124182 397352
rect 123206 349016 123262 349072
rect 122838 348472 122894 348528
rect 126242 374584 126298 374640
rect 125506 368600 125562 368656
rect 125506 368328 125562 368384
rect 125598 368192 125654 368248
rect 126886 368192 126942 368248
rect 124126 349016 124182 349072
rect 124126 347792 124182 347848
rect 123482 344256 123538 344312
rect 124034 343732 124090 343768
rect 124034 343712 124036 343732
rect 124036 343712 124088 343732
rect 124088 343712 124090 343732
rect 124862 350512 124918 350568
rect 124862 329976 124918 330032
rect 126886 367104 126942 367160
rect 187606 589348 187662 589384
rect 187606 589328 187608 589348
rect 187608 589328 187660 589348
rect 187660 589328 187662 589348
rect 129002 448568 129058 448624
rect 126978 366968 127034 367024
rect 127622 366968 127678 367024
rect 126978 366288 127034 366344
rect 127070 351872 127126 351928
rect 127714 351872 127770 351928
rect 133142 541048 133198 541104
rect 133142 536696 133198 536752
rect 131762 407768 131818 407824
rect 129738 353232 129794 353288
rect 129738 352008 129794 352064
rect 129002 345072 129058 345128
rect 134706 559544 134762 559600
rect 137926 545128 137982 545184
rect 133786 361664 133842 361720
rect 133694 354728 133750 354784
rect 130474 352008 130530 352064
rect 130474 342352 130530 342408
rect 131210 342352 131266 342408
rect 131118 338272 131174 338328
rect 131762 338408 131818 338464
rect 133878 352008 133934 352064
rect 134706 351056 134762 351112
rect 137282 364656 137338 364712
rect 136638 358808 136694 358864
rect 142066 542408 142122 542464
rect 141422 444896 141478 444952
rect 137926 358808 137982 358864
rect 140778 349288 140834 349344
rect 141422 349288 141478 349344
rect 148322 537104 148378 537160
rect 146942 535336 146998 535392
rect 143446 533976 143502 534032
rect 142802 533568 142858 533624
rect 143446 533568 143502 533624
rect 144182 391856 144238 391912
rect 142894 377304 142950 377360
rect 142802 341536 142858 341592
rect 144734 345616 144790 345672
rect 141882 331336 141938 331392
rect 148322 447072 148378 447128
rect 147586 363160 147642 363216
rect 146206 362208 146262 362264
rect 147586 355272 147642 355328
rect 146942 347928 146998 347984
rect 146758 334192 146814 334248
rect 147034 345072 147090 345128
rect 147034 337456 147090 337512
rect 155222 467880 155278 467936
rect 149702 355272 149758 355328
rect 150346 353504 150402 353560
rect 149058 334328 149114 334384
rect 152462 367648 152518 367704
rect 151082 334600 151138 334656
rect 152554 358672 152610 358728
rect 153106 358672 153162 358728
rect 153106 357720 153162 357776
rect 153014 339768 153070 339824
rect 153014 338680 153070 338736
rect 152646 329976 152702 330032
rect 155222 355952 155278 356008
rect 155222 353368 155278 353424
rect 155774 343984 155830 344040
rect 155130 341400 155186 341456
rect 155498 340992 155554 341048
rect 153842 339360 153898 339416
rect 155498 338000 155554 338056
rect 155774 336776 155830 336832
rect 159362 535744 159418 535800
rect 157982 444488 158038 444544
rect 156786 368600 156842 368656
rect 156694 367104 156750 367160
rect 154854 331880 154910 331936
rect 155866 334636 155868 334656
rect 155868 334636 155920 334656
rect 155920 334636 155922 334656
rect 155866 334600 155922 334636
rect 156786 329024 156842 329080
rect 157246 328480 157302 328536
rect 67822 308488 67878 308544
rect 159362 357992 159418 358048
rect 157430 331336 157486 331392
rect 157338 300328 157394 300384
rect 67730 296520 67786 296576
rect 156786 271088 156842 271144
rect 67822 270680 67878 270736
rect 67730 245656 67786 245712
rect 67638 228928 67694 228984
rect 80978 241984 81034 242040
rect 69754 241868 69810 241904
rect 69754 241848 69756 241868
rect 69756 241848 69808 241868
rect 69808 241848 69810 241868
rect 69662 241712 69718 241768
rect 69110 238448 69166 238504
rect 69754 217912 69810 217968
rect 71686 239400 71742 239456
rect 71778 238584 71834 238640
rect 71778 237360 71834 237416
rect 72422 237360 72478 237416
rect 77298 240080 77354 240136
rect 75826 210840 75882 210896
rect 78494 237224 78550 237280
rect 77298 214512 77354 214568
rect 79874 198600 79930 198656
rect 72422 195200 72478 195256
rect 80702 239536 80758 239592
rect 154670 241984 154726 242040
rect 83324 241440 83380 241496
rect 83554 241440 83610 241496
rect 81346 206216 81402 206272
rect 85118 239944 85174 240000
rect 86222 239400 86278 239456
rect 83462 230424 83518 230480
rect 82818 209616 82874 209672
rect 86774 208256 86830 208312
rect 87602 239536 87658 239592
rect 87142 212472 87198 212528
rect 87602 206760 87658 206816
rect 86866 197240 86922 197296
rect 88982 193840 89038 193896
rect 79966 192480 80022 192536
rect 89718 237224 89774 237280
rect 89718 236000 89774 236056
rect 90362 236000 90418 236056
rect 91006 216416 91062 216472
rect 92386 199280 92442 199336
rect 93950 235864 94006 235920
rect 95146 235864 95202 235920
rect 95146 235184 95202 235240
rect 93858 219272 93914 219328
rect 95146 219272 95202 219328
rect 93766 209480 93822 209536
rect 93122 193160 93178 193216
rect 96618 238176 96674 238232
rect 102782 228792 102838 228848
rect 103426 236680 103482 236736
rect 100942 224576 100998 224632
rect 102046 224576 102102 224632
rect 100666 212336 100722 212392
rect 97998 211112 98054 211168
rect 99286 211112 99342 211168
rect 99286 210704 99342 210760
rect 96526 206896 96582 206952
rect 102046 203496 102102 203552
rect 104806 190984 104862 191040
rect 107658 236680 107714 236736
rect 111062 221992 111118 222048
rect 112994 217640 113050 217696
rect 113638 239536 113694 239592
rect 114558 238312 114614 238368
rect 114650 235864 114706 235920
rect 117134 207576 117190 207632
rect 117410 233008 117466 233064
rect 118698 209344 118754 209400
rect 121366 240760 121422 240816
rect 121642 240216 121698 240272
rect 122286 239400 122342 239456
rect 121366 202816 121422 202872
rect 128358 210976 128414 211032
rect 129830 232872 129886 232928
rect 132590 233824 132646 233880
rect 135166 228656 135222 228712
rect 136454 215192 136510 215248
rect 131026 205536 131082 205592
rect 129646 202680 129702 202736
rect 136546 201184 136602 201240
rect 122746 196560 122802 196616
rect 107566 189624 107622 189680
rect 99286 186904 99342 186960
rect 95146 186224 95202 186280
rect 103426 183640 103482 183696
rect 99470 182144 99526 182200
rect 98458 180920 98514 180976
rect 97354 179424 97410 179480
rect 98458 177520 98514 177576
rect 97354 176840 97410 176896
rect 100758 180784 100814 180840
rect 100758 177520 100814 177576
rect 105910 177520 105966 177576
rect 107566 177520 107622 177576
rect 114374 179560 114430 179616
rect 114190 177556 114192 177576
rect 114192 177556 114244 177576
rect 114244 177556 114246 177576
rect 114190 177520 114246 177556
rect 138018 237224 138074 237280
rect 137282 226072 137338 226128
rect 139398 222128 139454 222184
rect 115846 182280 115902 182336
rect 115846 177520 115902 177576
rect 118606 177520 118662 177576
rect 121918 177520 121974 177576
rect 113086 177112 113142 177168
rect 114374 177112 114430 177168
rect 119894 177112 119950 177168
rect 125506 177520 125562 177576
rect 127990 177556 127992 177576
rect 127992 177556 128044 177576
rect 128044 177556 128046 177576
rect 127990 177520 128046 177556
rect 142986 237224 143042 237280
rect 142802 236544 142858 236600
rect 142986 235728 143042 235784
rect 143354 235184 143410 235240
rect 143538 237088 143594 237144
rect 143446 220632 143502 220688
rect 146804 241304 146860 241360
rect 147218 240216 147274 240272
rect 146850 236680 146906 236736
rect 146206 234368 146262 234424
rect 146850 231784 146906 231840
rect 144918 227432 144974 227488
rect 146942 226888 146998 226944
rect 147494 223488 147550 223544
rect 146942 216280 146998 216336
rect 146942 207032 146998 207088
rect 146942 206760 146998 206816
rect 147678 236952 147734 237008
rect 150438 235184 150494 235240
rect 150346 219000 150402 219056
rect 151910 240760 151966 240816
rect 154164 241440 154220 241496
rect 155130 241168 155186 241224
rect 152094 237224 152150 237280
rect 151726 204040 151782 204096
rect 142066 185544 142122 185600
rect 155222 240080 155278 240136
rect 155774 240080 155830 240136
rect 156694 241576 156750 241632
rect 158166 324944 158222 325000
rect 158810 343576 158866 343632
rect 158718 323176 158774 323232
rect 158718 322088 158774 322144
rect 158718 317736 158774 317792
rect 158718 316648 158774 316704
rect 158718 313404 158774 313440
rect 158718 313384 158720 313404
rect 158720 313384 158772 313404
rect 158772 313384 158774 313404
rect 158718 311208 158774 311264
rect 158902 328616 158958 328672
rect 160834 355952 160890 356008
rect 159454 342896 159510 342952
rect 158902 327528 158958 327584
rect 158994 326440 159050 326496
rect 159086 325352 159142 325408
rect 158902 324264 158958 324320
rect 159362 319368 159418 319424
rect 159270 318824 159326 318880
rect 158810 310120 158866 310176
rect 158718 307944 158774 308000
rect 158718 306856 158774 306912
rect 158718 305768 158774 305824
rect 158718 304680 158774 304736
rect 158810 303592 158866 303648
rect 158810 301416 158866 301472
rect 158810 298696 158866 298752
rect 158442 284824 158498 284880
rect 157982 264696 158038 264752
rect 157338 240760 157394 240816
rect 158442 261432 158498 261488
rect 158166 243480 158222 243536
rect 158074 236952 158130 237008
rect 158718 297064 158774 297120
rect 158718 295976 158774 296032
rect 158718 293800 158774 293856
rect 158718 291896 158774 291952
rect 158718 290808 158774 290864
rect 158810 289720 158866 289776
rect 158718 287544 158774 287600
rect 158718 286456 158774 286512
rect 158718 285368 158774 285424
rect 158718 284280 158774 284336
rect 158810 283192 158866 283248
rect 158718 282104 158774 282160
rect 158810 281016 158866 281072
rect 158718 279928 158774 279984
rect 158718 278840 158774 278896
rect 158718 276664 158774 276720
rect 158810 275576 158866 275632
rect 158718 274488 158774 274544
rect 158718 273400 158774 273456
rect 158718 269048 158774 269104
rect 158718 267980 158774 268016
rect 158718 267960 158720 267980
rect 158720 267960 158772 267980
rect 158772 267960 158774 267980
rect 158718 263628 158774 263664
rect 158718 263608 158720 263628
rect 158720 263608 158772 263628
rect 158772 263608 158774 263628
rect 158718 258168 158774 258224
rect 158810 256264 158866 256320
rect 158718 255212 158720 255232
rect 158720 255212 158772 255232
rect 158772 255212 158774 255232
rect 158718 255176 158774 255212
rect 158718 253000 158774 253056
rect 158810 249736 158866 249792
rect 158718 248648 158774 248704
rect 158626 245792 158682 245848
rect 158718 244316 158774 244352
rect 158718 244296 158720 244316
rect 158720 244296 158772 244316
rect 158772 244296 158774 244316
rect 158718 243208 158774 243264
rect 158810 241168 158866 241224
rect 159914 311072 159970 311128
rect 159454 300328 159510 300384
rect 159362 292984 159418 293040
rect 159638 298152 159694 298208
rect 159454 292440 159510 292496
rect 159362 282240 159418 282296
rect 159362 277752 159418 277808
rect 159362 271224 159418 271280
rect 159454 265784 159510 265840
rect 159362 261432 159418 261488
rect 159270 236000 159326 236056
rect 158626 233824 158682 233880
rect 155866 200640 155922 200696
rect 159914 259528 159970 259584
rect 159546 236000 159602 236056
rect 159362 221856 159418 221912
rect 159546 221448 159602 221504
rect 158626 199416 158682 199472
rect 154486 184184 154542 184240
rect 160006 254088 160062 254144
rect 160926 337456 160982 337512
rect 160926 328344 160982 328400
rect 160834 316648 160890 316704
rect 160834 311908 160890 311944
rect 160834 311888 160836 311908
rect 160836 311888 160888 311908
rect 160888 311888 160890 311908
rect 160834 262520 160890 262576
rect 160742 247152 160798 247208
rect 161202 251096 161258 251152
rect 160834 237224 160890 237280
rect 160742 220632 160798 220688
rect 161386 337320 161442 337376
rect 162214 355272 162270 355328
rect 162674 285640 162730 285696
rect 162122 269320 162178 269376
rect 161386 247152 161442 247208
rect 161294 244840 161350 244896
rect 162398 251776 162454 251832
rect 161202 209752 161258 209808
rect 162398 235728 162454 235784
rect 164146 313928 164202 313984
rect 163594 297336 163650 297392
rect 164698 356088 164754 356144
rect 164882 309712 164938 309768
rect 163594 279384 163650 279440
rect 162122 202680 162178 202736
rect 164146 266328 164202 266384
rect 164054 261432 164110 261488
rect 164146 237224 164202 237280
rect 164054 234640 164110 234696
rect 166354 364928 166410 364984
rect 165158 287680 165214 287736
rect 164974 251096 165030 251152
rect 164238 232872 164294 232928
rect 163594 230152 163650 230208
rect 165158 240760 165214 240816
rect 166446 332696 166502 332752
rect 166354 295160 166410 295216
rect 173162 536832 173218 536888
rect 169114 535608 169170 535664
rect 166906 272992 166962 273048
rect 166906 272448 166962 272504
rect 166446 245656 166502 245712
rect 166814 240080 166870 240136
rect 168194 355272 168250 355328
rect 166998 234640 167054 234696
rect 166814 223352 166870 223408
rect 166262 202136 166318 202192
rect 166354 201184 166410 201240
rect 169114 368328 169170 368384
rect 169022 334600 169078 334656
rect 168378 329704 168434 329760
rect 169758 385600 169814 385656
rect 169298 357584 169354 357640
rect 169666 357584 169722 357640
rect 169298 349696 169354 349752
rect 169022 301416 169078 301472
rect 169022 300192 169078 300248
rect 168654 268368 168710 268424
rect 167826 247560 167882 247616
rect 167826 241712 167882 241768
rect 168378 240760 168434 240816
rect 167826 232736 167882 232792
rect 159914 182824 159970 182880
rect 132406 177520 132462 177576
rect 133786 177520 133842 177576
rect 134798 177112 134854 177168
rect 99470 176704 99526 176760
rect 103426 176704 103482 176760
rect 123298 176704 123354 176760
rect 126794 176704 126850 176760
rect 129462 176704 129518 176760
rect 148230 176704 148286 176760
rect 158994 176740 158996 176760
rect 158996 176740 159048 176760
rect 159048 176740 159050 176760
rect 158994 176704 159050 176740
rect 128174 176432 128230 176488
rect 130750 175616 130806 175672
rect 135718 175616 135774 175672
rect 164882 178336 164938 178392
rect 166906 184320 166962 184376
rect 166262 179424 166318 179480
rect 167642 182144 167698 182200
rect 166446 179560 166502 179616
rect 166538 175480 166594 175536
rect 169298 303728 169354 303784
rect 169850 368328 169906 368384
rect 169850 325624 169906 325680
rect 169850 269184 169906 269240
rect 169850 222808 169906 222864
rect 170494 267552 170550 267608
rect 172610 349696 172666 349752
rect 173898 361528 173954 361584
rect 173254 330112 173310 330168
rect 172610 327120 172666 327176
rect 173162 311072 173218 311128
rect 172518 295296 172574 295352
rect 171874 273808 171930 273864
rect 175002 356768 175058 356824
rect 173346 319368 173402 319424
rect 175002 315968 175058 316024
rect 175002 315288 175058 315344
rect 174542 289040 174598 289096
rect 173254 283192 173310 283248
rect 173162 249736 173218 249792
rect 173162 246200 173218 246256
rect 172058 235728 172114 235784
rect 171782 226072 171838 226128
rect 169206 202816 169262 202872
rect 169390 202272 169446 202328
rect 169022 176840 169078 176896
rect 168286 175208 168342 175264
rect 167918 171536 167974 171592
rect 171782 178200 171838 178256
rect 170494 175344 170550 175400
rect 174542 276664 174598 276720
rect 173254 237088 173310 237144
rect 173806 233008 173862 233064
rect 173806 232600 173862 232656
rect 171874 175888 171930 175944
rect 67638 128016 67694 128072
rect 67730 100680 67786 100736
rect 107750 94696 107806 94752
rect 117134 94696 117190 94752
rect 95054 93472 95110 93528
rect 115846 93472 115902 93528
rect 103334 93200 103390 93256
rect 110326 93200 110382 93256
rect 86774 92384 86830 92440
rect 89074 92384 89130 92440
rect 86130 92248 86186 92304
rect 75734 91160 75790 91216
rect 85486 91160 85542 91216
rect 67638 82592 67694 82648
rect 67546 68176 67602 68232
rect 70306 62736 70362 62792
rect 68926 44784 68982 44840
rect 88062 91160 88118 91216
rect 86130 90344 86186 90400
rect 88062 86808 88118 86864
rect 75826 66952 75882 67008
rect 78586 65592 78642 65648
rect 79966 61512 80022 61568
rect 82726 26832 82782 26888
rect 89626 62872 89682 62928
rect 102046 92384 102102 92440
rect 97814 91296 97870 91352
rect 99286 91296 99342 91352
rect 101862 91296 101918 91352
rect 91006 91160 91062 91216
rect 93766 91160 93822 91216
rect 94686 91160 94742 91216
rect 96526 91160 96582 91216
rect 94686 85448 94742 85504
rect 96526 84088 96582 84144
rect 97906 91160 97962 91216
rect 99194 91160 99250 91216
rect 97814 82728 97870 82784
rect 95146 79600 95202 79656
rect 93766 76608 93822 76664
rect 100574 91160 100630 91216
rect 100574 87488 100630 87544
rect 101954 91160 102010 91216
rect 106922 91704 106978 91760
rect 106646 91568 106702 91624
rect 103426 91160 103482 91216
rect 104254 91160 104310 91216
rect 104806 91160 104862 91216
rect 105542 91160 105598 91216
rect 106094 91160 106150 91216
rect 105542 87896 105598 87952
rect 104806 78512 104862 78568
rect 104806 73888 104862 73944
rect 106646 89528 106702 89584
rect 106186 82048 106242 82104
rect 110234 91296 110290 91352
rect 108946 91160 109002 91216
rect 110142 91160 110198 91216
rect 108946 83952 109002 84008
rect 108946 76472 109002 76528
rect 162214 92520 162270 92576
rect 112350 92384 112406 92440
rect 111246 91296 111302 91352
rect 111706 91160 111762 91216
rect 111062 78376 111118 78432
rect 114374 91296 114430 91352
rect 112994 91160 113050 91216
rect 114466 91160 114522 91216
rect 111614 53080 111670 53136
rect 132406 92384 132462 92440
rect 134706 92384 134762 92440
rect 136086 92420 136088 92440
rect 136088 92420 136140 92440
rect 136140 92420 136142 92440
rect 136086 92384 136142 92420
rect 119710 91704 119766 91760
rect 121734 91704 121790 91760
rect 123758 91704 123814 91760
rect 115846 91160 115902 91216
rect 117226 91160 117282 91216
rect 118054 91160 118110 91216
rect 118606 91160 118662 91216
rect 118054 85312 118110 85368
rect 112442 11600 112498 11656
rect 119894 91160 119950 91216
rect 120446 91160 120502 91216
rect 120814 91160 120870 91216
rect 120078 86672 120134 86728
rect 120446 86536 120502 86592
rect 119986 80824 120042 80880
rect 124034 91432 124090 91488
rect 126794 91432 126850 91488
rect 123942 91160 123998 91216
rect 123758 89664 123814 89720
rect 123482 88984 123538 89040
rect 122746 74024 122802 74080
rect 125506 91296 125562 91352
rect 125414 91160 125470 91216
rect 126702 91160 126758 91216
rect 126242 84768 126298 84824
rect 126886 91296 126942 91352
rect 128266 91160 128322 91216
rect 130750 91160 130806 91216
rect 133786 91160 133842 91216
rect 130750 88032 130806 88088
rect 129002 87488 129058 87544
rect 151542 91432 151598 91488
rect 130382 69672 130438 69728
rect 151726 91296 151782 91352
rect 151634 91160 151690 91216
rect 151082 76744 151138 76800
rect 152094 91180 152150 91216
rect 152094 91160 152096 91180
rect 152096 91160 152148 91180
rect 152148 91160 152150 91180
rect 153106 91060 153108 91080
rect 153108 91060 153160 91080
rect 153160 91060 153162 91080
rect 153106 91024 153162 91060
rect 157982 90480 158038 90536
rect 160098 90344 160154 90400
rect 160098 88168 160154 88224
rect 132498 21256 132554 21312
rect 142802 20032 142858 20088
rect 125874 3440 125930 3496
rect 136454 11600 136510 11656
rect 162122 89800 162178 89856
rect 165526 94968 165582 95024
rect 165434 94152 165490 94208
rect 165526 92520 165582 92576
rect 165434 90480 165490 90536
rect 164974 90344 165030 90400
rect 162122 78512 162178 78568
rect 166538 88168 166594 88224
rect 167642 88032 167698 88088
rect 166446 86808 166502 86864
rect 167826 111732 167828 111752
rect 167828 111732 167880 111752
rect 167880 111732 167882 111752
rect 167826 111696 167882 111732
rect 168194 110064 168250 110120
rect 167918 108704 167974 108760
rect 167826 93880 167882 93936
rect 167918 85448 167974 85504
rect 169298 85312 169354 85368
rect 169114 82592 169170 82648
rect 171966 94424 172022 94480
rect 171874 89528 171930 89584
rect 170678 84088 170734 84144
rect 171782 81368 171838 81424
rect 172150 94152 172206 94208
rect 175186 332016 175242 332072
rect 177946 557504 178002 557560
rect 177394 538736 177450 538792
rect 177302 538056 177358 538112
rect 176014 504328 176070 504384
rect 176014 373224 176070 373280
rect 175738 297472 175794 297528
rect 175278 268368 175334 268424
rect 174726 250008 174782 250064
rect 174634 247288 174690 247344
rect 175186 232464 175242 232520
rect 175278 216008 175334 216064
rect 174726 195880 174782 195936
rect 176106 332832 176162 332888
rect 176014 292712 176070 292768
rect 176566 282240 176622 282296
rect 176474 252592 176530 252648
rect 176750 338000 176806 338056
rect 176750 337320 176806 337376
rect 177486 338272 177542 338328
rect 177946 337320 178002 337376
rect 178038 329976 178094 330032
rect 178038 324944 178094 325000
rect 178038 316648 178094 316704
rect 177302 249736 177358 249792
rect 177394 244976 177450 245032
rect 176566 243616 176622 243672
rect 177302 227704 177358 227760
rect 176474 217776 176530 217832
rect 176014 86536 176070 86592
rect 176198 94016 176254 94072
rect 175922 21256 175978 21312
rect 174542 19896 174598 19952
rect 178774 358944 178830 359000
rect 180706 373224 180762 373280
rect 180154 365744 180210 365800
rect 178866 347928 178922 347984
rect 178866 330384 178922 330440
rect 178866 285776 178922 285832
rect 180706 361392 180762 361448
rect 180338 331880 180394 331936
rect 180338 291760 180394 291816
rect 180246 287544 180302 287600
rect 180062 278024 180118 278080
rect 178774 241304 178830 241360
rect 178038 234368 178094 234424
rect 178038 234096 178094 234152
rect 178682 234096 178738 234152
rect 177946 228656 178002 228712
rect 177946 227704 178002 227760
rect 180246 257896 180302 257952
rect 180246 250416 180302 250472
rect 181442 360984 181498 361040
rect 180338 241576 180394 241632
rect 180614 241576 180670 241632
rect 180154 219136 180210 219192
rect 180062 203496 180118 203552
rect 178682 197920 178738 197976
rect 180338 238448 180394 238504
rect 180246 199552 180302 199608
rect 180154 182280 180210 182336
rect 184386 556144 184442 556200
rect 182822 539688 182878 539744
rect 181534 314064 181590 314120
rect 181718 247152 181774 247208
rect 181534 244840 181590 244896
rect 177578 92112 177634 92168
rect 177394 69672 177450 69728
rect 180154 86672 180210 86728
rect 184294 536968 184350 537024
rect 184386 369008 184442 369064
rect 184202 354728 184258 354784
rect 183190 349152 183246 349208
rect 183006 322224 183062 322280
rect 182270 245792 182326 245848
rect 183190 322088 183246 322144
rect 185398 365472 185454 365528
rect 186962 538192 187018 538248
rect 185582 361800 185638 361856
rect 184386 342352 184442 342408
rect 185766 377304 185822 377360
rect 186134 364384 186190 364440
rect 185674 314200 185730 314256
rect 184294 306992 184350 307048
rect 184202 298016 184258 298072
rect 186042 301416 186098 301472
rect 184846 298016 184902 298072
rect 184846 296792 184902 296848
rect 184294 293120 184350 293176
rect 184018 287680 184074 287736
rect 183098 273808 183154 273864
rect 183558 260888 183614 260944
rect 185674 287272 185730 287328
rect 185674 282240 185730 282296
rect 185582 278024 185638 278080
rect 183098 234368 183154 234424
rect 183282 213868 183284 213888
rect 183284 213868 183336 213888
rect 183336 213868 183338 213888
rect 183282 213832 183338 213868
rect 182822 199416 182878 199472
rect 181534 93064 181590 93120
rect 181442 83952 181498 84008
rect 183466 180648 183522 180704
rect 182822 30912 182878 30968
rect 184386 250416 184442 250472
rect 184754 241304 184810 241360
rect 184754 226244 184756 226264
rect 184756 226244 184808 226264
rect 184808 226244 184810 226264
rect 184754 226208 184810 226244
rect 184386 179968 184442 180024
rect 187514 554784 187570 554840
rect 187054 381112 187110 381168
rect 186962 347656 187018 347712
rect 186134 296112 186190 296168
rect 185674 244976 185730 245032
rect 185582 237088 185638 237144
rect 185674 219136 185730 219192
rect 186226 245792 186282 245848
rect 186226 241304 186282 241360
rect 186134 187040 186190 187096
rect 184570 180920 184626 180976
rect 185582 170312 185638 170368
rect 184386 93608 184442 93664
rect 184294 91024 184350 91080
rect 193218 559544 193274 559600
rect 193218 559000 193274 559056
rect 187606 374584 187662 374640
rect 188618 380976 188674 381032
rect 188526 357720 188582 357776
rect 188434 354048 188490 354104
rect 187238 291760 187294 291816
rect 187606 251776 187662 251832
rect 187146 243616 187202 243672
rect 188434 319368 188490 319424
rect 187698 216416 187754 216472
rect 187698 216008 187754 216064
rect 191102 547848 191158 547904
rect 190366 533432 190422 533488
rect 189722 335552 189778 335608
rect 188710 323584 188766 323640
rect 189078 320184 189134 320240
rect 188526 300192 188582 300248
rect 188526 291216 188582 291272
rect 187790 209344 187846 209400
rect 187790 208392 187846 208448
rect 188342 203496 188398 203552
rect 187238 87896 187294 87952
rect 188434 196696 188490 196752
rect 191194 545400 191250 545456
rect 191746 541320 191802 541376
rect 189906 339768 189962 339824
rect 190090 331744 190146 331800
rect 189078 260072 189134 260128
rect 190182 252456 190238 252512
rect 188802 216008 188858 216064
rect 189078 212472 189134 212528
rect 188618 208392 188674 208448
rect 188618 195336 188674 195392
rect 188526 180784 188582 180840
rect 191194 378392 191250 378448
rect 191746 373360 191802 373416
rect 192574 549480 192630 549536
rect 191654 353368 191710 353424
rect 191746 351056 191802 351112
rect 191194 338680 191250 338736
rect 191194 332016 191250 332072
rect 191194 294480 191250 294536
rect 191194 284008 191250 284064
rect 191194 252456 191250 252512
rect 190458 197104 190514 197160
rect 191286 236952 191342 237008
rect 192666 365744 192722 365800
rect 195334 547984 195390 548040
rect 193954 538328 194010 538384
rect 193954 382880 194010 382936
rect 193862 364520 193918 364576
rect 192482 320728 192538 320784
rect 191746 243480 191802 243536
rect 192574 289856 192630 289912
rect 192574 251096 192630 251152
rect 191746 236000 191802 236056
rect 191746 231512 191802 231568
rect 191654 210296 191710 210352
rect 189722 177384 189778 177440
rect 191102 142704 191158 142760
rect 189722 92248 189778 92304
rect 188434 28192 188490 28248
rect 188342 20032 188398 20088
rect 186962 14456 187018 14512
rect 193034 251096 193090 251152
rect 193954 305632 194010 305688
rect 195242 380160 195298 380216
rect 194598 379480 194654 379536
rect 195702 376488 195758 376544
rect 195242 373904 195298 373960
rect 195242 367784 195298 367840
rect 195702 351328 195758 351384
rect 195242 347112 195298 347168
rect 194138 328480 194194 328536
rect 193954 282104 194010 282160
rect 194506 279248 194562 279304
rect 194322 234232 194378 234288
rect 192574 200776 192630 200832
rect 192482 183640 192538 183696
rect 196622 542544 196678 542600
rect 196622 386960 196678 387016
rect 195886 375944 195942 376000
rect 196622 374720 196678 374776
rect 195794 300872 195850 300928
rect 195426 284280 195482 284336
rect 195334 267280 195390 267336
rect 195334 242800 195390 242856
rect 195334 232600 195390 232656
rect 195242 225664 195298 225720
rect 195334 225528 195390 225584
rect 195150 215872 195206 215928
rect 195150 213696 195206 213752
rect 194506 178744 194562 178800
rect 192666 177248 192722 177304
rect 193954 152360 194010 152416
rect 191194 91024 191250 91080
rect 192574 89664 192630 89720
rect 193954 119448 194010 119504
rect 191102 4800 191158 4856
rect 195334 207168 195390 207224
rect 196714 356904 196770 356960
rect 198002 535472 198058 535528
rect 197358 532208 197414 532264
rect 197358 529760 197414 529816
rect 197358 527312 197414 527368
rect 197450 524728 197506 524784
rect 197358 522280 197414 522336
rect 197358 519832 197414 519888
rect 197358 517384 197414 517440
rect 197358 510176 197414 510232
rect 197358 507592 197414 507648
rect 197358 500384 197414 500440
rect 197358 495508 197414 495544
rect 197358 495488 197360 495508
rect 197360 495488 197412 495508
rect 197412 495488 197414 495508
rect 197358 492904 197414 492960
rect 197358 490456 197414 490512
rect 197358 488008 197414 488064
rect 198002 483112 198058 483168
rect 197358 480664 197414 480720
rect 197358 478216 197414 478272
rect 197358 475768 197414 475824
rect 197358 473356 197360 473376
rect 197360 473356 197412 473376
rect 197412 473356 197414 473376
rect 197358 473320 197414 473356
rect 197634 470872 197690 470928
rect 197358 468424 197414 468480
rect 197358 465976 197414 466032
rect 197358 463256 197414 463312
rect 197358 460808 197414 460864
rect 197358 458360 197414 458416
rect 197358 448588 197414 448624
rect 197358 448568 197360 448588
rect 197360 448568 197412 448588
rect 197412 448568 197414 448588
rect 197358 446120 197414 446176
rect 197358 443692 197414 443728
rect 197358 443672 197360 443692
rect 197360 443672 197412 443692
rect 197412 443672 197414 443692
rect 197358 441360 197414 441416
rect 197358 433880 197414 433936
rect 197358 428984 197414 429040
rect 197358 426536 197414 426592
rect 197358 424088 197414 424144
rect 197358 419192 197414 419248
rect 197358 414296 197414 414352
rect 197358 411848 197414 411904
rect 197358 409536 197414 409592
rect 197358 406952 197414 407008
rect 197358 402056 197414 402112
rect 197358 399608 197414 399664
rect 197358 397160 197414 397216
rect 197358 394732 197414 394768
rect 197358 394712 197360 394732
rect 197360 394712 197412 394732
rect 197412 394712 197414 394732
rect 197358 392264 197414 392320
rect 197358 387368 197414 387424
rect 197266 384920 197322 384976
rect 197358 380024 197414 380080
rect 196714 292576 196770 292632
rect 198554 529760 198610 529816
rect 198738 530576 198794 530632
rect 198646 500384 198702 500440
rect 205638 545400 205694 545456
rect 206282 545400 206338 545456
rect 199106 505144 199162 505200
rect 198830 463256 198886 463312
rect 198830 458360 198886 458416
rect 198646 455912 198702 455968
rect 198554 453464 198610 453520
rect 198462 393372 198518 393408
rect 198462 393352 198464 393372
rect 198464 393352 198516 393372
rect 198516 393352 198518 393372
rect 198462 392264 198518 392320
rect 198002 325624 198058 325680
rect 197174 282920 197230 282976
rect 197358 282376 197414 282432
rect 198002 281560 198058 281616
rect 197358 280744 197414 280800
rect 198278 280492 198334 280528
rect 198278 280472 198280 280492
rect 198280 280472 198332 280492
rect 198332 280472 198334 280492
rect 197358 279520 197414 279576
rect 196622 253000 196678 253056
rect 197082 241576 197138 241632
rect 196990 240896 197046 240952
rect 197082 240760 197138 240816
rect 195518 191120 195574 191176
rect 195426 187584 195482 187640
rect 195426 183096 195482 183152
rect 195426 176976 195482 177032
rect 195426 160656 195482 160712
rect 195334 11600 195390 11656
rect 197082 199416 197138 199472
rect 196714 182960 196770 183016
rect 197358 278568 197414 278624
rect 197358 277208 197414 277264
rect 197358 276684 197414 276720
rect 197358 276664 197360 276684
rect 197360 276664 197412 276684
rect 197412 276664 197414 276684
rect 197450 275848 197506 275904
rect 197358 275032 197414 275088
rect 197358 274524 197360 274544
rect 197360 274524 197412 274544
rect 197412 274524 197414 274544
rect 197358 274488 197414 274524
rect 197358 273672 197414 273728
rect 197358 272856 197414 272912
rect 197450 272312 197506 272368
rect 197358 271496 197414 271552
rect 198370 270952 198426 271008
rect 197358 268776 197414 268832
rect 197450 267960 197506 268016
rect 197358 266600 197414 266656
rect 197450 265240 197506 265296
rect 197358 264424 197414 264480
rect 197358 263644 197360 263664
rect 197360 263644 197412 263664
rect 197412 263644 197414 263664
rect 197358 263608 197414 263644
rect 197358 261468 197360 261488
rect 197360 261468 197412 261488
rect 197412 261468 197414 261488
rect 197358 261432 197414 261468
rect 197358 260072 197414 260128
rect 197358 259256 197414 259312
rect 197450 258712 197506 258768
rect 197450 257896 197506 257952
rect 198094 257352 198150 257408
rect 197450 256536 197506 256592
rect 197358 255720 197414 255776
rect 197358 255212 197360 255232
rect 197360 255212 197412 255232
rect 197412 255212 197414 255232
rect 197358 255176 197414 255212
rect 197358 253544 197414 253600
rect 198002 251776 198058 251832
rect 197358 251640 197414 251696
rect 197910 250824 197966 250880
rect 197358 250008 197414 250064
rect 197358 249464 197414 249520
rect 197450 248684 197452 248704
rect 197452 248684 197504 248704
rect 197504 248684 197506 248704
rect 197450 248648 197506 248684
rect 197450 247832 197506 247888
rect 197358 245928 197414 245984
rect 197358 245112 197414 245168
rect 198922 416744 198978 416800
rect 199014 382472 199070 382528
rect 212538 553424 212594 553480
rect 213458 538464 213514 538520
rect 213458 538192 213514 538248
rect 230478 556144 230534 556200
rect 225326 552064 225382 552120
rect 218702 547984 218758 548040
rect 216586 538736 216642 538792
rect 203706 535472 203762 535528
rect 217138 538464 217194 538520
rect 216678 538228 216680 538248
rect 216680 538228 216732 538248
rect 216732 538228 216734 538248
rect 216678 538192 216734 538228
rect 222474 538328 222530 538384
rect 231950 549480 232006 549536
rect 241518 559000 241574 559056
rect 237378 557504 237434 557560
rect 235262 545264 235318 545320
rect 240230 554784 240286 554840
rect 238758 541320 238814 541376
rect 243542 547848 243598 547904
rect 248510 546624 248566 546680
rect 253938 542544 253994 542600
rect 255962 541592 256018 541648
rect 257342 541592 257398 541648
rect 262218 541184 262274 541240
rect 265530 538192 265586 538248
rect 268566 546488 268622 546544
rect 270866 543768 270922 543824
rect 278042 549344 278098 549400
rect 280618 539688 280674 539744
rect 284298 542952 284354 543008
rect 283470 542408 283526 542464
rect 295522 539688 295578 539744
rect 293866 537104 293922 537160
rect 303618 550704 303674 550760
rect 300030 545128 300086 545184
rect 302146 537104 302202 537160
rect 320178 545128 320234 545184
rect 318706 538192 318762 538248
rect 321558 543904 321614 543960
rect 323582 541048 323638 541104
rect 335450 536968 335506 537024
rect 333794 536832 333850 536888
rect 342074 539552 342130 539608
rect 348698 539824 348754 539880
rect 345386 539416 345442 539472
rect 347686 538736 347742 538792
rect 349158 539416 349214 539472
rect 350354 538328 350410 538384
rect 355322 538192 355378 538248
rect 313370 535744 313426 535800
rect 276018 535608 276074 535664
rect 276938 535608 276994 535664
rect 315670 535472 315726 535528
rect 201406 535336 201462 535392
rect 216586 535336 216642 535392
rect 199842 534928 199898 534984
rect 199842 533976 199898 534032
rect 357622 542952 357678 543008
rect 357438 522280 357494 522336
rect 357622 534656 357678 534712
rect 358726 532072 358782 532128
rect 358910 529624 358966 529680
rect 358726 527196 358782 527232
rect 358726 527176 358728 527196
rect 358728 527176 358780 527196
rect 358780 527176 358782 527196
rect 358726 524728 358782 524784
rect 358726 522300 358782 522336
rect 358726 522280 358728 522300
rect 358728 522280 358780 522300
rect 358780 522280 358782 522300
rect 357898 520004 357900 520024
rect 357900 520004 357952 520024
rect 357952 520004 357954 520024
rect 357898 519968 357954 520004
rect 358726 517384 358782 517440
rect 358634 514936 358690 514992
rect 357530 512624 357586 512680
rect 357622 510040 357678 510096
rect 358726 505164 358782 505200
rect 358726 505144 358728 505164
rect 358728 505144 358780 505164
rect 358780 505144 358782 505164
rect 358726 502696 358782 502752
rect 358726 500248 358782 500304
rect 199382 384784 199438 384840
rect 199842 378392 199898 378448
rect 199842 377168 199898 377224
rect 201406 377168 201462 377224
rect 200302 375264 200358 375320
rect 200302 374720 200358 374776
rect 200118 373360 200174 373416
rect 198830 366424 198886 366480
rect 199382 353504 199438 353560
rect 198830 296656 198886 296712
rect 198830 295976 198886 296032
rect 198830 284552 198886 284608
rect 200118 309712 200174 309768
rect 201406 338716 201408 338736
rect 201408 338716 201460 338736
rect 201460 338716 201462 338736
rect 201406 338680 201462 338716
rect 200762 309712 200818 309768
rect 202050 377304 202106 377360
rect 202234 377304 202290 377360
rect 204442 377576 204498 377632
rect 202234 312568 202290 312624
rect 201682 292576 201738 292632
rect 201406 288496 201462 288552
rect 200394 285776 200450 285832
rect 200302 284824 200358 284880
rect 200762 285640 200818 285696
rect 202234 291216 202290 291272
rect 203614 302776 203670 302832
rect 204902 375400 204958 375456
rect 207110 375944 207166 376000
rect 206650 375264 206706 375320
rect 204994 337456 205050 337512
rect 204442 290400 204498 290456
rect 203154 287272 203210 287328
rect 202878 285776 202934 285832
rect 205178 306448 205234 306504
rect 204258 284416 204314 284472
rect 203706 284280 203762 284336
rect 204902 285640 204958 285696
rect 206466 362208 206522 362264
rect 206558 330384 206614 330440
rect 206466 318008 206522 318064
rect 206466 295296 206522 295352
rect 206098 286048 206154 286104
rect 205546 285912 205602 285968
rect 207018 299376 207074 299432
rect 207754 299376 207810 299432
rect 207018 298288 207074 298344
rect 207570 285676 207572 285696
rect 207572 285676 207624 285696
rect 207624 285676 207626 285696
rect 207570 285640 207626 285676
rect 208122 289176 208178 289232
rect 208030 284280 208086 284336
rect 211066 342896 211122 342952
rect 209870 342216 209926 342272
rect 211066 342216 211122 342272
rect 209778 337592 209834 337648
rect 209226 317464 209282 317520
rect 209134 315288 209190 315344
rect 209410 317464 209466 317520
rect 214562 374040 214618 374096
rect 211986 358808 212042 358864
rect 211894 329024 211950 329080
rect 211066 295160 211122 295216
rect 211986 324944 212042 325000
rect 213274 316104 213330 316160
rect 213182 311208 213238 311264
rect 212906 296112 212962 296168
rect 211894 291080 211950 291136
rect 212446 291080 212502 291136
rect 211802 287408 211858 287464
rect 212354 284416 212410 284472
rect 217414 369008 217470 369064
rect 215942 345752 215998 345808
rect 216034 334056 216090 334112
rect 215390 328344 215446 328400
rect 214562 312432 214618 312488
rect 214746 285776 214802 285832
rect 214378 285640 214434 285696
rect 214746 284280 214802 284336
rect 215942 289176 215998 289232
rect 215390 285776 215446 285832
rect 215850 285640 215906 285696
rect 201406 284008 201462 284064
rect 218150 366424 218206 366480
rect 218702 362344 218758 362400
rect 217414 287272 217470 287328
rect 218702 302912 218758 302968
rect 222106 365744 222162 365800
rect 220818 365472 220874 365528
rect 222106 365472 222162 365528
rect 222934 369960 222990 370016
rect 219438 296248 219494 296304
rect 222842 337320 222898 337376
rect 221554 323584 221610 323640
rect 221186 293936 221242 293992
rect 218610 284552 218666 284608
rect 220082 287136 220138 287192
rect 220174 285776 220230 285832
rect 220634 285776 220690 285832
rect 223578 357992 223634 358048
rect 223026 357448 223082 357504
rect 221646 293936 221702 293992
rect 222842 293936 222898 293992
rect 223026 297472 223082 297528
rect 223026 295160 223082 295216
rect 222934 285912 222990 285968
rect 224314 320728 224370 320784
rect 223670 287272 223726 287328
rect 225142 303728 225198 303784
rect 224314 289992 224370 290048
rect 216034 284008 216090 284064
rect 201130 283872 201186 283928
rect 215942 283872 215998 283928
rect 219346 283872 219402 283928
rect 225142 285640 225198 285696
rect 226430 311072 226486 311128
rect 227166 312568 227222 312624
rect 226982 306992 227038 307048
rect 226890 289992 226946 290048
rect 226522 289720 226578 289776
rect 226522 288632 226578 288688
rect 229742 363160 229798 363216
rect 232502 351872 232558 351928
rect 229742 335416 229798 335472
rect 227718 305768 227774 305824
rect 228362 305768 228418 305824
rect 227166 289720 227222 289776
rect 227902 292440 227958 292496
rect 228638 305632 228694 305688
rect 227902 292032 227958 292088
rect 228454 292032 228510 292088
rect 228638 291216 228694 291272
rect 228914 291216 228970 291272
rect 224682 283872 224738 283928
rect 227994 283872 228050 283928
rect 230386 311208 230442 311264
rect 230754 287544 230810 287600
rect 229466 283872 229522 283928
rect 231030 283872 231086 283928
rect 233974 322088 234030 322144
rect 233882 319368 233938 319424
rect 232778 289856 232834 289912
rect 233146 287680 233202 287736
rect 233974 285640 234030 285696
rect 234618 302912 234674 302968
rect 235170 288360 235226 288416
rect 235170 287272 235226 287328
rect 239770 375264 239826 375320
rect 238022 357584 238078 357640
rect 236642 338680 236698 338736
rect 235906 288360 235962 288416
rect 240874 359352 240930 359408
rect 239402 329840 239458 329896
rect 238022 322088 238078 322144
rect 236642 287136 236698 287192
rect 236642 285640 236698 285696
rect 236734 283872 236790 283928
rect 239494 326304 239550 326360
rect 240874 351192 240930 351248
rect 238114 285912 238170 285968
rect 240138 305768 240194 305824
rect 239954 285640 240010 285696
rect 241426 298288 241482 298344
rect 240874 288360 240930 288416
rect 240874 287136 240930 287192
rect 243542 371864 243598 371920
rect 247038 376488 247094 376544
rect 248050 376488 248106 376544
rect 247038 368328 247094 368384
rect 243542 323584 243598 323640
rect 243910 313928 243966 313984
rect 242898 285912 242954 285968
rect 242346 284552 242402 284608
rect 238206 283872 238262 283928
rect 244094 300192 244150 300248
rect 244186 286048 244242 286104
rect 244186 283464 244242 283520
rect 251362 375264 251418 375320
rect 250442 353912 250498 353968
rect 248602 338136 248658 338192
rect 248418 334600 248474 334656
rect 247038 332560 247094 332616
rect 244278 278024 244334 278080
rect 200026 275848 200082 275904
rect 199474 270136 199530 270192
rect 199382 265784 199438 265840
rect 198646 263064 198702 263120
rect 198554 262248 198610 262304
rect 198462 244296 198518 244352
rect 198002 243752 198058 243808
rect 197450 243480 197506 243536
rect 197358 242936 197414 242992
rect 197818 242120 197874 242176
rect 198554 230288 198610 230344
rect 198462 211928 198518 211984
rect 198002 196560 198058 196616
rect 196714 100000 196770 100056
rect 244370 255176 244426 255232
rect 244278 250824 244334 250880
rect 199842 246200 199898 246256
rect 244002 244840 244058 244896
rect 199934 241712 199990 241768
rect 200026 241304 200082 241360
rect 199934 240080 199990 240136
rect 200578 240080 200634 240136
rect 199934 232600 199990 232656
rect 202602 240080 202658 240136
rect 202786 240116 202788 240136
rect 202788 240116 202840 240136
rect 202840 240116 202842 240136
rect 202786 240080 202842 240116
rect 201498 221992 201554 222048
rect 200762 192616 200818 192672
rect 202234 221992 202290 222048
rect 204258 238448 204314 238504
rect 204258 237360 204314 237416
rect 202970 234232 203026 234288
rect 203522 230288 203578 230344
rect 204166 234232 204222 234288
rect 203614 209072 203670 209128
rect 204442 235592 204498 235648
rect 205546 239536 205602 239592
rect 205822 238584 205878 238640
rect 205362 237360 205418 237416
rect 204994 222808 205050 222864
rect 204902 217368 204958 217424
rect 204166 181464 204222 181520
rect 203614 149232 203670 149288
rect 202234 113328 202290 113384
rect 200854 98368 200910 98424
rect 200762 43424 200818 43480
rect 205822 207032 205878 207088
rect 207018 237224 207074 237280
rect 207938 240080 207994 240136
rect 208214 240080 208270 240136
rect 207662 239536 207718 239592
rect 208306 239944 208362 240000
rect 207662 211928 207718 211984
rect 206466 207032 206522 207088
rect 208398 237224 208454 237280
rect 208398 235864 208454 235920
rect 209226 237224 209282 237280
rect 208858 235728 208914 235784
rect 208490 232600 208546 232656
rect 208398 231512 208454 231568
rect 208306 211928 208362 211984
rect 207754 209616 207810 209672
rect 210698 240080 210754 240136
rect 210330 237088 210386 237144
rect 209778 234504 209834 234560
rect 210974 234504 211030 234560
rect 210974 231104 211030 231160
rect 209778 219408 209834 219464
rect 209778 213560 209834 213616
rect 209686 211248 209742 211304
rect 206374 188536 206430 188592
rect 211894 234640 211950 234696
rect 211066 219408 211122 219464
rect 212722 235864 212778 235920
rect 212722 234640 212778 234696
rect 212170 228656 212226 228712
rect 212170 228248 212226 228304
rect 211342 215872 211398 215928
rect 213918 240116 213920 240136
rect 213920 240116 213972 240136
rect 213972 240116 213974 240136
rect 213918 240080 213974 240116
rect 214194 240080 214250 240136
rect 213826 239400 213882 239456
rect 213642 238584 213698 238640
rect 214194 238176 214250 238232
rect 213826 238040 213882 238096
rect 215298 234504 215354 234560
rect 216034 234504 216090 234560
rect 215298 231648 215354 231704
rect 211802 193160 211858 193216
rect 210422 181328 210478 181384
rect 207754 178064 207810 178120
rect 213274 215056 213330 215112
rect 213274 201320 213330 201376
rect 215114 222264 215170 222320
rect 215206 214512 215262 214568
rect 214562 207712 214618 207768
rect 216586 235728 216642 235784
rect 217506 240080 217562 240136
rect 217966 240080 218022 240136
rect 218426 240080 218482 240136
rect 218702 240080 218758 240136
rect 219530 238448 219586 238504
rect 218702 223488 218758 223544
rect 218058 204176 218114 204232
rect 217414 184456 217470 184512
rect 221370 240080 221426 240136
rect 221002 238312 221058 238368
rect 221462 234232 221518 234288
rect 223486 238584 223542 238640
rect 223302 233008 223358 233064
rect 220082 182960 220138 183016
rect 213826 178608 213882 178664
rect 213918 175616 213974 175672
rect 214562 175228 214618 175264
rect 214562 175208 214564 175228
rect 214564 175208 214616 175228
rect 214616 175208 214618 175228
rect 213918 174936 213974 174992
rect 214010 174256 214066 174312
rect 220266 210296 220322 210352
rect 220726 192480 220782 192536
rect 220726 185816 220782 185872
rect 223394 192480 223450 192536
rect 222842 181600 222898 181656
rect 226706 238312 226762 238368
rect 226706 238040 226762 238096
rect 226154 232464 226210 232520
rect 226246 180648 226302 180704
rect 224866 176840 224922 176896
rect 226338 176704 226394 176760
rect 228362 235592 228418 235648
rect 228178 234368 228234 234424
rect 227626 225936 227682 225992
rect 230570 240080 230626 240136
rect 230754 240080 230810 240136
rect 230202 235592 230258 235648
rect 228362 221856 228418 221912
rect 227718 219544 227774 219600
rect 226982 178880 227038 178936
rect 227718 178608 227774 178664
rect 226522 177384 226578 177440
rect 227718 177384 227774 177440
rect 229006 181192 229062 181248
rect 229190 178880 229246 178936
rect 229098 173712 229154 173768
rect 214930 173576 214986 173632
rect 213918 172896 213974 172952
rect 213918 172216 213974 172272
rect 214010 171536 214066 171592
rect 213918 171028 213920 171048
rect 213920 171028 213972 171048
rect 213972 171028 213974 171048
rect 213918 170992 213974 171028
rect 214010 170312 214066 170368
rect 214102 170176 214158 170232
rect 213918 169652 213974 169688
rect 213918 169632 213920 169652
rect 213920 169632 213972 169652
rect 213972 169632 213974 169652
rect 214010 168952 214066 169008
rect 213918 168292 213974 168328
rect 213918 168272 213920 168292
rect 213920 168272 213972 168292
rect 213972 168272 213974 168292
rect 214010 167592 214066 167648
rect 213918 166948 213920 166968
rect 213920 166948 213972 166968
rect 213972 166948 213974 166968
rect 213918 166912 213974 166948
rect 214102 166368 214158 166424
rect 214010 165688 214066 165744
rect 213918 165008 213974 165064
rect 214010 164328 214066 164384
rect 213918 163648 213974 163704
rect 214010 162968 214066 163024
rect 213918 162288 213974 162344
rect 204994 86128 205050 86184
rect 203614 82728 203670 82784
rect 214010 161744 214066 161800
rect 213918 161064 213974 161120
rect 214102 160656 214158 160712
rect 214010 160384 214066 160440
rect 213918 159704 213974 159760
rect 214102 159024 214158 159080
rect 213918 158344 213974 158400
rect 214010 157664 214066 157720
rect 213918 157120 213974 157176
rect 214010 156440 214066 156496
rect 213918 155796 213920 155816
rect 213920 155796 213972 155816
rect 213972 155796 213974 155816
rect 213918 155760 213974 155796
rect 214010 155080 214066 155136
rect 214010 154400 214066 154456
rect 213918 153720 213974 153776
rect 214010 153040 214066 153096
rect 214562 152496 214618 152552
rect 210514 119312 210570 119368
rect 209226 105168 209282 105224
rect 209134 91568 209190 91624
rect 213182 151816 213238 151872
rect 214010 151136 214066 151192
rect 213918 150492 213920 150512
rect 213920 150492 213972 150512
rect 213972 150492 213974 150512
rect 213918 150456 213974 150492
rect 214102 149096 214158 149152
rect 213918 148416 213974 148472
rect 213918 147872 213974 147928
rect 214010 147192 214066 147248
rect 213918 146512 213974 146568
rect 231950 240116 231952 240136
rect 231952 240116 232004 240136
rect 232004 240116 232006 240136
rect 231950 240080 232006 240116
rect 231214 237088 231270 237144
rect 232594 238448 232650 238504
rect 232962 234368 233018 234424
rect 231214 228928 231270 228984
rect 232962 228792 233018 228848
rect 231858 222128 231914 222184
rect 231122 219544 231178 219600
rect 230202 186224 230258 186280
rect 230662 184456 230718 184512
rect 229374 176976 229430 177032
rect 229374 175752 229430 175808
rect 229466 166096 229522 166152
rect 229190 155760 229246 155816
rect 229742 147872 229798 147928
rect 229098 146784 229154 146840
rect 215942 145832 215998 145888
rect 213918 145152 213974 145208
rect 214010 144472 214066 144528
rect 213918 143792 213974 143848
rect 213918 143248 213974 143304
rect 213918 141888 213974 141944
rect 214102 141208 214158 141264
rect 213918 140528 213974 140584
rect 214010 139848 214066 139904
rect 213918 138624 213974 138680
rect 214010 137944 214066 138000
rect 213366 136584 213422 136640
rect 213274 133864 213330 133920
rect 213182 119448 213238 119504
rect 210422 88984 210478 89040
rect 212446 94424 212502 94480
rect 211894 90344 211950 90400
rect 213918 135904 213974 135960
rect 213918 135260 213920 135280
rect 213920 135260 213972 135280
rect 213972 135260 213974 135280
rect 213918 135224 213974 135260
rect 213918 134544 213974 134600
rect 214838 139168 214894 139224
rect 214746 137264 214802 137320
rect 214010 133320 214066 133376
rect 213918 132640 213974 132696
rect 213918 131960 213974 132016
rect 214010 131280 214066 131336
rect 213918 130600 213974 130656
rect 214654 129920 214710 129976
rect 214562 129240 214618 129296
rect 213918 128696 213974 128752
rect 214010 128016 214066 128072
rect 213918 127336 213974 127392
rect 214010 126656 214066 126712
rect 213918 125976 213974 126032
rect 214010 125296 214066 125352
rect 213918 124616 213974 124672
rect 213918 124072 213974 124128
rect 214010 122712 214066 122768
rect 213918 122032 213974 122088
rect 214010 121352 214066 121408
rect 213918 120672 213974 120728
rect 214102 119992 214158 120048
rect 213918 119448 213974 119504
rect 214010 118788 214066 118824
rect 214010 118768 214012 118788
rect 214012 118768 214064 118788
rect 214064 118768 214066 118788
rect 214010 118088 214066 118144
rect 213918 117408 213974 117464
rect 214010 116728 214066 116784
rect 213918 116068 213974 116104
rect 213918 116048 213920 116068
rect 213920 116048 213972 116068
rect 213972 116048 213974 116068
rect 214010 115368 214066 115424
rect 213918 114824 213974 114880
rect 213918 114144 213974 114200
rect 214010 112784 214066 112840
rect 213918 112104 213974 112160
rect 214010 111424 214066 111480
rect 213918 110744 213974 110800
rect 214010 110200 214066 110256
rect 213918 109520 213974 109576
rect 214010 108840 214066 108896
rect 213918 108160 213974 108216
rect 214010 107480 214066 107536
rect 213918 106800 213974 106856
rect 214010 106120 214066 106176
rect 213918 104916 213974 104952
rect 213918 104896 213920 104916
rect 213920 104896 213972 104916
rect 213972 104896 213974 104916
rect 213918 104216 213974 104272
rect 213918 102856 213974 102912
rect 214010 102212 214012 102232
rect 214012 102212 214064 102232
rect 214064 102212 214066 102232
rect 214010 102176 214066 102212
rect 214010 101496 214066 101552
rect 213918 100952 213974 101008
rect 214102 100272 214158 100328
rect 214010 100000 214066 100056
rect 213918 99592 213974 99648
rect 213918 98232 213974 98288
rect 213918 97552 213974 97608
rect 213918 96328 213974 96384
rect 214654 96872 214710 96928
rect 213366 93744 213422 93800
rect 213182 22616 213238 22672
rect 216034 142568 216090 142624
rect 229834 145560 229890 145616
rect 229742 139168 229798 139224
rect 229742 135768 229798 135824
rect 216126 123392 216182 123448
rect 229098 97824 229154 97880
rect 229190 97144 229246 97200
rect 228362 95784 228418 95840
rect 225602 94424 225658 94480
rect 219346 93880 219402 93936
rect 222934 93200 222990 93256
rect 217230 87488 217286 87544
rect 198002 3984 198058 4040
rect 196622 3440 196678 3496
rect 177394 3304 177450 3360
rect 140042 2624 140098 2680
rect 142802 2624 142858 2680
rect 222934 64096 222990 64152
rect 226982 93880 227038 93936
rect 225694 79328 225750 79384
rect 230662 175616 230718 175672
rect 230570 169904 230626 169960
rect 230570 168952 230626 169008
rect 230754 172352 230810 172408
rect 233238 223524 233240 223544
rect 233240 223524 233292 223544
rect 233292 223524 233294 223544
rect 233238 223488 233294 223524
rect 231950 210976 232006 211032
rect 231122 185680 231178 185736
rect 231306 176024 231362 176080
rect 231306 175208 231362 175264
rect 231398 171808 231454 171864
rect 231306 171400 231362 171456
rect 231858 170448 231914 170504
rect 231122 168544 231178 168600
rect 230386 156576 230442 156632
rect 230570 153040 230626 153096
rect 230570 151544 230626 151600
rect 230386 148008 230442 148064
rect 230018 146240 230074 146296
rect 231030 163784 231086 163840
rect 230938 161880 230994 161936
rect 230846 157664 230902 157720
rect 231398 168036 231400 168056
rect 231400 168036 231452 168056
rect 231452 168036 231454 168056
rect 231398 168000 231454 168036
rect 231398 167084 231400 167104
rect 231400 167084 231452 167104
rect 231452 167084 231454 167104
rect 231398 167048 231454 167084
rect 231766 166676 231768 166696
rect 231768 166676 231820 166696
rect 231820 166676 231822 166696
rect 231766 166640 231822 166676
rect 231490 165180 231492 165200
rect 231492 165180 231544 165200
rect 231544 165180 231546 165200
rect 231490 165144 231546 165180
rect 231674 162832 231730 162888
rect 232042 164736 232098 164792
rect 231214 160520 231270 160576
rect 231398 159024 231454 159080
rect 231766 160012 231768 160032
rect 231768 160012 231820 160032
rect 231820 160012 231822 160032
rect 231766 159976 231822 160012
rect 231674 158616 231730 158672
rect 231214 158072 231270 158128
rect 231582 158072 231638 158128
rect 231490 155216 231546 155272
rect 231490 153312 231546 153368
rect 231490 152940 231492 152960
rect 231492 152940 231544 152960
rect 231544 152940 231546 152960
rect 231490 152904 231546 152940
rect 231674 157936 231730 157992
rect 231674 157120 231730 157176
rect 231766 156712 231822 156768
rect 231766 156168 231822 156224
rect 231674 154264 231730 154320
rect 231766 153856 231822 153912
rect 231582 151952 231638 152008
rect 231490 151000 231546 151056
rect 231766 151000 231822 151056
rect 231674 150592 231730 150648
rect 231490 148688 231546 148744
rect 231582 148280 231638 148336
rect 230754 139712 230810 139768
rect 229926 137808 229982 137864
rect 230570 135904 230626 135960
rect 229926 132776 229982 132832
rect 229834 106120 229890 106176
rect 230570 129784 230626 129840
rect 231122 142024 231178 142080
rect 231030 134408 231086 134464
rect 230846 133456 230902 133512
rect 230754 127336 230810 127392
rect 230570 126384 230626 126440
rect 230846 125976 230902 126032
rect 230018 123256 230074 123312
rect 229926 93880 229982 93936
rect 231766 148144 231822 148200
rect 233054 185000 233110 185056
rect 232226 174664 232282 174720
rect 236458 240080 236514 240136
rect 235906 238584 235962 238640
rect 237930 240080 237986 240136
rect 236826 227432 236882 227488
rect 236826 226888 236882 226944
rect 234986 224712 235042 224768
rect 237378 212472 237434 212528
rect 233514 194520 233570 194576
rect 232594 164872 232650 164928
rect 232502 159024 232558 159080
rect 231766 147056 231822 147112
rect 231674 144880 231730 144936
rect 231582 144336 231638 144392
rect 231766 143384 231822 143440
rect 231674 142976 231730 143032
rect 231766 140700 231768 140720
rect 231768 140700 231820 140720
rect 231820 140700 231822 140720
rect 231766 140664 231822 140700
rect 231490 138216 231546 138272
rect 231582 136856 231638 136912
rect 231490 135360 231546 135416
rect 231582 134000 231638 134056
rect 231766 133048 231822 133104
rect 231674 132504 231730 132560
rect 231306 131552 231362 131608
rect 231674 131144 231730 131200
rect 231214 130192 231270 130248
rect 231766 129240 231822 129296
rect 231674 128832 231730 128888
rect 231122 128288 231178 128344
rect 231766 127916 231768 127936
rect 231768 127916 231820 127936
rect 231820 127916 231822 127936
rect 231766 127880 231822 127916
rect 231122 127744 231178 127800
rect 230938 123120 230994 123176
rect 231306 127608 231362 127664
rect 231122 121624 231178 121680
rect 230754 120672 230810 120728
rect 230570 120264 230626 120320
rect 231214 119176 231270 119232
rect 230938 116456 230994 116512
rect 231122 116456 231178 116512
rect 230754 116048 230810 116104
rect 231030 114552 231086 114608
rect 230570 113192 230626 113248
rect 230570 110744 230626 110800
rect 230754 109792 230810 109848
rect 230662 101768 230718 101824
rect 230570 101360 230626 101416
rect 230662 100408 230718 100464
rect 230938 105168 230994 105224
rect 230938 104216 230994 104272
rect 231766 126948 231822 126984
rect 231766 126928 231768 126948
rect 231768 126928 231820 126948
rect 231820 126928 231822 126948
rect 231766 125024 231822 125080
rect 231490 124480 231546 124536
rect 231766 124108 231768 124128
rect 231768 124108 231820 124128
rect 231820 124108 231822 124128
rect 231766 124072 231822 124108
rect 231674 123528 231730 123584
rect 231766 122168 231822 122224
rect 231490 118904 231546 118960
rect 231398 117952 231454 118008
rect 231306 117136 231362 117192
rect 231214 115096 231270 115152
rect 231766 119992 231822 120048
rect 231766 119312 231822 119368
rect 233422 164328 233478 164384
rect 236090 191120 236146 191176
rect 234710 181600 234766 181656
rect 233974 154944 234030 155000
rect 232594 125432 232650 125488
rect 232778 124616 232834 124672
rect 232502 118360 232558 118416
rect 231766 117408 231822 117464
rect 231766 115504 231822 115560
rect 231582 113600 231638 113656
rect 232686 113464 232742 113520
rect 231766 112648 231822 112704
rect 232502 112376 232558 112432
rect 231674 112240 231730 112296
rect 231398 111288 231454 111344
rect 231766 109384 231822 109440
rect 231766 108432 231822 108488
rect 231490 107888 231546 107944
rect 231766 107072 231822 107128
rect 231490 106528 231546 106584
rect 231766 105576 231822 105632
rect 231306 103672 231362 103728
rect 231766 102720 231822 102776
rect 231490 102312 231546 102368
rect 231306 101496 231362 101552
rect 231122 98912 231178 98968
rect 230754 97552 230810 97608
rect 231122 97008 231178 97064
rect 230570 96600 230626 96656
rect 230478 96192 230534 96248
rect 230570 90888 230626 90944
rect 229742 76608 229798 76664
rect 231674 100816 231730 100872
rect 231674 100680 231730 100736
rect 231674 99864 231730 99920
rect 231766 99456 231822 99512
rect 233882 140664 233938 140720
rect 232686 54440 232742 54496
rect 234066 145424 234122 145480
rect 233974 105304 234030 105360
rect 234250 153720 234306 153776
rect 234802 180240 234858 180296
rect 235998 180104 236054 180160
rect 235446 175072 235502 175128
rect 235354 166368 235410 166424
rect 236182 175752 236238 175808
rect 236090 175208 236146 175264
rect 236182 167048 236238 167104
rect 234158 117816 234214 117872
rect 234066 103264 234122 103320
rect 235262 115912 235318 115968
rect 236642 128696 236698 128752
rect 235538 73888 235594 73944
rect 235262 58520 235318 58576
rect 239218 239944 239274 240000
rect 239402 235864 239458 235920
rect 239218 235592 239274 235648
rect 238022 117408 238078 117464
rect 236734 59880 236790 59936
rect 236642 36488 236698 36544
rect 241242 239400 241298 239456
rect 240690 235864 240746 235920
rect 239770 230424 239826 230480
rect 240138 213832 240194 213888
rect 238850 165688 238906 165744
rect 238114 105440 238170 105496
rect 238206 103944 238262 104000
rect 239402 137128 239458 137184
rect 241426 215872 241482 215928
rect 240874 213832 240930 213888
rect 240782 204040 240838 204096
rect 240230 186904 240286 186960
rect 240322 183096 240378 183152
rect 240230 175208 240286 175264
rect 239678 166232 239734 166288
rect 240414 177384 240470 177440
rect 240322 163376 240378 163432
rect 240966 170312 241022 170368
rect 239678 124752 239734 124808
rect 239586 116456 239642 116512
rect 240782 122032 240838 122088
rect 239494 66952 239550 67008
rect 242714 236952 242770 237008
rect 243542 238448 243598 238504
rect 242254 180104 242310 180160
rect 244554 270952 244610 271008
rect 244462 253816 244518 253872
rect 246026 297336 246082 297392
rect 245842 289040 245898 289096
rect 245934 283772 245936 283792
rect 245936 283772 245988 283792
rect 245988 283772 245990 283792
rect 245934 283736 245990 283772
rect 245750 281560 245806 281616
rect 245658 281016 245714 281072
rect 245658 280200 245714 280256
rect 245658 280064 245714 280120
rect 245474 253852 245476 253872
rect 245476 253852 245528 253872
rect 245528 253852 245530 253872
rect 245474 253816 245530 253852
rect 244646 253000 244702 253056
rect 245474 253000 245530 253056
rect 244462 247288 244518 247344
rect 245750 278840 245806 278896
rect 245750 277480 245806 277536
rect 245934 282376 245990 282432
rect 245934 279420 245936 279440
rect 245936 279420 245988 279440
rect 245988 279420 245990 279440
rect 245934 279384 245990 279420
rect 245842 275848 245898 275904
rect 246946 283192 247002 283248
rect 246118 276684 246174 276720
rect 246118 276664 246120 276684
rect 246120 276664 246172 276684
rect 246172 276664 246174 276684
rect 245934 274488 245990 274544
rect 245934 273672 245990 273728
rect 245842 272312 245898 272368
rect 246946 273128 247002 273184
rect 245750 270136 245806 270192
rect 245842 269592 245898 269648
rect 246210 267960 246266 268016
rect 245934 267416 245990 267472
rect 245934 266328 245990 266384
rect 246210 266192 246266 266248
rect 245934 265784 245990 265840
rect 246762 265240 246818 265296
rect 245842 263880 245898 263936
rect 245750 263064 245806 263120
rect 245934 262268 245990 262304
rect 245934 262248 245936 262268
rect 245936 262248 245988 262268
rect 245988 262248 245990 262268
rect 246394 260888 246450 260944
rect 245842 260072 245898 260128
rect 245934 259528 245990 259584
rect 245934 258712 245990 258768
rect 245842 258168 245898 258224
rect 245750 250280 245806 250336
rect 245658 246472 245714 246528
rect 245750 245928 245806 245984
rect 245658 245656 245714 245712
rect 245750 244568 245806 244624
rect 245658 240760 245714 240816
rect 244462 233144 244518 233200
rect 244186 192616 244242 192672
rect 243910 189080 243966 189136
rect 242346 173848 242402 173904
rect 242254 162832 242310 162888
rect 242162 143928 242218 143984
rect 241518 140120 241574 140176
rect 242162 136856 242218 136912
rect 241058 94424 241114 94480
rect 240874 77832 240930 77888
rect 242346 143928 242402 143984
rect 242438 142704 242494 142760
rect 243542 116048 243598 116104
rect 242438 104624 242494 104680
rect 242346 69672 242402 69728
rect 246026 257352 246082 257408
rect 245934 256536 245990 256592
rect 245934 254360 245990 254416
rect 245934 251640 245990 251696
rect 245934 249500 245936 249520
rect 245936 249500 245988 249520
rect 245988 249500 245990 249520
rect 245934 249464 245990 249500
rect 245934 248668 245990 248704
rect 245934 248648 245936 248668
rect 245936 248648 245988 248668
rect 245988 248648 245990 248668
rect 246946 248104 247002 248160
rect 246118 245656 246174 245712
rect 245934 240216 245990 240272
rect 246394 242392 246450 242448
rect 246302 241440 246358 241496
rect 245934 227568 245990 227624
rect 244462 166368 244518 166424
rect 244554 146920 244610 146976
rect 243910 127744 243966 127800
rect 245198 146920 245254 146976
rect 244922 91840 244978 91896
rect 243634 62872 243690 62928
rect 242898 9016 242954 9072
rect 239310 5616 239366 5672
rect 244094 7520 244150 7576
rect 245106 109384 245162 109440
rect 246026 197104 246082 197160
rect 246302 150456 246358 150512
rect 245658 136312 245714 136368
rect 245198 108840 245254 108896
rect 244922 5616 244978 5672
rect 246394 139440 246450 139496
rect 247130 273128 247186 273184
rect 247222 271496 247278 271552
rect 247130 264424 247186 264480
rect 247222 235592 247278 235648
rect 247038 153720 247094 153776
rect 246670 140664 246726 140720
rect 248602 249872 248658 249928
rect 250074 328616 250130 328672
rect 249982 295976 250038 296032
rect 249982 278724 250038 278760
rect 249982 278704 249984 278724
rect 249984 278704 250036 278724
rect 250036 278704 250038 278724
rect 248510 160928 248566 160984
rect 246486 102176 246542 102232
rect 248694 176024 248750 176080
rect 248602 147736 248658 147792
rect 247866 119176 247922 119232
rect 249154 135904 249210 135960
rect 249062 111696 249118 111752
rect 249062 99728 249118 99784
rect 247958 88984 248014 89040
rect 247866 74024 247922 74080
rect 248418 71168 248474 71224
rect 247590 3440 247646 3496
rect 249890 215056 249946 215112
rect 250718 171536 250774 171592
rect 249798 170312 249854 170368
rect 250442 160384 250498 160440
rect 249338 127608 249394 127664
rect 249338 110608 249394 110664
rect 250442 128968 250498 129024
rect 250626 148416 250682 148472
rect 249338 76472 249394 76528
rect 249246 61512 249302 61568
rect 250534 107888 250590 107944
rect 252558 358944 252614 359000
rect 251822 268776 251878 268832
rect 251362 217912 251418 217968
rect 253294 358944 253350 359000
rect 256698 375264 256754 375320
rect 255318 289992 255374 290048
rect 254030 261160 254086 261216
rect 251270 158072 251326 158128
rect 251178 148280 251234 148336
rect 250718 141480 250774 141536
rect 250626 107480 250682 107536
rect 253478 168408 253534 168464
rect 253202 161472 253258 161528
rect 251914 156440 251970 156496
rect 251822 120128 251878 120184
rect 250718 101496 250774 101552
rect 250626 76744 250682 76800
rect 251914 99592 251970 99648
rect 253294 131552 253350 131608
rect 253202 112104 253258 112160
rect 252006 69536 252062 69592
rect 253938 162424 253994 162480
rect 253386 100816 253442 100872
rect 254858 167592 254914 167648
rect 254766 142840 254822 142896
rect 253294 72528 253350 72584
rect 254858 131008 254914 131064
rect 254766 98640 254822 98696
rect 255594 280064 255650 280120
rect 255502 234232 255558 234288
rect 258722 376624 258778 376680
rect 258078 331200 258134 331256
rect 256882 300056 256938 300112
rect 256698 203496 256754 203552
rect 259458 366288 259514 366344
rect 259734 366288 259790 366344
rect 258722 297472 258778 297528
rect 258722 268368 258778 268424
rect 258262 266464 258318 266520
rect 259366 266464 259422 266520
rect 259366 264152 259422 264208
rect 259550 288496 259606 288552
rect 259734 287680 259790 287736
rect 260102 287272 260158 287328
rect 259642 239944 259698 240000
rect 260194 238448 260250 238504
rect 259458 215192 259514 215248
rect 260746 215192 260802 215248
rect 257342 174256 257398 174312
rect 255318 96464 255374 96520
rect 255870 96464 255926 96520
rect 254674 73752 254730 73808
rect 257618 172760 257674 172816
rect 257342 141344 257398 141400
rect 256054 106528 256110 106584
rect 256146 79600 256202 79656
rect 257526 149640 257582 149696
rect 257434 119992 257490 120048
rect 257342 68312 257398 68368
rect 257618 75248 257674 75304
rect 257434 55800 257490 55856
rect 256054 33904 256110 33960
rect 253202 22616 253258 22672
rect 252374 3304 252430 3360
rect 253938 22072 253994 22128
rect 253478 3440 253534 3496
rect 260102 167048 260158 167104
rect 258722 151952 258778 152008
rect 258722 110336 258778 110392
rect 262494 377440 262550 377496
rect 264978 348472 265034 348528
rect 264978 347792 265034 347848
rect 263598 343848 263654 343904
rect 264242 343848 264298 343904
rect 262218 291760 262274 291816
rect 262862 239400 262918 239456
rect 263598 235728 263654 235784
rect 262954 233008 263010 233064
rect 267002 301008 267058 301064
rect 266358 296112 266414 296168
rect 266266 283464 266322 283520
rect 266358 244196 266360 244216
rect 266360 244196 266412 244216
rect 266412 244196 266414 244216
rect 266358 244160 266414 244196
rect 266358 219136 266414 219192
rect 268382 285640 268438 285696
rect 269026 285640 269082 285696
rect 267830 266192 267886 266248
rect 269762 317464 269818 317520
rect 269026 266192 269082 266248
rect 269026 265512 269082 265568
rect 268474 229744 268530 229800
rect 268382 216280 268438 216336
rect 267830 195880 267886 195936
rect 268382 195880 268438 195936
rect 266266 190304 266322 190360
rect 266266 189760 266322 189816
rect 269026 216280 269082 216336
rect 269026 215872 269082 215928
rect 270038 266328 270094 266384
rect 270406 266328 270462 266384
rect 270038 224848 270094 224904
rect 270406 224848 270462 224904
rect 270406 224168 270462 224224
rect 269854 183096 269910 183152
rect 268474 180104 268530 180160
rect 264978 177248 265034 177304
rect 271142 288632 271198 288688
rect 272614 234368 272670 234424
rect 273994 200776 274050 200832
rect 281354 376624 281410 376680
rect 276754 294072 276810 294128
rect 273994 180240 274050 180296
rect 273258 179968 273314 180024
rect 271142 178744 271198 178800
rect 276018 178880 276074 178936
rect 273258 177248 273314 177304
rect 280894 374584 280950 374640
rect 279422 300872 279478 300928
rect 276754 177384 276810 177440
rect 279514 224168 279570 224224
rect 279422 211928 279478 211984
rect 279330 192480 279386 192536
rect 279238 182960 279294 183016
rect 264978 175616 265034 175672
rect 265622 175208 265678 175264
rect 264978 174800 265034 174856
rect 265070 174004 265126 174040
rect 265070 173984 265072 174004
rect 265072 173984 265124 174004
rect 265124 173984 265126 174004
rect 264242 173576 264298 173632
rect 260838 173304 260894 173360
rect 260378 162696 260434 162752
rect 260194 157936 260250 157992
rect 260286 155216 260342 155272
rect 259366 109112 259422 109168
rect 258906 65456 258962 65512
rect 262770 135904 262826 135960
rect 262770 135360 262826 135416
rect 260286 114416 260342 114472
rect 260470 112376 260526 112432
rect 260286 105712 260342 105768
rect 260286 62736 260342 62792
rect 262770 125024 262826 125080
rect 262770 124616 262826 124672
rect 262862 121352 262918 121408
rect 262862 118904 262918 118960
rect 262126 107752 262182 107808
rect 261574 80824 261630 80880
rect 261482 48864 261538 48920
rect 259458 28192 259514 28248
rect 260838 21256 260894 21312
rect 264978 172624 265034 172680
rect 265070 172216 265126 172272
rect 264978 171400 265034 171456
rect 265070 170992 265126 171048
rect 264978 170040 265034 170096
rect 265162 170448 265218 170504
rect 264978 169632 265034 169688
rect 265070 168816 265126 168872
rect 265070 167864 265126 167920
rect 264978 167456 265034 167512
rect 265254 169224 265310 169280
rect 265162 167592 265218 167648
rect 265070 166640 265126 166696
rect 264978 166232 265034 166288
rect 265254 166368 265310 166424
rect 265162 165824 265218 165880
rect 265070 165280 265126 165336
rect 264978 164872 265034 164928
rect 265162 165008 265218 165064
rect 265254 164464 265310 164520
rect 264978 164056 265034 164112
rect 265070 163648 265126 163704
rect 265162 163240 265218 163296
rect 264978 162288 265034 162344
rect 265070 161880 265126 161936
rect 265070 161064 265126 161120
rect 264978 160248 265034 160304
rect 265070 159704 265126 159760
rect 264978 158888 265034 158944
rect 265070 158480 265126 158536
rect 264978 158072 265034 158128
rect 264334 157392 264390 157448
rect 265254 162696 265310 162752
rect 265346 157664 265402 157720
rect 265162 157392 265218 157448
rect 265070 157120 265126 157176
rect 264978 156304 265034 156360
rect 265162 155896 265218 155952
rect 264978 154536 265034 154592
rect 265070 153720 265126 153776
rect 264978 153332 265034 153368
rect 264978 153312 264980 153332
rect 264980 153312 265032 153332
rect 265032 153312 265034 153332
rect 264978 152904 265034 152960
rect 265254 152496 265310 152552
rect 265070 151544 265126 151600
rect 264978 151136 265034 151192
rect 264978 149912 265034 149968
rect 265070 149504 265126 149560
rect 265070 148416 265126 148472
rect 265254 150728 265310 150784
rect 265162 148144 265218 148200
rect 264978 147736 265034 147792
rect 264978 147328 265034 147384
rect 265070 146396 265126 146432
rect 265070 146376 265072 146396
rect 265072 146376 265124 146396
rect 265124 146376 265126 146396
rect 265070 145968 265126 146024
rect 264978 145152 265034 145208
rect 280158 184320 280214 184376
rect 279514 182960 279570 183016
rect 279330 172216 279386 172272
rect 281354 307672 281410 307728
rect 280894 291080 280950 291136
rect 280986 287136 281042 287192
rect 280894 284552 280950 284608
rect 280894 182008 280950 182064
rect 280250 168680 280306 168736
rect 280158 162560 280214 162616
rect 265714 154128 265770 154184
rect 265254 146920 265310 146976
rect 265438 146920 265494 146976
rect 265162 145560 265218 145616
rect 264610 144744 264666 144800
rect 264426 140800 264482 140856
rect 264334 122712 264390 122768
rect 264242 119312 264298 119368
rect 263046 83408 263102 83464
rect 263598 17312 263654 17368
rect 264334 109928 264390 109984
rect 264978 143792 265034 143848
rect 264978 143384 265034 143440
rect 265438 142704 265494 142760
rect 265162 142568 265218 142624
rect 265070 141208 265126 141264
rect 264978 139168 265034 139224
rect 265622 142160 265678 142216
rect 265162 139984 265218 140040
rect 265346 139984 265402 140040
rect 265070 138624 265126 138680
rect 264978 137808 265034 137864
rect 265070 136584 265126 136640
rect 264978 135632 265034 135688
rect 264978 134000 265034 134056
rect 264978 132640 265034 132696
rect 264978 132232 265034 132288
rect 264978 131008 265034 131064
rect 265070 130464 265126 130520
rect 264978 129240 265034 129296
rect 264978 127472 265034 127528
rect 265162 129648 265218 129704
rect 265070 126520 265126 126576
rect 264978 125840 265034 125896
rect 279330 155896 279386 155952
rect 267094 148960 267150 149016
rect 265806 148552 265862 148608
rect 264978 124480 265034 124536
rect 264978 123664 265034 123720
rect 265622 122848 265678 122904
rect 264978 121896 265034 121952
rect 265070 121524 265072 121544
rect 265072 121524 265124 121544
rect 265124 121524 265126 121544
rect 265070 121488 265126 121524
rect 264978 121080 265034 121136
rect 265070 120672 265126 120728
rect 264978 119720 265034 119776
rect 264978 118496 265034 118552
rect 265070 117136 265126 117192
rect 264978 116728 265034 116784
rect 265070 115096 265126 115152
rect 264978 114572 265034 114608
rect 264978 114552 264980 114572
rect 264980 114552 265032 114572
rect 265032 114552 265034 114572
rect 265070 113736 265126 113792
rect 264978 113328 265034 113384
rect 264978 112512 265034 112568
rect 264978 111560 265034 111616
rect 265070 110336 265126 110392
rect 264978 108976 265034 109032
rect 265346 108568 265402 108624
rect 264978 107344 265034 107400
rect 264886 106392 264942 106448
rect 264978 105168 265034 105224
rect 264978 104352 265034 104408
rect 265070 103400 265126 103456
rect 264978 102584 265034 102640
rect 264978 101768 265034 101824
rect 265070 101224 265126 101280
rect 265070 99184 265126 99240
rect 264978 98640 265034 98696
rect 265070 97824 265126 97880
rect 264978 96600 265034 96656
rect 264978 96192 265034 96248
rect 267002 138216 267058 138272
rect 265806 127880 265862 127936
rect 265898 126248 265954 126304
rect 265990 111968 266046 112024
rect 265806 98776 265862 98832
rect 265990 98232 266046 98288
rect 265714 97416 265770 97472
rect 265622 84768 265678 84824
rect 265714 80688 265770 80744
rect 265990 79464 266046 79520
rect 279330 148280 279386 148336
rect 280066 148280 280122 148336
rect 283562 374040 283618 374096
rect 283562 360848 283618 360904
rect 281630 202272 281686 202328
rect 280986 166368 281042 166424
rect 280894 145832 280950 145888
rect 279422 144744 279478 144800
rect 267094 134408 267150 134464
rect 267186 124072 267242 124128
rect 281906 178880 281962 178936
rect 281722 175480 281778 175536
rect 281630 163240 281686 163296
rect 282182 173984 282238 174040
rect 282458 172488 282514 172544
rect 282274 170892 282276 170912
rect 282276 170892 282328 170912
rect 282328 170892 282330 170912
rect 282274 170856 282330 170892
rect 282826 169360 282882 169416
rect 282274 167864 282330 167920
rect 282826 165552 282882 165608
rect 283102 207712 283158 207768
rect 283010 182008 283066 182064
rect 281906 164872 281962 164928
rect 282826 164056 282882 164112
rect 282826 161744 282882 161800
rect 282826 161064 282882 161120
rect 281722 160248 281778 160304
rect 281906 159432 281962 159488
rect 282366 158752 282422 158808
rect 282826 157936 282882 157992
rect 281630 154944 281686 155000
rect 281630 154128 281686 154184
rect 281630 152632 281686 152688
rect 282182 153720 282238 153776
rect 281722 151816 281778 151872
rect 281630 151136 281686 151192
rect 281630 150356 281632 150376
rect 281632 150356 281684 150376
rect 281684 150356 281686 150376
rect 281630 150320 281686 150356
rect 281722 149640 281778 149696
rect 281814 148824 281870 148880
rect 281630 148008 281686 148064
rect 282090 141208 282146 141264
rect 284942 298288 284998 298344
rect 284298 198600 284354 198656
rect 283102 153448 283158 153504
rect 282826 147328 282882 147384
rect 282366 145016 282422 145072
rect 282826 142704 282882 142760
rect 282826 142044 282882 142080
rect 282826 142024 282828 142044
rect 282828 142024 282880 142044
rect 282880 142024 282882 142044
rect 282826 139712 282882 139768
rect 282826 138896 282882 138952
rect 282826 138216 282882 138272
rect 282826 137400 282882 137456
rect 282826 136604 282882 136640
rect 282826 136584 282828 136604
rect 282828 136584 282880 136604
rect 282880 136584 282882 136604
rect 282826 136312 282882 136368
rect 282458 134408 282514 134464
rect 282826 133592 282882 133648
rect 282734 132776 282790 132832
rect 282182 132096 282238 132152
rect 282826 131280 282882 131336
rect 282826 130600 282882 130656
rect 282734 129784 282790 129840
rect 281814 128968 281870 129024
rect 282826 128308 282882 128344
rect 282826 128288 282828 128308
rect 282828 128288 282880 128308
rect 282880 128288 282882 128308
rect 282734 127472 282790 127528
rect 282366 125976 282422 126032
rect 282826 125160 282882 125216
rect 282734 124480 282790 124536
rect 282826 123684 282882 123720
rect 282826 123664 282828 123684
rect 282828 123664 282880 123684
rect 282880 123664 282882 123684
rect 282090 122984 282146 123040
rect 282090 120672 282146 120728
rect 281538 119176 281594 119232
rect 267738 111152 267794 111208
rect 267646 100408 267702 100464
rect 267186 82048 267242 82104
rect 267094 65592 267150 65648
rect 282826 122168 282882 122224
rect 282826 121388 282828 121408
rect 282828 121388 282880 121408
rect 282880 121388 282882 121408
rect 282826 121352 282882 121388
rect 282826 119856 282882 119912
rect 282826 118360 282882 118416
rect 282734 117952 282790 118008
rect 282826 117544 282882 117600
rect 282826 116864 282882 116920
rect 282734 116048 282790 116104
rect 282826 115368 282882 115424
rect 282642 114552 282698 114608
rect 282826 113736 282882 113792
rect 282826 113092 282828 113112
rect 282828 113092 282880 113112
rect 282880 113092 282882 113112
rect 282826 113056 282882 113092
rect 282182 112240 282238 112296
rect 282090 111596 282092 111616
rect 282092 111596 282144 111616
rect 282144 111596 282146 111616
rect 282090 111560 282146 111596
rect 282826 110744 282882 110800
rect 281722 109928 281778 109984
rect 282642 109248 282698 109304
rect 281722 108432 281778 108488
rect 282826 107752 282882 107808
rect 282826 106956 282882 106992
rect 282826 106936 282828 106956
rect 282828 106936 282880 106956
rect 282880 106936 282882 106956
rect 282826 106120 282882 106176
rect 282826 105440 282882 105496
rect 282826 104624 282882 104680
rect 281538 103944 281594 104000
rect 282090 103128 282146 103184
rect 282274 101632 282330 101688
rect 281538 100816 281594 100872
rect 279330 100544 279386 100600
rect 279330 98096 279386 98152
rect 269118 92520 269174 92576
rect 267002 53080 267058 53136
rect 266358 37168 266414 37224
rect 264978 22616 265034 22672
rect 268382 43424 268438 43480
rect 268290 12960 268346 13016
rect 267738 3984 267794 4040
rect 270590 94968 270646 95024
rect 270498 93200 270554 93256
rect 269210 51720 269266 51776
rect 278778 95784 278834 95840
rect 278778 95104 278834 95160
rect 273258 91704 273314 91760
rect 269118 30912 269174 30968
rect 268474 10240 268530 10296
rect 268474 3984 268530 4040
rect 270774 11600 270830 11656
rect 276018 91024 276074 91080
rect 276754 91024 276810 91080
rect 281630 99340 281686 99376
rect 281630 99320 281632 99340
rect 281632 99320 281684 99340
rect 281684 99320 281686 99340
rect 285770 270544 285826 270600
rect 286046 270544 286102 270600
rect 285678 222944 285734 223000
rect 285034 215872 285090 215928
rect 285034 176840 285090 176896
rect 289634 375264 289690 375320
rect 287058 369824 287114 369880
rect 287702 369824 287758 369880
rect 285862 238312 285918 238368
rect 291198 219408 291254 219464
rect 289910 209072 289966 209128
rect 289818 153720 289874 153776
rect 290094 176704 290150 176760
rect 290646 117292 290702 117328
rect 290646 117272 290648 117292
rect 290648 117272 290700 117292
rect 290700 117272 290702 117292
rect 291474 195336 291530 195392
rect 295982 355408 296038 355464
rect 296810 296792 296866 296848
rect 294142 181328 294198 181384
rect 281998 97824 282054 97880
rect 281538 88168 281594 88224
rect 277398 87488 277454 87544
rect 276110 68176 276166 68232
rect 276110 67496 276166 67552
rect 277306 67496 277362 67552
rect 277122 3440 277178 3496
rect 280158 86128 280214 86184
rect 278778 37848 278834 37904
rect 280802 19896 280858 19952
rect 277306 3304 277362 3360
rect 281906 4800 281962 4856
rect 285678 93064 285734 93120
rect 289818 19896 289874 19952
rect 284298 3304 284354 3360
rect 285402 3304 285458 3360
rect 287794 3440 287850 3496
rect 296718 204992 296774 205048
rect 291382 3440 291438 3496
rect 293682 3440 293738 3496
rect 298742 295976 298798 296032
rect 298190 291216 298246 291272
rect 298098 216008 298154 216064
rect 299570 293936 299626 293992
rect 299478 241440 299534 241496
rect 298742 235728 298798 235784
rect 302238 342080 302294 342136
rect 302238 340856 302294 340912
rect 300122 200640 300178 200696
rect 302146 226888 302202 226944
rect 301042 187040 301098 187096
rect 307022 375264 307078 375320
rect 304538 374584 304594 374640
rect 304262 349016 304318 349072
rect 304262 348336 304318 348392
rect 303710 310392 303766 310448
rect 304262 310392 304318 310448
rect 303710 309712 303766 309768
rect 303618 211792 303674 211848
rect 302514 189760 302570 189816
rect 302330 117952 302386 118008
rect 305734 349016 305790 349072
rect 308402 364928 308458 364984
rect 307022 342080 307078 342136
rect 305734 206216 305790 206272
rect 302882 14456 302938 14512
rect 298466 4800 298522 4856
rect 300766 3440 300822 3496
rect 307758 66816 307814 66872
rect 309874 237088 309930 237144
rect 309874 220088 309930 220144
rect 312818 375264 312874 375320
rect 311898 369008 311954 369064
rect 311898 368464 311954 368520
rect 313278 355272 313334 355328
rect 313278 202136 313334 202192
rect 316038 184184 316094 184240
rect 316774 302232 316830 302288
rect 316682 190984 316738 191040
rect 318798 376896 318854 376952
rect 319626 376896 319682 376952
rect 320178 361664 320234 361720
rect 318798 352552 318854 352608
rect 317510 237224 317566 237280
rect 317510 199416 317566 199472
rect 317510 75112 317566 75168
rect 322202 308352 322258 308408
rect 325698 368600 325754 368656
rect 326342 368600 326398 368656
rect 324318 356768 324374 356824
rect 322938 193840 322994 193896
rect 317326 3304 317382 3360
rect 324318 188264 324374 188320
rect 327078 353368 327134 353424
rect 328458 363024 328514 363080
rect 329102 363024 329158 363080
rect 331862 324944 331918 325000
rect 326342 6840 326398 6896
rect 326802 6840 326858 6896
rect 330390 3304 330446 3360
rect 333978 345072 334034 345128
rect 332598 311072 332654 311128
rect 332598 185544 332654 185600
rect 340234 375944 340290 376000
rect 338762 362208 338818 362264
rect 335358 209752 335414 209808
rect 342350 374584 342406 374640
rect 346122 375264 346178 375320
rect 349158 375264 349214 375320
rect 347042 349696 347098 349752
rect 345018 312432 345074 312488
rect 342350 235864 342406 235920
rect 340970 208936 341026 208992
rect 338854 185544 338910 185600
rect 338762 18536 338818 18592
rect 342902 206352 342958 206408
rect 342258 72392 342314 72448
rect 342994 3984 343050 4040
rect 352562 375264 352618 375320
rect 351090 374720 351146 374776
rect 354126 377440 354182 377496
rect 353298 361528 353354 361584
rect 351918 195200 351974 195256
rect 346950 3984 347006 4040
rect 354678 376352 354734 376408
rect 354678 373224 354734 373280
rect 354126 367648 354182 367704
rect 356242 492632 356298 492688
rect 358082 497800 358138 497856
rect 357162 495488 357218 495544
rect 356610 490320 356666 490376
rect 357438 482840 357494 482896
rect 356794 465704 356850 465760
rect 358634 493040 358690 493096
rect 358726 487736 358782 487792
rect 358726 485288 358782 485344
rect 358726 477944 358782 478000
rect 358726 475496 358782 475552
rect 358726 473048 358782 473104
rect 358726 470620 358782 470656
rect 358726 470600 358728 470620
rect 358728 470600 358780 470620
rect 358780 470600 358782 470620
rect 358726 468152 358782 468208
rect 358726 463256 358782 463312
rect 358450 460808 358506 460864
rect 358726 455912 358782 455968
rect 358726 453464 358782 453520
rect 358726 451016 358782 451072
rect 358726 448588 358782 448624
rect 358726 448568 358728 448588
rect 358728 448568 358780 448588
rect 358780 448568 358782 448588
rect 357530 446120 357586 446176
rect 358726 443672 358782 443728
rect 358726 441224 358782 441280
rect 358726 438932 358782 438968
rect 358726 438912 358728 438932
rect 358728 438912 358780 438932
rect 358780 438912 358782 438932
rect 358726 436328 358782 436384
rect 358726 433880 358782 433936
rect 358726 431432 358782 431488
rect 358726 428984 358782 429040
rect 357530 426536 357586 426592
rect 358726 424088 358782 424144
rect 358726 421640 358782 421696
rect 358726 419192 358782 419248
rect 357622 416744 357678 416800
rect 358726 414296 358782 414352
rect 358726 411848 358782 411904
rect 358726 409400 358782 409456
rect 358726 404232 358782 404288
rect 358726 401784 358782 401840
rect 357990 399336 358046 399392
rect 358726 396888 358782 396944
rect 357714 391992 357770 392048
rect 358818 382336 358874 382392
rect 357898 379752 357954 379808
rect 358358 377984 358414 378040
rect 358818 374720 358874 374776
rect 359002 406952 359058 407008
rect 359002 377440 359058 377496
rect 363602 542952 363658 543008
rect 361578 538328 361634 538384
rect 360382 535472 360438 535528
rect 360474 348472 360530 348528
rect 361854 373904 361910 373960
rect 361762 346976 361818 347032
rect 374090 539552 374146 539608
rect 371238 538192 371294 538248
rect 364614 345616 364670 345672
rect 360290 182824 360346 182880
rect 367374 377304 367430 377360
rect 370134 369008 370190 369064
rect 370042 365608 370098 365664
rect 371422 335960 371478 336016
rect 371238 184184 371294 184240
rect 374642 376488 374698 376544
rect 375562 351056 375618 351112
rect 375470 207576 375526 207632
rect 381542 284416 381598 284472
rect 380898 219272 380954 219328
rect 382922 374584 382978 374640
rect 582470 697176 582526 697232
rect 582378 564304 582434 564360
rect 580170 537784 580226 537840
rect 582378 524456 582434 524512
rect 582378 511264 582434 511320
rect 580262 484608 580318 484664
rect 582562 683848 582618 683904
rect 583206 670656 583262 670712
rect 582746 644000 582802 644056
rect 582654 577632 582710 577688
rect 582378 418240 582434 418296
rect 582378 378392 582434 378448
rect 583022 630808 583078 630864
rect 582930 590960 582986 591016
rect 583114 617480 583170 617536
rect 583114 541592 583170 541648
rect 582930 471416 582986 471472
rect 582838 458088 582894 458144
rect 582838 431568 582894 431624
rect 582746 404912 582802 404968
rect 582654 376896 582710 376952
rect 583206 376624 583262 376680
rect 582378 365064 582434 365120
rect 580170 351872 580226 351928
rect 582378 342896 582434 342952
rect 580722 298696 580778 298752
rect 580722 296656 580778 296712
rect 579802 272176 579858 272232
rect 580262 261432 580318 261488
rect 580170 258848 580226 258904
rect 580170 245520 580226 245576
rect 574742 234504 574798 234560
rect 574742 228248 574798 228304
rect 385038 6840 385094 6896
rect 580262 179152 580318 179208
rect 580170 165824 580226 165880
rect 582930 325216 582986 325272
rect 582654 292576 582710 292632
rect 582654 192480 582710 192536
rect 582562 72936 582618 72992
rect 583022 312024 583078 312080
rect 583574 287680 583630 287736
rect 583206 284280 583262 284336
rect 583022 264152 583078 264208
rect 582930 231104 582986 231160
rect 582838 112784 582894 112840
rect 583206 219000 583262 219056
rect 583482 265512 583538 265568
rect 583482 232872 583538 232928
rect 583482 213152 583538 213208
rect 583390 152632 583446 152688
rect 583298 139304 583354 139360
rect 583114 125976 583170 126032
rect 583022 99456 583078 99512
rect 582930 59608 582986 59664
rect 582746 46280 582802 46336
rect 583390 33108 583446 33144
rect 583390 33088 583392 33108
rect 583392 33088 583444 33108
rect 583444 33088 583446 33108
rect 582470 19760 582526 19816
rect 580170 6568 580226 6624
rect 353298 3304 353354 3360
rect 583758 225528 583814 225584
rect 583666 222808 583722 222864
rect 583574 206216 583630 206272
rect 583574 204856 583630 204912
rect 583758 86672 583814 86728
<< metal3 >>
rect 69606 702476 69612 702540
rect 69676 702538 69682 702540
rect 154113 702538 154179 702541
rect 69676 702536 154179 702538
rect 69676 702480 154118 702536
rect 154174 702480 154179 702536
rect 69676 702478 154179 702480
rect 69676 702476 69682 702478
rect 154113 702475 154179 702478
rect -960 697220 480 697460
rect 582465 697234 582531 697237
rect 583520 697234 584960 697324
rect 582465 697232 584960 697234
rect 582465 697176 582470 697232
rect 582526 697176 584960 697232
rect 582465 697174 584960 697176
rect 582465 697171 582531 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 3417 684314 3483 684317
rect -960 684312 3483 684314
rect -960 684256 3422 684312
rect 3478 684256 3483 684312
rect -960 684254 3483 684256
rect -960 684164 480 684254
rect 3417 684251 3483 684254
rect 582557 683906 582623 683909
rect 583520 683906 584960 683996
rect 582557 683904 584960 683906
rect 582557 683848 582562 683904
rect 582618 683848 584960 683904
rect 582557 683846 584960 683848
rect 582557 683843 582623 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3509 671258 3575 671261
rect -960 671256 3575 671258
rect -960 671200 3514 671256
rect 3570 671200 3575 671256
rect -960 671198 3575 671200
rect -960 671108 480 671198
rect 3509 671195 3575 671198
rect 583201 670714 583267 670717
rect 583520 670714 584960 670804
rect 583201 670712 584960 670714
rect 583201 670656 583206 670712
rect 583262 670656 584960 670712
rect 583201 670654 584960 670656
rect 583201 670651 583267 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 3417 658202 3483 658205
rect -960 658200 3483 658202
rect -960 658144 3422 658200
rect 3478 658144 3483 658200
rect -960 658142 3483 658144
rect -960 658052 480 658142
rect 3417 658139 3483 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 582741 644058 582807 644061
rect 583520 644058 584960 644148
rect 582741 644056 584960 644058
rect 582741 644000 582746 644056
rect 582802 644000 584960 644056
rect 582741 643998 584960 644000
rect 582741 643995 582807 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 3417 632090 3483 632093
rect -960 632088 3483 632090
rect -960 632032 3422 632088
rect 3478 632032 3483 632088
rect -960 632030 3483 632032
rect -960 631940 480 632030
rect 3417 632027 3483 632030
rect 583017 630866 583083 630869
rect 583520 630866 584960 630956
rect 583017 630864 584960 630866
rect 583017 630808 583022 630864
rect 583078 630808 584960 630864
rect 583017 630806 584960 630808
rect 583017 630803 583083 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 3141 619170 3207 619173
rect -960 619168 3207 619170
rect -960 619112 3146 619168
rect 3202 619112 3207 619168
rect -960 619110 3207 619112
rect -960 619020 480 619110
rect 3141 619107 3207 619110
rect 583109 617538 583175 617541
rect 583520 617538 584960 617628
rect 583109 617536 584960 617538
rect 583109 617480 583114 617536
rect 583170 617480 584960 617536
rect 583109 617478 584960 617480
rect 583109 617475 583175 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 3233 606114 3299 606117
rect -960 606112 3299 606114
rect -960 606056 3238 606112
rect 3294 606056 3299 606112
rect -960 606054 3299 606056
rect -960 605964 480 606054
rect 3233 606051 3299 606054
rect 583520 604060 584960 604300
rect 72877 595506 72943 595509
rect 87597 595506 87663 595509
rect 72877 595504 87663 595506
rect 72877 595448 72882 595504
rect 72938 595448 87602 595504
rect 87658 595448 87663 595504
rect 72877 595446 87663 595448
rect 72877 595443 72943 595446
rect 87597 595443 87663 595446
rect -960 592908 480 593148
rect 78581 592106 78647 592109
rect 103513 592106 103579 592109
rect 78581 592104 103579 592106
rect 78581 592048 78586 592104
rect 78642 592048 103518 592104
rect 103574 592048 103579 592104
rect 78581 592046 103579 592048
rect 78581 592043 78647 592046
rect 103513 592043 103579 592046
rect 83181 591018 83247 591021
rect 100753 591018 100819 591021
rect 83181 591016 100819 591018
rect 83181 590960 83186 591016
rect 83242 590960 100758 591016
rect 100814 590960 100819 591016
rect 83181 590958 100819 590960
rect 83181 590955 83247 590958
rect 100753 590955 100819 590958
rect 582925 591018 582991 591021
rect 583520 591018 584960 591108
rect 582925 591016 584960 591018
rect 582925 590960 582930 591016
rect 582986 590960 584960 591016
rect 582925 590958 584960 590960
rect 582925 590955 582991 590958
rect 583520 590868 584960 590958
rect 66069 590746 66135 590749
rect 70301 590746 70367 590749
rect 71129 590746 71195 590749
rect 66069 590744 71195 590746
rect 66069 590688 66074 590744
rect 66130 590688 70306 590744
rect 70362 590688 71134 590744
rect 71190 590688 71195 590744
rect 66069 590686 71195 590688
rect 66069 590683 66135 590686
rect 70301 590683 70367 590686
rect 71129 590683 71195 590686
rect 82261 590746 82327 590749
rect 88006 590746 88012 590748
rect 82261 590744 88012 590746
rect 82261 590688 82266 590744
rect 82322 590688 88012 590744
rect 82261 590686 88012 590688
rect 82261 590683 82327 590686
rect 88006 590684 88012 590686
rect 88076 590684 88082 590748
rect 73153 589930 73219 589933
rect 90357 589930 90423 589933
rect 73153 589928 90423 589930
rect 73153 589872 73158 589928
rect 73214 589872 90362 589928
rect 90418 589872 90423 589928
rect 73153 589870 90423 589872
rect 73153 589867 73219 589870
rect 90357 589867 90423 589870
rect 77661 589522 77727 589525
rect 100845 589522 100911 589525
rect 77661 589520 100911 589522
rect 77661 589464 77666 589520
rect 77722 589464 100850 589520
rect 100906 589464 100911 589520
rect 77661 589462 100911 589464
rect 77661 589459 77727 589462
rect 100845 589459 100911 589462
rect 81341 589386 81407 589389
rect 93761 589386 93827 589389
rect 187601 589386 187667 589389
rect 81341 589384 187667 589386
rect 81341 589328 81346 589384
rect 81402 589328 93766 589384
rect 93822 589328 187606 589384
rect 187662 589328 187667 589384
rect 81341 589326 187667 589328
rect 81341 589323 81407 589326
rect 93761 589323 93827 589326
rect 187601 589323 187667 589326
rect 81709 588706 81775 588709
rect 93894 588706 93900 588708
rect 81709 588704 93900 588706
rect 81709 588648 81714 588704
rect 81770 588648 93900 588704
rect 81709 588646 93900 588648
rect 81709 588643 81775 588646
rect 93894 588644 93900 588646
rect 93964 588644 93970 588708
rect 88057 588570 88123 588573
rect 88190 588570 88196 588572
rect 88057 588568 88196 588570
rect 88057 588512 88062 588568
rect 88118 588512 88196 588568
rect 88057 588510 88196 588512
rect 88057 588507 88123 588510
rect 88190 588508 88196 588510
rect 88260 588508 88266 588572
rect 66805 588434 66871 588437
rect 66805 588432 68908 588434
rect 66805 588376 66810 588432
rect 66866 588376 68908 588432
rect 66805 588374 68908 588376
rect 66805 588371 66871 588374
rect 91737 587618 91803 587621
rect 88596 587616 91803 587618
rect 88596 587560 91742 587616
rect 91798 587560 91803 587616
rect 88596 587558 91803 587560
rect 91737 587555 91803 587558
rect 66253 586530 66319 586533
rect 66253 586528 66362 586530
rect 66253 586472 66258 586528
rect 66314 586472 66362 586528
rect 66253 586467 66362 586472
rect 66302 586394 66362 586467
rect 68878 586394 68938 587044
rect 66302 586334 68938 586394
rect 89713 586258 89779 586261
rect 88596 586256 89779 586258
rect 88596 586200 89718 586256
rect 89774 586200 89779 586256
rect 88596 586198 89779 586200
rect 89713 586195 89779 586198
rect 66805 585714 66871 585717
rect 66805 585712 68908 585714
rect 66805 585656 66810 585712
rect 66866 585656 68908 585712
rect 66805 585654 68908 585656
rect 66805 585651 66871 585654
rect 88190 585652 88196 585716
rect 88260 585714 88266 585716
rect 118693 585714 118759 585717
rect 88260 585712 118759 585714
rect 88260 585656 118698 585712
rect 118754 585656 118759 585712
rect 88260 585654 118759 585656
rect 88260 585652 88266 585654
rect 118693 585651 118759 585654
rect 91369 584898 91435 584901
rect 88596 584896 91435 584898
rect 88596 584840 91374 584896
rect 91430 584840 91435 584896
rect 88596 584838 91435 584840
rect 91369 584835 91435 584838
rect 67633 584354 67699 584357
rect 67633 584352 68908 584354
rect 67633 584296 67638 584352
rect 67694 584296 68908 584352
rect 67633 584294 68908 584296
rect 67633 584291 67699 584294
rect 91185 583674 91251 583677
rect 88596 583672 91251 583674
rect 88596 583616 91190 583672
rect 91246 583616 91251 583672
rect 88596 583614 91251 583616
rect 91185 583611 91251 583614
rect 66805 582994 66871 582997
rect 109033 582994 109099 582997
rect 66805 582992 68908 582994
rect 66805 582936 66810 582992
rect 66866 582936 68908 582992
rect 66805 582934 68908 582936
rect 89670 582992 109099 582994
rect 89670 582936 109038 582992
rect 109094 582936 109099 582992
rect 89670 582934 109099 582936
rect 66805 582931 66871 582934
rect 88190 582796 88196 582860
rect 88260 582858 88266 582860
rect 89670 582858 89730 582934
rect 109033 582931 109099 582934
rect 88260 582798 89730 582858
rect 88260 582796 88266 582798
rect 69422 582252 69428 582316
rect 69492 582252 69498 582316
rect 66437 581770 66503 581773
rect 69430 581770 69490 582252
rect 91737 582178 91803 582181
rect 88596 582176 91803 582178
rect 88596 582120 91742 582176
rect 91798 582120 91803 582176
rect 88596 582118 91803 582120
rect 91737 582115 91803 582118
rect 66437 581768 69490 581770
rect 66437 581712 66442 581768
rect 66498 581740 69490 581768
rect 66498 581712 69460 581740
rect 66437 581710 69460 581712
rect 66437 581707 66503 581710
rect 91737 580818 91803 580821
rect 88596 580816 91803 580818
rect 88596 580760 91742 580816
rect 91798 580760 91803 580816
rect 88596 580758 91803 580760
rect 91737 580755 91803 580758
rect 66805 580274 66871 580277
rect 66805 580272 68908 580274
rect 66805 580216 66810 580272
rect 66866 580216 68908 580272
rect 66805 580214 68908 580216
rect 66805 580211 66871 580214
rect -960 580002 480 580092
rect 3417 580002 3483 580005
rect -960 580000 3483 580002
rect -960 579944 3422 580000
rect 3478 579944 3483 580000
rect -960 579942 3483 579944
rect -960 579852 480 579942
rect 3417 579939 3483 579942
rect 91737 579458 91803 579461
rect 88596 579456 91803 579458
rect 88596 579400 91742 579456
rect 91798 579400 91803 579456
rect 88596 579398 91803 579400
rect 91737 579395 91803 579398
rect 67725 578914 67791 578917
rect 67725 578912 68908 578914
rect 67725 578856 67730 578912
rect 67786 578856 68908 578912
rect 67725 578854 68908 578856
rect 67725 578851 67791 578854
rect 91502 578098 91508 578100
rect 88596 578038 91508 578098
rect 91502 578036 91508 578038
rect 91572 578036 91578 578100
rect 582649 577690 582715 577693
rect 583520 577690 584960 577780
rect 582649 577688 584960 577690
rect 582649 577632 582654 577688
rect 582710 577632 584960 577688
rect 582649 577630 584960 577632
rect 582649 577627 582715 577630
rect 67265 577554 67331 577557
rect 88885 577554 88951 577557
rect 124254 577554 124260 577556
rect 67265 577552 68908 577554
rect 67265 577496 67270 577552
rect 67326 577496 68908 577552
rect 67265 577494 68908 577496
rect 88885 577552 124260 577554
rect 88885 577496 88890 577552
rect 88946 577496 124260 577552
rect 88885 577494 124260 577496
rect 67265 577491 67331 577494
rect 88885 577491 88951 577494
rect 124254 577492 124260 577494
rect 124324 577492 124330 577556
rect 583520 577540 584960 577630
rect 91093 576738 91159 576741
rect 88596 576736 91159 576738
rect 88596 576680 91098 576736
rect 91154 576680 91159 576736
rect 88596 576678 91159 576680
rect 91093 576675 91159 576678
rect 67357 576194 67423 576197
rect 67357 576192 68908 576194
rect 67357 576136 67362 576192
rect 67418 576136 68908 576192
rect 67357 576134 68908 576136
rect 67357 576131 67423 576134
rect 91093 575378 91159 575381
rect 88596 575376 91159 575378
rect 88596 575320 91098 575376
rect 91154 575320 91159 575376
rect 88596 575318 91159 575320
rect 91093 575315 91159 575318
rect 67081 574834 67147 574837
rect 67541 574834 67607 574837
rect 67081 574832 68908 574834
rect 67081 574776 67086 574832
rect 67142 574776 67546 574832
rect 67602 574776 68908 574832
rect 67081 574774 68908 574776
rect 67081 574771 67147 574774
rect 67541 574771 67607 574774
rect 65885 573474 65951 573477
rect 65885 573472 68908 573474
rect 65885 573416 65890 573472
rect 65946 573416 68908 573472
rect 65885 573414 68908 573416
rect 65885 573411 65951 573414
rect 88566 573338 88626 573988
rect 88566 573278 93870 573338
rect 93810 572794 93870 573278
rect 121678 572794 121684 572796
rect 93810 572734 121684 572794
rect 121678 572732 121684 572734
rect 121748 572732 121754 572796
rect 91093 572658 91159 572661
rect 88596 572656 91159 572658
rect 88596 572600 91098 572656
rect 91154 572600 91159 572656
rect 88596 572598 91159 572600
rect 91093 572595 91159 572598
rect 66805 572114 66871 572117
rect 66805 572112 68908 572114
rect 66805 572056 66810 572112
rect 66866 572056 68908 572112
rect 66805 572054 68908 572056
rect 66805 572051 66871 572054
rect 91185 571434 91251 571437
rect 88596 571432 91251 571434
rect 88596 571376 91190 571432
rect 91246 571376 91251 571432
rect 88596 571374 91251 571376
rect 91185 571371 91251 571374
rect 67173 570754 67239 570757
rect 67173 570752 68908 570754
rect 67173 570696 67178 570752
rect 67234 570696 68908 570752
rect 67173 570694 68908 570696
rect 67173 570691 67239 570694
rect 91093 570074 91159 570077
rect 88596 570072 91159 570074
rect 88596 570016 91098 570072
rect 91154 570016 91159 570072
rect 88596 570014 91159 570016
rect 91093 570011 91159 570014
rect 66805 569394 66871 569397
rect 66805 569392 68908 569394
rect 66805 569336 66810 569392
rect 66866 569336 68908 569392
rect 66805 569334 68908 569336
rect 66805 569331 66871 569334
rect 91093 568714 91159 568717
rect 88596 568712 91159 568714
rect 88596 568656 91098 568712
rect 91154 568656 91159 568712
rect 88596 568654 91159 568656
rect 91093 568651 91159 568654
rect 66713 568034 66779 568037
rect 66713 568032 68908 568034
rect 66713 567976 66718 568032
rect 66774 567976 68908 568032
rect 66713 567974 68908 567976
rect 66713 567971 66779 567974
rect 89805 567354 89871 567357
rect 88596 567352 89871 567354
rect 88596 567296 89810 567352
rect 89866 567296 89871 567352
rect 88596 567294 89871 567296
rect 89805 567291 89871 567294
rect -960 566946 480 567036
rect 3417 566946 3483 566949
rect -960 566944 3483 566946
rect -960 566888 3422 566944
rect 3478 566888 3483 566944
rect -960 566886 3483 566888
rect -960 566796 480 566886
rect 3417 566883 3483 566886
rect 67449 566810 67515 566813
rect 67449 566808 68908 566810
rect 67449 566752 67454 566808
rect 67510 566752 68908 566808
rect 67449 566750 68908 566752
rect 67449 566747 67515 566750
rect 91369 565858 91435 565861
rect 88596 565856 91435 565858
rect 88596 565800 91374 565856
rect 91430 565800 91435 565856
rect 88596 565798 91435 565800
rect 91369 565795 91435 565798
rect 66805 565042 66871 565045
rect 66805 565040 68908 565042
rect 66805 564984 66810 565040
rect 66866 564984 68908 565040
rect 66805 564982 68908 564984
rect 66805 564979 66871 564982
rect 91369 564498 91435 564501
rect 88596 564496 91435 564498
rect 88596 564440 91374 564496
rect 91430 564440 91435 564496
rect 88596 564438 91435 564440
rect 91369 564435 91435 564438
rect 582373 564362 582439 564365
rect 583520 564362 584960 564452
rect 582373 564360 584960 564362
rect 582373 564304 582378 564360
rect 582434 564304 584960 564360
rect 582373 564302 584960 564304
rect 582373 564299 582439 564302
rect 583520 564212 584960 564302
rect 66805 563682 66871 563685
rect 66805 563680 68908 563682
rect 66805 563624 66810 563680
rect 66866 563624 68908 563680
rect 66805 563622 68908 563624
rect 66805 563619 66871 563622
rect 91369 563138 91435 563141
rect 88596 563136 91435 563138
rect 88596 563080 91374 563136
rect 91430 563080 91435 563136
rect 88596 563078 91435 563080
rect 91369 563075 91435 563078
rect 66805 562322 66871 562325
rect 66805 562320 68908 562322
rect 66805 562264 66810 562320
rect 66866 562264 68908 562320
rect 66805 562262 68908 562264
rect 66805 562259 66871 562262
rect 91093 561506 91159 561509
rect 88596 561504 91159 561506
rect 88596 561448 91098 561504
rect 91154 561448 91159 561504
rect 88596 561446 91159 561448
rect 91093 561443 91159 561446
rect 66805 560962 66871 560965
rect 66805 560960 68908 560962
rect 66805 560904 66810 560960
rect 66866 560904 68908 560960
rect 66805 560902 68908 560904
rect 66805 560899 66871 560902
rect 88885 560146 88951 560149
rect 89621 560146 89687 560149
rect 88596 560144 89687 560146
rect 88596 560088 88890 560144
rect 88946 560088 89626 560144
rect 89682 560088 89687 560144
rect 88596 560086 89687 560088
rect 88885 560083 88951 560086
rect 89621 560083 89687 560086
rect 66805 559602 66871 559605
rect 134701 559602 134767 559605
rect 193213 559602 193279 559605
rect 66805 559600 68908 559602
rect 66805 559544 66810 559600
rect 66866 559544 68908 559600
rect 66805 559542 68908 559544
rect 134701 559600 193279 559602
rect 134701 559544 134706 559600
rect 134762 559544 193218 559600
rect 193274 559544 193279 559600
rect 134701 559542 193279 559544
rect 66805 559539 66871 559542
rect 134701 559539 134767 559542
rect 193213 559539 193279 559542
rect 193213 559058 193279 559061
rect 241513 559058 241579 559061
rect 193213 559056 241579 559058
rect 193213 559000 193218 559056
rect 193274 559000 241518 559056
rect 241574 559000 241579 559056
rect 193213 558998 241579 559000
rect 193213 558995 193279 558998
rect 241513 558995 241579 558998
rect 92381 558786 92447 558789
rect 88596 558784 92447 558786
rect 88596 558728 92386 558784
rect 92442 558728 92447 558784
rect 88596 558726 92447 558728
rect 92381 558723 92447 558726
rect 66805 558242 66871 558245
rect 66805 558240 68908 558242
rect 66805 558184 66810 558240
rect 66866 558184 68908 558240
rect 66805 558182 68908 558184
rect 66805 558179 66871 558182
rect 177941 557562 178007 557565
rect 237373 557562 237439 557565
rect 177941 557560 237439 557562
rect 177941 557504 177946 557560
rect 178002 557504 237378 557560
rect 237434 557504 237439 557560
rect 177941 557502 237439 557504
rect 177941 557499 178007 557502
rect 237373 557499 237439 557502
rect 91185 557426 91251 557429
rect 88596 557424 91251 557426
rect 88596 557368 91190 557424
rect 91246 557368 91251 557424
rect 88596 557366 91251 557368
rect 91185 557363 91251 557366
rect 67398 556820 67404 556884
rect 67468 556882 67474 556884
rect 67468 556822 68908 556882
rect 67468 556820 67474 556822
rect 184381 556202 184447 556205
rect 230473 556202 230539 556205
rect 184381 556200 230539 556202
rect 184381 556144 184386 556200
rect 184442 556144 230478 556200
rect 230534 556144 230539 556200
rect 184381 556142 230539 556144
rect 184381 556139 184447 556142
rect 230473 556139 230539 556142
rect 91737 556066 91803 556069
rect 88596 556064 91803 556066
rect 88596 556008 91742 556064
rect 91798 556008 91803 556064
rect 88596 556006 91803 556008
rect 91737 556003 91803 556006
rect 66805 555522 66871 555525
rect 66805 555520 68908 555522
rect 66805 555464 66810 555520
rect 66866 555464 68908 555520
rect 66805 555462 68908 555464
rect 66805 555459 66871 555462
rect 187509 554842 187575 554845
rect 240225 554842 240291 554845
rect 187509 554840 240291 554842
rect 187509 554784 187514 554840
rect 187570 554784 240230 554840
rect 240286 554784 240291 554840
rect 187509 554782 240291 554784
rect 187509 554779 187575 554782
rect 240225 554779 240291 554782
rect 91737 554706 91803 554709
rect 88596 554704 91803 554706
rect 88596 554648 91742 554704
rect 91798 554648 91803 554704
rect 88596 554646 91803 554648
rect 91737 554643 91803 554646
rect 66529 554162 66595 554165
rect 66529 554160 68908 554162
rect 66529 554104 66534 554160
rect 66590 554104 68908 554160
rect 66529 554102 68908 554104
rect 66529 554099 66595 554102
rect -960 553890 480 553980
rect 3417 553890 3483 553893
rect -960 553888 3483 553890
rect -960 553832 3422 553888
rect 3478 553832 3483 553888
rect -960 553830 3483 553832
rect -960 553740 480 553830
rect 3417 553827 3483 553830
rect 117957 553482 118023 553485
rect 118601 553482 118667 553485
rect 212533 553482 212599 553485
rect 117957 553480 212599 553482
rect 117957 553424 117962 553480
rect 118018 553424 118606 553480
rect 118662 553424 212538 553480
rect 212594 553424 212599 553480
rect 117957 553422 212599 553424
rect 117957 553419 118023 553422
rect 118601 553419 118667 553422
rect 212533 553419 212599 553422
rect 91737 553346 91803 553349
rect 88596 553344 91803 553346
rect 88596 553288 91742 553344
rect 91798 553288 91803 553344
rect 88596 553286 91803 553288
rect 91737 553283 91803 553286
rect 67449 552802 67515 552805
rect 67449 552800 68908 552802
rect 67449 552744 67454 552800
rect 67510 552744 68908 552800
rect 67449 552742 68908 552744
rect 67449 552739 67515 552742
rect 91185 552122 91251 552125
rect 88596 552120 91251 552122
rect 88596 552064 91190 552120
rect 91246 552064 91251 552120
rect 88596 552062 91251 552064
rect 91185 552059 91251 552062
rect 170254 552060 170260 552124
rect 170324 552122 170330 552124
rect 225321 552122 225387 552125
rect 170324 552120 225387 552122
rect 170324 552064 225326 552120
rect 225382 552064 225387 552120
rect 170324 552062 225387 552064
rect 170324 552060 170330 552062
rect 225321 552059 225387 552062
rect 66662 551380 66668 551444
rect 66732 551442 66738 551444
rect 66732 551382 68908 551442
rect 66732 551380 66738 551382
rect 583520 551020 584960 551260
rect 91185 550762 91251 550765
rect 88596 550760 91251 550762
rect 88596 550704 91190 550760
rect 91246 550704 91251 550760
rect 88596 550702 91251 550704
rect 91185 550699 91251 550702
rect 173014 550700 173020 550764
rect 173084 550762 173090 550764
rect 303613 550762 303679 550765
rect 173084 550760 303679 550762
rect 173084 550704 303618 550760
rect 303674 550704 303679 550760
rect 173084 550702 303679 550704
rect 173084 550700 173090 550702
rect 303613 550699 303679 550702
rect 66437 550082 66503 550085
rect 66437 550080 68908 550082
rect 66437 550024 66442 550080
rect 66498 550024 68908 550080
rect 66437 550022 68908 550024
rect 66437 550019 66503 550022
rect 192569 549538 192635 549541
rect 231945 549538 232011 549541
rect 192569 549536 232011 549538
rect 192569 549480 192574 549536
rect 192630 549480 231950 549536
rect 232006 549480 232011 549536
rect 192569 549478 232011 549480
rect 192569 549475 192635 549478
rect 231945 549475 232011 549478
rect 95141 549402 95207 549405
rect 278037 549402 278103 549405
rect 88596 549400 278103 549402
rect 88596 549344 95146 549400
rect 95202 549344 278042 549400
rect 278098 549344 278103 549400
rect 88596 549342 278103 549344
rect 95141 549339 95207 549342
rect 278037 549339 278103 549342
rect 66437 548722 66503 548725
rect 66437 548720 68908 548722
rect 66437 548664 66442 548720
rect 66498 548664 68908 548720
rect 66437 548662 68908 548664
rect 66437 548659 66503 548662
rect 195329 548042 195395 548045
rect 218697 548042 218763 548045
rect 195329 548040 218763 548042
rect 195329 547984 195334 548040
rect 195390 547984 218702 548040
rect 218758 547984 218763 548040
rect 195329 547982 218763 547984
rect 195329 547979 195395 547982
rect 218697 547979 218763 547982
rect 91461 547906 91527 547909
rect 88596 547904 91527 547906
rect 88596 547848 91466 547904
rect 91522 547848 91527 547904
rect 88596 547846 91527 547848
rect 91461 547843 91527 547846
rect 191097 547906 191163 547909
rect 243537 547906 243603 547909
rect 191097 547904 243603 547906
rect 191097 547848 191102 547904
rect 191158 547848 243542 547904
rect 243598 547848 243603 547904
rect 191097 547846 243603 547848
rect 191097 547843 191163 547846
rect 243537 547843 243603 547846
rect 66161 547362 66227 547365
rect 66161 547360 68908 547362
rect 66161 547304 66166 547360
rect 66222 547304 68908 547360
rect 66161 547302 68908 547304
rect 66161 547299 66227 547302
rect 197854 546620 197860 546684
rect 197924 546682 197930 546684
rect 248505 546682 248571 546685
rect 197924 546680 248571 546682
rect 197924 546624 248510 546680
rect 248566 546624 248571 546680
rect 197924 546622 248571 546624
rect 197924 546620 197930 546622
rect 248505 546619 248571 546622
rect 91185 546546 91251 546549
rect 88596 546544 91251 546546
rect 88596 546488 91190 546544
rect 91246 546488 91251 546544
rect 88596 546486 91251 546488
rect 91185 546483 91251 546486
rect 199510 546484 199516 546548
rect 199580 546546 199586 546548
rect 268561 546546 268627 546549
rect 199580 546544 268627 546546
rect 199580 546488 268566 546544
rect 268622 546488 268627 546544
rect 199580 546486 268627 546488
rect 199580 546484 199586 546486
rect 268561 546483 268627 546486
rect 67766 545940 67772 546004
rect 67836 546002 67842 546004
rect 67836 545942 68908 546002
rect 67836 545940 67842 545942
rect 191189 545458 191255 545461
rect 205633 545458 205699 545461
rect 206277 545458 206343 545461
rect 191189 545456 206343 545458
rect 191189 545400 191194 545456
rect 191250 545400 205638 545456
rect 205694 545400 206282 545456
rect 206338 545400 206343 545456
rect 191189 545398 206343 545400
rect 191189 545395 191255 545398
rect 205633 545395 205699 545398
rect 206277 545395 206343 545398
rect 200614 545260 200620 545324
rect 200684 545322 200690 545324
rect 235257 545322 235323 545325
rect 200684 545320 235323 545322
rect 200684 545264 235262 545320
rect 235318 545264 235323 545320
rect 200684 545262 235323 545264
rect 200684 545260 200690 545262
rect 235257 545259 235323 545262
rect 66805 545186 66871 545189
rect 67766 545186 67772 545188
rect 66805 545184 67772 545186
rect 66805 545128 66810 545184
rect 66866 545128 67772 545184
rect 66805 545126 67772 545128
rect 66805 545123 66871 545126
rect 67766 545124 67772 545126
rect 67836 545124 67842 545188
rect 91185 545186 91251 545189
rect 88596 545184 91251 545186
rect 88596 545128 91190 545184
rect 91246 545128 91251 545184
rect 88596 545126 91251 545128
rect 91185 545123 91251 545126
rect 137921 545186 137987 545189
rect 300025 545186 300091 545189
rect 137921 545184 300091 545186
rect 137921 545128 137926 545184
rect 137982 545128 300030 545184
rect 300086 545128 300091 545184
rect 137921 545126 300091 545128
rect 137921 545123 137987 545126
rect 300025 545123 300091 545126
rect 320173 545186 320239 545189
rect 353334 545186 353340 545188
rect 320173 545184 353340 545186
rect 320173 545128 320178 545184
rect 320234 545128 353340 545184
rect 320173 545126 353340 545128
rect 320173 545123 320239 545126
rect 353334 545124 353340 545126
rect 353404 545124 353410 545188
rect 66805 544642 66871 544645
rect 66805 544640 68908 544642
rect 66805 544584 66810 544640
rect 66866 544584 68908 544640
rect 66805 544582 68908 544584
rect 66805 544579 66871 544582
rect 91829 543962 91895 543965
rect 88596 543960 91895 543962
rect 88596 543904 91834 543960
rect 91890 543904 91895 543960
rect 88596 543902 91895 543904
rect 91829 543899 91895 543902
rect 161974 543900 161980 543964
rect 162044 543962 162050 543964
rect 321553 543962 321619 543965
rect 162044 543960 321619 543962
rect 162044 543904 321558 543960
rect 321614 543904 321619 543960
rect 162044 543902 321619 543904
rect 162044 543900 162050 543902
rect 321553 543899 321619 543902
rect 89621 543826 89687 543829
rect 270861 543826 270927 543829
rect 89621 543824 270927 543826
rect 89621 543768 89626 543824
rect 89682 543768 270866 543824
rect 270922 543768 270927 543824
rect 89621 543766 270927 543768
rect 89621 543763 89687 543766
rect 270861 543763 270927 543766
rect 66805 543282 66871 543285
rect 66805 543280 68908 543282
rect 66805 543224 66810 543280
rect 66866 543224 68908 543280
rect 66805 543222 68908 543224
rect 66805 543219 66871 543222
rect 284293 543010 284359 543013
rect 357617 543010 357683 543013
rect 363597 543010 363663 543013
rect 284293 543008 363663 543010
rect 284293 542952 284298 543008
rect 284354 542952 357622 543008
rect 357678 542952 363602 543008
rect 363658 542952 363663 543008
rect 284293 542950 363663 542952
rect 284293 542947 284359 542950
rect 357617 542947 357683 542950
rect 363597 542947 363663 542950
rect 196617 542602 196683 542605
rect 253933 542602 253999 542605
rect 196617 542600 253999 542602
rect 196617 542544 196622 542600
rect 196678 542544 253938 542600
rect 253994 542544 253999 542600
rect 196617 542542 253999 542544
rect 196617 542539 196683 542542
rect 253933 542539 253999 542542
rect 91185 542466 91251 542469
rect 88596 542464 91251 542466
rect 88596 542408 91190 542464
rect 91246 542408 91251 542464
rect 88596 542406 91251 542408
rect 91185 542403 91251 542406
rect 142061 542466 142127 542469
rect 283465 542466 283531 542469
rect 142061 542464 283531 542466
rect 142061 542408 142066 542464
rect 142122 542408 283470 542464
rect 283526 542408 283531 542464
rect 142061 542406 283531 542408
rect 142061 542403 142127 542406
rect 283465 542403 283531 542406
rect 65885 542330 65951 542333
rect 69422 542330 69428 542332
rect 65885 542328 69428 542330
rect 65885 542272 65890 542328
rect 65946 542272 69428 542328
rect 65885 542270 69428 542272
rect 65885 542267 65951 542270
rect 69422 542268 69428 542270
rect 69492 542268 69498 542332
rect 67081 541922 67147 541925
rect 67081 541920 68908 541922
rect 67081 541864 67086 541920
rect 67142 541864 68908 541920
rect 67081 541862 68908 541864
rect 67081 541859 67147 541862
rect 255957 541650 256023 541653
rect 257337 541650 257403 541653
rect 583109 541650 583175 541653
rect 255957 541648 583175 541650
rect 255957 541592 255962 541648
rect 256018 541592 257342 541648
rect 257398 541592 583114 541648
rect 583170 541592 583175 541648
rect 255957 541590 583175 541592
rect 255957 541587 256023 541590
rect 257337 541587 257403 541590
rect 583109 541587 583175 541590
rect 191741 541378 191807 541381
rect 238753 541378 238819 541381
rect 191741 541376 238819 541378
rect 191741 541320 191746 541376
rect 191802 541320 238758 541376
rect 238814 541320 238819 541376
rect 191741 541318 238819 541320
rect 191741 541315 191807 541318
rect 238753 541315 238819 541318
rect 91185 541242 91251 541245
rect 88596 541240 91251 541242
rect 88596 541184 91190 541240
rect 91246 541184 91251 541240
rect 88596 541182 91251 541184
rect 91185 541179 91251 541182
rect 188838 541180 188844 541244
rect 188908 541242 188914 541244
rect 262213 541242 262279 541245
rect 188908 541240 262279 541242
rect 188908 541184 262218 541240
rect 262274 541184 262279 541240
rect 188908 541182 262279 541184
rect 188908 541180 188914 541182
rect 262213 541179 262279 541182
rect 133137 541106 133203 541109
rect 323577 541106 323643 541109
rect 133137 541104 323643 541106
rect 133137 541048 133142 541104
rect 133198 541048 323582 541104
rect 323638 541048 323643 541104
rect 133137 541046 323643 541048
rect 133137 541043 133203 541046
rect 323577 541043 323643 541046
rect -960 540684 480 540924
rect 67541 539610 67607 539613
rect 69430 539610 69490 540532
rect 160686 539820 160692 539884
rect 160756 539882 160762 539884
rect 348693 539882 348759 539885
rect 160756 539880 348759 539882
rect 160756 539824 348698 539880
rect 348754 539824 348759 539880
rect 160756 539822 348759 539824
rect 160756 539820 160762 539822
rect 348693 539819 348759 539822
rect 92381 539746 92447 539749
rect 88596 539744 92447 539746
rect 88596 539688 92386 539744
rect 92442 539688 92447 539744
rect 88596 539686 92447 539688
rect 92381 539683 92447 539686
rect 182817 539746 182883 539749
rect 280613 539746 280679 539749
rect 182817 539744 280679 539746
rect 182817 539688 182822 539744
rect 182878 539688 280618 539744
rect 280674 539688 280679 539744
rect 182817 539686 280679 539688
rect 182817 539683 182883 539686
rect 280613 539683 280679 539686
rect 295517 539746 295583 539749
rect 362902 539746 362908 539748
rect 295517 539744 362908 539746
rect 295517 539688 295522 539744
rect 295578 539688 362908 539744
rect 295517 539686 362908 539688
rect 295517 539683 295583 539686
rect 362902 539684 362908 539686
rect 362972 539684 362978 539748
rect 342069 539610 342135 539613
rect 374085 539610 374151 539613
rect 67541 539608 74550 539610
rect 67541 539552 67546 539608
rect 67602 539552 74550 539608
rect 67541 539550 74550 539552
rect 67541 539547 67607 539550
rect 74490 538794 74550 539550
rect 342069 539608 374151 539610
rect 342069 539552 342074 539608
rect 342130 539552 374090 539608
rect 374146 539552 374151 539608
rect 342069 539550 374151 539552
rect 342069 539547 342135 539550
rect 374085 539547 374151 539550
rect 345381 539474 345447 539477
rect 349153 539474 349219 539477
rect 345381 539472 349219 539474
rect 345381 539416 345386 539472
rect 345442 539416 349158 539472
rect 349214 539416 349219 539472
rect 345381 539414 349219 539416
rect 345381 539411 345447 539414
rect 349153 539411 349219 539414
rect 177389 538794 177455 538797
rect 74490 538792 177455 538794
rect 74490 538736 177394 538792
rect 177450 538736 177455 538792
rect 74490 538734 177455 538736
rect 177389 538731 177455 538734
rect 216581 538794 216647 538797
rect 347681 538794 347747 538797
rect 216581 538792 347747 538794
rect 216581 538736 216586 538792
rect 216642 538736 347686 538792
rect 347742 538736 347747 538792
rect 216581 538734 347747 538736
rect 216581 538731 216647 538734
rect 347681 538731 347747 538734
rect 213453 538522 213519 538525
rect 217133 538522 217199 538525
rect 213453 538520 217199 538522
rect 213453 538464 213458 538520
rect 213514 538464 217138 538520
rect 217194 538464 217199 538520
rect 213453 538462 217199 538464
rect 213453 538459 213519 538462
rect 217133 538459 217199 538462
rect 193949 538386 194015 538389
rect 222469 538386 222535 538389
rect 193949 538384 222535 538386
rect 193949 538328 193954 538384
rect 194010 538328 222474 538384
rect 222530 538328 222535 538384
rect 193949 538326 222535 538328
rect 193949 538323 194015 538326
rect 222469 538323 222535 538326
rect 350349 538386 350415 538389
rect 361573 538386 361639 538389
rect 350349 538384 361639 538386
rect 350349 538328 350354 538384
rect 350410 538328 361578 538384
rect 361634 538328 361639 538384
rect 350349 538326 361639 538328
rect 350349 538323 350415 538326
rect 361573 538323 361639 538326
rect 186957 538250 187023 538253
rect 213453 538250 213519 538253
rect 186957 538248 213519 538250
rect 186957 538192 186962 538248
rect 187018 538192 213458 538248
rect 213514 538192 213519 538248
rect 186957 538190 213519 538192
rect 186957 538187 187023 538190
rect 213453 538187 213519 538190
rect 216673 538250 216739 538253
rect 265525 538250 265591 538253
rect 216673 538248 265591 538250
rect 216673 538192 216678 538248
rect 216734 538192 265530 538248
rect 265586 538192 265591 538248
rect 216673 538190 265591 538192
rect 216673 538187 216739 538190
rect 265525 538187 265591 538190
rect 318701 538250 318767 538253
rect 352046 538250 352052 538252
rect 318701 538248 352052 538250
rect 318701 538192 318706 538248
rect 318762 538192 352052 538248
rect 318701 538190 352052 538192
rect 318701 538187 318767 538190
rect 352046 538188 352052 538190
rect 352116 538188 352122 538252
rect 355317 538250 355383 538253
rect 371233 538250 371299 538253
rect 355317 538248 371299 538250
rect 355317 538192 355322 538248
rect 355378 538192 371238 538248
rect 371294 538192 371299 538248
rect 355317 538190 371299 538192
rect 355317 538187 355383 538190
rect 371233 538187 371299 538190
rect 67357 538114 67423 538117
rect 177297 538114 177363 538117
rect 67357 538112 177363 538114
rect 67357 538056 67362 538112
rect 67418 538056 177302 538112
rect 177358 538056 177363 538112
rect 67357 538054 177363 538056
rect 67357 538051 67423 538054
rect 177297 538051 177363 538054
rect 580165 537842 580231 537845
rect 583520 537842 584960 537932
rect 580165 537840 584960 537842
rect 580165 537784 580170 537840
rect 580226 537784 584960 537840
rect 580165 537782 584960 537784
rect 580165 537779 580231 537782
rect 583520 537692 584960 537782
rect 67081 537434 67147 537437
rect 67398 537434 67404 537436
rect 67081 537432 67404 537434
rect 67081 537376 67086 537432
rect 67142 537376 67404 537432
rect 67081 537374 67404 537376
rect 67081 537371 67147 537374
rect 67398 537372 67404 537374
rect 67468 537372 67474 537436
rect 148317 537162 148383 537165
rect 293861 537162 293927 537165
rect 148317 537160 293927 537162
rect 148317 537104 148322 537160
rect 148378 537104 293866 537160
rect 293922 537104 293927 537160
rect 148317 537102 293927 537104
rect 148317 537099 148383 537102
rect 293861 537099 293927 537102
rect 302141 537162 302207 537165
rect 357566 537162 357572 537164
rect 302141 537160 357572 537162
rect 302141 537104 302146 537160
rect 302202 537104 357572 537160
rect 302141 537102 357572 537104
rect 302141 537099 302207 537102
rect 357566 537100 357572 537102
rect 357636 537100 357642 537164
rect 184289 537026 184355 537029
rect 335445 537026 335511 537029
rect 184289 537024 335511 537026
rect 184289 536968 184294 537024
rect 184350 536968 335450 537024
rect 335506 536968 335511 537024
rect 184289 536966 335511 536968
rect 184289 536963 184355 536966
rect 335445 536963 335511 536966
rect 173157 536890 173223 536893
rect 333789 536890 333855 536893
rect 173157 536888 333855 536890
rect 173157 536832 173162 536888
rect 173218 536832 333794 536888
rect 333850 536832 333855 536888
rect 173157 536830 333855 536832
rect 173157 536827 173223 536830
rect 333789 536827 333855 536830
rect 72417 536754 72483 536757
rect 133137 536754 133203 536757
rect 72417 536752 133203 536754
rect 72417 536696 72422 536752
rect 72478 536696 133142 536752
rect 133198 536696 133203 536752
rect 72417 536694 133203 536696
rect 72417 536691 72483 536694
rect 133137 536691 133203 536694
rect 68645 536618 68711 536621
rect 88149 536618 88215 536621
rect 68645 536616 88215 536618
rect 68645 536560 68650 536616
rect 68706 536560 88154 536616
rect 88210 536560 88215 536616
rect 68645 536558 88215 536560
rect 68645 536555 68711 536558
rect 88149 536555 88215 536558
rect 159357 535802 159423 535805
rect 313365 535802 313431 535805
rect 159357 535800 313431 535802
rect 159357 535744 159362 535800
rect 159418 535744 313370 535800
rect 313426 535744 313431 535800
rect 159357 535742 313431 535744
rect 159357 535739 159423 535742
rect 313365 535739 313431 535742
rect 169109 535666 169175 535669
rect 276013 535666 276079 535669
rect 276933 535666 276999 535669
rect 169109 535664 276999 535666
rect 169109 535608 169114 535664
rect 169170 535608 276018 535664
rect 276074 535608 276938 535664
rect 276994 535608 276999 535664
rect 169109 535606 276999 535608
rect 169109 535603 169175 535606
rect 276013 535603 276079 535606
rect 276933 535603 276999 535606
rect 68134 535468 68140 535532
rect 68204 535530 68210 535532
rect 68645 535530 68711 535533
rect 69565 535532 69631 535533
rect 69565 535530 69612 535532
rect 68204 535528 68711 535530
rect 68204 535472 68650 535528
rect 68706 535472 68711 535528
rect 68204 535470 68711 535472
rect 69520 535528 69612 535530
rect 69520 535472 69570 535528
rect 69520 535470 69612 535472
rect 68204 535468 68210 535470
rect 68645 535467 68711 535470
rect 69565 535468 69612 535470
rect 69676 535468 69682 535532
rect 197997 535530 198063 535533
rect 203701 535530 203767 535533
rect 197997 535528 203767 535530
rect 197997 535472 198002 535528
rect 198058 535472 203706 535528
rect 203762 535472 203767 535528
rect 197997 535470 203767 535472
rect 69565 535467 69631 535468
rect 197997 535467 198063 535470
rect 203701 535467 203767 535470
rect 315665 535530 315731 535533
rect 360377 535530 360443 535533
rect 315665 535528 360443 535530
rect 315665 535472 315670 535528
rect 315726 535472 360382 535528
rect 360438 535472 360443 535528
rect 315665 535470 360443 535472
rect 315665 535467 315731 535470
rect 360377 535467 360443 535470
rect 67766 535332 67772 535396
rect 67836 535394 67842 535396
rect 146937 535394 147003 535397
rect 67836 535392 147003 535394
rect 67836 535336 146942 535392
rect 146998 535336 147003 535392
rect 67836 535334 147003 535336
rect 67836 535332 67842 535334
rect 146937 535331 147003 535334
rect 191598 535332 191604 535396
rect 191668 535394 191674 535396
rect 201401 535394 201467 535397
rect 216581 535394 216647 535397
rect 191668 535392 201467 535394
rect 191668 535336 201406 535392
rect 201462 535336 201467 535392
rect 191668 535334 201467 535336
rect 191668 535332 191674 535334
rect 201401 535331 201467 535334
rect 209730 535392 216647 535394
rect 209730 535336 216586 535392
rect 216642 535336 216647 535392
rect 209730 535334 216647 535336
rect 199837 534986 199903 534989
rect 209730 534986 209790 535334
rect 216581 535331 216647 535334
rect 199837 534984 209790 534986
rect 199837 534928 199842 534984
rect 199898 534928 209790 534984
rect 199837 534926 209790 534928
rect 199837 534923 199903 534926
rect 93669 534714 93735 534717
rect 106406 534714 106412 534716
rect 93669 534712 106412 534714
rect 93669 534656 93674 534712
rect 93730 534656 106412 534712
rect 93669 534654 106412 534656
rect 93669 534651 93735 534654
rect 106406 534652 106412 534654
rect 106476 534652 106482 534716
rect 357617 534714 357683 534717
rect 356132 534712 357683 534714
rect 356132 534656 357622 534712
rect 357678 534656 357683 534712
rect 356132 534654 357683 534656
rect 357617 534651 357683 534654
rect 183318 534108 183324 534172
rect 183388 534170 183394 534172
rect 200070 534170 200130 534548
rect 183388 534110 200130 534170
rect 183388 534108 183394 534110
rect 143441 534034 143507 534037
rect 199837 534034 199903 534037
rect 143441 534032 199903 534034
rect 143441 533976 143446 534032
rect 143502 533976 199842 534032
rect 199898 533976 199903 534032
rect 143441 533974 199903 533976
rect 143441 533971 143507 533974
rect 199837 533971 199903 533974
rect 142797 533626 142863 533629
rect 143441 533626 143507 533629
rect 142797 533624 143507 533626
rect 142797 533568 142802 533624
rect 142858 533568 143446 533624
rect 143502 533568 143507 533624
rect 142797 533566 143507 533568
rect 142797 533563 142863 533566
rect 143441 533563 143507 533566
rect 190361 533490 190427 533493
rect 200062 533490 200068 533492
rect 190361 533488 200068 533490
rect 190361 533432 190366 533488
rect 190422 533432 200068 533488
rect 190361 533430 200068 533432
rect 190361 533427 190427 533430
rect 200062 533428 200068 533430
rect 200132 533428 200138 533492
rect 197353 532266 197419 532269
rect 197353 532264 200100 532266
rect 197353 532208 197358 532264
rect 197414 532208 200100 532264
rect 197353 532206 200100 532208
rect 197353 532203 197419 532206
rect 358721 532130 358787 532133
rect 356132 532128 358787 532130
rect 356132 532072 358726 532128
rect 358782 532072 358787 532128
rect 356132 532070 358787 532072
rect 358721 532067 358787 532070
rect 179270 530572 179276 530636
rect 179340 530634 179346 530636
rect 198733 530634 198799 530637
rect 179340 530632 198799 530634
rect 179340 530576 198738 530632
rect 198794 530576 198799 530632
rect 179340 530574 198799 530576
rect 179340 530572 179346 530574
rect 198733 530571 198799 530574
rect 197353 529818 197419 529821
rect 198549 529818 198615 529821
rect 197353 529816 200100 529818
rect 197353 529760 197358 529816
rect 197414 529760 198554 529816
rect 198610 529760 200100 529816
rect 197353 529758 200100 529760
rect 197353 529755 197419 529758
rect 198549 529755 198615 529758
rect 358905 529682 358971 529685
rect 356132 529680 358971 529682
rect 356132 529624 358910 529680
rect 358966 529624 358971 529680
rect 356132 529622 358971 529624
rect 358905 529619 358971 529622
rect -960 527914 480 528004
rect 3417 527914 3483 527917
rect -960 527912 3483 527914
rect -960 527856 3422 527912
rect 3478 527856 3483 527912
rect -960 527854 3483 527856
rect -960 527764 480 527854
rect 3417 527851 3483 527854
rect 197353 527370 197419 527373
rect 197353 527368 200100 527370
rect 197353 527312 197358 527368
rect 197414 527312 200100 527368
rect 197353 527310 200100 527312
rect 197353 527307 197419 527310
rect 358721 527234 358787 527237
rect 356132 527232 358787 527234
rect 356132 527176 358726 527232
rect 358782 527176 358787 527232
rect 356132 527174 358787 527176
rect 358721 527171 358787 527174
rect 35801 526418 35867 526421
rect 197854 526418 197860 526420
rect 35801 526416 197860 526418
rect 35801 526360 35806 526416
rect 35862 526360 197860 526416
rect 35801 526358 197860 526360
rect 35801 526355 35867 526358
rect 197854 526356 197860 526358
rect 197924 526356 197930 526420
rect 197445 524786 197511 524789
rect 358721 524786 358787 524789
rect 197445 524784 200100 524786
rect 197445 524728 197450 524784
rect 197506 524728 200100 524784
rect 197445 524726 200100 524728
rect 356132 524784 358787 524786
rect 356132 524728 358726 524784
rect 358782 524728 358787 524784
rect 356132 524726 358787 524728
rect 197445 524723 197511 524726
rect 358721 524723 358787 524726
rect 582373 524514 582439 524517
rect 583520 524514 584960 524604
rect 582373 524512 584960 524514
rect 582373 524456 582378 524512
rect 582434 524456 584960 524512
rect 582373 524454 584960 524456
rect 582373 524451 582439 524454
rect 583520 524364 584960 524454
rect 66478 523772 66484 523836
rect 66548 523834 66554 523836
rect 66897 523834 66963 523837
rect 66548 523832 66963 523834
rect 66548 523776 66902 523832
rect 66958 523776 66963 523832
rect 66548 523774 66963 523776
rect 66548 523772 66554 523774
rect 66897 523771 66963 523774
rect 66662 523636 66668 523700
rect 66732 523698 66738 523700
rect 67081 523698 67147 523701
rect 66732 523696 67147 523698
rect 66732 523640 67086 523696
rect 67142 523640 67147 523696
rect 66732 523638 67147 523640
rect 66732 523636 66738 523638
rect 67081 523635 67147 523638
rect 197353 522338 197419 522341
rect 357433 522338 357499 522341
rect 358721 522338 358787 522341
rect 197353 522336 200100 522338
rect 197353 522280 197358 522336
rect 197414 522280 200100 522336
rect 197353 522278 200100 522280
rect 356132 522336 358787 522338
rect 356132 522280 357438 522336
rect 357494 522280 358726 522336
rect 358782 522280 358787 522336
rect 356132 522278 358787 522280
rect 197353 522275 197419 522278
rect 357433 522275 357499 522278
rect 358721 522275 358787 522278
rect 357893 520026 357959 520029
rect 356132 520024 357959 520026
rect 356132 519968 357898 520024
rect 357954 519968 357959 520024
rect 356132 519966 357959 519968
rect 357893 519963 357959 519966
rect 197353 519890 197419 519893
rect 197353 519888 200100 519890
rect 197353 519832 197358 519888
rect 197414 519832 200100 519888
rect 197353 519830 200100 519832
rect 197353 519827 197419 519830
rect 197353 517442 197419 517445
rect 358721 517442 358787 517445
rect 197353 517440 200100 517442
rect 197353 517384 197358 517440
rect 197414 517384 200100 517440
rect 197353 517382 200100 517384
rect 356132 517440 358787 517442
rect 356132 517384 358726 517440
rect 358782 517384 358787 517440
rect 356132 517382 358787 517384
rect 197353 517379 197419 517382
rect 358721 517379 358787 517382
rect -960 514858 480 514948
rect 195094 514932 195100 514996
rect 195164 514994 195170 514996
rect 358629 514994 358695 514997
rect 195164 514934 200100 514994
rect 356132 514992 358695 514994
rect 356132 514936 358634 514992
rect 358690 514936 358695 514992
rect 356132 514934 358695 514936
rect 195164 514932 195170 514934
rect 358629 514931 358695 514934
rect 2773 514858 2839 514861
rect -960 514856 2839 514858
rect -960 514800 2778 514856
rect 2834 514800 2839 514856
rect -960 514798 2839 514800
rect -960 514708 480 514798
rect 2773 514795 2839 514798
rect 357525 512682 357591 512685
rect 356132 512680 357591 512682
rect 356132 512624 357530 512680
rect 357586 512624 357591 512680
rect 356132 512622 357591 512624
rect 357525 512619 357591 512622
rect 198590 512484 198596 512548
rect 198660 512546 198666 512548
rect 198660 512486 200100 512546
rect 198660 512484 198666 512486
rect 582373 511322 582439 511325
rect 583520 511322 584960 511412
rect 582373 511320 584960 511322
rect 582373 511264 582378 511320
rect 582434 511264 584960 511320
rect 582373 511262 584960 511264
rect 582373 511259 582439 511262
rect 583520 511172 584960 511262
rect 197353 510234 197419 510237
rect 197353 510232 200100 510234
rect 197353 510176 197358 510232
rect 197414 510176 200100 510232
rect 197353 510174 200100 510176
rect 197353 510171 197419 510174
rect 357617 510098 357683 510101
rect 356132 510096 357683 510098
rect 356132 510040 357622 510096
rect 357678 510040 357683 510096
rect 356132 510038 357683 510040
rect 357617 510035 357683 510038
rect 197353 507650 197419 507653
rect 197353 507648 200100 507650
rect 197353 507592 197358 507648
rect 197414 507592 200100 507648
rect 197353 507590 200100 507592
rect 197353 507587 197419 507590
rect 356102 507106 356162 507620
rect 356278 507106 356284 507108
rect 356102 507046 356284 507106
rect 356278 507044 356284 507046
rect 356348 507044 356354 507108
rect 199101 505202 199167 505205
rect 358721 505202 358787 505205
rect 199101 505200 200100 505202
rect 199101 505144 199106 505200
rect 199162 505144 200100 505200
rect 199101 505142 200100 505144
rect 356132 505200 358787 505202
rect 356132 505144 358726 505200
rect 358782 505144 358787 505200
rect 356132 505142 358787 505144
rect 199101 505139 199167 505142
rect 358721 505139 358787 505142
rect 155718 504324 155724 504388
rect 155788 504386 155794 504388
rect 176009 504386 176075 504389
rect 155788 504384 176075 504386
rect 155788 504328 176014 504384
rect 176070 504328 176075 504384
rect 155788 504326 176075 504328
rect 155788 504324 155794 504326
rect 176009 504323 176075 504326
rect 358721 502754 358787 502757
rect 356132 502752 358787 502754
rect 184790 502420 184796 502484
rect 184860 502482 184866 502484
rect 200070 502482 200130 502724
rect 356132 502696 358726 502752
rect 358782 502696 358787 502752
rect 356132 502694 358787 502696
rect 358721 502691 358787 502694
rect 184860 502422 200130 502482
rect 184860 502420 184866 502422
rect -960 501802 480 501892
rect 3509 501802 3575 501805
rect -960 501800 3575 501802
rect -960 501744 3514 501800
rect 3570 501744 3575 501800
rect -960 501742 3575 501744
rect -960 501652 480 501742
rect 3509 501739 3575 501742
rect 197353 500442 197419 500445
rect 198641 500442 198707 500445
rect 197353 500440 200100 500442
rect 197353 500384 197358 500440
rect 197414 500384 198646 500440
rect 198702 500384 200100 500440
rect 197353 500382 200100 500384
rect 197353 500379 197419 500382
rect 198641 500379 198707 500382
rect 358721 500306 358787 500309
rect 356132 500304 358787 500306
rect 356132 500248 358726 500304
rect 358782 500248 358787 500304
rect 356132 500246 358787 500248
rect 358721 500243 358787 500246
rect 358077 497858 358143 497861
rect 356132 497856 358143 497858
rect 177798 496844 177804 496908
rect 177868 496906 177874 496908
rect 200070 496906 200130 497828
rect 356132 497800 358082 497856
rect 358138 497800 358143 497856
rect 583520 497844 584960 498084
rect 356132 497798 358143 497800
rect 358077 497795 358143 497798
rect 177868 496846 200130 496906
rect 177868 496844 177874 496846
rect 197353 495546 197419 495549
rect 357157 495546 357223 495549
rect 197353 495544 200100 495546
rect 197353 495488 197358 495544
rect 197414 495488 200100 495544
rect 197353 495486 200100 495488
rect 356132 495544 357223 495546
rect 356132 495488 357162 495544
rect 357218 495488 357223 495544
rect 356132 495486 357223 495488
rect 197353 495483 197419 495486
rect 357157 495483 357223 495486
rect 358629 493098 358695 493101
rect 356132 493096 358695 493098
rect 356132 493068 358634 493096
rect 356102 493040 358634 493068
rect 358690 493040 358695 493096
rect 356102 493038 358695 493040
rect 197353 492962 197419 492965
rect 197353 492960 200100 492962
rect 197353 492904 197358 492960
rect 197414 492904 200100 492960
rect 197353 492902 200100 492904
rect 197353 492899 197419 492902
rect 356102 492690 356162 493038
rect 358629 493035 358695 493038
rect 356237 492690 356303 492693
rect 356102 492688 356303 492690
rect 356102 492632 356242 492688
rect 356298 492632 356303 492688
rect 356102 492630 356303 492632
rect 356237 492627 356303 492630
rect 197353 490514 197419 490517
rect 197353 490512 200100 490514
rect 197353 490456 197358 490512
rect 197414 490456 200100 490512
rect 197353 490454 200100 490456
rect 197353 490451 197419 490454
rect 356605 490378 356671 490381
rect 356132 490376 356671 490378
rect 356132 490320 356610 490376
rect 356666 490320 356671 490376
rect 356132 490318 356671 490320
rect 356605 490315 356671 490318
rect -960 488596 480 488836
rect 197353 488066 197419 488069
rect 197353 488064 200100 488066
rect 197353 488008 197358 488064
rect 197414 488008 200100 488064
rect 197353 488006 200100 488008
rect 197353 488003 197419 488006
rect 358721 487794 358787 487797
rect 356132 487792 358787 487794
rect 356132 487736 358726 487792
rect 358782 487736 358787 487792
rect 356132 487734 358787 487736
rect 358721 487731 358787 487734
rect 198774 485556 198780 485620
rect 198844 485618 198850 485620
rect 198844 485558 200100 485618
rect 198844 485556 198850 485558
rect 358721 485346 358787 485349
rect 356132 485344 358787 485346
rect 356132 485288 358726 485344
rect 358782 485288 358787 485344
rect 356132 485286 358787 485288
rect 358721 485283 358787 485286
rect 580257 484666 580323 484669
rect 583520 484666 584960 484756
rect 580257 484664 584960 484666
rect 580257 484608 580262 484664
rect 580318 484608 584960 484664
rect 580257 484606 584960 484608
rect 580257 484603 580323 484606
rect 583520 484516 584960 484606
rect 197997 483170 198063 483173
rect 197997 483168 200100 483170
rect 197997 483112 198002 483168
rect 198058 483112 200100 483168
rect 197997 483110 200100 483112
rect 197997 483107 198063 483110
rect 357433 482898 357499 482901
rect 356132 482896 357499 482898
rect 356132 482840 357438 482896
rect 357494 482840 357499 482896
rect 356132 482838 357499 482840
rect 357433 482835 357499 482838
rect 197353 480722 197419 480725
rect 197353 480720 200100 480722
rect 197353 480664 197358 480720
rect 197414 480664 200100 480720
rect 197353 480662 200100 480664
rect 197353 480659 197419 480662
rect 360142 480450 360148 480452
rect 356132 480390 360148 480450
rect 360142 480388 360148 480390
rect 360212 480388 360218 480452
rect 107009 479498 107075 479501
rect 122598 479498 122604 479500
rect 107009 479496 122604 479498
rect 107009 479440 107014 479496
rect 107070 479440 122604 479496
rect 107009 479438 122604 479440
rect 107009 479435 107075 479438
rect 122598 479436 122604 479438
rect 122668 479436 122674 479500
rect 197353 478274 197419 478277
rect 197353 478272 200100 478274
rect 197353 478216 197358 478272
rect 197414 478216 200100 478272
rect 197353 478214 200100 478216
rect 197353 478211 197419 478214
rect 358721 478002 358787 478005
rect 356132 478000 358787 478002
rect 356132 477944 358726 478000
rect 358782 477944 358787 478000
rect 356132 477942 358787 477944
rect 358721 477939 358787 477942
rect 197353 475826 197419 475829
rect 197353 475824 200100 475826
rect -960 475690 480 475780
rect 197353 475768 197358 475824
rect 197414 475768 200100 475824
rect 197353 475766 200100 475768
rect 197353 475763 197419 475766
rect 3325 475690 3391 475693
rect -960 475688 3391 475690
rect -960 475632 3330 475688
rect 3386 475632 3391 475688
rect -960 475630 3391 475632
rect -960 475540 480 475630
rect 3325 475627 3391 475630
rect 358721 475554 358787 475557
rect 356132 475552 358787 475554
rect 356132 475496 358726 475552
rect 358782 475496 358787 475552
rect 356132 475494 358787 475496
rect 358721 475491 358787 475494
rect 100109 474058 100175 474061
rect 115974 474058 115980 474060
rect 100109 474056 115980 474058
rect 100109 474000 100114 474056
rect 100170 474000 115980 474056
rect 100109 473998 115980 474000
rect 100109 473995 100175 473998
rect 115974 473996 115980 473998
rect 116044 473996 116050 474060
rect 197353 473378 197419 473381
rect 197353 473376 200100 473378
rect 197353 473320 197358 473376
rect 197414 473320 200100 473376
rect 197353 473318 200100 473320
rect 197353 473315 197419 473318
rect 358721 473106 358787 473109
rect 356132 473104 358787 473106
rect 356132 473048 358726 473104
rect 358782 473048 358787 473104
rect 356132 473046 358787 473048
rect 358721 473043 358787 473046
rect 582925 471474 582991 471477
rect 583520 471474 584960 471564
rect 582925 471472 584960 471474
rect 582925 471416 582930 471472
rect 582986 471416 584960 471472
rect 582925 471414 584960 471416
rect 582925 471411 582991 471414
rect 583520 471324 584960 471414
rect 197629 470930 197695 470933
rect 197629 470928 200100 470930
rect 197629 470872 197634 470928
rect 197690 470872 200100 470928
rect 197629 470870 200100 470872
rect 197629 470867 197695 470870
rect 98729 470658 98795 470661
rect 104934 470658 104940 470660
rect 98729 470656 104940 470658
rect 98729 470600 98734 470656
rect 98790 470600 104940 470656
rect 98729 470598 104940 470600
rect 98729 470595 98795 470598
rect 104934 470596 104940 470598
rect 105004 470596 105010 470660
rect 358721 470658 358787 470661
rect 356132 470656 358787 470658
rect 356132 470600 358726 470656
rect 358782 470600 358787 470656
rect 356132 470598 358787 470600
rect 358721 470595 358787 470598
rect 97349 469842 97415 469845
rect 118182 469842 118188 469844
rect 97349 469840 118188 469842
rect 97349 469784 97354 469840
rect 97410 469784 118188 469840
rect 97349 469782 118188 469784
rect 97349 469779 97415 469782
rect 118182 469780 118188 469782
rect 118252 469780 118258 469844
rect 197353 468482 197419 468485
rect 197353 468480 200100 468482
rect 197353 468424 197358 468480
rect 197414 468424 200100 468480
rect 197353 468422 200100 468424
rect 197353 468419 197419 468422
rect 358721 468210 358787 468213
rect 356132 468208 358787 468210
rect 356132 468152 358726 468208
rect 358782 468152 358787 468208
rect 356132 468150 358787 468152
rect 358721 468147 358787 468150
rect 70158 467876 70164 467940
rect 70228 467938 70234 467940
rect 155217 467938 155283 467941
rect 70228 467936 155283 467938
rect 70228 467880 155222 467936
rect 155278 467880 155283 467936
rect 70228 467878 155283 467880
rect 70228 467876 70234 467878
rect 155217 467875 155283 467878
rect 108941 467802 109007 467805
rect 113214 467802 113220 467804
rect 108941 467800 113220 467802
rect 108941 467744 108946 467800
rect 109002 467744 113220 467800
rect 108941 467742 113220 467744
rect 108941 467739 109007 467742
rect 113214 467740 113220 467742
rect 113284 467740 113290 467804
rect 94497 467122 94563 467125
rect 107694 467122 107700 467124
rect 94497 467120 107700 467122
rect 94497 467064 94502 467120
rect 94558 467064 107700 467120
rect 94497 467062 107700 467064
rect 94497 467059 94563 467062
rect 107694 467060 107700 467062
rect 107764 467060 107770 467124
rect 197353 466034 197419 466037
rect 197353 466032 200100 466034
rect 197353 465976 197358 466032
rect 197414 465976 200100 466032
rect 197353 465974 200100 465976
rect 197353 465971 197419 465974
rect 356789 465762 356855 465765
rect 356132 465760 356855 465762
rect 356132 465704 356794 465760
rect 356850 465704 356855 465760
rect 356132 465702 356855 465704
rect 356789 465699 356855 465702
rect 93209 464402 93275 464405
rect 102174 464402 102180 464404
rect 93209 464400 102180 464402
rect 93209 464344 93214 464400
rect 93270 464344 102180 464400
rect 93209 464342 102180 464344
rect 93209 464339 93275 464342
rect 102174 464340 102180 464342
rect 102244 464340 102250 464404
rect 197353 463314 197419 463317
rect 198825 463314 198891 463317
rect 358721 463314 358787 463317
rect 197353 463312 200100 463314
rect 197353 463256 197358 463312
rect 197414 463256 198830 463312
rect 198886 463256 200100 463312
rect 197353 463254 200100 463256
rect 356132 463312 358787 463314
rect 356132 463256 358726 463312
rect 358782 463256 358787 463312
rect 356132 463254 358787 463256
rect 197353 463251 197419 463254
rect 198825 463251 198891 463254
rect 358721 463251 358787 463254
rect 61837 462906 61903 462909
rect 71814 462906 71820 462908
rect 61837 462904 71820 462906
rect 61837 462848 61842 462904
rect 61898 462848 71820 462904
rect 61837 462846 71820 462848
rect 61837 462843 61903 462846
rect 71814 462844 71820 462846
rect 71884 462844 71890 462908
rect 82813 462906 82879 462909
rect 92974 462906 92980 462908
rect 82813 462904 92980 462906
rect 82813 462848 82818 462904
rect 82874 462848 92980 462904
rect 82813 462846 92980 462848
rect 82813 462843 82879 462846
rect 92974 462844 92980 462846
rect 93044 462844 93050 462908
rect -960 462634 480 462724
rect 3509 462634 3575 462637
rect -960 462632 3575 462634
rect -960 462576 3514 462632
rect 3570 462576 3575 462632
rect -960 462574 3575 462576
rect -960 462484 480 462574
rect 3509 462571 3575 462574
rect 197353 460866 197419 460869
rect 358445 460866 358511 460869
rect 197353 460864 200100 460866
rect 197353 460808 197358 460864
rect 197414 460808 200100 460864
rect 197353 460806 200100 460808
rect 356132 460864 358511 460866
rect 356132 460808 358450 460864
rect 358506 460808 358511 460864
rect 356132 460806 358511 460808
rect 197353 460803 197419 460806
rect 358445 460803 358511 460806
rect 83457 460186 83523 460189
rect 89662 460186 89668 460188
rect 83457 460184 89668 460186
rect 83457 460128 83462 460184
rect 83518 460128 89668 460184
rect 83457 460126 89668 460128
rect 83457 460123 83523 460126
rect 89662 460124 89668 460126
rect 89732 460124 89738 460188
rect 95141 460186 95207 460189
rect 111742 460186 111748 460188
rect 95141 460184 111748 460186
rect 95141 460128 95146 460184
rect 95202 460128 111748 460184
rect 95141 460126 111748 460128
rect 95141 460123 95207 460126
rect 111742 460124 111748 460126
rect 111812 460124 111818 460188
rect 89069 459642 89135 459645
rect 94078 459642 94084 459644
rect 89069 459640 94084 459642
rect 89069 459584 89074 459640
rect 89130 459584 94084 459640
rect 89069 459582 94084 459584
rect 89069 459579 89135 459582
rect 94078 459580 94084 459582
rect 94148 459580 94154 459644
rect 112437 458826 112503 458829
rect 118734 458826 118740 458828
rect 112437 458824 118740 458826
rect 112437 458768 112442 458824
rect 112498 458768 118740 458824
rect 112437 458766 118740 458768
rect 112437 458763 112503 458766
rect 118734 458764 118740 458766
rect 118804 458764 118810 458828
rect 197353 458418 197419 458421
rect 198825 458418 198891 458421
rect 358854 458418 358860 458420
rect 197353 458416 200100 458418
rect 197353 458360 197358 458416
rect 197414 458360 198830 458416
rect 198886 458360 200100 458416
rect 197353 458358 200100 458360
rect 356132 458358 358860 458418
rect 197353 458355 197419 458358
rect 198825 458355 198891 458358
rect 358854 458356 358860 458358
rect 358924 458356 358930 458420
rect 582833 458146 582899 458149
rect 583520 458146 584960 458236
rect 582833 458144 584960 458146
rect 582833 458088 582838 458144
rect 582894 458088 584960 458144
rect 582833 458086 584960 458088
rect 582833 458083 582899 458086
rect 583520 457996 584960 458086
rect 86861 457466 86927 457469
rect 96654 457466 96660 457468
rect 86861 457464 96660 457466
rect 86861 457408 86866 457464
rect 86922 457408 96660 457464
rect 86861 457406 96660 457408
rect 86861 457403 86927 457406
rect 96654 457404 96660 457406
rect 96724 457404 96730 457468
rect 97257 457466 97323 457469
rect 108982 457466 108988 457468
rect 97257 457464 108988 457466
rect 97257 457408 97262 457464
rect 97318 457408 108988 457464
rect 97257 457406 108988 457408
rect 97257 457403 97323 457406
rect 108982 457404 108988 457406
rect 109052 457404 109058 457468
rect 97993 456922 98059 456925
rect 98637 456922 98703 456925
rect 172462 456922 172468 456924
rect 97993 456920 172468 456922
rect 97993 456864 97998 456920
rect 98054 456864 98642 456920
rect 98698 456864 172468 456920
rect 97993 456862 172468 456864
rect 97993 456859 98059 456862
rect 98637 456859 98703 456862
rect 172462 456860 172468 456862
rect 172532 456860 172538 456924
rect 81433 456242 81499 456245
rect 90214 456242 90220 456244
rect 81433 456240 90220 456242
rect 81433 456184 81438 456240
rect 81494 456184 90220 456240
rect 81433 456182 90220 456184
rect 81433 456179 81499 456182
rect 90214 456180 90220 456182
rect 90284 456180 90290 456244
rect 90449 456106 90515 456109
rect 100702 456106 100708 456108
rect 90449 456104 100708 456106
rect 90449 456048 90454 456104
rect 90510 456048 100708 456104
rect 90449 456046 100708 456048
rect 90449 456043 90515 456046
rect 100702 456044 100708 456046
rect 100772 456044 100778 456108
rect 198641 455970 198707 455973
rect 358721 455970 358787 455973
rect 198641 455968 200100 455970
rect 198641 455912 198646 455968
rect 198702 455912 200100 455968
rect 198641 455910 200100 455912
rect 356132 455968 358787 455970
rect 356132 455912 358726 455968
rect 358782 455912 358787 455968
rect 356132 455910 358787 455912
rect 198641 455907 198707 455910
rect 358721 455907 358787 455910
rect 86953 454746 87019 454749
rect 98126 454746 98132 454748
rect 86953 454744 98132 454746
rect 86953 454688 86958 454744
rect 87014 454688 98132 454744
rect 86953 454686 98132 454688
rect 86953 454683 87019 454686
rect 98126 454684 98132 454686
rect 98196 454684 98202 454748
rect 198549 453522 198615 453525
rect 358721 453522 358787 453525
rect 198549 453520 200100 453522
rect 198549 453464 198554 453520
rect 198610 453464 200100 453520
rect 198549 453462 200100 453464
rect 356132 453520 358787 453522
rect 356132 453464 358726 453520
rect 358782 453464 358787 453520
rect 356132 453462 358787 453464
rect 198549 453459 198615 453462
rect 358721 453459 358787 453462
rect 104157 453250 104223 453253
rect 122966 453250 122972 453252
rect 104157 453248 122972 453250
rect 104157 453192 104162 453248
rect 104218 453192 122972 453248
rect 104157 453190 122972 453192
rect 104157 453187 104223 453190
rect 122966 453188 122972 453190
rect 123036 453188 123042 453252
rect 100017 451890 100083 451893
rect 123569 451890 123635 451893
rect 100017 451888 123635 451890
rect 100017 451832 100022 451888
rect 100078 451832 123574 451888
rect 123630 451832 123635 451888
rect 100017 451830 123635 451832
rect 100017 451827 100083 451830
rect 123569 451827 123635 451830
rect 358721 451074 358787 451077
rect 356132 451072 358787 451074
rect 91502 450468 91508 450532
rect 91572 450530 91578 450532
rect 120022 450530 120028 450532
rect 91572 450470 120028 450530
rect 91572 450468 91578 450470
rect 120022 450468 120028 450470
rect 120092 450468 120098 450532
rect 172094 449924 172100 449988
rect 172164 449986 172170 449988
rect 200070 449986 200130 451044
rect 356132 451016 358726 451072
rect 358782 451016 358787 451072
rect 356132 451014 358787 451016
rect 358721 451011 358787 451014
rect 172164 449926 200130 449986
rect 172164 449924 172170 449926
rect -960 449578 480 449668
rect 3141 449578 3207 449581
rect -960 449576 3207 449578
rect -960 449520 3146 449576
rect 3202 449520 3207 449576
rect -960 449518 3207 449520
rect -960 449428 480 449518
rect 3141 449515 3207 449518
rect 78029 448626 78095 448629
rect 128997 448626 129063 448629
rect 78029 448624 129063 448626
rect 78029 448568 78034 448624
rect 78090 448568 129002 448624
rect 129058 448568 129063 448624
rect 78029 448566 129063 448568
rect 78029 448563 78095 448566
rect 128997 448563 129063 448566
rect 197353 448626 197419 448629
rect 358721 448626 358787 448629
rect 197353 448624 200100 448626
rect 197353 448568 197358 448624
rect 197414 448568 200100 448624
rect 197353 448566 200100 448568
rect 356132 448624 358787 448626
rect 356132 448568 358726 448624
rect 358782 448568 358787 448624
rect 356132 448566 358787 448568
rect 197353 448563 197419 448566
rect 358721 448563 358787 448566
rect 84193 447266 84259 447269
rect 91502 447266 91508 447268
rect 84193 447264 91508 447266
rect 84193 447208 84198 447264
rect 84254 447208 91508 447264
rect 84193 447206 91508 447208
rect 84193 447203 84259 447206
rect 91502 447204 91508 447206
rect 91572 447204 91578 447268
rect 115289 447266 115355 447269
rect 115790 447266 115796 447268
rect 115289 447264 115796 447266
rect 115289 447208 115294 447264
rect 115350 447208 115796 447264
rect 115289 447206 115796 447208
rect 115289 447203 115355 447206
rect 115790 447204 115796 447206
rect 115860 447266 115866 447268
rect 124305 447266 124371 447269
rect 115860 447264 124371 447266
rect 115860 447208 124310 447264
rect 124366 447208 124371 447264
rect 115860 447206 124371 447208
rect 115860 447204 115866 447206
rect 124305 447203 124371 447206
rect 70209 447132 70275 447133
rect 70158 447130 70164 447132
rect 70118 447070 70164 447130
rect 70228 447128 70275 447132
rect 70270 447072 70275 447128
rect 70158 447068 70164 447070
rect 70228 447068 70275 447072
rect 70209 447067 70275 447068
rect 109033 447130 109099 447133
rect 148317 447130 148383 447133
rect 109033 447128 148383 447130
rect 109033 447072 109038 447128
rect 109094 447072 148322 447128
rect 148378 447072 148383 447128
rect 109033 447070 148383 447072
rect 109033 447067 109099 447070
rect 148317 447067 148383 447070
rect 70393 446450 70459 446453
rect 72366 446450 72372 446452
rect 70393 446448 72372 446450
rect 70393 446392 70398 446448
rect 70454 446392 72372 446448
rect 70393 446390 72372 446392
rect 70393 446387 70459 446390
rect 72366 446388 72372 446390
rect 72436 446388 72442 446452
rect 197353 446178 197419 446181
rect 357525 446178 357591 446181
rect 197353 446176 200100 446178
rect 197353 446120 197358 446176
rect 197414 446120 200100 446176
rect 197353 446118 200100 446120
rect 356132 446176 357591 446178
rect 356132 446120 357530 446176
rect 357586 446120 357591 446176
rect 356132 446118 357591 446120
rect 197353 446115 197419 446118
rect 357525 446115 357591 446118
rect 60641 445906 60707 445909
rect 68318 445906 68324 445908
rect 60641 445904 68324 445906
rect 60641 445848 60646 445904
rect 60702 445848 68324 445904
rect 60641 445846 68324 445848
rect 60641 445843 60707 445846
rect 68318 445844 68324 445846
rect 68388 445906 68394 445908
rect 68737 445906 68803 445909
rect 71773 445908 71839 445909
rect 71773 445906 71820 445908
rect 68388 445904 68803 445906
rect 68388 445848 68742 445904
rect 68798 445848 68803 445904
rect 68388 445846 68803 445848
rect 71728 445904 71820 445906
rect 71884 445906 71890 445908
rect 72734 445906 72740 445908
rect 71728 445848 71778 445904
rect 71728 445846 71820 445848
rect 68388 445844 68394 445846
rect 68737 445843 68803 445846
rect 71773 445844 71820 445846
rect 71884 445846 72740 445906
rect 71884 445844 71890 445846
rect 72734 445844 72740 445846
rect 72804 445844 72810 445908
rect 71773 445843 71839 445844
rect 55029 445770 55095 445773
rect 85573 445770 85639 445773
rect 55029 445768 85639 445770
rect 55029 445712 55034 445768
rect 55090 445712 85578 445768
rect 85634 445712 85639 445768
rect 55029 445710 85639 445712
rect 55029 445707 55095 445710
rect 85573 445707 85639 445710
rect 93894 445708 93900 445772
rect 93964 445770 93970 445772
rect 94773 445770 94839 445773
rect 93964 445768 94839 445770
rect 93964 445712 94778 445768
rect 94834 445712 94839 445768
rect 93964 445710 94839 445712
rect 93964 445708 93970 445710
rect 94773 445707 94839 445710
rect 96286 445708 96292 445772
rect 96356 445770 96362 445772
rect 96613 445770 96679 445773
rect 97625 445770 97691 445773
rect 96356 445768 97691 445770
rect 96356 445712 96618 445768
rect 96674 445712 97630 445768
rect 97686 445712 97691 445768
rect 96356 445710 97691 445712
rect 96356 445708 96362 445710
rect 96613 445707 96679 445710
rect 97625 445707 97691 445710
rect 100518 445708 100524 445772
rect 100588 445770 100594 445772
rect 100845 445770 100911 445773
rect 100588 445768 100911 445770
rect 100588 445712 100850 445768
rect 100906 445712 100911 445768
rect 100588 445710 100911 445712
rect 100588 445708 100594 445710
rect 100845 445707 100911 445710
rect 113173 445770 113239 445773
rect 114369 445772 114435 445773
rect 114318 445770 114324 445772
rect 113173 445768 114324 445770
rect 114388 445768 114435 445772
rect 113173 445712 113178 445768
rect 113234 445712 114324 445768
rect 114430 445712 114435 445768
rect 113173 445710 114324 445712
rect 113173 445707 113239 445710
rect 114318 445708 114324 445710
rect 114388 445708 114435 445712
rect 114369 445707 114435 445708
rect 117589 445770 117655 445773
rect 117998 445770 118004 445772
rect 117589 445768 118004 445770
rect 117589 445712 117594 445768
rect 117650 445712 118004 445768
rect 117589 445710 118004 445712
rect 117589 445707 117655 445710
rect 117998 445708 118004 445710
rect 118068 445770 118074 445772
rect 118601 445770 118667 445773
rect 118068 445768 118667 445770
rect 118068 445712 118606 445768
rect 118662 445712 118667 445768
rect 118068 445710 118667 445712
rect 118068 445708 118074 445710
rect 118601 445707 118667 445710
rect 96521 444954 96587 444957
rect 141417 444954 141483 444957
rect 96521 444952 141483 444954
rect 96521 444896 96526 444952
rect 96582 444896 141422 444952
rect 141478 444896 141483 444952
rect 96521 444894 141483 444896
rect 96521 444891 96587 444894
rect 141417 444891 141483 444894
rect 124857 444818 124923 444821
rect 103470 444816 124923 444818
rect 103470 444760 124862 444816
rect 124918 444760 124923 444816
rect 103470 444758 124923 444760
rect 87045 444682 87111 444685
rect 103470 444682 103530 444758
rect 124857 444755 124923 444758
rect 87045 444680 103530 444682
rect 87045 444624 87050 444680
rect 87106 444624 103530 444680
rect 87045 444622 103530 444624
rect 87045 444619 87111 444622
rect 108798 444620 108804 444684
rect 108868 444682 108874 444684
rect 109033 444682 109099 444685
rect 108868 444680 109099 444682
rect 108868 444624 109038 444680
rect 109094 444624 109099 444680
rect 108868 444622 109099 444624
rect 108868 444620 108874 444622
rect 109033 444619 109099 444622
rect 111558 444620 111564 444684
rect 111628 444682 111634 444684
rect 111701 444682 111767 444685
rect 111628 444680 111767 444682
rect 111628 444624 111706 444680
rect 111762 444624 111767 444680
rect 583520 444668 584960 444908
rect 111628 444622 111767 444624
rect 111628 444620 111634 444622
rect 111701 444619 111767 444622
rect 53741 444546 53807 444549
rect 79409 444546 79475 444549
rect 53741 444544 79475 444546
rect 53741 444488 53746 444544
rect 53802 444488 79414 444544
rect 79470 444488 79475 444544
rect 53741 444486 79475 444488
rect 53741 444483 53807 444486
rect 79409 444483 79475 444486
rect 83825 444546 83891 444549
rect 157977 444546 158043 444549
rect 83825 444544 158043 444546
rect 83825 444488 83830 444544
rect 83886 444488 157982 444544
rect 158038 444488 158043 444544
rect 83825 444486 158043 444488
rect 83825 444483 83891 444486
rect 157977 444483 158043 444486
rect 120582 443866 120642 444244
rect 124254 443866 124260 443868
rect 120582 443806 124260 443866
rect 124254 443804 124260 443806
rect 124324 443866 124330 443868
rect 125501 443866 125567 443869
rect 124324 443864 125567 443866
rect 124324 443808 125506 443864
rect 125562 443808 125567 443864
rect 124324 443806 125567 443808
rect 124324 443804 124330 443806
rect 125501 443803 125567 443806
rect 197353 443730 197419 443733
rect 358721 443730 358787 443733
rect 197353 443728 200100 443730
rect 197353 443672 197358 443728
rect 197414 443672 200100 443728
rect 197353 443670 200100 443672
rect 356132 443728 358787 443730
rect 356132 443672 358726 443728
rect 358782 443672 358787 443728
rect 356132 443670 358787 443672
rect 197353 443667 197419 443670
rect 358721 443667 358787 443670
rect 67817 442234 67883 442237
rect 121637 442234 121703 442237
rect 154062 442234 154068 442236
rect 67817 442232 68908 442234
rect 67817 442176 67822 442232
rect 67878 442176 68908 442232
rect 67817 442174 68908 442176
rect 121637 442232 154068 442234
rect 121637 442176 121642 442232
rect 121698 442176 154068 442232
rect 121637 442174 154068 442176
rect 67817 442171 67883 442174
rect 121637 442171 121703 442174
rect 154062 442172 154068 442174
rect 154132 442172 154138 442236
rect 124121 442098 124187 442101
rect 120612 442096 124187 442098
rect 120612 442040 124126 442096
rect 124182 442040 124187 442096
rect 120612 442038 124187 442040
rect 124121 442035 124187 442038
rect 197353 441418 197419 441421
rect 197353 441416 200100 441418
rect 197353 441360 197358 441416
rect 197414 441360 200100 441416
rect 197353 441358 200100 441360
rect 197353 441355 197419 441358
rect 358721 441282 358787 441285
rect 356132 441280 358787 441282
rect 356132 441224 358726 441280
rect 358782 441224 358787 441280
rect 356132 441222 358787 441224
rect 358721 441219 358787 441222
rect 121545 440058 121611 440061
rect 120612 440056 121611 440058
rect 120612 440000 121550 440056
rect 121606 440000 121611 440056
rect 120612 439998 121611 440000
rect 121545 439995 121611 439998
rect 67633 439922 67699 439925
rect 67633 439920 68908 439922
rect 67633 439864 67638 439920
rect 67694 439864 68908 439920
rect 67633 439862 68908 439864
rect 67633 439859 67699 439862
rect 197118 438908 197124 438972
rect 197188 438970 197194 438972
rect 358721 438970 358787 438973
rect 197188 438910 200100 438970
rect 356132 438968 358787 438970
rect 356132 438912 358726 438968
rect 358782 438912 358787 438968
rect 356132 438910 358787 438912
rect 197188 438908 197194 438910
rect 358721 438907 358787 438910
rect 66805 437882 66871 437885
rect 124121 437882 124187 437885
rect 66805 437880 68908 437882
rect 66805 437824 66810 437880
rect 66866 437824 68908 437880
rect 66805 437822 68908 437824
rect 120612 437880 124187 437882
rect 120612 437824 124126 437880
rect 124182 437824 124187 437880
rect 120612 437822 124187 437824
rect 66805 437819 66871 437822
rect 124121 437819 124187 437822
rect -960 436508 480 436748
rect 358721 436386 358787 436389
rect 356132 436384 358787 436386
rect 160870 436052 160876 436116
rect 160940 436114 160946 436116
rect 200070 436114 200130 436356
rect 356132 436328 358726 436384
rect 358782 436328 358787 436384
rect 356132 436326 358787 436328
rect 358721 436323 358787 436326
rect 160940 436054 200130 436114
rect 160940 436052 160946 436054
rect 66713 435434 66779 435437
rect 121545 435434 121611 435437
rect 122966 435434 122972 435436
rect 66713 435432 68908 435434
rect 66713 435376 66718 435432
rect 66774 435376 68908 435432
rect 66713 435374 68908 435376
rect 120612 435432 122972 435434
rect 120612 435376 121550 435432
rect 121606 435376 122972 435432
rect 120612 435374 122972 435376
rect 66713 435371 66779 435374
rect 121545 435371 121611 435374
rect 122966 435372 122972 435374
rect 123036 435372 123042 435436
rect 197353 433938 197419 433941
rect 358721 433938 358787 433941
rect 197353 433936 200100 433938
rect 197353 433880 197358 433936
rect 197414 433880 200100 433936
rect 197353 433878 200100 433880
rect 356132 433936 358787 433938
rect 356132 433880 358726 433936
rect 358782 433880 358787 433936
rect 356132 433878 358787 433880
rect 197353 433875 197419 433878
rect 358721 433875 358787 433878
rect 66805 433122 66871 433125
rect 124121 433122 124187 433125
rect 66805 433120 68908 433122
rect 66805 433064 66810 433120
rect 66866 433064 68908 433120
rect 66805 433062 68908 433064
rect 120612 433120 124187 433122
rect 120612 433064 124126 433120
rect 124182 433064 124187 433120
rect 120612 433062 124187 433064
rect 66805 433059 66871 433062
rect 124121 433059 124187 433062
rect 582833 431626 582899 431629
rect 583520 431626 584960 431716
rect 582833 431624 584960 431626
rect 582833 431568 582838 431624
rect 582894 431568 584960 431624
rect 582833 431566 584960 431568
rect 582833 431563 582899 431566
rect 358721 431490 358787 431493
rect 356132 431488 358787 431490
rect 66805 431082 66871 431085
rect 124121 431082 124187 431085
rect 66805 431080 68908 431082
rect 66805 431024 66810 431080
rect 66866 431024 68908 431080
rect 66805 431022 68908 431024
rect 120612 431080 124187 431082
rect 120612 431024 124126 431080
rect 124182 431024 124187 431080
rect 120612 431022 124187 431024
rect 66805 431019 66871 431022
rect 124121 431019 124187 431022
rect 186814 430612 186820 430676
rect 186884 430674 186890 430676
rect 200070 430674 200130 431460
rect 356132 431432 358726 431488
rect 358782 431432 358787 431488
rect 583520 431476 584960 431566
rect 356132 431430 358787 431432
rect 358721 431427 358787 431430
rect 186884 430614 200130 430674
rect 186884 430612 186890 430614
rect 120717 429314 120783 429317
rect 120582 429312 120783 429314
rect 120582 429256 120722 429312
rect 120778 429256 120783 429312
rect 120582 429254 120783 429256
rect 66805 428634 66871 428637
rect 66805 428632 68908 428634
rect 66805 428576 66810 428632
rect 66866 428576 68908 428632
rect 66805 428574 68908 428576
rect 66805 428571 66871 428574
rect 120582 428498 120642 429254
rect 120717 429251 120783 429254
rect 197353 429042 197419 429045
rect 358721 429042 358787 429045
rect 197353 429040 200100 429042
rect 197353 428984 197358 429040
rect 197414 428984 200100 429040
rect 197353 428982 200100 428984
rect 356132 429040 358787 429042
rect 356132 428984 358726 429040
rect 358782 428984 358787 429040
rect 356132 428982 358787 428984
rect 197353 428979 197419 428982
rect 358721 428979 358787 428982
rect 122741 428498 122807 428501
rect 120582 428496 122807 428498
rect 120582 428468 122746 428496
rect 120612 428440 122746 428468
rect 122802 428440 122807 428496
rect 120612 428438 122807 428440
rect 122741 428435 122807 428438
rect 197353 426594 197419 426597
rect 357525 426594 357591 426597
rect 197353 426592 200100 426594
rect 197353 426536 197358 426592
rect 197414 426536 200100 426592
rect 197353 426534 200100 426536
rect 356132 426592 357591 426594
rect 356132 426536 357530 426592
rect 357586 426536 357591 426592
rect 356132 426534 357591 426536
rect 197353 426531 197419 426534
rect 357525 426531 357591 426534
rect 66713 426322 66779 426325
rect 66713 426320 68908 426322
rect 66713 426264 66718 426320
rect 66774 426264 68908 426320
rect 66713 426262 68908 426264
rect 66713 426259 66779 426262
rect 120030 426052 120090 426292
rect 120022 425988 120028 426052
rect 120092 426050 120098 426052
rect 123477 426050 123543 426053
rect 120092 426048 123543 426050
rect 120092 425992 123482 426048
rect 123538 425992 123543 426048
rect 120092 425990 123543 425992
rect 120092 425988 120098 425990
rect 123477 425987 123543 425990
rect 66805 424146 66871 424149
rect 123017 424146 123083 424149
rect 66805 424144 68908 424146
rect 66805 424088 66810 424144
rect 66866 424088 68908 424144
rect 66805 424086 68908 424088
rect 120612 424144 123083 424146
rect 120612 424088 123022 424144
rect 123078 424088 123083 424144
rect 120612 424086 123083 424088
rect 66805 424083 66871 424086
rect 123017 424083 123083 424086
rect 197353 424146 197419 424149
rect 358721 424146 358787 424149
rect 197353 424144 200100 424146
rect 197353 424088 197358 424144
rect 197414 424088 200100 424144
rect 197353 424086 200100 424088
rect 356132 424144 358787 424146
rect 356132 424088 358726 424144
rect 358782 424088 358787 424144
rect 356132 424086 358787 424088
rect 197353 424083 197419 424086
rect 358721 424083 358787 424086
rect -960 423602 480 423692
rect 3417 423602 3483 423605
rect -960 423600 3483 423602
rect -960 423544 3422 423600
rect 3478 423544 3483 423600
rect -960 423542 3483 423544
rect -960 423452 480 423542
rect 3417 423539 3483 423542
rect 66253 421970 66319 421973
rect 122925 421970 122991 421973
rect 66253 421968 68908 421970
rect 66253 421912 66258 421968
rect 66314 421912 68908 421968
rect 66253 421910 68908 421912
rect 120612 421968 122991 421970
rect 120612 421912 122930 421968
rect 122986 421912 122991 421968
rect 120612 421910 122991 421912
rect 66253 421907 66319 421910
rect 122925 421907 122991 421910
rect 197854 421636 197860 421700
rect 197924 421698 197930 421700
rect 358721 421698 358787 421701
rect 197924 421638 200100 421698
rect 356132 421696 358787 421698
rect 356132 421640 358726 421696
rect 358782 421640 358787 421696
rect 356132 421638 358787 421640
rect 197924 421636 197930 421638
rect 358721 421635 358787 421638
rect 121494 420820 121500 420884
rect 121564 420882 121570 420884
rect 124121 420882 124187 420885
rect 121564 420880 124187 420882
rect 121564 420824 124126 420880
rect 124182 420824 124187 420880
rect 121564 420822 124187 420824
rect 121564 420820 121570 420822
rect 124121 420819 124187 420822
rect 66662 419596 66668 419660
rect 66732 419658 66738 419660
rect 67725 419658 67791 419661
rect 121494 419658 121500 419660
rect 66732 419656 68908 419658
rect 66732 419600 67730 419656
rect 67786 419600 68908 419656
rect 66732 419598 68908 419600
rect 120612 419598 121500 419658
rect 66732 419596 66738 419598
rect 67725 419595 67791 419598
rect 121494 419596 121500 419598
rect 121564 419596 121570 419660
rect 197353 419250 197419 419253
rect 358721 419250 358787 419253
rect 197353 419248 200100 419250
rect 197353 419192 197358 419248
rect 197414 419192 200100 419248
rect 197353 419190 200100 419192
rect 356132 419248 358787 419250
rect 356132 419192 358726 419248
rect 358782 419192 358787 419248
rect 356132 419190 358787 419192
rect 197353 419187 197419 419190
rect 358721 419187 358787 419190
rect 582373 418298 582439 418301
rect 583520 418298 584960 418388
rect 582373 418296 584960 418298
rect 582373 418240 582378 418296
rect 582434 418240 584960 418296
rect 582373 418238 584960 418240
rect 582373 418235 582439 418238
rect 583520 418148 584960 418238
rect 68878 416802 68938 417316
rect 120582 417074 120642 417316
rect 120717 417074 120783 417077
rect 120582 417072 120783 417074
rect 120582 417016 120722 417072
rect 120778 417016 120783 417072
rect 120582 417014 120783 417016
rect 120717 417011 120783 417014
rect 66854 416742 68938 416802
rect 198917 416802 198983 416805
rect 357617 416802 357683 416805
rect 198917 416800 200100 416802
rect 198917 416744 198922 416800
rect 198978 416744 200100 416800
rect 198917 416742 200100 416744
rect 356132 416800 357683 416802
rect 356132 416744 357622 416800
rect 357678 416744 357683 416800
rect 356132 416742 357683 416744
rect 62849 416666 62915 416669
rect 66854 416666 66914 416742
rect 198917 416739 198983 416742
rect 357617 416739 357683 416742
rect 62849 416664 66914 416666
rect 62849 416608 62854 416664
rect 62910 416608 66914 416664
rect 62849 416606 66914 416608
rect 62849 416603 62915 416606
rect 41321 415442 41387 415445
rect 53649 415442 53715 415445
rect 62849 415442 62915 415445
rect 63401 415442 63467 415445
rect 41321 415440 63467 415442
rect 41321 415384 41326 415440
rect 41382 415384 53654 415440
rect 53710 415384 62854 415440
rect 62910 415384 63406 415440
rect 63462 415384 63467 415440
rect 41321 415382 63467 415384
rect 41321 415379 41387 415382
rect 53649 415379 53715 415382
rect 62849 415379 62915 415382
rect 63401 415379 63467 415382
rect 121177 415306 121243 415309
rect 120612 415304 121243 415306
rect 120612 415276 121182 415304
rect 120582 415248 121182 415276
rect 121238 415248 121243 415304
rect 120582 415246 121243 415248
rect 66805 415170 66871 415173
rect 66805 415168 68908 415170
rect 66805 415112 66810 415168
rect 66866 415112 68908 415168
rect 66805 415110 68908 415112
rect 66805 415107 66871 415110
rect 120582 414629 120642 415246
rect 121177 415243 121243 415246
rect 120582 414624 120691 414629
rect 120582 414568 120630 414624
rect 120686 414568 120691 414624
rect 120582 414566 120691 414568
rect 120625 414563 120691 414566
rect 197353 414354 197419 414357
rect 358721 414354 358787 414357
rect 197353 414352 200100 414354
rect 197353 414296 197358 414352
rect 197414 414296 200100 414352
rect 197353 414294 200100 414296
rect 356132 414352 358787 414354
rect 356132 414296 358726 414352
rect 358782 414296 358787 414352
rect 356132 414294 358787 414296
rect 197353 414291 197419 414294
rect 358721 414291 358787 414294
rect 67449 412858 67515 412861
rect 123845 412858 123911 412861
rect 67449 412856 68908 412858
rect 67449 412800 67454 412856
rect 67510 412800 68908 412856
rect 67449 412798 68908 412800
rect 120612 412856 123911 412858
rect 120612 412800 123850 412856
rect 123906 412800 123911 412856
rect 120612 412798 123911 412800
rect 67449 412795 67515 412798
rect 123845 412795 123911 412798
rect 197353 411906 197419 411909
rect 358721 411906 358787 411909
rect 197353 411904 200100 411906
rect 197353 411848 197358 411904
rect 197414 411848 200100 411904
rect 197353 411846 200100 411848
rect 356132 411904 358787 411906
rect 356132 411848 358726 411904
rect 358782 411848 358787 411904
rect 356132 411846 358787 411848
rect 197353 411843 197419 411846
rect 358721 411843 358787 411846
rect 66897 410682 66963 410685
rect 123569 410682 123635 410685
rect 66897 410680 68908 410682
rect -960 410546 480 410636
rect 66897 410624 66902 410680
rect 66958 410624 68908 410680
rect 66897 410622 68908 410624
rect 120612 410680 123635 410682
rect 120612 410624 123574 410680
rect 123630 410624 123635 410680
rect 120612 410622 123635 410624
rect 66897 410619 66963 410622
rect 123569 410619 123635 410622
rect 3417 410546 3483 410549
rect -960 410544 3483 410546
rect -960 410488 3422 410544
rect 3478 410488 3483 410544
rect -960 410486 3483 410488
rect -960 410396 480 410486
rect 3417 410483 3483 410486
rect 197353 409594 197419 409597
rect 197353 409592 200100 409594
rect 197353 409536 197358 409592
rect 197414 409536 200100 409592
rect 197353 409534 200100 409536
rect 197353 409531 197419 409534
rect 358721 409458 358787 409461
rect 356132 409456 358787 409458
rect 356132 409400 358726 409456
rect 358782 409400 358787 409456
rect 356132 409398 358787 409400
rect 358721 409395 358787 409398
rect 124121 408370 124187 408373
rect 120612 408368 124187 408370
rect 69246 407828 69306 408340
rect 120612 408312 124126 408368
rect 124182 408312 124187 408368
rect 120612 408310 124187 408312
rect 124121 408307 124187 408310
rect 69238 407764 69244 407828
rect 69308 407764 69314 407828
rect 131757 407826 131823 407829
rect 165654 407826 165660 407828
rect 131757 407824 165660 407826
rect 131757 407768 131762 407824
rect 131818 407768 165660 407824
rect 131757 407766 165660 407768
rect 131757 407763 131823 407766
rect 165654 407764 165660 407766
rect 165724 407764 165730 407828
rect 56501 407146 56567 407149
rect 69238 407146 69244 407148
rect 56501 407144 69244 407146
rect 56501 407088 56506 407144
rect 56562 407088 69244 407144
rect 56501 407086 69244 407088
rect 56501 407083 56567 407086
rect 69238 407084 69244 407086
rect 69308 407084 69314 407148
rect 197353 407010 197419 407013
rect 358997 407010 359063 407013
rect 197353 407008 200100 407010
rect 197353 406952 197358 407008
rect 197414 406952 200100 407008
rect 197353 406950 200100 406952
rect 356132 407008 359063 407010
rect 356132 406952 359002 407008
rect 359058 406952 359063 407008
rect 356132 406950 359063 406952
rect 197353 406947 197419 406950
rect 358997 406947 359063 406950
rect 66253 406194 66319 406197
rect 124121 406194 124187 406197
rect 66253 406192 68908 406194
rect 66253 406136 66258 406192
rect 66314 406136 68908 406192
rect 66253 406134 68908 406136
rect 120612 406192 124187 406194
rect 120612 406136 124126 406192
rect 124182 406136 124187 406192
rect 120612 406134 124187 406136
rect 66253 406131 66319 406134
rect 124121 406131 124187 406134
rect 582741 404970 582807 404973
rect 583520 404970 584960 405060
rect 582741 404968 584960 404970
rect 582741 404912 582746 404968
rect 582802 404912 584960 404968
rect 582741 404910 584960 404912
rect 582741 404907 582807 404910
rect 583520 404820 584960 404910
rect 192702 404500 192708 404564
rect 192772 404562 192778 404564
rect 192772 404502 200100 404562
rect 192772 404500 192778 404502
rect 358721 404290 358787 404293
rect 356132 404288 358787 404290
rect 356132 404232 358726 404288
rect 358782 404232 358787 404288
rect 356132 404230 358787 404232
rect 358721 404227 358787 404230
rect 66253 403746 66319 403749
rect 122598 403746 122604 403748
rect 66253 403744 68908 403746
rect 66253 403688 66258 403744
rect 66314 403688 68908 403744
rect 66253 403686 68908 403688
rect 120612 403686 122604 403746
rect 66253 403683 66319 403686
rect 122598 403684 122604 403686
rect 122668 403746 122674 403748
rect 123753 403746 123819 403749
rect 122668 403744 123819 403746
rect 122668 403688 123758 403744
rect 123814 403688 123819 403744
rect 122668 403686 123819 403688
rect 122668 403684 122674 403686
rect 123753 403683 123819 403686
rect 197353 402114 197419 402117
rect 197353 402112 200100 402114
rect 197353 402056 197358 402112
rect 197414 402056 200100 402112
rect 197353 402054 200100 402056
rect 197353 402051 197419 402054
rect 358721 401842 358787 401845
rect 356132 401840 358787 401842
rect 356132 401784 358726 401840
rect 358782 401784 358787 401840
rect 356132 401782 358787 401784
rect 358721 401779 358787 401782
rect 66253 401570 66319 401573
rect 124121 401570 124187 401573
rect 66253 401568 68908 401570
rect 66253 401512 66258 401568
rect 66314 401512 68908 401568
rect 66253 401510 68908 401512
rect 120612 401568 124187 401570
rect 120612 401512 124126 401568
rect 124182 401512 124187 401568
rect 120612 401510 124187 401512
rect 66253 401507 66319 401510
rect 124121 401507 124187 401510
rect 197353 399666 197419 399669
rect 197353 399664 200100 399666
rect 197353 399608 197358 399664
rect 197414 399608 200100 399664
rect 197353 399606 200100 399608
rect 197353 399603 197419 399606
rect 66253 399530 66319 399533
rect 124121 399530 124187 399533
rect 66253 399528 68908 399530
rect 66253 399472 66258 399528
rect 66314 399472 68908 399528
rect 66253 399470 68908 399472
rect 120612 399528 124187 399530
rect 120612 399472 124126 399528
rect 124182 399472 124187 399528
rect 120612 399470 124187 399472
rect 66253 399467 66319 399470
rect 124121 399467 124187 399470
rect 357985 399394 358051 399397
rect 356132 399392 358051 399394
rect 356132 399336 357990 399392
rect 358046 399336 358051 399392
rect 356132 399334 358051 399336
rect 357985 399331 358051 399334
rect -960 397490 480 397580
rect 2773 397490 2839 397493
rect -960 397488 2839 397490
rect -960 397432 2778 397488
rect 2834 397432 2839 397488
rect -960 397430 2839 397432
rect -960 397340 480 397430
rect 2773 397427 2839 397430
rect 123017 397354 123083 397357
rect 124121 397354 124187 397357
rect 120582 397352 124187 397354
rect 120582 397296 123022 397352
rect 123078 397296 124126 397352
rect 124182 397296 124187 397352
rect 120582 397294 124187 397296
rect 120582 397052 120642 397294
rect 123017 397291 123083 397294
rect 124121 397291 124187 397294
rect 197353 397218 197419 397221
rect 197353 397216 200100 397218
rect 197353 397160 197358 397216
rect 197414 397160 200100 397216
rect 197353 397158 200100 397160
rect 197353 397155 197419 397158
rect 66989 396946 67055 396949
rect 358721 396946 358787 396949
rect 66989 396944 68908 396946
rect 66989 396888 66994 396944
rect 67050 396888 68908 396944
rect 66989 396886 68908 396888
rect 356132 396944 358787 396946
rect 356132 396888 358726 396944
rect 358782 396888 358787 396944
rect 356132 396886 358787 396888
rect 66989 396883 67055 396886
rect 358721 396883 358787 396886
rect 67541 394906 67607 394909
rect 67541 394904 68908 394906
rect 67541 394848 67546 394904
rect 67602 394848 68908 394904
rect 67541 394846 68908 394848
rect 67541 394843 67607 394846
rect 122925 394770 122991 394773
rect 120612 394768 122991 394770
rect 120612 394712 122930 394768
rect 122986 394712 122991 394768
rect 120612 394710 122991 394712
rect 122925 394707 122991 394710
rect 197353 394770 197419 394773
rect 197353 394768 200100 394770
rect 197353 394712 197358 394768
rect 197414 394712 200100 394768
rect 197353 394710 200100 394712
rect 197353 394707 197419 394710
rect 356462 394498 356468 394500
rect 356132 394438 356468 394498
rect 356462 394436 356468 394438
rect 356532 394436 356538 394500
rect 198457 393410 198523 393413
rect 198590 393410 198596 393412
rect 198457 393408 198596 393410
rect 198457 393352 198462 393408
rect 198518 393352 198596 393408
rect 198457 393350 198596 393352
rect 198457 393347 198523 393350
rect 198590 393348 198596 393350
rect 198660 393348 198666 393412
rect 121453 392730 121519 392733
rect 120612 392728 121519 392730
rect 120612 392672 121458 392728
rect 121514 392672 121519 392728
rect 120612 392670 121519 392672
rect 121453 392667 121519 392670
rect 66621 392594 66687 392597
rect 66621 392592 68908 392594
rect 66621 392536 66626 392592
rect 66682 392536 68908 392592
rect 66621 392534 68908 392536
rect 66621 392531 66687 392534
rect 197353 392322 197419 392325
rect 198457 392322 198523 392325
rect 197353 392320 200100 392322
rect 197353 392264 197358 392320
rect 197414 392264 198462 392320
rect 198518 392264 200100 392320
rect 197353 392262 200100 392264
rect 197353 392259 197419 392262
rect 198457 392259 198523 392262
rect 357709 392050 357775 392053
rect 356132 392048 357775 392050
rect 356132 391992 357714 392048
rect 357770 391992 357775 392048
rect 356132 391990 357775 391992
rect 357709 391987 357775 391990
rect 72366 391852 72372 391916
rect 72436 391914 72442 391916
rect 73102 391914 73108 391916
rect 72436 391854 73108 391914
rect 72436 391852 72442 391854
rect 73102 391852 73108 391854
rect 73172 391914 73178 391916
rect 144177 391914 144243 391917
rect 73172 391912 144243 391914
rect 73172 391856 144182 391912
rect 144238 391856 144243 391912
rect 73172 391854 144243 391856
rect 73172 391852 73178 391854
rect 144177 391851 144243 391854
rect 583520 391628 584960 391868
rect 64781 391234 64847 391237
rect 64781 391232 64890 391234
rect 64781 391176 64786 391232
rect 64842 391176 64890 391232
rect 64781 391171 64890 391176
rect 64830 391098 64890 391171
rect 77661 391098 77727 391101
rect 92933 391100 92999 391101
rect 92933 391098 92980 391100
rect 64830 391096 77727 391098
rect 64830 391040 77666 391096
rect 77722 391040 77727 391096
rect 64830 391038 77727 391040
rect 92888 391096 92980 391098
rect 92888 391040 92938 391096
rect 92888 391038 92980 391040
rect 77661 391035 77727 391038
rect 92933 391036 92980 391038
rect 93044 391036 93050 391100
rect 92933 391035 92999 391036
rect 115749 390690 115815 390693
rect 121494 390690 121500 390692
rect 115749 390688 121500 390690
rect 115749 390632 115754 390688
rect 115810 390632 121500 390688
rect 115749 390630 121500 390632
rect 115749 390627 115815 390630
rect 121494 390628 121500 390630
rect 121564 390628 121570 390692
rect 69606 390356 69612 390420
rect 69676 390418 69682 390420
rect 69933 390418 69999 390421
rect 69676 390416 69999 390418
rect 69676 390360 69938 390416
rect 69994 390360 69999 390416
rect 69676 390358 69999 390360
rect 69676 390356 69682 390358
rect 69933 390355 69999 390358
rect 89662 390356 89668 390420
rect 89732 390418 89738 390420
rect 89805 390418 89871 390421
rect 89732 390416 89871 390418
rect 89732 390360 89810 390416
rect 89866 390360 89871 390416
rect 89732 390358 89871 390360
rect 89732 390356 89738 390358
rect 89805 390355 89871 390358
rect 94078 390356 94084 390420
rect 94148 390418 94154 390420
rect 94221 390418 94287 390421
rect 94148 390416 94287 390418
rect 94148 390360 94226 390416
rect 94282 390360 94287 390416
rect 94148 390358 94287 390360
rect 94148 390356 94154 390358
rect 94221 390355 94287 390358
rect 96654 390356 96660 390420
rect 96724 390418 96730 390420
rect 97349 390418 97415 390421
rect 96724 390416 97415 390418
rect 96724 390360 97354 390416
rect 97410 390360 97415 390416
rect 96724 390358 97415 390360
rect 96724 390356 96730 390358
rect 97349 390355 97415 390358
rect 98126 390356 98132 390420
rect 98196 390418 98202 390420
rect 98821 390418 98887 390421
rect 98196 390416 98887 390418
rect 98196 390360 98826 390416
rect 98882 390360 98887 390416
rect 98196 390358 98887 390360
rect 98196 390356 98202 390358
rect 98821 390355 98887 390358
rect 102133 390420 102199 390421
rect 104985 390420 105051 390421
rect 102133 390416 102180 390420
rect 102244 390418 102250 390420
rect 104934 390418 104940 390420
rect 102133 390360 102138 390416
rect 102133 390356 102180 390360
rect 102244 390358 102290 390418
rect 104894 390358 104940 390418
rect 105004 390416 105051 390420
rect 105046 390360 105051 390416
rect 102244 390356 102250 390358
rect 104934 390356 104940 390358
rect 105004 390356 105051 390360
rect 106406 390356 106412 390420
rect 106476 390418 106482 390420
rect 106549 390418 106615 390421
rect 106476 390416 106615 390418
rect 106476 390360 106554 390416
rect 106610 390360 106615 390416
rect 106476 390358 106615 390360
rect 106476 390356 106482 390358
rect 102133 390355 102199 390356
rect 104985 390355 105051 390356
rect 106549 390355 106615 390358
rect 107694 390356 107700 390420
rect 107764 390418 107770 390420
rect 108021 390418 108087 390421
rect 107764 390416 108087 390418
rect 107764 390360 108026 390416
rect 108082 390360 108087 390416
rect 107764 390358 108087 390360
rect 107764 390356 107770 390358
rect 108021 390355 108087 390358
rect 108982 390356 108988 390420
rect 109052 390418 109058 390420
rect 109493 390418 109559 390421
rect 109052 390416 109559 390418
rect 109052 390360 109498 390416
rect 109554 390360 109559 390416
rect 109052 390358 109559 390360
rect 109052 390356 109058 390358
rect 109493 390355 109559 390358
rect 115933 390420 115999 390421
rect 115933 390416 115980 390420
rect 116044 390418 116050 390420
rect 117865 390418 117931 390421
rect 118785 390420 118851 390421
rect 118182 390418 118188 390420
rect 115933 390360 115938 390416
rect 115933 390356 115980 390360
rect 116044 390358 116090 390418
rect 117865 390416 118188 390418
rect 117865 390360 117870 390416
rect 117926 390360 118188 390416
rect 117865 390358 118188 390360
rect 116044 390356 116050 390358
rect 115933 390355 115999 390356
rect 117865 390355 117931 390358
rect 118182 390356 118188 390358
rect 118252 390356 118258 390420
rect 118734 390418 118740 390420
rect 118694 390358 118740 390418
rect 118804 390416 118851 390420
rect 118846 390360 118851 390416
rect 118734 390356 118740 390358
rect 118804 390356 118851 390360
rect 118785 390355 118851 390356
rect 100753 390284 100819 390285
rect 100702 390282 100708 390284
rect 100662 390222 100708 390282
rect 100772 390280 100819 390284
rect 100814 390224 100819 390280
rect 100702 390220 100708 390222
rect 100772 390220 100819 390224
rect 100753 390219 100819 390220
rect 68645 389330 68711 389333
rect 70894 389330 70900 389332
rect 68645 389328 70900 389330
rect 68645 389272 68650 389328
rect 68706 389272 70900 389328
rect 68645 389270 70900 389272
rect 68645 389267 68711 389270
rect 70894 389268 70900 389270
rect 70964 389268 70970 389332
rect 108389 389330 108455 389333
rect 169702 389330 169708 389332
rect 108389 389328 169708 389330
rect 108389 389272 108394 389328
rect 108450 389272 169708 389328
rect 108389 389270 169708 389272
rect 108389 389267 108455 389270
rect 169702 389268 169708 389270
rect 169772 389268 169778 389332
rect 63401 389194 63467 389197
rect 200070 389194 200130 389844
rect 356102 389332 356162 389572
rect 356094 389268 356100 389332
rect 356164 389268 356170 389332
rect 63401 389192 200130 389194
rect 63401 389136 63406 389192
rect 63462 389136 200130 389192
rect 63401 389134 200130 389136
rect 63401 389131 63467 389134
rect 65793 389058 65859 389061
rect 68134 389058 68140 389060
rect 65793 389056 68140 389058
rect 65793 389000 65798 389056
rect 65854 389000 68140 389056
rect 65793 388998 68140 389000
rect 65793 388995 65859 388998
rect 68134 388996 68140 388998
rect 68204 389058 68210 389060
rect 68737 389058 68803 389061
rect 68204 389056 68803 389058
rect 68204 389000 68742 389056
rect 68798 389000 68803 389056
rect 68204 388998 68803 389000
rect 68204 388996 68210 388998
rect 68737 388995 68803 388998
rect 71773 389058 71839 389061
rect 73061 389060 73127 389061
rect 73061 389058 73108 389060
rect 71773 389056 73108 389058
rect 73172 389058 73178 389060
rect 81433 389058 81499 389061
rect 71773 389000 71778 389056
rect 71834 389000 73066 389056
rect 71773 388998 73108 389000
rect 71773 388995 71839 388998
rect 73061 388996 73108 388998
rect 73172 388998 73254 389058
rect 81433 389056 84210 389058
rect 81433 389000 81438 389056
rect 81494 389000 84210 389056
rect 81433 388998 84210 389000
rect 73172 388996 73178 388998
rect 73061 388995 73127 388996
rect 81433 388995 81499 388998
rect 65885 388922 65951 388925
rect 73153 388922 73219 388925
rect 73797 388922 73863 388925
rect 65885 388920 73863 388922
rect 65885 388864 65890 388920
rect 65946 388864 73158 388920
rect 73214 388864 73802 388920
rect 73858 388864 73863 388920
rect 65885 388862 73863 388864
rect 84150 388922 84210 388998
rect 90214 388996 90220 389060
rect 90284 389058 90290 389060
rect 91645 389058 91711 389061
rect 95233 389058 95299 389061
rect 96245 389058 96311 389061
rect 90284 389056 91711 389058
rect 90284 389000 91650 389056
rect 91706 389000 91711 389056
rect 90284 388998 91711 389000
rect 90284 388996 90290 388998
rect 91645 388995 91711 388998
rect 93810 389056 96311 389058
rect 93810 389000 95238 389056
rect 95294 389000 96250 389056
rect 96306 389000 96311 389056
rect 93810 388998 96311 389000
rect 90449 388922 90515 388925
rect 84150 388920 90515 388922
rect 84150 388864 90454 388920
rect 90510 388864 90515 388920
rect 84150 388862 90515 388864
rect 65885 388859 65951 388862
rect 73153 388859 73219 388862
rect 73797 388859 73863 388862
rect 90449 388859 90515 388862
rect 91502 388860 91508 388924
rect 91572 388922 91578 388924
rect 93810 388922 93870 388998
rect 95233 388995 95299 388998
rect 96245 388995 96311 388998
rect 99189 389058 99255 389061
rect 100753 389058 100819 389061
rect 99189 389056 100819 389058
rect 99189 389000 99194 389056
rect 99250 389000 100758 389056
rect 100814 389000 100819 389056
rect 99189 388998 100819 389000
rect 99189 388995 99255 388998
rect 100753 388995 100819 388998
rect 102317 389058 102383 389061
rect 103329 389058 103395 389061
rect 102317 389056 103395 389058
rect 102317 389000 102322 389056
rect 102378 389000 103334 389056
rect 103390 389000 103395 389056
rect 102317 388998 103395 389000
rect 102317 388995 102383 388998
rect 103329 388995 103395 388998
rect 111742 388996 111748 389060
rect 111812 389058 111818 389060
rect 112897 389058 112963 389061
rect 111812 389056 112963 389058
rect 111812 389000 112902 389056
rect 112958 389000 112963 389056
rect 111812 388998 112963 389000
rect 111812 388996 111818 388998
rect 112897 388995 112963 388998
rect 113173 389060 113239 389061
rect 113173 389056 113220 389060
rect 113284 389058 113290 389060
rect 114369 389058 114435 389061
rect 113284 389056 114435 389058
rect 113173 389000 113178 389056
rect 113284 389000 114374 389056
rect 114430 389000 114435 389056
rect 113173 388996 113220 389000
rect 113284 388998 114435 389000
rect 113284 388996 113290 388998
rect 113173 388995 113239 388996
rect 114369 388995 114435 388998
rect 91572 388862 93870 388922
rect 91572 388860 91578 388862
rect 65609 388786 65675 388789
rect 79501 388786 79567 388789
rect 65609 388784 79567 388786
rect 65609 388728 65614 388784
rect 65670 388728 79506 388784
rect 79562 388728 79567 388784
rect 65609 388726 79567 388728
rect 65609 388723 65675 388726
rect 79501 388723 79567 388726
rect 93025 388786 93091 388789
rect 101397 388786 101463 388789
rect 93025 388784 101463 388786
rect 93025 388728 93030 388784
rect 93086 388728 101402 388784
rect 101458 388728 101463 388784
rect 93025 388726 101463 388728
rect 93025 388723 93091 388726
rect 101397 388723 101463 388726
rect 106917 388378 106983 388381
rect 120441 388378 120507 388381
rect 106917 388376 120507 388378
rect 106917 388320 106922 388376
rect 106978 388320 120446 388376
rect 120502 388320 120507 388376
rect 106917 388318 120507 388320
rect 106917 388315 106983 388318
rect 120441 388315 120507 388318
rect 197353 387426 197419 387429
rect 197353 387424 200100 387426
rect 197353 387368 197358 387424
rect 197414 387368 200100 387424
rect 197353 387366 200100 387368
rect 197353 387363 197419 387366
rect 63309 387018 63375 387021
rect 79961 387018 80027 387021
rect 80881 387018 80947 387021
rect 63309 387016 80947 387018
rect 63309 386960 63314 387016
rect 63370 386960 79966 387016
rect 80022 386960 80886 387016
rect 80942 386960 80947 387016
rect 63309 386958 80947 386960
rect 63309 386955 63375 386958
rect 79961 386955 80027 386958
rect 80881 386955 80947 386958
rect 120717 387018 120783 387021
rect 196617 387018 196683 387021
rect 120717 387016 196683 387018
rect 120717 386960 120722 387016
rect 120778 386960 196622 387016
rect 196678 386960 196683 387016
rect 120717 386958 196683 386960
rect 120717 386955 120783 386958
rect 196617 386955 196683 386958
rect 356102 386612 356162 387124
rect 356094 386548 356100 386612
rect 356164 386548 356170 386612
rect 76373 385658 76439 385661
rect 169753 385658 169819 385661
rect 76373 385656 169819 385658
rect 76373 385600 76378 385656
rect 76434 385600 169758 385656
rect 169814 385600 169819 385656
rect 76373 385598 169819 385600
rect 76373 385595 76439 385598
rect 169753 385595 169819 385598
rect 197261 384978 197327 384981
rect 197261 384976 200100 384978
rect 197261 384920 197266 384976
rect 197322 384920 200100 384976
rect 197261 384918 200100 384920
rect 197261 384915 197327 384918
rect 195830 384780 195836 384844
rect 195900 384842 195906 384844
rect 199377 384842 199443 384845
rect 195900 384840 199443 384842
rect 195900 384784 199382 384840
rect 199438 384784 199443 384840
rect 195900 384782 199443 384784
rect 195900 384780 195906 384782
rect 199377 384779 199443 384782
rect 363086 384706 363092 384708
rect 356132 384646 363092 384706
rect 363086 384644 363092 384646
rect 363156 384644 363162 384708
rect -960 384284 480 384524
rect 39849 384298 39915 384301
rect 122925 384298 122991 384301
rect 39849 384296 122991 384298
rect 39849 384240 39854 384296
rect 39910 384240 122930 384296
rect 122986 384240 122991 384296
rect 39849 384238 122991 384240
rect 39849 384235 39915 384238
rect 122925 384235 122991 384238
rect 356278 383964 356284 384028
rect 356348 383964 356354 384028
rect 15837 383754 15903 383757
rect 119337 383754 119403 383757
rect 356286 383756 356346 383964
rect 15837 383752 119403 383754
rect 15837 383696 15842 383752
rect 15898 383696 119342 383752
rect 119398 383696 119403 383752
rect 15837 383694 119403 383696
rect 15837 383691 15903 383694
rect 119337 383691 119403 383694
rect 356278 383692 356284 383756
rect 356348 383692 356354 383756
rect 75821 382938 75887 382941
rect 193949 382938 194015 382941
rect 75821 382936 194015 382938
rect 75821 382880 75826 382936
rect 75882 382880 193954 382936
rect 194010 382880 194015 382936
rect 75821 382878 194015 382880
rect 75821 382875 75887 382878
rect 193949 382875 194015 382878
rect 199009 382530 199075 382533
rect 199009 382528 200100 382530
rect 199009 382472 199014 382528
rect 199070 382472 200100 382528
rect 199009 382470 200100 382472
rect 199009 382467 199075 382470
rect 358813 382394 358879 382397
rect 356132 382392 358879 382394
rect 356132 382336 358818 382392
rect 358874 382336 358879 382392
rect 356132 382334 358879 382336
rect 358813 382331 358879 382334
rect 106181 381578 106247 381581
rect 121545 381578 121611 381581
rect 106181 381576 121611 381578
rect 106181 381520 106186 381576
rect 106242 381520 121550 381576
rect 121606 381520 121611 381576
rect 106181 381518 121611 381520
rect 106181 381515 106247 381518
rect 121545 381515 121611 381518
rect 356094 381516 356100 381580
rect 356164 381578 356170 381580
rect 356462 381578 356468 381580
rect 356164 381518 356468 381578
rect 356164 381516 356170 381518
rect 356462 381516 356468 381518
rect 356532 381516 356538 381580
rect 187049 381170 187115 381173
rect 200062 381170 200068 381172
rect 187049 381168 200068 381170
rect 187049 381112 187054 381168
rect 187110 381112 200068 381168
rect 187049 381110 200068 381112
rect 187049 381107 187115 381110
rect 200062 381108 200068 381110
rect 200132 381108 200138 381172
rect 4797 381034 4863 381037
rect 104985 381034 105051 381037
rect 105537 381034 105603 381037
rect 4797 381032 105603 381034
rect 4797 380976 4802 381032
rect 4858 380976 104990 381032
rect 105046 380976 105542 381032
rect 105598 380976 105603 381032
rect 4797 380974 105603 380976
rect 4797 380971 4863 380974
rect 104985 380971 105051 380974
rect 105537 380971 105603 380974
rect 111057 381034 111123 381037
rect 111558 381034 111564 381036
rect 111057 381032 111564 381034
rect 111057 380976 111062 381032
rect 111118 380976 111564 381032
rect 111057 380974 111564 380976
rect 111057 380971 111123 380974
rect 111558 380972 111564 380974
rect 111628 381034 111634 381036
rect 188613 381034 188679 381037
rect 111628 381032 188679 381034
rect 111628 380976 188618 381032
rect 188674 380976 188679 381032
rect 111628 380974 188679 380976
rect 111628 380972 111634 380974
rect 188613 380971 188679 380974
rect 69657 380218 69723 380221
rect 195237 380218 195303 380221
rect 69657 380216 195303 380218
rect 69657 380160 69662 380216
rect 69718 380160 195242 380216
rect 195298 380160 195303 380216
rect 69657 380158 195303 380160
rect 69657 380155 69723 380158
rect 195237 380155 195303 380158
rect 197353 380082 197419 380085
rect 197353 380080 200100 380082
rect 197353 380024 197358 380080
rect 197414 380024 200100 380080
rect 197353 380022 200100 380024
rect 197353 380019 197419 380022
rect 357893 379810 357959 379813
rect 356132 379808 357959 379810
rect 356132 379752 357898 379808
rect 357954 379752 357959 379808
rect 356132 379750 357959 379752
rect 357893 379747 357959 379750
rect 73797 379538 73863 379541
rect 194593 379538 194659 379541
rect 73797 379536 194659 379538
rect 73797 379480 73802 379536
rect 73858 379480 194598 379536
rect 194654 379480 194659 379536
rect 73797 379478 194659 379480
rect 73797 379475 73863 379478
rect 194593 379475 194659 379478
rect 115657 379266 115723 379269
rect 115790 379266 115796 379268
rect 115657 379264 115796 379266
rect 115657 379208 115662 379264
rect 115718 379208 115796 379264
rect 115657 379206 115796 379208
rect 115657 379203 115723 379206
rect 115790 379204 115796 379206
rect 115860 379204 115866 379268
rect 63309 378722 63375 378725
rect 111742 378722 111748 378724
rect 63309 378720 111748 378722
rect 63309 378664 63314 378720
rect 63370 378664 111748 378720
rect 63309 378662 111748 378664
rect 63309 378659 63375 378662
rect 111742 378660 111748 378662
rect 111812 378660 111818 378724
rect 191189 378450 191255 378453
rect 199837 378450 199903 378453
rect 191189 378448 199903 378450
rect 191189 378392 191194 378448
rect 191250 378392 199842 378448
rect 199898 378392 199903 378448
rect 191189 378390 199903 378392
rect 191189 378387 191255 378390
rect 199837 378387 199903 378390
rect 582373 378450 582439 378453
rect 583520 378450 584960 378540
rect 582373 378448 584960 378450
rect 582373 378392 582378 378448
rect 582434 378392 584960 378448
rect 582373 378390 584960 378392
rect 582373 378387 582439 378390
rect 115657 378314 115723 378317
rect 115657 378312 122850 378314
rect 115657 378256 115662 378312
rect 115718 378256 122850 378312
rect 583520 378300 584960 378390
rect 115657 378254 122850 378256
rect 115657 378251 115723 378254
rect 114318 378116 114324 378180
rect 114388 378178 114394 378180
rect 119981 378178 120047 378181
rect 114388 378176 120047 378178
rect 114388 378120 119986 378176
rect 120042 378120 120047 378176
rect 114388 378118 120047 378120
rect 122790 378178 122850 378254
rect 196566 378178 196572 378180
rect 122790 378118 196572 378178
rect 114388 378116 114394 378118
rect 119981 378115 120047 378118
rect 196566 378116 196572 378118
rect 196636 378116 196642 378180
rect 357566 377980 357572 378044
rect 357636 378042 357642 378044
rect 358353 378042 358419 378045
rect 357636 378040 358419 378042
rect 357636 377984 358358 378040
rect 358414 377984 358419 378040
rect 357636 377982 358419 377984
rect 357636 377980 357642 377982
rect 358353 377979 358419 377982
rect 198774 377572 198780 377636
rect 198844 377634 198850 377636
rect 204437 377634 204503 377637
rect 198844 377632 204503 377634
rect 198844 377576 204442 377632
rect 204498 377576 204503 377632
rect 198844 377574 204503 377576
rect 198844 377572 198850 377574
rect 204437 377571 204503 377574
rect 67766 377436 67772 377500
rect 67836 377498 67842 377500
rect 116485 377498 116551 377501
rect 262489 377498 262555 377501
rect 67836 377496 262555 377498
rect 67836 377440 116490 377496
rect 116546 377440 262494 377496
rect 262550 377440 262555 377496
rect 67836 377438 262555 377440
rect 67836 377436 67842 377438
rect 116485 377435 116551 377438
rect 262489 377435 262555 377438
rect 354121 377498 354187 377501
rect 358997 377498 359063 377501
rect 354121 377496 359063 377498
rect 354121 377440 354126 377496
rect 354182 377440 359002 377496
rect 359058 377440 359063 377496
rect 354121 377438 359063 377440
rect 354121 377435 354187 377438
rect 358997 377435 359063 377438
rect 68318 377300 68324 377364
rect 68388 377362 68394 377364
rect 142889 377362 142955 377365
rect 68388 377360 142955 377362
rect 68388 377304 142894 377360
rect 142950 377304 142955 377360
rect 68388 377302 142955 377304
rect 68388 377300 68394 377302
rect 142889 377299 142955 377302
rect 185761 377362 185827 377365
rect 202045 377362 202111 377365
rect 185761 377360 202111 377362
rect 185761 377304 185766 377360
rect 185822 377304 202050 377360
rect 202106 377304 202111 377360
rect 185761 377302 202111 377304
rect 185761 377299 185827 377302
rect 202045 377299 202111 377302
rect 202229 377362 202295 377365
rect 367369 377362 367435 377365
rect 202229 377360 367435 377362
rect 202229 377304 202234 377360
rect 202290 377304 367374 377360
rect 367430 377304 367435 377360
rect 202229 377302 367435 377304
rect 202229 377299 202295 377302
rect 367369 377299 367435 377302
rect 199837 377226 199903 377229
rect 201401 377226 201467 377229
rect 199837 377224 201467 377226
rect 199837 377168 199842 377224
rect 199898 377168 201406 377224
rect 201462 377168 201467 377224
rect 199837 377166 201467 377168
rect 199837 377163 199903 377166
rect 201401 377163 201467 377166
rect 318793 376954 318859 376957
rect 319621 376954 319687 376957
rect 582649 376954 582715 376957
rect 318793 376952 582715 376954
rect 318793 376896 318798 376952
rect 318854 376896 319626 376952
rect 319682 376896 582654 376952
rect 582710 376896 582715 376952
rect 318793 376894 582715 376896
rect 318793 376891 318859 376894
rect 319621 376891 319687 376894
rect 582649 376891 582715 376894
rect 64689 376682 64755 376685
rect 258717 376682 258783 376685
rect 64689 376680 258783 376682
rect 64689 376624 64694 376680
rect 64750 376624 258722 376680
rect 258778 376624 258783 376680
rect 64689 376622 258783 376624
rect 64689 376619 64755 376622
rect 258717 376619 258783 376622
rect 281349 376682 281415 376685
rect 583201 376682 583267 376685
rect 281349 376680 583267 376682
rect 281349 376624 281354 376680
rect 281410 376624 583206 376680
rect 583262 376624 583267 376680
rect 281349 376622 583267 376624
rect 281349 376619 281415 376622
rect 583201 376619 583267 376622
rect 114553 376546 114619 376549
rect 115749 376546 115815 376549
rect 114553 376544 115815 376546
rect 114553 376488 114558 376544
rect 114614 376488 115754 376544
rect 115810 376488 115815 376544
rect 114553 376486 115815 376488
rect 114553 376483 114619 376486
rect 115749 376483 115815 376486
rect 195697 376546 195763 376549
rect 195830 376546 195836 376548
rect 195697 376544 195836 376546
rect 195697 376488 195702 376544
rect 195758 376488 195836 376544
rect 195697 376486 195836 376488
rect 195697 376483 195763 376486
rect 195830 376484 195836 376486
rect 195900 376484 195906 376548
rect 247033 376546 247099 376549
rect 248045 376546 248111 376549
rect 374637 376546 374703 376549
rect 247033 376544 374703 376546
rect 247033 376488 247038 376544
rect 247094 376488 248050 376544
rect 248106 376488 374642 376544
rect 374698 376488 374703 376544
rect 247033 376486 374703 376488
rect 247033 376483 247099 376486
rect 248045 376483 248111 376486
rect 374637 376483 374703 376486
rect 354673 376410 354739 376413
rect 354806 376410 354812 376412
rect 354673 376408 354812 376410
rect 354673 376352 354678 376408
rect 354734 376352 354812 376408
rect 354673 376350 354812 376352
rect 354673 376347 354739 376350
rect 354806 376348 354812 376350
rect 354876 376348 354882 376412
rect 195881 376002 195947 376005
rect 207105 376002 207171 376005
rect 195881 376000 207171 376002
rect 195881 375944 195886 376000
rect 195942 375944 207110 376000
rect 207166 375944 207171 376000
rect 195881 375942 207171 375944
rect 195881 375939 195947 375942
rect 207105 375939 207171 375942
rect 340229 376002 340295 376005
rect 353334 376002 353340 376004
rect 340229 376000 353340 376002
rect 340229 375944 340234 376000
rect 340290 375944 353340 376000
rect 340229 375942 353340 375944
rect 340229 375939 340295 375942
rect 353334 375940 353340 375942
rect 353404 375940 353410 376004
rect 115749 375458 115815 375461
rect 204897 375458 204963 375461
rect 115749 375456 204963 375458
rect 115749 375400 115754 375456
rect 115810 375400 204902 375456
rect 204958 375400 204963 375456
rect 115749 375398 204963 375400
rect 115749 375395 115815 375398
rect 204897 375395 204963 375398
rect 200297 375322 200363 375325
rect 206645 375322 206711 375325
rect 200297 375320 206711 375322
rect 200297 375264 200302 375320
rect 200358 375264 206650 375320
rect 206706 375264 206711 375320
rect 200297 375262 206711 375264
rect 200297 375259 200363 375262
rect 206645 375259 206711 375262
rect 239765 375322 239831 375325
rect 241646 375322 241652 375324
rect 239765 375320 241652 375322
rect 239765 375264 239770 375320
rect 239826 375264 241652 375320
rect 239765 375262 241652 375264
rect 239765 375259 239831 375262
rect 241646 375260 241652 375262
rect 241716 375260 241722 375324
rect 251357 375322 251423 375325
rect 256693 375322 256759 375325
rect 251357 375320 256759 375322
rect 251357 375264 251362 375320
rect 251418 375264 256698 375320
rect 256754 375264 256759 375320
rect 251357 375262 256759 375264
rect 251357 375259 251423 375262
rect 256693 375259 256759 375262
rect 288382 375260 288388 375324
rect 288452 375322 288458 375324
rect 289629 375322 289695 375325
rect 288452 375320 289695 375322
rect 288452 375264 289634 375320
rect 289690 375264 289695 375320
rect 288452 375262 289695 375264
rect 288452 375260 288458 375262
rect 289629 375259 289695 375262
rect 307017 375322 307083 375325
rect 312813 375322 312879 375325
rect 307017 375320 312879 375322
rect 307017 375264 307022 375320
rect 307078 375264 312818 375320
rect 312874 375264 312879 375320
rect 307017 375262 312879 375264
rect 307017 375259 307083 375262
rect 312813 375259 312879 375262
rect 346117 375322 346183 375325
rect 349153 375322 349219 375325
rect 346117 375320 349219 375322
rect 346117 375264 346122 375320
rect 346178 375264 349158 375320
rect 349214 375264 349219 375320
rect 346117 375262 349219 375264
rect 346117 375259 346183 375262
rect 349153 375259 349219 375262
rect 352557 375322 352623 375325
rect 354438 375322 354444 375324
rect 352557 375320 354444 375322
rect 352557 375264 352562 375320
rect 352618 375264 354444 375320
rect 352557 375262 354444 375264
rect 352557 375259 352623 375262
rect 354438 375260 354444 375262
rect 354508 375260 354514 375324
rect 196617 374778 196683 374781
rect 200297 374778 200363 374781
rect 196617 374776 200363 374778
rect 196617 374720 196622 374776
rect 196678 374720 200302 374776
rect 200358 374720 200363 374776
rect 196617 374718 200363 374720
rect 196617 374715 196683 374718
rect 200297 374715 200363 374718
rect 351085 374778 351151 374781
rect 358813 374778 358879 374781
rect 351085 374776 358879 374778
rect 351085 374720 351090 374776
rect 351146 374720 358818 374776
rect 358874 374720 358879 374776
rect 351085 374718 358879 374720
rect 351085 374715 351151 374718
rect 358813 374715 358879 374718
rect 97257 374642 97323 374645
rect 126237 374642 126303 374645
rect 97257 374640 126303 374642
rect 97257 374584 97262 374640
rect 97318 374584 126242 374640
rect 126298 374584 126303 374640
rect 97257 374582 126303 374584
rect 97257 374579 97323 374582
rect 126237 374579 126303 374582
rect 187601 374642 187667 374645
rect 244774 374642 244780 374644
rect 187601 374640 244780 374642
rect 187601 374584 187606 374640
rect 187662 374584 244780 374640
rect 187601 374582 244780 374584
rect 187601 374579 187667 374582
rect 244774 374580 244780 374582
rect 244844 374580 244850 374644
rect 280889 374642 280955 374645
rect 304533 374642 304599 374645
rect 280889 374640 304599 374642
rect 280889 374584 280894 374640
rect 280950 374584 304538 374640
rect 304594 374584 304599 374640
rect 280889 374582 304599 374584
rect 280889 374579 280955 374582
rect 304533 374579 304599 374582
rect 342345 374642 342411 374645
rect 382917 374642 382983 374645
rect 342345 374640 382983 374642
rect 342345 374584 342350 374640
rect 342406 374584 382922 374640
rect 382978 374584 382983 374640
rect 342345 374582 382983 374584
rect 342345 374579 342411 374582
rect 382917 374579 382983 374582
rect 59169 374098 59235 374101
rect 214557 374098 214623 374101
rect 59169 374096 214623 374098
rect 59169 374040 59174 374096
rect 59230 374040 214562 374096
rect 214618 374040 214623 374096
rect 59169 374038 214623 374040
rect 59169 374035 59235 374038
rect 214557 374035 214623 374038
rect 283557 374098 283623 374101
rect 303654 374098 303660 374100
rect 283557 374096 303660 374098
rect 283557 374040 283562 374096
rect 283618 374040 303660 374096
rect 283557 374038 303660 374040
rect 283557 374035 283623 374038
rect 303654 374036 303660 374038
rect 303724 374036 303730 374100
rect 195237 373962 195303 373965
rect 361849 373962 361915 373965
rect 195237 373960 361915 373962
rect 195237 373904 195242 373960
rect 195298 373904 361854 373960
rect 361910 373904 361915 373960
rect 195237 373902 361915 373904
rect 195237 373899 195303 373902
rect 361849 373899 361915 373902
rect 81341 373418 81407 373421
rect 96286 373418 96292 373420
rect 81341 373416 96292 373418
rect 81341 373360 81346 373416
rect 81402 373360 96292 373416
rect 81341 373358 96292 373360
rect 81341 373355 81407 373358
rect 96286 373356 96292 373358
rect 96356 373356 96362 373420
rect 191741 373418 191807 373421
rect 200113 373418 200179 373421
rect 191741 373416 200179 373418
rect 191741 373360 191746 373416
rect 191802 373360 200118 373416
rect 200174 373360 200179 373416
rect 191741 373358 200179 373360
rect 191741 373355 191807 373358
rect 200113 373355 200179 373358
rect 54937 373282 55003 373285
rect 176009 373282 176075 373285
rect 54937 373280 176075 373282
rect 54937 373224 54942 373280
rect 54998 373224 176014 373280
rect 176070 373224 176075 373280
rect 54937 373222 176075 373224
rect 54937 373219 55003 373222
rect 176009 373219 176075 373222
rect 180701 373282 180767 373285
rect 354673 373282 354739 373285
rect 180701 373280 354739 373282
rect 180701 373224 180706 373280
rect 180762 373224 354678 373280
rect 354734 373224 354739 373280
rect 180701 373222 354739 373224
rect 180701 373219 180767 373222
rect 354673 373219 354739 373222
rect 99281 371922 99347 371925
rect 243537 371922 243603 371925
rect 99281 371920 243603 371922
rect 99281 371864 99286 371920
rect 99342 371864 243542 371920
rect 243598 371864 243603 371920
rect 99281 371862 243603 371864
rect 99281 371859 99347 371862
rect 243537 371859 243603 371862
rect -960 371378 480 371468
rect 3509 371378 3575 371381
rect -960 371376 3575 371378
rect -960 371320 3514 371376
rect 3570 371320 3575 371376
rect -960 371318 3575 371320
rect -960 371228 480 371318
rect 3509 371315 3575 371318
rect 89621 371378 89687 371381
rect 356094 371378 356100 371380
rect 89621 371376 356100 371378
rect 89621 371320 89626 371376
rect 89682 371320 356100 371376
rect 89621 371318 356100 371320
rect 89621 371315 89687 371318
rect 356094 371316 356100 371318
rect 356164 371316 356170 371380
rect 69790 370500 69796 370564
rect 69860 370562 69866 370564
rect 87597 370562 87663 370565
rect 69860 370560 87663 370562
rect 69860 370504 87602 370560
rect 87658 370504 87663 370560
rect 69860 370502 87663 370504
rect 69860 370500 69866 370502
rect 87597 370499 87663 370502
rect 100017 370018 100083 370021
rect 100518 370018 100524 370020
rect 100017 370016 100524 370018
rect 100017 369960 100022 370016
rect 100078 369960 100524 370016
rect 100017 369958 100524 369960
rect 100017 369955 100083 369958
rect 100518 369956 100524 369958
rect 100588 370018 100594 370020
rect 222929 370018 222995 370021
rect 100588 370016 222995 370018
rect 100588 369960 222934 370016
rect 222990 369960 222995 370016
rect 100588 369958 222995 369960
rect 100588 369956 100594 369958
rect 222929 369955 222995 369958
rect 93117 369882 93183 369885
rect 287053 369882 287119 369885
rect 287697 369882 287763 369885
rect 93117 369880 287763 369882
rect 93117 369824 93122 369880
rect 93178 369824 287058 369880
rect 287114 369824 287702 369880
rect 287758 369824 287763 369880
rect 93117 369822 287763 369824
rect 93117 369819 93183 369822
rect 287053 369819 287119 369822
rect 287697 369819 287763 369822
rect 184381 369066 184447 369069
rect 217409 369066 217475 369069
rect 184381 369064 217475 369066
rect 184381 369008 184386 369064
rect 184442 369008 217414 369064
rect 217470 369008 217475 369064
rect 184381 369006 217475 369008
rect 184381 369003 184447 369006
rect 217409 369003 217475 369006
rect 311893 369066 311959 369069
rect 370129 369066 370195 369069
rect 311893 369064 370195 369066
rect 311893 369008 311898 369064
rect 311954 369008 370134 369064
rect 370190 369008 370195 369064
rect 311893 369006 370195 369008
rect 311893 369003 311959 369006
rect 370129 369003 370195 369006
rect 125501 368658 125567 368661
rect 156781 368658 156847 368661
rect 125501 368656 156847 368658
rect 125501 368600 125506 368656
rect 125562 368600 156786 368656
rect 156842 368600 156847 368656
rect 125501 368598 156847 368600
rect 125501 368595 125567 368598
rect 156781 368595 156847 368598
rect 195278 368596 195284 368660
rect 195348 368658 195354 368660
rect 325693 368658 325759 368661
rect 326337 368658 326403 368661
rect 195348 368656 326403 368658
rect 195348 368600 325698 368656
rect 325754 368600 326342 368656
rect 326398 368600 326403 368656
rect 195348 368598 326403 368600
rect 195348 368596 195354 368598
rect 325693 368595 325759 368598
rect 326337 368595 326403 368598
rect 69606 368460 69612 368524
rect 69676 368522 69682 368524
rect 311893 368522 311959 368525
rect 69676 368520 311959 368522
rect 69676 368464 311898 368520
rect 311954 368464 311959 368520
rect 69676 368462 311959 368464
rect 69676 368460 69682 368462
rect 311893 368459 311959 368462
rect 55029 368386 55095 368389
rect 125501 368386 125567 368389
rect 55029 368384 125567 368386
rect 55029 368328 55034 368384
rect 55090 368328 125506 368384
rect 125562 368328 125567 368384
rect 55029 368326 125567 368328
rect 55029 368323 55095 368326
rect 125501 368323 125567 368326
rect 169109 368386 169175 368389
rect 169845 368386 169911 368389
rect 247033 368386 247099 368389
rect 169109 368384 247099 368386
rect 169109 368328 169114 368384
rect 169170 368328 169850 368384
rect 169906 368328 247038 368384
rect 247094 368328 247099 368384
rect 169109 368326 247099 368328
rect 169109 368323 169175 368326
rect 169845 368323 169911 368326
rect 247033 368323 247099 368326
rect 125593 368250 125659 368253
rect 126881 368250 126947 368253
rect 125593 368248 126947 368250
rect 125593 368192 125598 368248
rect 125654 368192 126886 368248
rect 126942 368192 126947 368248
rect 125593 368190 126947 368192
rect 125593 368187 125659 368190
rect 126881 368187 126947 368190
rect 195237 367842 195303 367845
rect 224902 367842 224908 367844
rect 195237 367840 224908 367842
rect 195237 367784 195242 367840
rect 195298 367784 224908 367840
rect 195237 367782 224908 367784
rect 195237 367779 195303 367782
rect 224902 367780 224908 367782
rect 224972 367780 224978 367844
rect 116577 367706 116643 367709
rect 152457 367706 152523 367709
rect 116577 367704 152523 367706
rect 116577 367648 116582 367704
rect 116638 367648 152462 367704
rect 152518 367648 152523 367704
rect 116577 367646 152523 367648
rect 116577 367643 116643 367646
rect 152457 367643 152523 367646
rect 157926 367644 157932 367708
rect 157996 367706 158002 367708
rect 354121 367706 354187 367709
rect 157996 367704 354187 367706
rect 157996 367648 354126 367704
rect 354182 367648 354187 367704
rect 157996 367646 354187 367648
rect 157996 367644 158002 367646
rect 354121 367643 354187 367646
rect 126881 367162 126947 367165
rect 156689 367162 156755 367165
rect 126881 367160 156755 367162
rect 126881 367104 126886 367160
rect 126942 367104 156694 367160
rect 156750 367104 156755 367160
rect 126881 367102 156755 367104
rect 126881 367099 126947 367102
rect 156689 367099 156755 367102
rect 126973 367026 127039 367029
rect 127617 367026 127683 367029
rect 126973 367024 127683 367026
rect 126973 366968 126978 367024
rect 127034 366968 127622 367024
rect 127678 366968 127683 367024
rect 126973 366966 127683 366968
rect 126973 366963 127039 366966
rect 127617 366963 127683 366966
rect 198825 366482 198891 366485
rect 218145 366482 218211 366485
rect 198825 366480 218211 366482
rect 198825 366424 198830 366480
rect 198886 366424 218150 366480
rect 218206 366424 218211 366480
rect 198825 366422 218211 366424
rect 198825 366419 198891 366422
rect 218145 366419 218211 366422
rect 126973 366346 127039 366349
rect 259453 366346 259519 366349
rect 259729 366346 259795 366349
rect 126973 366344 259795 366346
rect 126973 366288 126978 366344
rect 127034 366288 259458 366344
rect 259514 366288 259734 366344
rect 259790 366288 259795 366344
rect 126973 366286 259795 366288
rect 126973 366283 127039 366286
rect 259453 366283 259519 366286
rect 259729 366283 259795 366286
rect 73061 365802 73127 365805
rect 180149 365802 180215 365805
rect 73061 365800 180215 365802
rect 73061 365744 73066 365800
rect 73122 365744 180154 365800
rect 180210 365744 180215 365800
rect 73061 365742 180215 365744
rect 73061 365739 73127 365742
rect 180149 365739 180215 365742
rect 192661 365802 192727 365805
rect 222101 365802 222167 365805
rect 285622 365802 285628 365804
rect 192661 365800 200130 365802
rect 192661 365744 192666 365800
rect 192722 365744 200130 365800
rect 192661 365742 200130 365744
rect 192661 365739 192727 365742
rect 200070 365666 200130 365742
rect 222101 365800 285628 365802
rect 222101 365744 222106 365800
rect 222162 365744 285628 365800
rect 222101 365742 285628 365744
rect 222101 365739 222167 365742
rect 285622 365740 285628 365742
rect 285692 365740 285698 365804
rect 370037 365666 370103 365669
rect 200070 365664 370103 365666
rect 200070 365608 370042 365664
rect 370098 365608 370103 365664
rect 200070 365606 370103 365608
rect 370037 365603 370103 365606
rect 185393 365530 185459 365533
rect 220813 365530 220879 365533
rect 222101 365530 222167 365533
rect 185393 365528 222167 365530
rect 185393 365472 185398 365528
rect 185454 365472 220818 365528
rect 220874 365472 222106 365528
rect 222162 365472 222167 365528
rect 185393 365470 222167 365472
rect 185393 365467 185459 365470
rect 220813 365467 220879 365470
rect 222101 365467 222167 365470
rect 582373 365122 582439 365125
rect 583520 365122 584960 365212
rect 582373 365120 584960 365122
rect 582373 365064 582378 365120
rect 582434 365064 584960 365120
rect 582373 365062 584960 365064
rect 582373 365059 582439 365062
rect 166349 364986 166415 364989
rect 308397 364986 308463 364989
rect 166349 364984 308463 364986
rect 166349 364928 166354 364984
rect 166410 364928 308402 364984
rect 308458 364928 308463 364984
rect 583520 364972 584960 365062
rect 166349 364926 308463 364928
rect 166349 364923 166415 364926
rect 308397 364923 308463 364926
rect 64638 364652 64644 364716
rect 64708 364714 64714 364716
rect 137277 364714 137343 364717
rect 64708 364712 137343 364714
rect 64708 364656 137282 364712
rect 137338 364656 137343 364712
rect 64708 364654 137343 364656
rect 64708 364652 64714 364654
rect 137277 364651 137343 364654
rect 116669 364578 116735 364581
rect 193857 364578 193923 364581
rect 116669 364576 193923 364578
rect 116669 364520 116674 364576
rect 116730 364520 193862 364576
rect 193918 364520 193923 364576
rect 116669 364518 193923 364520
rect 116669 364515 116735 364518
rect 193857 364515 193923 364518
rect 93853 364442 93919 364445
rect 95141 364442 95207 364445
rect 186129 364442 186195 364445
rect 93853 364440 186195 364442
rect 93853 364384 93858 364440
rect 93914 364384 95146 364440
rect 95202 364384 186134 364440
rect 186190 364384 186195 364440
rect 93853 364382 186195 364384
rect 93853 364379 93919 364382
rect 95141 364379 95207 364382
rect 186129 364379 186195 364382
rect 147581 363218 147647 363221
rect 229737 363218 229803 363221
rect 147581 363216 229803 363218
rect 147581 363160 147586 363216
rect 147642 363160 229742 363216
rect 229798 363160 229803 363216
rect 147581 363158 229803 363160
rect 147581 363155 147647 363158
rect 229737 363155 229803 363158
rect 61929 363082 61995 363085
rect 328453 363082 328519 363085
rect 329097 363082 329163 363085
rect 61929 363080 329163 363082
rect 61929 363024 61934 363080
rect 61990 363024 328458 363080
rect 328514 363024 329102 363080
rect 329158 363024 329163 363080
rect 61929 363022 329163 363024
rect 61929 363019 61995 363022
rect 328453 363019 328519 363022
rect 329097 363019 329163 363022
rect 196566 362340 196572 362404
rect 196636 362402 196642 362404
rect 218697 362402 218763 362405
rect 196636 362400 218763 362402
rect 196636 362344 218702 362400
rect 218758 362344 218763 362400
rect 196636 362342 218763 362344
rect 196636 362340 196642 362342
rect 218697 362339 218763 362342
rect 146201 362266 146267 362269
rect 206461 362266 206527 362269
rect 146201 362264 206527 362266
rect 146201 362208 146206 362264
rect 146262 362208 206466 362264
rect 206522 362208 206527 362264
rect 146201 362206 206527 362208
rect 146201 362203 146267 362206
rect 206461 362203 206527 362206
rect 338757 362266 338823 362269
rect 357566 362266 357572 362268
rect 338757 362264 357572 362266
rect 338757 362208 338762 362264
rect 338818 362208 357572 362264
rect 338757 362206 357572 362208
rect 338757 362203 338823 362206
rect 357566 362204 357572 362206
rect 357636 362204 357642 362268
rect 71078 361796 71084 361860
rect 71148 361858 71154 361860
rect 185577 361858 185643 361861
rect 71148 361856 185643 361858
rect 71148 361800 185582 361856
rect 185638 361800 185643 361856
rect 71148 361798 185643 361800
rect 71148 361796 71154 361798
rect 185577 361795 185643 361798
rect 133781 361722 133847 361725
rect 320173 361722 320239 361725
rect 133781 361720 320239 361722
rect 133781 361664 133786 361720
rect 133842 361664 320178 361720
rect 320234 361664 320239 361720
rect 133781 361662 320239 361664
rect 133781 361659 133847 361662
rect 320173 361659 320239 361662
rect 173893 361586 173959 361589
rect 353293 361586 353359 361589
rect 173893 361584 353359 361586
rect 173893 361528 173898 361584
rect 173954 361528 353298 361584
rect 353354 361528 353359 361584
rect 173893 361526 353359 361528
rect 173893 361523 173959 361526
rect 353293 361523 353359 361526
rect 180701 361450 180767 361453
rect 180701 361448 180810 361450
rect 180701 361392 180706 361448
rect 180762 361392 180810 361448
rect 180701 361387 180810 361392
rect 115841 361042 115907 361045
rect 180750 361042 180810 361387
rect 181437 361042 181503 361045
rect 115841 361040 181503 361042
rect 115841 360984 115846 361040
rect 115902 360984 181442 361040
rect 181498 360984 181503 361040
rect 115841 360982 181503 360984
rect 115841 360979 115907 360982
rect 181437 360979 181503 360982
rect 66069 360906 66135 360909
rect 283557 360906 283623 360909
rect 66069 360904 283623 360906
rect 66069 360848 66074 360904
rect 66130 360848 283562 360904
rect 283618 360848 283623 360904
rect 66069 360846 283623 360848
rect 66069 360843 66135 360846
rect 283557 360843 283623 360846
rect 97809 360090 97875 360093
rect 157742 360090 157748 360092
rect 97809 360088 157748 360090
rect 97809 360032 97814 360088
rect 97870 360032 157748 360088
rect 97809 360030 157748 360032
rect 97809 360027 97875 360030
rect 157742 360028 157748 360030
rect 157812 360028 157818 360092
rect 240869 359410 240935 359413
rect 356278 359410 356284 359412
rect 240869 359408 356284 359410
rect 240869 359352 240874 359408
rect 240930 359352 356284 359408
rect 240869 359350 356284 359352
rect 240869 359347 240935 359350
rect 356278 359348 356284 359350
rect 356348 359348 356354 359412
rect 178769 359002 178835 359005
rect 252553 359002 252619 359005
rect 253289 359002 253355 359005
rect 178769 359000 253355 359002
rect 178769 358944 178774 359000
rect 178830 358944 252558 359000
rect 252614 358944 253294 359000
rect 253350 358944 253355 359000
rect 178769 358942 253355 358944
rect 178769 358939 178835 358942
rect 252553 358939 252619 358942
rect 253289 358939 253355 358942
rect 136633 358866 136699 358869
rect 137921 358866 137987 358869
rect 211981 358866 212047 358869
rect 136633 358864 212047 358866
rect 136633 358808 136638 358864
rect 136694 358808 137926 358864
rect 137982 358808 211986 358864
rect 212042 358808 212047 358864
rect 136633 358806 212047 358808
rect 136633 358803 136699 358806
rect 137921 358803 137987 358806
rect 211981 358803 212047 358806
rect 152549 358730 152615 358733
rect 153101 358730 153167 358733
rect 152549 358728 153167 358730
rect 152549 358672 152554 358728
rect 152610 358672 153106 358728
rect 153162 358672 153167 358728
rect 152549 358670 153167 358672
rect 152549 358667 152615 358670
rect 153101 358667 153167 358670
rect -960 358458 480 358548
rect 3325 358458 3391 358461
rect -960 358456 3391 358458
rect -960 358400 3330 358456
rect 3386 358400 3391 358456
rect -960 358398 3391 358400
rect -960 358308 480 358398
rect 3325 358395 3391 358398
rect 121453 358050 121519 358053
rect 159357 358050 159423 358053
rect 223573 358050 223639 358053
rect 121453 358048 159423 358050
rect 121453 357992 121458 358048
rect 121514 357992 159362 358048
rect 159418 357992 159423 358048
rect 121453 357990 159423 357992
rect 121453 357987 121519 357990
rect 159357 357987 159423 357990
rect 190410 358048 223639 358050
rect 190410 357992 223578 358048
rect 223634 357992 223639 358048
rect 190410 357990 223639 357992
rect 153101 357778 153167 357781
rect 188521 357778 188587 357781
rect 190410 357778 190470 357990
rect 223573 357987 223639 357990
rect 153101 357776 190470 357778
rect 153101 357720 153106 357776
rect 153162 357720 188526 357776
rect 188582 357720 190470 357776
rect 153101 357718 190470 357720
rect 153101 357715 153167 357718
rect 188521 357715 188587 357718
rect 169293 357642 169359 357645
rect 169661 357642 169727 357645
rect 238017 357642 238083 357645
rect 169293 357640 238083 357642
rect 169293 357584 169298 357640
rect 169354 357584 169666 357640
rect 169722 357584 238022 357640
rect 238078 357584 238083 357640
rect 169293 357582 238083 357584
rect 169293 357579 169359 357582
rect 169661 357579 169727 357582
rect 238017 357579 238083 357582
rect 110229 357506 110295 357509
rect 223021 357506 223087 357509
rect 110229 357504 223087 357506
rect 110229 357448 110234 357504
rect 110290 357448 223026 357504
rect 223082 357448 223087 357504
rect 110229 357446 223087 357448
rect 110229 357443 110295 357446
rect 223021 357443 223087 357446
rect 98821 356962 98887 356965
rect 99189 356962 99255 356965
rect 196709 356962 196775 356965
rect 98821 356960 196775 356962
rect 98821 356904 98826 356960
rect 98882 356904 99194 356960
rect 99250 356904 196714 356960
rect 196770 356904 196775 356960
rect 98821 356902 196775 356904
rect 98821 356899 98887 356902
rect 99189 356899 99255 356902
rect 196709 356899 196775 356902
rect 174997 356826 175063 356829
rect 324313 356826 324379 356829
rect 174997 356824 324379 356826
rect 174997 356768 175002 356824
rect 175058 356768 324318 356824
rect 324374 356768 324379 356824
rect 174997 356766 324379 356768
rect 174997 356763 175063 356766
rect 324313 356763 324379 356766
rect 159950 356628 159956 356692
rect 160020 356690 160026 356692
rect 358854 356690 358860 356692
rect 160020 356630 358860 356690
rect 160020 356628 160026 356630
rect 358854 356628 358860 356630
rect 358924 356628 358930 356692
rect 96521 356146 96587 356149
rect 164693 356146 164759 356149
rect 96521 356144 164759 356146
rect 96521 356088 96526 356144
rect 96582 356088 164698 356144
rect 164754 356088 164759 356144
rect 96521 356086 164759 356088
rect 96521 356083 96587 356086
rect 164693 356083 164759 356086
rect 155217 356010 155283 356013
rect 160829 356010 160895 356013
rect 155217 356008 160895 356010
rect 155217 355952 155222 356008
rect 155278 355952 160834 356008
rect 160890 355952 160895 356008
rect 155217 355950 160895 355952
rect 155217 355947 155283 355950
rect 160829 355947 160895 355950
rect 295977 355466 296043 355469
rect 352046 355466 352052 355468
rect 295977 355464 352052 355466
rect 295977 355408 295982 355464
rect 296038 355408 352052 355464
rect 295977 355406 352052 355408
rect 295977 355403 296043 355406
rect 352046 355404 352052 355406
rect 352116 355404 352122 355468
rect 103329 355330 103395 355333
rect 147581 355330 147647 355333
rect 103329 355328 147647 355330
rect 103329 355272 103334 355328
rect 103390 355272 147586 355328
rect 147642 355272 147647 355328
rect 103329 355270 147647 355272
rect 103329 355267 103395 355270
rect 147581 355267 147647 355270
rect 149697 355330 149763 355333
rect 162209 355330 162275 355333
rect 149697 355328 162275 355330
rect 149697 355272 149702 355328
rect 149758 355272 162214 355328
rect 162270 355272 162275 355328
rect 149697 355270 162275 355272
rect 149697 355267 149763 355270
rect 162209 355267 162275 355270
rect 168189 355330 168255 355333
rect 313273 355330 313339 355333
rect 168189 355328 313339 355330
rect 168189 355272 168194 355328
rect 168250 355272 313278 355328
rect 313334 355272 313339 355328
rect 168189 355270 313339 355272
rect 168189 355267 168255 355270
rect 313273 355267 313339 355270
rect 133689 354786 133755 354789
rect 184197 354786 184263 354789
rect 133689 354784 184263 354786
rect 133689 354728 133694 354784
rect 133750 354728 184202 354784
rect 184258 354728 184263 354784
rect 133689 354726 184263 354728
rect 133689 354723 133755 354726
rect 184197 354723 184263 354726
rect 180558 354044 180564 354108
rect 180628 354106 180634 354108
rect 188429 354106 188495 354109
rect 180628 354104 188495 354106
rect 180628 354048 188434 354104
rect 188490 354048 188495 354104
rect 180628 354046 188495 354048
rect 180628 354044 180634 354046
rect 188429 354043 188495 354046
rect 121729 353970 121795 353973
rect 250437 353970 250503 353973
rect 121729 353968 250503 353970
rect 121729 353912 121734 353968
rect 121790 353912 250442 353968
rect 250498 353912 250503 353968
rect 121729 353910 250503 353912
rect 121729 353907 121795 353910
rect 250437 353907 250503 353910
rect 150341 353562 150407 353565
rect 180558 353562 180564 353564
rect 150341 353560 180564 353562
rect 150341 353504 150346 353560
rect 150402 353504 180564 353560
rect 150341 353502 180564 353504
rect 150341 353499 150407 353502
rect 180558 353500 180564 353502
rect 180628 353500 180634 353564
rect 199377 353562 199443 353565
rect 199510 353562 199516 353564
rect 199377 353560 199516 353562
rect 199377 353504 199382 353560
rect 199438 353504 199516 353560
rect 199377 353502 199516 353504
rect 199377 353499 199443 353502
rect 199510 353500 199516 353502
rect 199580 353500 199586 353564
rect 76741 353426 76807 353429
rect 113173 353426 113239 353429
rect 113817 353426 113883 353429
rect 76741 353424 113883 353426
rect 76741 353368 76746 353424
rect 76802 353368 113178 353424
rect 113234 353368 113822 353424
rect 113878 353368 113883 353424
rect 76741 353366 113883 353368
rect 76741 353363 76807 353366
rect 113173 353363 113239 353366
rect 113817 353363 113883 353366
rect 118601 353426 118667 353429
rect 155217 353426 155283 353429
rect 118601 353424 155283 353426
rect 118601 353368 118606 353424
rect 118662 353368 155222 353424
rect 155278 353368 155283 353424
rect 118601 353366 155283 353368
rect 118601 353363 118667 353366
rect 155217 353363 155283 353366
rect 191649 353426 191715 353429
rect 327073 353426 327139 353429
rect 191649 353424 327139 353426
rect 191649 353368 191654 353424
rect 191710 353368 327078 353424
rect 327134 353368 327139 353424
rect 191649 353366 327139 353368
rect 191649 353363 191715 353366
rect 327073 353363 327139 353366
rect 90357 353290 90423 353293
rect 129733 353290 129799 353293
rect 90357 353288 129799 353290
rect 90357 353232 90362 353288
rect 90418 353232 129738 353288
rect 129794 353232 129799 353288
rect 90357 353230 129799 353232
rect 90357 353227 90423 353230
rect 129733 353227 129799 353230
rect 234470 352610 234476 352612
rect 219390 352550 234476 352610
rect 129733 352066 129799 352069
rect 130469 352066 130535 352069
rect 129733 352064 130535 352066
rect 129733 352008 129738 352064
rect 129794 352008 130474 352064
rect 130530 352008 130535 352064
rect 129733 352006 130535 352008
rect 129733 352003 129799 352006
rect 130469 352003 130535 352006
rect 133873 352066 133939 352069
rect 219390 352066 219450 352550
rect 234470 352548 234476 352550
rect 234540 352610 234546 352612
rect 318793 352610 318859 352613
rect 234540 352608 318859 352610
rect 234540 352552 318798 352608
rect 318854 352552 318859 352608
rect 234540 352550 318859 352552
rect 234540 352548 234546 352550
rect 318793 352547 318859 352550
rect 133873 352064 219450 352066
rect 133873 352008 133878 352064
rect 133934 352008 219450 352064
rect 133873 352006 219450 352008
rect 133873 352003 133939 352006
rect 127065 351930 127131 351933
rect 127709 351930 127775 351933
rect 232497 351930 232563 351933
rect 127065 351928 232563 351930
rect 127065 351872 127070 351928
rect 127126 351872 127714 351928
rect 127770 351872 232502 351928
rect 232558 351872 232563 351928
rect 127065 351870 232563 351872
rect 127065 351867 127131 351870
rect 127709 351867 127775 351870
rect 232497 351867 232563 351870
rect 580165 351930 580231 351933
rect 583520 351930 584960 352020
rect 580165 351928 584960 351930
rect 580165 351872 580170 351928
rect 580226 351872 584960 351928
rect 580165 351870 584960 351872
rect 580165 351867 580231 351870
rect 583520 351780 584960 351870
rect 195697 351386 195763 351389
rect 211654 351386 211660 351388
rect 195697 351384 211660 351386
rect 195697 351328 195702 351384
rect 195758 351328 211660 351384
rect 195697 351326 211660 351328
rect 195697 351323 195763 351326
rect 211654 351324 211660 351326
rect 211724 351324 211730 351388
rect 107745 351250 107811 351253
rect 240726 351250 240732 351252
rect 107745 351248 240732 351250
rect 107745 351192 107750 351248
rect 107806 351192 240732 351248
rect 107745 351190 240732 351192
rect 107745 351187 107811 351190
rect 240726 351188 240732 351190
rect 240796 351250 240802 351252
rect 240869 351250 240935 351253
rect 240796 351248 240935 351250
rect 240796 351192 240874 351248
rect 240930 351192 240935 351248
rect 240796 351190 240935 351192
rect 240796 351188 240802 351190
rect 240869 351187 240935 351190
rect 91001 351114 91067 351117
rect 134701 351114 134767 351117
rect 191741 351114 191807 351117
rect 375557 351114 375623 351117
rect 91001 351112 134767 351114
rect 91001 351056 91006 351112
rect 91062 351056 134706 351112
rect 134762 351056 134767 351112
rect 91001 351054 134767 351056
rect 91001 351051 91067 351054
rect 134701 351051 134767 351054
rect 180750 351112 375623 351114
rect 180750 351056 191746 351112
rect 191802 351056 375562 351112
rect 375618 351056 375623 351112
rect 180750 351054 375623 351056
rect 124857 350570 124923 350573
rect 180750 350570 180810 351054
rect 191741 351051 191807 351054
rect 375557 351051 375623 351054
rect 124857 350568 180810 350570
rect 124857 350512 124862 350568
rect 124918 350512 180810 350568
rect 124857 350510 180810 350512
rect 124857 350507 124923 350510
rect 100661 349754 100727 349757
rect 169293 349754 169359 349757
rect 172605 349754 172671 349757
rect 347037 349754 347103 349757
rect 100661 349752 169359 349754
rect 100661 349696 100666 349752
rect 100722 349696 169298 349752
rect 169354 349696 169359 349752
rect 100661 349694 169359 349696
rect 100661 349691 100727 349694
rect 169293 349691 169359 349694
rect 171090 349752 347103 349754
rect 171090 349696 172610 349752
rect 172666 349696 347042 349752
rect 347098 349696 347103 349752
rect 171090 349694 347103 349696
rect 140773 349346 140839 349349
rect 141417 349346 141483 349349
rect 171090 349346 171150 349694
rect 172605 349691 172671 349694
rect 347037 349691 347103 349694
rect 140773 349344 171150 349346
rect 140773 349288 140778 349344
rect 140834 349288 141422 349344
rect 141478 349288 171150 349344
rect 140773 349286 171150 349288
rect 140773 349283 140839 349286
rect 141417 349283 141483 349286
rect 108481 349210 108547 349213
rect 108798 349210 108804 349212
rect 108481 349208 108804 349210
rect 108481 349152 108486 349208
rect 108542 349152 108804 349208
rect 108481 349150 108804 349152
rect 108481 349147 108547 349150
rect 108798 349148 108804 349150
rect 108868 349210 108874 349212
rect 183185 349210 183251 349213
rect 108868 349208 183251 349210
rect 108868 349152 183190 349208
rect 183246 349152 183251 349208
rect 108868 349150 183251 349152
rect 108868 349148 108874 349150
rect 183185 349147 183251 349150
rect 72734 349012 72740 349076
rect 72804 349074 72810 349076
rect 123201 349074 123267 349077
rect 124121 349074 124187 349077
rect 72804 349072 124187 349074
rect 72804 349016 123206 349072
rect 123262 349016 124126 349072
rect 124182 349016 124187 349072
rect 72804 349014 124187 349016
rect 72804 349012 72810 349014
rect 123201 349011 123267 349014
rect 124121 349011 124187 349014
rect 304257 349074 304323 349077
rect 305729 349074 305795 349077
rect 304257 349072 305795 349074
rect 304257 349016 304262 349072
rect 304318 349016 305734 349072
rect 305790 349016 305795 349072
rect 304257 349014 305795 349016
rect 304257 349011 304323 349014
rect 305729 349011 305795 349014
rect 68870 348468 68876 348532
rect 68940 348530 68946 348532
rect 122833 348530 122899 348533
rect 68940 348528 122899 348530
rect 68940 348472 122838 348528
rect 122894 348472 122899 348528
rect 68940 348470 122899 348472
rect 68940 348468 68946 348470
rect 122833 348467 122899 348470
rect 264973 348530 265039 348533
rect 360469 348530 360535 348533
rect 264973 348528 360535 348530
rect 264973 348472 264978 348528
rect 265034 348472 360474 348528
rect 360530 348472 360535 348528
rect 264973 348470 360535 348472
rect 264973 348467 265039 348470
rect 360469 348467 360535 348470
rect 111701 348394 111767 348397
rect 304257 348394 304323 348397
rect 111701 348392 304323 348394
rect 111701 348336 111706 348392
rect 111762 348336 304262 348392
rect 304318 348336 304323 348392
rect 111701 348334 304323 348336
rect 111701 348331 111767 348334
rect 304257 348331 304323 348334
rect 146937 347986 147003 347989
rect 178861 347986 178927 347989
rect 146937 347984 178927 347986
rect 146937 347928 146942 347984
rect 146998 347928 178866 347984
rect 178922 347928 178927 347984
rect 146937 347926 178927 347928
rect 146937 347923 147003 347926
rect 178861 347923 178927 347926
rect 124121 347850 124187 347853
rect 264973 347850 265039 347853
rect 124121 347848 265039 347850
rect 124121 347792 124126 347848
rect 124182 347792 264978 347848
rect 265034 347792 265039 347848
rect 124121 347790 265039 347792
rect 124121 347787 124187 347790
rect 264973 347787 265039 347790
rect 186957 347716 187023 347717
rect 186957 347712 187004 347716
rect 187068 347714 187074 347716
rect 186957 347656 186962 347712
rect 186957 347652 187004 347656
rect 187068 347654 187114 347714
rect 187068 347652 187074 347654
rect 186957 347651 187023 347652
rect 195237 347170 195303 347173
rect 248454 347170 248460 347172
rect 195237 347168 248460 347170
rect 195237 347112 195242 347168
rect 195298 347112 248460 347168
rect 195237 347110 248460 347112
rect 195237 347107 195303 347110
rect 248454 347108 248460 347110
rect 248524 347108 248530 347172
rect 66662 346972 66668 347036
rect 66732 347034 66738 347036
rect 361757 347034 361823 347037
rect 66732 347032 361823 347034
rect 66732 346976 361762 347032
rect 361818 346976 361823 347032
rect 66732 346974 361823 346976
rect 66732 346972 66738 346974
rect 361757 346971 361823 346974
rect 100569 346490 100635 346493
rect 186998 346490 187004 346492
rect 100569 346488 187004 346490
rect 100569 346432 100574 346488
rect 100630 346432 187004 346488
rect 100569 346430 187004 346432
rect 100569 346427 100635 346430
rect 186998 346428 187004 346430
rect 187068 346428 187074 346492
rect 104985 346354 105051 346357
rect 106181 346354 106247 346357
rect 104985 346352 106247 346354
rect 104985 346296 104990 346352
rect 105046 346296 106186 346352
rect 106242 346296 106247 346352
rect 104985 346294 106247 346296
rect 104985 346291 105051 346294
rect 106181 346291 106247 346294
rect 106181 345810 106247 345813
rect 215937 345810 216003 345813
rect 245694 345810 245700 345812
rect 106181 345808 245700 345810
rect 106181 345752 106186 345808
rect 106242 345752 215942 345808
rect 215998 345752 245700 345808
rect 106181 345750 245700 345752
rect 106181 345747 106247 345750
rect 215937 345747 216003 345750
rect 245694 345748 245700 345750
rect 245764 345748 245770 345812
rect 67357 345674 67423 345677
rect 121545 345674 121611 345677
rect 67357 345672 121611 345674
rect 67357 345616 67362 345672
rect 67418 345616 121550 345672
rect 121606 345616 121611 345672
rect 67357 345614 121611 345616
rect 67357 345611 67423 345614
rect 121545 345611 121611 345614
rect 144729 345674 144795 345677
rect 364609 345674 364675 345677
rect 144729 345672 364675 345674
rect 144729 345616 144734 345672
rect 144790 345616 364614 345672
rect 364670 345616 364675 345672
rect 144729 345614 364675 345616
rect 144729 345611 144795 345614
rect 364609 345611 364675 345614
rect -960 345402 480 345492
rect 2773 345402 2839 345405
rect -960 345400 2839 345402
rect -960 345344 2778 345400
rect 2834 345344 2839 345400
rect -960 345342 2839 345344
rect -960 345252 480 345342
rect 2773 345339 2839 345342
rect 128997 345130 129063 345133
rect 147029 345130 147095 345133
rect 128997 345128 147095 345130
rect 128997 345072 129002 345128
rect 129058 345072 147034 345128
rect 147090 345072 147095 345128
rect 128997 345070 147095 345072
rect 128997 345067 129063 345070
rect 147029 345067 147095 345070
rect 155718 345068 155724 345132
rect 155788 345130 155794 345132
rect 333973 345130 334039 345133
rect 155788 345128 334039 345130
rect 155788 345072 333978 345128
rect 334034 345072 334039 345128
rect 155788 345070 334039 345072
rect 155788 345068 155794 345070
rect 333973 345067 334039 345070
rect 69841 344314 69907 344317
rect 123477 344314 123543 344317
rect 360142 344314 360148 344316
rect 69841 344312 123543 344314
rect 69841 344256 69846 344312
rect 69902 344256 123482 344312
rect 123538 344256 123543 344312
rect 69841 344254 123543 344256
rect 69841 344251 69907 344254
rect 123477 344251 123543 344254
rect 296670 344254 360148 344314
rect 102041 344042 102107 344045
rect 155769 344042 155835 344045
rect 102041 344040 155835 344042
rect 102041 343984 102046 344040
rect 102102 343984 155774 344040
rect 155830 343984 155835 344040
rect 102041 343982 155835 343984
rect 102041 343979 102107 343982
rect 155769 343979 155835 343982
rect 119889 343906 119955 343909
rect 263593 343906 263659 343909
rect 264237 343906 264303 343909
rect 119889 343904 264303 343906
rect 119889 343848 119894 343904
rect 119950 343848 263598 343904
rect 263654 343848 264242 343904
rect 264298 343848 264303 343904
rect 119889 343846 264303 343848
rect 119889 343843 119955 343846
rect 263593 343843 263659 343846
rect 264237 343843 264303 343846
rect 124029 343770 124095 343773
rect 295374 343770 295380 343772
rect 124029 343768 295380 343770
rect 124029 343712 124034 343768
rect 124090 343712 295380 343768
rect 124029 343710 295380 343712
rect 124029 343707 124095 343710
rect 295374 343708 295380 343710
rect 295444 343770 295450 343772
rect 296670 343770 296730 344254
rect 360142 344252 360148 344254
rect 360212 344252 360218 344316
rect 295444 343710 296730 343770
rect 295444 343708 295450 343710
rect 113817 343634 113883 343637
rect 158805 343634 158871 343637
rect 113817 343632 158871 343634
rect 113817 343576 113822 343632
rect 113878 343576 158810 343632
rect 158866 343576 158871 343632
rect 113817 343574 158871 343576
rect 113817 343571 113883 343574
rect 158805 343571 158871 343574
rect 159449 342954 159515 342957
rect 168966 342954 168972 342956
rect 159449 342952 168972 342954
rect 159449 342896 159454 342952
rect 159510 342896 168972 342952
rect 159449 342894 168972 342896
rect 159449 342891 159515 342894
rect 168966 342892 168972 342894
rect 169036 342892 169042 342956
rect 211061 342954 211127 342957
rect 582373 342954 582439 342957
rect 211061 342952 582439 342954
rect 211061 342896 211066 342952
rect 211122 342896 582378 342952
rect 582434 342896 582439 342952
rect 211061 342894 582439 342896
rect 211061 342891 211127 342894
rect 582373 342891 582439 342894
rect 130469 342410 130535 342413
rect 131205 342410 131271 342413
rect 184381 342410 184447 342413
rect 130469 342408 184447 342410
rect 130469 342352 130474 342408
rect 130530 342352 131210 342408
rect 131266 342352 184386 342408
rect 184442 342352 184447 342408
rect 130469 342350 184447 342352
rect 130469 342347 130535 342350
rect 131205 342347 131271 342350
rect 184381 342347 184447 342350
rect 87137 342274 87203 342277
rect 209865 342274 209931 342277
rect 211061 342274 211127 342277
rect 87137 342272 211127 342274
rect 87137 342216 87142 342272
rect 87198 342216 209870 342272
rect 209926 342216 211066 342272
rect 211122 342216 211127 342272
rect 87137 342214 211127 342216
rect 87137 342211 87203 342214
rect 209865 342211 209931 342214
rect 211061 342211 211127 342214
rect 302233 342138 302299 342141
rect 307017 342138 307083 342141
rect 302233 342136 307083 342138
rect 302233 342080 302238 342136
rect 302294 342080 307022 342136
rect 307078 342080 307083 342136
rect 302233 342078 307083 342080
rect 302233 342075 302299 342078
rect 307017 342075 307083 342078
rect 142797 341594 142863 341597
rect 159398 341594 159404 341596
rect 142797 341592 159404 341594
rect 142797 341536 142802 341592
rect 142858 341536 159404 341592
rect 142797 341534 159404 341536
rect 142797 341531 142863 341534
rect 159398 341532 159404 341534
rect 159468 341532 159474 341596
rect 78438 341396 78444 341460
rect 78508 341458 78514 341460
rect 97257 341458 97323 341461
rect 78508 341456 97323 341458
rect 78508 341400 97262 341456
rect 97318 341400 97323 341456
rect 78508 341398 97323 341400
rect 78508 341396 78514 341398
rect 97257 341395 97323 341398
rect 155125 341458 155191 341461
rect 251766 341458 251772 341460
rect 155125 341456 251772 341458
rect 155125 341400 155130 341456
rect 155186 341400 251772 341456
rect 155125 341398 251772 341400
rect 155125 341395 155191 341398
rect 251766 341396 251772 341398
rect 251836 341396 251842 341460
rect 89529 341050 89595 341053
rect 155493 341050 155559 341053
rect 89529 341048 155559 341050
rect 89529 340992 89534 341048
rect 89590 340992 155498 341048
rect 155554 340992 155559 341048
rect 89529 340990 155559 340992
rect 89529 340987 89595 340990
rect 155493 340987 155559 340990
rect 111609 340914 111675 340917
rect 302233 340914 302299 340917
rect 111609 340912 302299 340914
rect 111609 340856 111614 340912
rect 111670 340856 302238 340912
rect 302294 340856 302299 340912
rect 111609 340854 302299 340856
rect 111609 340851 111675 340854
rect 302233 340851 302299 340854
rect 73470 340036 73476 340100
rect 73540 340098 73546 340100
rect 104157 340098 104223 340101
rect 73540 340096 104223 340098
rect 73540 340040 104162 340096
rect 104218 340040 104223 340096
rect 73540 340038 104223 340040
rect 73540 340036 73546 340038
rect 104157 340035 104223 340038
rect 153009 339826 153075 339829
rect 189901 339826 189967 339829
rect 153009 339824 189967 339826
rect 153009 339768 153014 339824
rect 153070 339768 189906 339824
rect 189962 339768 189967 339824
rect 153009 339766 189967 339768
rect 153009 339763 153075 339766
rect 189901 339763 189967 339766
rect 112345 339690 112411 339693
rect 212574 339690 212580 339692
rect 112345 339688 212580 339690
rect 112345 339632 112350 339688
rect 112406 339632 212580 339688
rect 112345 339630 212580 339632
rect 112345 339627 112411 339630
rect 212574 339628 212580 339630
rect 212644 339628 212650 339692
rect 81433 339554 81499 339557
rect 230422 339554 230428 339556
rect 81433 339552 230428 339554
rect 81433 339496 81438 339552
rect 81494 339496 230428 339552
rect 81433 339494 230428 339496
rect 81433 339491 81499 339494
rect 230422 339492 230428 339494
rect 230492 339492 230498 339556
rect 67950 339356 67956 339420
rect 68020 339418 68026 339420
rect 68870 339418 68876 339420
rect 68020 339358 68876 339418
rect 68020 339356 68026 339358
rect 68870 339356 68876 339358
rect 68940 339356 68946 339420
rect 117998 339356 118004 339420
rect 118068 339418 118074 339420
rect 118509 339418 118575 339421
rect 118068 339416 118575 339418
rect 118068 339360 118514 339416
rect 118570 339360 118575 339416
rect 118068 339358 118575 339360
rect 118068 339356 118074 339358
rect 118509 339355 118575 339358
rect 153837 339418 153903 339421
rect 156638 339418 156644 339420
rect 153837 339416 156644 339418
rect 153837 339360 153842 339416
rect 153898 339360 156644 339416
rect 153837 339358 156644 339360
rect 153837 339355 153903 339358
rect 156638 339356 156644 339358
rect 156708 339356 156714 339420
rect 57697 338738 57763 338741
rect 153009 338738 153075 338741
rect 57697 338736 153075 338738
rect 57697 338680 57702 338736
rect 57758 338680 153014 338736
rect 153070 338680 153075 338736
rect 57697 338678 153075 338680
rect 57697 338675 57763 338678
rect 153009 338675 153075 338678
rect 191189 338738 191255 338741
rect 201401 338738 201467 338741
rect 191189 338736 201467 338738
rect 191189 338680 191194 338736
rect 191250 338680 201406 338736
rect 201462 338680 201467 338736
rect 191189 338678 201467 338680
rect 191189 338675 191255 338678
rect 201401 338675 201467 338678
rect 210734 338676 210740 338740
rect 210804 338738 210810 338740
rect 236637 338738 236703 338741
rect 210804 338736 236703 338738
rect 210804 338680 236642 338736
rect 236698 338680 236703 338736
rect 210804 338678 236703 338680
rect 210804 338676 210810 338678
rect 236637 338675 236703 338678
rect 131757 338466 131823 338469
rect 122790 338464 131823 338466
rect 122790 338408 131762 338464
rect 131818 338408 131823 338464
rect 583520 338452 584960 338692
rect 122790 338406 131823 338408
rect 67950 338268 67956 338332
rect 68020 338330 68026 338332
rect 122790 338330 122850 338406
rect 131757 338403 131823 338406
rect 68020 338270 122850 338330
rect 131113 338330 131179 338333
rect 177481 338330 177547 338333
rect 131113 338328 177547 338330
rect 131113 338272 131118 338328
rect 131174 338272 177486 338328
rect 177542 338272 177547 338328
rect 131113 338270 177547 338272
rect 68020 338268 68026 338270
rect 131113 338267 131179 338270
rect 177481 338267 177547 338270
rect 85665 338194 85731 338197
rect 248597 338194 248663 338197
rect 85665 338192 248663 338194
rect 85665 338136 85670 338192
rect 85726 338136 248602 338192
rect 248658 338136 248663 338192
rect 85665 338134 248663 338136
rect 85665 338131 85731 338134
rect 248597 338131 248663 338134
rect 155493 338058 155559 338061
rect 176745 338058 176811 338061
rect 155493 338056 176811 338058
rect 155493 338000 155498 338056
rect 155554 338000 176750 338056
rect 176806 338000 176811 338056
rect 155493 337998 176811 338000
rect 155493 337995 155559 337998
rect 176745 337995 176811 337998
rect 202638 337588 202644 337652
rect 202708 337650 202714 337652
rect 209773 337650 209839 337653
rect 202708 337648 209839 337650
rect 202708 337592 209778 337648
rect 209834 337592 209839 337648
rect 202708 337590 209839 337592
rect 202708 337588 202714 337590
rect 209773 337587 209839 337590
rect 83958 337452 83964 337516
rect 84028 337514 84034 337516
rect 101397 337514 101463 337517
rect 84028 337512 101463 337514
rect 84028 337456 101402 337512
rect 101458 337456 101463 337512
rect 84028 337454 101463 337456
rect 84028 337452 84034 337454
rect 101397 337451 101463 337454
rect 147029 337514 147095 337517
rect 160921 337514 160987 337517
rect 204989 337514 205055 337517
rect 147029 337512 160987 337514
rect 147029 337456 147034 337512
rect 147090 337456 160926 337512
rect 160982 337456 160987 337512
rect 147029 337454 160987 337456
rect 147029 337451 147095 337454
rect 160921 337451 160987 337454
rect 161430 337512 205055 337514
rect 161430 337456 204994 337512
rect 205050 337456 205055 337512
rect 161430 337454 205055 337456
rect 161430 337381 161490 337454
rect 204989 337451 205055 337454
rect 77109 337378 77175 337381
rect 161381 337378 161490 337381
rect 77109 337376 161490 337378
rect 77109 337320 77114 337376
rect 77170 337320 161386 337376
rect 161442 337320 161490 337376
rect 77109 337318 161490 337320
rect 176745 337378 176811 337381
rect 177941 337378 178007 337381
rect 222837 337378 222903 337381
rect 176745 337376 222903 337378
rect 176745 337320 176750 337376
rect 176806 337320 177946 337376
rect 178002 337320 222842 337376
rect 222898 337320 222903 337376
rect 176745 337318 222903 337320
rect 77109 337315 77175 337318
rect 161381 337315 161447 337318
rect 176745 337315 176811 337318
rect 177941 337315 178007 337318
rect 222837 337315 222903 337318
rect 65885 336834 65951 336837
rect 155769 336834 155835 336837
rect 65885 336832 155835 336834
rect 65885 336776 65890 336832
rect 65946 336776 155774 336832
rect 155830 336776 155835 336832
rect 65885 336774 155835 336776
rect 65885 336771 65951 336774
rect 155769 336771 155835 336774
rect 81014 335956 81020 336020
rect 81084 336018 81090 336020
rect 371417 336018 371483 336021
rect 81084 336016 371483 336018
rect 81084 335960 371422 336016
rect 371478 335960 371483 336016
rect 81084 335958 371483 335960
rect 81084 335956 81090 335958
rect 371417 335955 371483 335958
rect 57605 335610 57671 335613
rect 189717 335610 189783 335613
rect 57605 335608 189783 335610
rect 57605 335552 57610 335608
rect 57666 335552 189722 335608
rect 189778 335552 189783 335608
rect 57605 335550 189783 335552
rect 57605 335547 57671 335550
rect 189717 335547 189783 335550
rect 69790 335412 69796 335476
rect 69860 335474 69866 335476
rect 229737 335474 229803 335477
rect 69860 335472 229803 335474
rect 69860 335416 229742 335472
rect 229798 335416 229803 335472
rect 69860 335414 229803 335416
rect 69860 335412 69866 335414
rect 229737 335411 229803 335414
rect 151077 334658 151143 334661
rect 154614 334658 154620 334660
rect 151077 334656 154620 334658
rect 151077 334600 151082 334656
rect 151138 334600 154620 334656
rect 151077 334598 154620 334600
rect 151077 334595 151143 334598
rect 154614 334596 154620 334598
rect 154684 334596 154690 334660
rect 155861 334658 155927 334661
rect 169017 334658 169083 334661
rect 155861 334656 169083 334658
rect 155861 334600 155866 334656
rect 155922 334600 169022 334656
rect 169078 334600 169083 334656
rect 155861 334598 169083 334600
rect 155861 334595 155927 334598
rect 169017 334595 169083 334598
rect 214414 334596 214420 334660
rect 214484 334658 214490 334660
rect 248413 334658 248479 334661
rect 214484 334656 248479 334658
rect 214484 334600 248418 334656
rect 248474 334600 248479 334656
rect 214484 334598 248479 334600
rect 214484 334596 214490 334598
rect 248413 334595 248479 334598
rect 59261 334386 59327 334389
rect 149053 334386 149119 334389
rect 59261 334384 149119 334386
rect 59261 334328 59266 334384
rect 59322 334328 149058 334384
rect 149114 334328 149119 334384
rect 59261 334326 149119 334328
rect 59261 334323 59327 334326
rect 149053 334323 149119 334326
rect 146753 334250 146819 334253
rect 222326 334250 222332 334252
rect 146753 334248 222332 334250
rect 146753 334192 146758 334248
rect 146814 334192 222332 334248
rect 146753 334190 222332 334192
rect 146753 334187 146819 334190
rect 222326 334188 222332 334190
rect 222396 334188 222402 334252
rect 72233 334114 72299 334117
rect 216029 334114 216095 334117
rect 72233 334112 216095 334114
rect 72233 334056 72238 334112
rect 72294 334056 216034 334112
rect 216090 334056 216095 334112
rect 72233 334054 216095 334056
rect 72233 334051 72299 334054
rect 216029 334051 216095 334054
rect 97809 332890 97875 332893
rect 176101 332890 176167 332893
rect 97809 332888 176167 332890
rect 97809 332832 97814 332888
rect 97870 332832 176106 332888
rect 176162 332832 176167 332888
rect 97809 332830 176167 332832
rect 97809 332827 97875 332830
rect 176101 332827 176167 332830
rect 63217 332754 63283 332757
rect 166441 332754 166507 332757
rect 63217 332752 166507 332754
rect 63217 332696 63222 332752
rect 63278 332696 166446 332752
rect 166502 332696 166507 332752
rect 63217 332694 166507 332696
rect 63217 332691 63283 332694
rect 166441 332691 166507 332694
rect 117037 332618 117103 332621
rect 247033 332618 247099 332621
rect 117037 332616 247099 332618
rect 117037 332560 117042 332616
rect 117098 332560 247038 332616
rect 247094 332560 247099 332616
rect 117037 332558 247099 332560
rect 117037 332555 117103 332558
rect 247033 332555 247099 332558
rect -960 332196 480 332436
rect 175181 332074 175247 332077
rect 191189 332074 191255 332077
rect 161430 332072 191255 332074
rect 161430 332016 175186 332072
rect 175242 332016 191194 332072
rect 191250 332016 191255 332072
rect 161430 332014 191255 332016
rect 154849 331938 154915 331941
rect 155718 331938 155724 331940
rect 154849 331936 155724 331938
rect 154849 331880 154854 331936
rect 154910 331880 155724 331936
rect 154849 331878 155724 331880
rect 154849 331875 154915 331878
rect 155718 331876 155724 331878
rect 155788 331876 155794 331940
rect 70025 331802 70091 331805
rect 161430 331802 161490 332014
rect 175181 332011 175247 332014
rect 191189 332011 191255 332014
rect 180333 331938 180399 331941
rect 189942 331938 189948 331940
rect 180333 331936 189948 331938
rect 180333 331880 180338 331936
rect 180394 331880 189948 331936
rect 180333 331878 189948 331880
rect 180333 331875 180399 331878
rect 189942 331876 189948 331878
rect 190012 331876 190018 331940
rect 70025 331800 161490 331802
rect 70025 331744 70030 331800
rect 70086 331744 161490 331800
rect 70025 331742 161490 331744
rect 190085 331802 190151 331805
rect 232078 331802 232084 331804
rect 190085 331800 232084 331802
rect 190085 331744 190090 331800
rect 190146 331744 232084 331800
rect 190085 331742 232084 331744
rect 70025 331739 70091 331742
rect 190085 331739 190151 331742
rect 232078 331740 232084 331742
rect 232148 331740 232154 331804
rect 141877 331394 141943 331397
rect 156822 331394 156828 331396
rect 141877 331392 156828 331394
rect 141877 331336 141882 331392
rect 141938 331336 156828 331392
rect 141877 331334 156828 331336
rect 141877 331331 141943 331334
rect 156822 331332 156828 331334
rect 156892 331332 156898 331396
rect 157425 331394 157491 331397
rect 158478 331394 158484 331396
rect 157425 331392 158484 331394
rect 157425 331336 157430 331392
rect 157486 331336 158484 331392
rect 157425 331334 158484 331336
rect 157425 331331 157491 331334
rect 158478 331332 158484 331334
rect 158548 331332 158554 331396
rect 75177 331258 75243 331261
rect 75678 331258 75684 331260
rect 75177 331256 75684 331258
rect 75177 331200 75182 331256
rect 75238 331200 75684 331256
rect 75177 331198 75684 331200
rect 75177 331195 75243 331198
rect 75678 331196 75684 331198
rect 75748 331258 75754 331260
rect 75821 331258 75887 331261
rect 75748 331256 75887 331258
rect 75748 331200 75826 331256
rect 75882 331200 75887 331256
rect 75748 331198 75887 331200
rect 75748 331196 75754 331198
rect 75821 331195 75887 331198
rect 114461 331258 114527 331261
rect 258073 331258 258139 331261
rect 114461 331256 258139 331258
rect 114461 331200 114466 331256
rect 114522 331200 258078 331256
rect 258134 331200 258139 331256
rect 114461 331198 258139 331200
rect 114461 331195 114527 331198
rect 258073 331195 258139 331198
rect 178861 330442 178927 330445
rect 206553 330442 206619 330445
rect 178861 330440 206619 330442
rect 178861 330384 178866 330440
rect 178922 330384 206558 330440
rect 206614 330384 206619 330440
rect 178861 330382 206619 330384
rect 178861 330379 178927 330382
rect 206553 330379 206619 330382
rect 91921 330170 91987 330173
rect 93894 330170 93900 330172
rect 91921 330168 93900 330170
rect 91921 330112 91926 330168
rect 91982 330112 93900 330168
rect 91921 330110 93900 330112
rect 91921 330107 91987 330110
rect 93894 330108 93900 330110
rect 93964 330170 93970 330172
rect 173249 330170 173315 330173
rect 93964 330168 173315 330170
rect 93964 330112 173254 330168
rect 173310 330112 173315 330168
rect 93964 330110 173315 330112
rect 93964 330108 93970 330110
rect 173249 330107 173315 330110
rect 17217 330034 17283 330037
rect 124857 330034 124923 330037
rect 17217 330032 124923 330034
rect 17217 329976 17222 330032
rect 17278 329976 124862 330032
rect 124918 329976 124923 330032
rect 17217 329974 124923 329976
rect 17217 329971 17283 329974
rect 124857 329971 124923 329974
rect 152641 330034 152707 330037
rect 178033 330034 178099 330037
rect 152641 330032 178099 330034
rect 152641 329976 152646 330032
rect 152702 329976 178038 330032
rect 178094 329976 178099 330032
rect 152641 329974 178099 329976
rect 152641 329971 152707 329974
rect 178033 329971 178099 329974
rect 76649 329898 76715 329901
rect 239397 329898 239463 329901
rect 76649 329896 239463 329898
rect 76649 329840 76654 329896
rect 76710 329840 239402 329896
rect 239458 329840 239463 329896
rect 76649 329838 239463 329840
rect 76649 329835 76715 329838
rect 239397 329835 239463 329838
rect 168230 329700 168236 329764
rect 168300 329762 168306 329764
rect 168373 329762 168439 329765
rect 168300 329760 168439 329762
rect 168300 329704 168378 329760
rect 168434 329704 168439 329760
rect 168300 329702 168439 329704
rect 168300 329700 168306 329702
rect 168373 329699 168439 329702
rect 69841 329626 69907 329629
rect 69246 329624 69907 329626
rect 69246 329568 69846 329624
rect 69902 329568 69907 329624
rect 69246 329566 69907 329568
rect 66621 328946 66687 328949
rect 69246 328946 69306 329566
rect 69841 329563 69907 329566
rect 69422 329156 69428 329220
rect 69492 329218 69498 329220
rect 71078 329218 71084 329220
rect 69492 329158 71084 329218
rect 69492 329156 69498 329158
rect 71078 329156 71084 329158
rect 71148 329156 71154 329220
rect 77150 329156 77156 329220
rect 77220 329218 77226 329220
rect 77477 329218 77543 329221
rect 77220 329216 77543 329218
rect 77220 329160 77482 329216
rect 77538 329160 77543 329216
rect 77220 329158 77543 329160
rect 77220 329156 77226 329158
rect 77477 329155 77543 329158
rect 82670 329156 82676 329220
rect 82740 329218 82746 329220
rect 83181 329218 83247 329221
rect 82740 329216 83247 329218
rect 82740 329160 83186 329216
rect 83242 329160 83247 329216
rect 82740 329158 83247 329160
rect 82740 329156 82746 329158
rect 83181 329155 83247 329158
rect 156781 329082 156847 329085
rect 211889 329082 211955 329085
rect 156781 329080 211955 329082
rect 156781 329024 156786 329080
rect 156842 329024 211894 329080
rect 211950 329024 211955 329080
rect 156781 329022 211955 329024
rect 156781 329019 156847 329022
rect 211889 329019 211955 329022
rect 66621 328944 69306 328946
rect 66621 328888 66626 328944
rect 66682 328916 69306 328944
rect 66682 328888 69276 328916
rect 66621 328886 69276 328888
rect 66621 328883 66687 328886
rect 158897 328674 158963 328677
rect 250069 328674 250135 328677
rect 156676 328672 158963 328674
rect 156676 328616 158902 328672
rect 158958 328616 158963 328672
rect 156676 328614 158963 328616
rect 158897 328611 158963 328614
rect 161430 328672 250135 328674
rect 161430 328616 250074 328672
rect 250130 328616 250135 328672
rect 161430 328614 250135 328616
rect 157241 328538 157307 328541
rect 161430 328538 161490 328614
rect 250069 328611 250135 328614
rect 157241 328536 161490 328538
rect 157241 328480 157246 328536
rect 157302 328480 161490 328536
rect 157241 328478 161490 328480
rect 194133 328538 194199 328541
rect 255262 328538 255268 328540
rect 194133 328536 255268 328538
rect 194133 328480 194138 328536
rect 194194 328480 255268 328536
rect 194133 328478 255268 328480
rect 157241 328475 157307 328478
rect 194133 328475 194199 328478
rect 255262 328476 255268 328478
rect 255332 328476 255338 328540
rect 69422 328340 69428 328404
rect 69492 328340 69498 328404
rect 160921 328402 160987 328405
rect 215385 328402 215451 328405
rect 160921 328400 215451 328402
rect 160921 328344 160926 328400
rect 160982 328344 215390 328400
rect 215446 328344 215451 328400
rect 160921 328342 215451 328344
rect 69430 327828 69490 328340
rect 160921 328339 160987 328342
rect 215385 328339 215451 328342
rect 158897 327586 158963 327589
rect 156676 327584 158963 327586
rect 156676 327528 158902 327584
rect 158958 327528 158963 327584
rect 156676 327526 158963 327528
rect 158897 327523 158963 327526
rect 169518 327116 169524 327180
rect 169588 327178 169594 327180
rect 172605 327178 172671 327181
rect 169588 327176 172671 327178
rect 169588 327120 172610 327176
rect 172666 327120 172671 327176
rect 169588 327118 172671 327120
rect 169588 327116 169594 327118
rect 172605 327115 172671 327118
rect 68878 326090 68938 326740
rect 158989 326498 159055 326501
rect 156676 326496 159055 326498
rect 156676 326440 158994 326496
rect 159050 326440 159055 326496
rect 156676 326438 159055 326440
rect 158989 326435 159055 326438
rect 156822 326300 156828 326364
rect 156892 326362 156898 326364
rect 239489 326362 239555 326365
rect 156892 326360 239555 326362
rect 156892 326304 239494 326360
rect 239550 326304 239555 326360
rect 156892 326302 239555 326304
rect 156892 326300 156898 326302
rect 239489 326299 239555 326302
rect 64830 326030 68938 326090
rect 61878 325756 61884 325820
rect 61948 325818 61954 325820
rect 64830 325818 64890 326030
rect 61948 325758 64890 325818
rect 61948 325756 61954 325758
rect 169845 325682 169911 325685
rect 197997 325682 198063 325685
rect 169845 325680 198063 325682
rect 69430 325548 69490 325652
rect 169845 325624 169850 325680
rect 169906 325624 198002 325680
rect 198058 325624 198063 325680
rect 169845 325622 198063 325624
rect 169845 325619 169911 325622
rect 197997 325619 198063 325622
rect 69422 325484 69428 325548
rect 69492 325484 69498 325548
rect 159081 325410 159147 325413
rect 156676 325408 159147 325410
rect 156676 325352 159086 325408
rect 159142 325352 159147 325408
rect 156676 325350 159147 325352
rect 159081 325347 159147 325350
rect 582925 325274 582991 325277
rect 583520 325274 584960 325364
rect 582925 325272 584960 325274
rect 582925 325216 582930 325272
rect 582986 325216 584960 325272
rect 582925 325214 584960 325216
rect 582925 325211 582991 325214
rect 583520 325124 584960 325214
rect 158161 325002 158227 325005
rect 178033 325002 178099 325005
rect 158161 325000 178099 325002
rect 158161 324944 158166 325000
rect 158222 324944 178038 325000
rect 178094 324944 178099 325000
rect 158161 324942 178099 324944
rect 158161 324939 158227 324942
rect 178033 324939 178099 324942
rect 211981 325002 212047 325005
rect 331857 325002 331923 325005
rect 211981 325000 331923 325002
rect 211981 324944 211986 325000
rect 212042 324944 331862 325000
rect 331918 324944 331923 325000
rect 211981 324942 331923 324944
rect 211981 324939 212047 324942
rect 331857 324939 331923 324942
rect 67265 324594 67331 324597
rect 67265 324592 68908 324594
rect 67265 324536 67270 324592
rect 67326 324536 68908 324592
rect 67265 324534 68908 324536
rect 67265 324531 67331 324534
rect 158897 324322 158963 324325
rect 156676 324320 158963 324322
rect 156676 324264 158902 324320
rect 158958 324264 158963 324320
rect 156676 324262 158963 324264
rect 158897 324259 158963 324262
rect 69422 323988 69428 324052
rect 69492 323988 69498 324052
rect 69430 323476 69490 323988
rect 188705 323642 188771 323645
rect 221549 323642 221615 323645
rect 188705 323640 221615 323642
rect 188705 323584 188710 323640
rect 188766 323584 221554 323640
rect 221610 323584 221615 323640
rect 188705 323582 221615 323584
rect 188705 323579 188771 323582
rect 221549 323579 221615 323582
rect 243537 323642 243603 323645
rect 291142 323642 291148 323644
rect 243537 323640 291148 323642
rect 243537 323584 243542 323640
rect 243598 323584 291148 323640
rect 243537 323582 291148 323584
rect 243537 323579 243603 323582
rect 291142 323580 291148 323582
rect 291212 323580 291218 323644
rect 158713 323234 158779 323237
rect 156676 323232 158779 323234
rect 156676 323176 158718 323232
rect 158774 323176 158779 323232
rect 156676 323174 158779 323176
rect 158713 323171 158779 323174
rect 65793 322418 65859 322421
rect 65977 322418 66043 322421
rect 65793 322416 68908 322418
rect 65793 322360 65798 322416
rect 65854 322360 65982 322416
rect 66038 322360 68908 322416
rect 65793 322358 68908 322360
rect 65793 322355 65859 322358
rect 65977 322355 66043 322358
rect 183001 322282 183067 322285
rect 195094 322282 195100 322284
rect 183001 322280 195100 322282
rect 183001 322224 183006 322280
rect 183062 322224 195100 322280
rect 183001 322222 195100 322224
rect 183001 322219 183067 322222
rect 195094 322220 195100 322222
rect 195164 322220 195170 322284
rect 158713 322146 158779 322149
rect 156676 322144 158779 322146
rect 156676 322088 158718 322144
rect 158774 322088 158779 322144
rect 156676 322086 158779 322088
rect 158713 322083 158779 322086
rect 183185 322146 183251 322149
rect 233969 322146 234035 322149
rect 183185 322144 234035 322146
rect 183185 322088 183190 322144
rect 183246 322088 233974 322144
rect 234030 322088 234035 322144
rect 183185 322086 234035 322088
rect 183185 322083 183251 322086
rect 233969 322083 234035 322086
rect 238017 322146 238083 322149
rect 253054 322146 253060 322148
rect 238017 322144 253060 322146
rect 238017 322088 238022 322144
rect 238078 322088 253060 322144
rect 238017 322086 253060 322088
rect 238017 322083 238083 322086
rect 253054 322084 253060 322086
rect 253124 322084 253130 322148
rect 66805 321330 66871 321333
rect 66805 321328 68908 321330
rect 66805 321272 66810 321328
rect 66866 321272 68908 321328
rect 66805 321270 68908 321272
rect 66805 321267 66871 321270
rect 156646 320378 156706 321028
rect 192477 320786 192543 320789
rect 224309 320786 224375 320789
rect 192477 320784 224375 320786
rect 192477 320728 192482 320784
rect 192538 320728 224314 320784
rect 224370 320728 224375 320784
rect 192477 320726 224375 320728
rect 192477 320723 192543 320726
rect 224309 320723 224375 320726
rect 156646 320318 161490 320378
rect 66897 320242 66963 320245
rect 161430 320242 161490 320318
rect 189073 320242 189139 320245
rect 66897 320240 68908 320242
rect 66897 320184 66902 320240
rect 66958 320184 68908 320240
rect 66897 320182 68908 320184
rect 161430 320240 189139 320242
rect 161430 320184 189078 320240
rect 189134 320184 189139 320240
rect 161430 320182 189139 320184
rect 66897 320179 66963 320182
rect 189073 320179 189139 320182
rect 156646 319426 156706 319940
rect 159357 319426 159423 319429
rect 173341 319426 173407 319429
rect 156646 319424 173407 319426
rect -960 319290 480 319380
rect 156646 319368 159362 319424
rect 159418 319368 173346 319424
rect 173402 319368 173407 319424
rect 156646 319366 173407 319368
rect 159357 319363 159423 319366
rect 173341 319363 173407 319366
rect 188429 319426 188495 319429
rect 233877 319426 233943 319429
rect 188429 319424 233943 319426
rect 188429 319368 188434 319424
rect 188490 319368 233882 319424
rect 233938 319368 233943 319424
rect 188429 319366 233943 319368
rect 188429 319363 188495 319366
rect 233877 319363 233943 319366
rect 4061 319290 4127 319293
rect -960 319288 4127 319290
rect -960 319232 4066 319288
rect 4122 319232 4127 319288
rect -960 319230 4127 319232
rect -960 319140 480 319230
rect 4061 319227 4127 319230
rect 66897 319154 66963 319157
rect 66897 319152 68908 319154
rect 66897 319096 66902 319152
rect 66958 319096 68908 319152
rect 66897 319094 68908 319096
rect 66897 319091 66963 319094
rect 159265 318882 159331 318885
rect 156676 318880 159331 318882
rect 156676 318824 159270 318880
rect 159326 318824 159331 318880
rect 156676 318822 159331 318824
rect 159265 318819 159331 318822
rect 66805 318066 66871 318069
rect 66805 318064 68908 318066
rect 66805 318008 66810 318064
rect 66866 318008 68908 318064
rect 66805 318006 68908 318008
rect 66805 318003 66871 318006
rect 176510 318004 176516 318068
rect 176580 318066 176586 318068
rect 206461 318066 206527 318069
rect 176580 318064 206527 318066
rect 176580 318008 206466 318064
rect 206522 318008 206527 318064
rect 176580 318006 206527 318008
rect 176580 318004 176586 318006
rect 206461 318003 206527 318006
rect 158713 317794 158779 317797
rect 156676 317792 158779 317794
rect 156676 317736 158718 317792
rect 158774 317736 158779 317792
rect 156676 317734 158779 317736
rect 158713 317731 158779 317734
rect 209221 317522 209287 317525
rect 209405 317522 209471 317525
rect 269757 317522 269823 317525
rect 209221 317520 269823 317522
rect 209221 317464 209226 317520
rect 209282 317464 209410 317520
rect 209466 317464 269762 317520
rect 269818 317464 269823 317520
rect 209221 317462 269823 317464
rect 209221 317459 209287 317462
rect 209405 317459 209471 317462
rect 269757 317459 269823 317462
rect 67357 316978 67423 316981
rect 67357 316976 68908 316978
rect 67357 316920 67362 316976
rect 67418 316920 68908 316976
rect 67357 316918 68908 316920
rect 67357 316915 67423 316918
rect 158713 316706 158779 316709
rect 156676 316704 158779 316706
rect 156676 316648 158718 316704
rect 158774 316648 158779 316704
rect 156676 316646 158779 316648
rect 158713 316643 158779 316646
rect 160829 316706 160895 316709
rect 178033 316706 178099 316709
rect 160829 316704 180810 316706
rect 160829 316648 160834 316704
rect 160890 316648 178038 316704
rect 178094 316648 180810 316704
rect 160829 316646 180810 316648
rect 160829 316643 160895 316646
rect 178033 316643 178099 316646
rect 180750 316162 180810 316646
rect 213269 316162 213335 316165
rect 180750 316160 213335 316162
rect 180750 316104 213274 316160
rect 213330 316104 213335 316160
rect 180750 316102 213335 316104
rect 213269 316099 213335 316102
rect 174997 316026 175063 316029
rect 156646 316024 175063 316026
rect 156646 315968 175002 316024
rect 175058 315968 175063 316024
rect 156646 315966 175063 315968
rect 66253 315890 66319 315893
rect 66253 315888 68908 315890
rect 66253 315832 66258 315888
rect 66314 315832 68908 315888
rect 66253 315830 68908 315832
rect 66253 315827 66319 315830
rect 156646 315588 156706 315966
rect 174997 315963 175063 315966
rect 174997 315346 175063 315349
rect 185342 315346 185348 315348
rect 174997 315344 185348 315346
rect 174997 315288 175002 315344
rect 175058 315288 185348 315344
rect 174997 315286 185348 315288
rect 174997 315283 175063 315286
rect 185342 315284 185348 315286
rect 185412 315284 185418 315348
rect 209129 315346 209195 315349
rect 249742 315346 249748 315348
rect 209129 315344 249748 315346
rect 209129 315288 209134 315344
rect 209190 315288 249748 315344
rect 209129 315286 249748 315288
rect 209129 315283 209195 315286
rect 249742 315284 249748 315286
rect 249812 315284 249818 315348
rect 52269 314938 52335 314941
rect 52269 314936 68938 314938
rect 52269 314880 52274 314936
rect 52330 314880 68938 314936
rect 52269 314878 68938 314880
rect 52269 314875 52335 314878
rect 68878 314772 68938 314878
rect 198590 314740 198596 314804
rect 198660 314802 198666 314804
rect 277894 314802 277900 314804
rect 198660 314742 277900 314802
rect 198660 314740 198666 314742
rect 277894 314740 277900 314742
rect 277964 314740 277970 314804
rect 66805 313986 66871 313989
rect 156646 313986 156706 314500
rect 174670 314196 174676 314260
rect 174740 314258 174746 314260
rect 185669 314258 185735 314261
rect 174740 314256 185735 314258
rect 174740 314200 185674 314256
rect 185730 314200 185735 314256
rect 174740 314198 185735 314200
rect 174740 314196 174746 314198
rect 185669 314195 185735 314198
rect 181529 314122 181595 314125
rect 215334 314122 215340 314124
rect 181529 314120 215340 314122
rect 181529 314064 181534 314120
rect 181590 314064 215340 314120
rect 181529 314062 215340 314064
rect 181529 314059 181595 314062
rect 215334 314060 215340 314062
rect 215404 314060 215410 314124
rect 164141 313986 164207 313989
rect 243905 313986 243971 313989
rect 66805 313984 68908 313986
rect 66805 313928 66810 313984
rect 66866 313928 68908 313984
rect 66805 313926 68908 313928
rect 156646 313984 243971 313986
rect 156646 313928 164146 313984
rect 164202 313928 243910 313984
rect 243966 313928 243971 313984
rect 156646 313926 243971 313928
rect 66805 313923 66871 313926
rect 164141 313923 164207 313926
rect 243905 313923 243971 313926
rect 158713 313442 158779 313445
rect 156676 313440 158779 313442
rect 156676 313384 158718 313440
rect 158774 313384 158779 313440
rect 156676 313382 158779 313384
rect 158713 313379 158779 313382
rect 66437 312898 66503 312901
rect 66437 312896 68908 312898
rect 66437 312840 66442 312896
rect 66498 312840 68908 312896
rect 66437 312838 68908 312840
rect 66437 312835 66503 312838
rect 202229 312626 202295 312629
rect 227161 312626 227227 312629
rect 202229 312624 227227 312626
rect 202229 312568 202234 312624
rect 202290 312568 227166 312624
rect 227222 312568 227227 312624
rect 202229 312566 227227 312568
rect 202229 312563 202295 312566
rect 227161 312563 227227 312566
rect 200614 312428 200620 312492
rect 200684 312490 200690 312492
rect 213862 312490 213868 312492
rect 200684 312430 213868 312490
rect 200684 312428 200690 312430
rect 213862 312428 213868 312430
rect 213932 312428 213938 312492
rect 214557 312490 214623 312493
rect 345013 312490 345079 312493
rect 214557 312488 345079 312490
rect 214557 312432 214562 312488
rect 214618 312432 345018 312488
rect 345074 312432 345079 312488
rect 214557 312430 345079 312432
rect 214557 312427 214623 312430
rect 345013 312427 345079 312430
rect 156646 311946 156706 312324
rect 583017 312082 583083 312085
rect 583520 312082 584960 312172
rect 583017 312080 584960 312082
rect 583017 312024 583022 312080
rect 583078 312024 584960 312080
rect 583017 312022 584960 312024
rect 583017 312019 583083 312022
rect 160686 311946 160692 311948
rect 156646 311886 160692 311946
rect 160686 311884 160692 311886
rect 160756 311946 160762 311948
rect 160829 311946 160895 311949
rect 160756 311944 160895 311946
rect 160756 311888 160834 311944
rect 160890 311888 160895 311944
rect 583520 311932 584960 312022
rect 160756 311886 160895 311888
rect 160756 311884 160762 311886
rect 160829 311883 160895 311886
rect 66989 311810 67055 311813
rect 66989 311808 68908 311810
rect 66989 311752 66994 311808
rect 67050 311752 68908 311808
rect 66989 311750 68908 311752
rect 66989 311747 67055 311750
rect 158713 311266 158779 311269
rect 156676 311264 158779 311266
rect 156676 311208 158718 311264
rect 158774 311208 158779 311264
rect 156676 311206 158779 311208
rect 158713 311203 158779 311206
rect 213177 311266 213243 311269
rect 230381 311266 230447 311269
rect 213177 311264 230447 311266
rect 213177 311208 213182 311264
rect 213238 311208 230386 311264
rect 230442 311208 230447 311264
rect 213177 311206 230447 311208
rect 213177 311203 213243 311206
rect 230381 311203 230447 311206
rect 159909 311130 159975 311133
rect 173157 311130 173223 311133
rect 159909 311128 173223 311130
rect 159909 311072 159914 311128
rect 159970 311072 173162 311128
rect 173218 311072 173223 311128
rect 159909 311070 173223 311072
rect 159909 311067 159975 311070
rect 173157 311067 173223 311070
rect 226425 311130 226491 311133
rect 332593 311130 332659 311133
rect 226425 311128 332659 311130
rect 226425 311072 226430 311128
rect 226486 311072 332598 311128
rect 332654 311072 332659 311128
rect 226425 311070 332659 311072
rect 226425 311067 226491 311070
rect 332593 311067 332659 311070
rect 67449 310722 67515 310725
rect 67633 310722 67699 310725
rect 67449 310720 68908 310722
rect 67449 310664 67454 310720
rect 67510 310664 67638 310720
rect 67694 310664 68908 310720
rect 67449 310662 68908 310664
rect 67449 310659 67515 310662
rect 67633 310659 67699 310662
rect 303705 310450 303771 310453
rect 304257 310450 304323 310453
rect 303705 310448 304323 310450
rect 303705 310392 303710 310448
rect 303766 310392 304262 310448
rect 304318 310392 304323 310448
rect 303705 310390 304323 310392
rect 303705 310387 303771 310390
rect 304257 310387 304323 310390
rect 158805 310178 158871 310181
rect 156676 310176 158871 310178
rect 156676 310120 158810 310176
rect 158866 310120 158871 310176
rect 156676 310118 158871 310120
rect 158805 310115 158871 310118
rect 159214 309708 159220 309772
rect 159284 309770 159290 309772
rect 164877 309770 164943 309773
rect 159284 309768 164943 309770
rect 159284 309712 164882 309768
rect 164938 309712 164943 309768
rect 159284 309710 164943 309712
rect 159284 309708 159290 309710
rect 164877 309707 164943 309710
rect 200113 309770 200179 309773
rect 200757 309770 200823 309773
rect 303705 309770 303771 309773
rect 200113 309768 303771 309770
rect 200113 309712 200118 309768
rect 200174 309712 200762 309768
rect 200818 309712 303710 309768
rect 303766 309712 303771 309768
rect 200113 309710 303771 309712
rect 200113 309707 200179 309710
rect 200757 309707 200823 309710
rect 303705 309707 303771 309710
rect 66805 309634 66871 309637
rect 66805 309632 68908 309634
rect 66805 309576 66810 309632
rect 66866 309576 68908 309632
rect 66805 309574 68908 309576
rect 66805 309571 66871 309574
rect 159950 309090 159956 309092
rect 156676 309030 159956 309090
rect 159950 309028 159956 309030
rect 160020 309028 160026 309092
rect 67817 308546 67883 308549
rect 67817 308544 68908 308546
rect 67817 308488 67822 308544
rect 67878 308488 68908 308544
rect 67817 308486 68908 308488
rect 67817 308483 67883 308486
rect 159950 308348 159956 308412
rect 160020 308410 160026 308412
rect 322197 308410 322263 308413
rect 160020 308408 322263 308410
rect 160020 308352 322202 308408
rect 322258 308352 322263 308408
rect 160020 308350 322263 308352
rect 160020 308348 160026 308350
rect 322197 308347 322263 308350
rect 158713 308002 158779 308005
rect 156676 308000 158779 308002
rect 156676 307944 158718 308000
rect 158774 307944 158779 308000
rect 156676 307942 158779 307944
rect 158713 307939 158779 307942
rect 281349 307730 281415 307733
rect 281574 307730 281580 307732
rect 281349 307728 281580 307730
rect 281349 307672 281354 307728
rect 281410 307672 281580 307728
rect 281349 307670 281580 307672
rect 281349 307667 281415 307670
rect 281574 307668 281580 307670
rect 281644 307668 281650 307732
rect 66897 307458 66963 307461
rect 66897 307456 68908 307458
rect 66897 307400 66902 307456
rect 66958 307400 68908 307456
rect 66897 307398 68908 307400
rect 66897 307395 66963 307398
rect 184289 307050 184355 307053
rect 226977 307050 227043 307053
rect 184289 307048 227043 307050
rect 184289 306992 184294 307048
rect 184350 306992 226982 307048
rect 227038 306992 227043 307048
rect 184289 306990 227043 306992
rect 184289 306987 184355 306990
rect 226977 306987 227043 306990
rect 158713 306914 158779 306917
rect 156676 306912 158779 306914
rect 156676 306856 158718 306912
rect 158774 306856 158779 306912
rect 156676 306854 158779 306856
rect 158713 306851 158779 306854
rect 205173 306506 205239 306509
rect 263542 306506 263548 306508
rect 205173 306504 263548 306506
rect 205173 306448 205178 306504
rect 205234 306448 263548 306504
rect 205173 306446 263548 306448
rect 205173 306443 205239 306446
rect 263542 306444 263548 306446
rect 263612 306444 263618 306508
rect 67081 306370 67147 306373
rect 67081 306368 68908 306370
rect -960 306234 480 306324
rect 67081 306312 67086 306368
rect 67142 306312 68908 306368
rect 67081 306310 68908 306312
rect 67081 306307 67147 306310
rect 3509 306234 3575 306237
rect -960 306232 3575 306234
rect -960 306176 3514 306232
rect 3570 306176 3575 306232
rect -960 306174 3575 306176
rect -960 306084 480 306174
rect 3509 306171 3575 306174
rect 158713 305826 158779 305829
rect 156676 305824 158779 305826
rect 156676 305768 158718 305824
rect 158774 305768 158779 305824
rect 156676 305766 158779 305768
rect 158713 305763 158779 305766
rect 207974 305764 207980 305828
rect 208044 305826 208050 305828
rect 227713 305826 227779 305829
rect 208044 305824 227779 305826
rect 208044 305768 227718 305824
rect 227774 305768 227779 305824
rect 208044 305766 227779 305768
rect 208044 305764 208050 305766
rect 227713 305763 227779 305766
rect 228357 305826 228423 305829
rect 240133 305826 240199 305829
rect 228357 305824 240199 305826
rect 228357 305768 228362 305824
rect 228418 305768 240138 305824
rect 240194 305768 240199 305824
rect 228357 305766 240199 305768
rect 228357 305763 228423 305766
rect 240133 305763 240199 305766
rect 193949 305690 194015 305693
rect 228633 305690 228699 305693
rect 193949 305688 228699 305690
rect 193949 305632 193954 305688
rect 194010 305632 228638 305688
rect 228694 305632 228699 305688
rect 193949 305630 228699 305632
rect 193949 305627 194015 305630
rect 228633 305627 228699 305630
rect 66805 305282 66871 305285
rect 66805 305280 68908 305282
rect 66805 305224 66810 305280
rect 66866 305224 68908 305280
rect 66805 305222 68908 305224
rect 66805 305219 66871 305222
rect 158713 304738 158779 304741
rect 156676 304736 158779 304738
rect 156676 304680 158718 304736
rect 158774 304680 158779 304736
rect 156676 304678 158779 304680
rect 158713 304675 158779 304678
rect 66805 304194 66871 304197
rect 66805 304192 68908 304194
rect 66805 304136 66810 304192
rect 66866 304136 68908 304192
rect 66805 304134 68908 304136
rect 66805 304131 66871 304134
rect 159398 303724 159404 303788
rect 159468 303786 159474 303788
rect 159468 303726 161490 303786
rect 159468 303724 159474 303726
rect 158805 303650 158871 303653
rect 156676 303648 158871 303650
rect 156676 303592 158810 303648
rect 158866 303592 158871 303648
rect 156676 303590 158871 303592
rect 161430 303650 161490 303726
rect 168966 303724 168972 303788
rect 169036 303786 169042 303788
rect 169293 303786 169359 303789
rect 225137 303786 225203 303789
rect 169036 303784 225203 303786
rect 169036 303728 169298 303784
rect 169354 303728 225142 303784
rect 225198 303728 225203 303784
rect 169036 303726 225203 303728
rect 169036 303724 169042 303726
rect 169293 303723 169359 303726
rect 225137 303723 225203 303726
rect 247718 303650 247724 303652
rect 161430 303590 247724 303650
rect 158805 303587 158871 303590
rect 247718 303588 247724 303590
rect 247788 303588 247794 303652
rect 65885 303106 65951 303109
rect 65885 303104 68908 303106
rect 65885 303048 65890 303104
rect 65946 303048 68908 303104
rect 65885 303046 68908 303048
rect 65885 303043 65951 303046
rect 218697 302970 218763 302973
rect 234613 302970 234679 302973
rect 218697 302968 234679 302970
rect 218697 302912 218702 302968
rect 218758 302912 234618 302968
rect 234674 302912 234679 302968
rect 218697 302910 234679 302912
rect 218697 302907 218763 302910
rect 234613 302907 234679 302910
rect 203609 302834 203675 302837
rect 227662 302834 227668 302836
rect 203609 302832 227668 302834
rect 203609 302776 203614 302832
rect 203670 302776 227668 302832
rect 203609 302774 227668 302776
rect 203609 302771 203675 302774
rect 227662 302772 227668 302774
rect 227732 302772 227738 302836
rect 156646 302290 156706 302532
rect 316769 302290 316835 302293
rect 156646 302288 316835 302290
rect 156646 302232 316774 302288
rect 316830 302232 316835 302288
rect 156646 302230 316835 302232
rect 316769 302227 316835 302230
rect 66805 302018 66871 302021
rect 66805 302016 68908 302018
rect 66805 301960 66810 302016
rect 66866 301960 68908 302016
rect 66805 301958 68908 301960
rect 66805 301955 66871 301958
rect 158805 301474 158871 301477
rect 156676 301472 158871 301474
rect 156676 301416 158810 301472
rect 158866 301416 158871 301472
rect 156676 301414 158871 301416
rect 158805 301411 158871 301414
rect 169017 301474 169083 301477
rect 186037 301474 186103 301477
rect 169017 301472 190470 301474
rect 169017 301416 169022 301472
rect 169078 301416 186042 301472
rect 186098 301416 190470 301472
rect 169017 301414 190470 301416
rect 169017 301411 169083 301414
rect 186037 301411 186103 301414
rect 190410 301066 190470 301414
rect 266997 301066 267063 301069
rect 190410 301064 267063 301066
rect 190410 301008 267002 301064
rect 267058 301008 267063 301064
rect 190410 301006 267063 301008
rect 266997 301003 267063 301006
rect 66897 300930 66963 300933
rect 195789 300932 195855 300933
rect 195789 300930 195836 300932
rect 66897 300928 68908 300930
rect 66897 300872 66902 300928
rect 66958 300872 68908 300928
rect 66897 300870 68908 300872
rect 195708 300928 195836 300930
rect 195900 300930 195906 300932
rect 279417 300930 279483 300933
rect 195900 300928 279483 300930
rect 195708 300872 195794 300928
rect 195900 300872 279422 300928
rect 279478 300872 279483 300928
rect 195708 300870 195836 300872
rect 66897 300867 66963 300870
rect 195789 300868 195836 300870
rect 195900 300870 279483 300872
rect 195900 300868 195906 300870
rect 195789 300867 195855 300868
rect 279417 300867 279483 300870
rect 157333 300386 157399 300389
rect 159449 300386 159515 300389
rect 156676 300384 159515 300386
rect 156676 300328 157338 300384
rect 157394 300328 159454 300384
rect 159510 300328 159515 300384
rect 156676 300326 159515 300328
rect 157333 300323 157399 300326
rect 159449 300323 159515 300326
rect 169017 300250 169083 300253
rect 188521 300250 188587 300253
rect 244089 300250 244155 300253
rect 169017 300248 244155 300250
rect 169017 300192 169022 300248
rect 169078 300192 188526 300248
rect 188582 300192 244094 300248
rect 244150 300192 244155 300248
rect 169017 300190 244155 300192
rect 169017 300187 169083 300190
rect 188521 300187 188587 300190
rect 244089 300187 244155 300190
rect 157926 300052 157932 300116
rect 157996 300114 158002 300116
rect 158478 300114 158484 300116
rect 157996 300054 158484 300114
rect 157996 300052 158002 300054
rect 158478 300052 158484 300054
rect 158548 300114 158554 300116
rect 256877 300114 256943 300117
rect 158548 300112 256943 300114
rect 158548 300056 256882 300112
rect 256938 300056 256943 300112
rect 158548 300054 256943 300056
rect 158548 300052 158554 300054
rect 256877 300051 256943 300054
rect 67541 299842 67607 299845
rect 67541 299840 68908 299842
rect 67541 299784 67546 299840
rect 67602 299784 68908 299840
rect 67541 299782 68908 299784
rect 67541 299779 67607 299782
rect 207013 299434 207079 299437
rect 207749 299434 207815 299437
rect 207013 299432 207815 299434
rect 207013 299376 207018 299432
rect 207074 299376 207754 299432
rect 207810 299376 207815 299432
rect 207013 299374 207815 299376
rect 207013 299371 207079 299374
rect 207749 299371 207815 299374
rect 66621 298756 66687 298757
rect 66621 298754 66668 298756
rect 66540 298752 66668 298754
rect 66732 298754 66738 298756
rect 66540 298696 66626 298752
rect 66540 298694 66668 298696
rect 66621 298692 66668 298694
rect 66732 298694 68908 298754
rect 66732 298692 66738 298694
rect 66621 298691 66687 298692
rect 156646 298618 156706 299268
rect 158805 298754 158871 298757
rect 242934 298754 242940 298756
rect 158805 298752 242940 298754
rect 158805 298696 158810 298752
rect 158866 298696 242940 298752
rect 158805 298694 242940 298696
rect 158805 298691 158871 298694
rect 242934 298692 242940 298694
rect 243004 298692 243010 298756
rect 580717 298754 580783 298757
rect 583520 298754 584960 298844
rect 580717 298752 584960 298754
rect 580717 298696 580722 298752
rect 580778 298696 584960 298752
rect 580717 298694 584960 298696
rect 580717 298691 580783 298694
rect 156646 298558 161490 298618
rect 583520 298604 584960 298694
rect 159633 298210 159699 298213
rect 156676 298208 159699 298210
rect 156676 298152 159638 298208
rect 159694 298152 159699 298208
rect 156676 298150 159699 298152
rect 161430 298210 161490 298558
rect 240358 298482 240364 298484
rect 219390 298422 240364 298482
rect 207013 298346 207079 298349
rect 219390 298346 219450 298422
rect 240358 298420 240364 298422
rect 240428 298420 240434 298484
rect 207013 298344 219450 298346
rect 207013 298288 207018 298344
rect 207074 298288 219450 298344
rect 207013 298286 219450 298288
rect 241421 298346 241487 298349
rect 284937 298346 285003 298349
rect 241421 298344 285003 298346
rect 241421 298288 241426 298344
rect 241482 298288 284942 298344
rect 284998 298288 285003 298344
rect 241421 298286 285003 298288
rect 207013 298283 207079 298286
rect 241421 298283 241487 298286
rect 284937 298283 285003 298286
rect 244406 298210 244412 298212
rect 161430 298150 244412 298210
rect 159633 298147 159699 298150
rect 244406 298148 244412 298150
rect 244476 298148 244482 298212
rect 184197 298074 184263 298077
rect 184841 298074 184907 298077
rect 184197 298072 184907 298074
rect 184197 298016 184202 298072
rect 184258 298016 184846 298072
rect 184902 298016 184907 298072
rect 184197 298014 184907 298016
rect 184197 298011 184263 298014
rect 184841 298011 184907 298014
rect 66805 297666 66871 297669
rect 66805 297664 68908 297666
rect 66805 297608 66810 297664
rect 66866 297608 68908 297664
rect 66805 297606 68908 297608
rect 66805 297603 66871 297606
rect 175733 297530 175799 297533
rect 184054 297530 184060 297532
rect 175733 297528 184060 297530
rect 175733 297472 175738 297528
rect 175794 297472 184060 297528
rect 175733 297470 184060 297472
rect 175733 297467 175799 297470
rect 184054 297468 184060 297470
rect 184124 297468 184130 297532
rect 223021 297530 223087 297533
rect 258717 297530 258783 297533
rect 223021 297528 258783 297530
rect 223021 297472 223026 297528
rect 223082 297472 258722 297528
rect 258778 297472 258783 297528
rect 223021 297470 258783 297472
rect 223021 297467 223087 297470
rect 258717 297467 258783 297470
rect 163589 297394 163655 297397
rect 246021 297394 246087 297397
rect 163589 297392 246087 297394
rect 163589 297336 163594 297392
rect 163650 297336 246026 297392
rect 246082 297336 246087 297392
rect 163589 297334 246087 297336
rect 163589 297331 163655 297334
rect 246021 297331 246087 297334
rect 158713 297122 158779 297125
rect 156676 297120 158779 297122
rect 156676 297064 158718 297120
rect 158774 297064 158779 297120
rect 156676 297062 158779 297064
rect 158713 297059 158779 297062
rect 184841 296850 184907 296853
rect 296805 296850 296871 296853
rect 184841 296848 296871 296850
rect 184841 296792 184846 296848
rect 184902 296792 296810 296848
rect 296866 296792 296871 296848
rect 184841 296790 296871 296792
rect 184841 296787 184907 296790
rect 296805 296787 296871 296790
rect 172462 296652 172468 296716
rect 172532 296714 172538 296716
rect 198825 296714 198891 296717
rect 172532 296712 198891 296714
rect 172532 296656 198830 296712
rect 198886 296656 198891 296712
rect 172532 296654 198891 296656
rect 172532 296652 172538 296654
rect 198825 296651 198891 296654
rect 357566 296652 357572 296716
rect 357636 296714 357642 296716
rect 580717 296714 580783 296717
rect 357636 296712 580783 296714
rect 357636 296656 580722 296712
rect 580778 296656 580783 296712
rect 357636 296654 580783 296656
rect 357636 296652 357642 296654
rect 580717 296651 580783 296654
rect 67725 296578 67791 296581
rect 67725 296576 68908 296578
rect 67725 296520 67730 296576
rect 67786 296520 68908 296576
rect 67725 296518 68908 296520
rect 67725 296515 67791 296518
rect 157006 296244 157012 296308
rect 157076 296306 157082 296308
rect 172462 296306 172468 296308
rect 157076 296246 172468 296306
rect 157076 296244 157082 296246
rect 172462 296244 172468 296246
rect 172532 296244 172538 296308
rect 206870 296244 206876 296308
rect 206940 296306 206946 296308
rect 219433 296306 219499 296309
rect 206940 296304 219499 296306
rect 206940 296248 219438 296304
rect 219494 296248 219499 296304
rect 206940 296246 219499 296248
rect 206940 296244 206946 296246
rect 219433 296243 219499 296246
rect 186129 296170 186195 296173
rect 212901 296170 212967 296173
rect 186129 296168 212967 296170
rect 186129 296112 186134 296168
rect 186190 296112 212906 296168
rect 212962 296112 212967 296168
rect 186129 296110 212967 296112
rect 186129 296107 186195 296110
rect 212901 296107 212967 296110
rect 219198 296108 219204 296172
rect 219268 296170 219274 296172
rect 266353 296170 266419 296173
rect 219268 296168 266419 296170
rect 219268 296112 266358 296168
rect 266414 296112 266419 296168
rect 219268 296110 266419 296112
rect 219268 296108 219274 296110
rect 266353 296107 266419 296110
rect 158713 296034 158779 296037
rect 156676 296032 158779 296034
rect 156676 295976 158718 296032
rect 158774 295976 158779 296032
rect 156676 295974 158779 295976
rect 158713 295971 158779 295974
rect 198825 296034 198891 296037
rect 249977 296034 250043 296037
rect 198825 296032 250043 296034
rect 198825 295976 198830 296032
rect 198886 295976 249982 296032
rect 250038 295976 250043 296032
rect 198825 295974 250043 295976
rect 198825 295971 198891 295974
rect 249977 295971 250043 295974
rect 298737 296034 298803 296037
rect 357566 296034 357572 296036
rect 298737 296032 357572 296034
rect 298737 295976 298742 296032
rect 298798 295976 357572 296032
rect 298737 295974 357572 295976
rect 298737 295971 298803 295974
rect 357566 295972 357572 295974
rect 357636 295972 357642 296036
rect 66713 295490 66779 295493
rect 66713 295488 68908 295490
rect 66713 295432 66718 295488
rect 66774 295432 68908 295488
rect 66713 295430 68908 295432
rect 66713 295427 66779 295430
rect 172513 295354 172579 295357
rect 173750 295354 173756 295356
rect 172513 295352 173756 295354
rect 172513 295296 172518 295352
rect 172574 295296 173756 295352
rect 172513 295294 173756 295296
rect 172513 295291 172579 295294
rect 173750 295292 173756 295294
rect 173820 295292 173826 295356
rect 203190 295292 203196 295356
rect 203260 295354 203266 295356
rect 206461 295354 206527 295357
rect 203260 295352 206527 295354
rect 203260 295296 206466 295352
rect 206522 295296 206527 295352
rect 203260 295294 206527 295296
rect 203260 295292 203266 295294
rect 206461 295291 206527 295294
rect 166349 295218 166415 295221
rect 156646 295216 166415 295218
rect 156646 295160 166354 295216
rect 166410 295160 166415 295216
rect 156646 295158 166415 295160
rect 156646 294916 156706 295158
rect 166349 295155 166415 295158
rect 211061 295218 211127 295221
rect 223021 295218 223087 295221
rect 211061 295216 223087 295218
rect 211061 295160 211066 295216
rect 211122 295160 223026 295216
rect 223082 295160 223087 295216
rect 211061 295158 223087 295160
rect 211061 295155 211127 295158
rect 223021 295155 223087 295158
rect 191189 294538 191255 294541
rect 200614 294538 200620 294540
rect 191189 294536 200620 294538
rect 191189 294480 191194 294536
rect 191250 294480 200620 294536
rect 191189 294478 200620 294480
rect 191189 294475 191255 294478
rect 200614 294476 200620 294478
rect 200684 294476 200690 294540
rect 66805 294402 66871 294405
rect 66805 294400 68908 294402
rect 66805 294344 66810 294400
rect 66866 294344 68908 294400
rect 66805 294342 68908 294344
rect 66805 294339 66871 294342
rect 276749 294130 276815 294133
rect 222702 294128 276815 294130
rect 222702 294072 276754 294128
rect 276810 294072 276815 294128
rect 222702 294070 276815 294072
rect 221181 293994 221247 293997
rect 221641 293994 221707 293997
rect 222702 293994 222762 294070
rect 276749 294067 276815 294070
rect 221181 293992 222762 293994
rect 221181 293936 221186 293992
rect 221242 293936 221646 293992
rect 221702 293936 222762 293992
rect 221181 293934 222762 293936
rect 222837 293994 222903 293997
rect 299565 293994 299631 293997
rect 222837 293992 299631 293994
rect 222837 293936 222842 293992
rect 222898 293936 299570 293992
rect 299626 293936 299631 293992
rect 222837 293934 299631 293936
rect 221181 293931 221247 293934
rect 221641 293931 221707 293934
rect 222837 293931 222903 293934
rect 299565 293931 299631 293934
rect 158713 293858 158779 293861
rect 156676 293856 158779 293858
rect 156676 293800 158718 293856
rect 158774 293800 158779 293856
rect 156676 293798 158779 293800
rect 158713 293795 158779 293798
rect 66805 293314 66871 293317
rect 66805 293312 68908 293314
rect -960 293178 480 293268
rect 66805 293256 66810 293312
rect 66866 293256 68908 293312
rect 66805 293254 68908 293256
rect 66805 293251 66871 293254
rect 3509 293178 3575 293181
rect -960 293176 3575 293178
rect -960 293120 3514 293176
rect 3570 293120 3575 293176
rect -960 293118 3575 293120
rect -960 293028 480 293118
rect 3509 293115 3575 293118
rect 163446 293116 163452 293180
rect 163516 293178 163522 293180
rect 184289 293178 184355 293181
rect 163516 293176 184355 293178
rect 163516 293120 184294 293176
rect 184350 293120 184355 293176
rect 163516 293118 184355 293120
rect 163516 293116 163522 293118
rect 184289 293115 184355 293118
rect 159357 293042 159423 293045
rect 156676 293040 159423 293042
rect 156676 292984 159362 293040
rect 159418 292984 159423 293040
rect 156676 292982 159423 292984
rect 159357 292979 159423 292982
rect 176009 292770 176075 292773
rect 249926 292770 249932 292772
rect 176009 292768 249932 292770
rect 176009 292712 176014 292768
rect 176070 292712 249932 292768
rect 176009 292710 249932 292712
rect 176009 292707 176075 292710
rect 249926 292708 249932 292710
rect 249996 292708 250002 292772
rect 196709 292634 196775 292637
rect 201677 292634 201743 292637
rect 582649 292634 582715 292637
rect 196709 292632 582715 292634
rect 196709 292576 196714 292632
rect 196770 292576 201682 292632
rect 201738 292576 582654 292632
rect 582710 292576 582715 292632
rect 196709 292574 582715 292576
rect 196709 292571 196775 292574
rect 201677 292571 201743 292574
rect 582649 292571 582715 292574
rect 159449 292498 159515 292501
rect 227897 292498 227963 292501
rect 159449 292496 227963 292498
rect 159449 292440 159454 292496
rect 159510 292440 227902 292496
rect 227958 292440 227963 292496
rect 159449 292438 227963 292440
rect 159449 292435 159515 292438
rect 227897 292435 227963 292438
rect 66805 292226 66871 292229
rect 66805 292224 68908 292226
rect 66805 292168 66810 292224
rect 66866 292168 68908 292224
rect 66805 292166 68908 292168
rect 66805 292163 66871 292166
rect 227897 292090 227963 292093
rect 228449 292090 228515 292093
rect 227897 292088 228515 292090
rect 227897 292032 227902 292088
rect 227958 292032 228454 292088
rect 228510 292032 228515 292088
rect 227897 292030 228515 292032
rect 227897 292027 227963 292030
rect 228449 292027 228515 292030
rect 158713 291954 158779 291957
rect 156676 291952 158779 291954
rect 156676 291896 158718 291952
rect 158774 291896 158779 291952
rect 156676 291894 158779 291896
rect 158713 291891 158779 291894
rect 180333 291818 180399 291821
rect 187233 291818 187299 291821
rect 180333 291816 187299 291818
rect 180333 291760 180338 291816
rect 180394 291760 187238 291816
rect 187294 291760 187299 291816
rect 180333 291758 187299 291760
rect 180333 291755 180399 291758
rect 187233 291755 187299 291758
rect 217542 291756 217548 291820
rect 217612 291818 217618 291820
rect 262213 291818 262279 291821
rect 217612 291816 262279 291818
rect 217612 291760 262218 291816
rect 262274 291760 262279 291816
rect 217612 291758 262279 291760
rect 217612 291756 217618 291758
rect 262213 291755 262279 291758
rect 188521 291274 188587 291277
rect 202229 291274 202295 291277
rect 188521 291272 202295 291274
rect 188521 291216 188526 291272
rect 188582 291216 202234 291272
rect 202290 291216 202295 291272
rect 188521 291214 202295 291216
rect 188521 291211 188587 291214
rect 202229 291211 202295 291214
rect 228633 291274 228699 291277
rect 228909 291274 228975 291277
rect 298185 291274 298251 291277
rect 228633 291272 298251 291274
rect 228633 291216 228638 291272
rect 228694 291216 228914 291272
rect 228970 291216 298190 291272
rect 298246 291216 298251 291272
rect 228633 291214 298251 291216
rect 228633 291211 228699 291214
rect 228909 291211 228975 291214
rect 298185 291211 298251 291214
rect 66805 291138 66871 291141
rect 211889 291138 211955 291141
rect 212441 291138 212507 291141
rect 280889 291138 280955 291141
rect 66805 291136 68908 291138
rect 66805 291080 66810 291136
rect 66866 291080 68908 291136
rect 66805 291078 68908 291080
rect 211889 291136 280955 291138
rect 211889 291080 211894 291136
rect 211950 291080 212446 291136
rect 212502 291080 280894 291136
rect 280950 291080 280955 291136
rect 211889 291078 280955 291080
rect 66805 291075 66871 291078
rect 211889 291075 211955 291078
rect 212441 291075 212507 291078
rect 280889 291075 280955 291078
rect 158713 290866 158779 290869
rect 156676 290864 158779 290866
rect 156676 290808 158718 290864
rect 158774 290808 158779 290864
rect 156676 290806 158779 290808
rect 158713 290803 158779 290806
rect 196934 290396 196940 290460
rect 197004 290458 197010 290460
rect 204437 290458 204503 290461
rect 197004 290456 204503 290458
rect 197004 290400 204442 290456
rect 204498 290400 204503 290456
rect 197004 290398 204503 290400
rect 197004 290396 197010 290398
rect 204437 290395 204503 290398
rect 66897 290050 66963 290053
rect 224309 290050 224375 290053
rect 226885 290050 226951 290053
rect 255313 290050 255379 290053
rect 66897 290048 68908 290050
rect 66897 289992 66902 290048
rect 66958 289992 68908 290048
rect 66897 289990 68908 289992
rect 224309 290048 255379 290050
rect 224309 289992 224314 290048
rect 224370 289992 226890 290048
rect 226946 289992 255318 290048
rect 255374 289992 255379 290048
rect 224309 289990 255379 289992
rect 66897 289987 66963 289990
rect 224309 289987 224375 289990
rect 226885 289987 226951 289990
rect 255313 289987 255379 289990
rect 192569 289914 192635 289917
rect 232773 289914 232839 289917
rect 192569 289912 232839 289914
rect 192569 289856 192574 289912
rect 192630 289856 232778 289912
rect 232834 289856 232839 289912
rect 192569 289854 232839 289856
rect 192569 289851 192635 289854
rect 232773 289851 232839 289854
rect 158805 289778 158871 289781
rect 156676 289776 158871 289778
rect 156676 289720 158810 289776
rect 158866 289720 158871 289776
rect 156676 289718 158871 289720
rect 158805 289715 158871 289718
rect 226517 289778 226583 289781
rect 227161 289778 227227 289781
rect 226517 289776 227227 289778
rect 226517 289720 226522 289776
rect 226578 289720 227166 289776
rect 227222 289720 227227 289776
rect 226517 289718 227227 289720
rect 226517 289715 226583 289718
rect 227161 289715 227227 289718
rect 156822 289172 156828 289236
rect 156892 289234 156898 289236
rect 208117 289234 208183 289237
rect 215937 289234 216003 289237
rect 156892 289232 216003 289234
rect 156892 289176 208122 289232
rect 208178 289176 215942 289232
rect 215998 289176 216003 289232
rect 156892 289174 216003 289176
rect 156892 289172 156898 289174
rect 208117 289171 208183 289174
rect 215937 289171 216003 289174
rect 174537 289098 174603 289101
rect 245837 289098 245903 289101
rect 174537 289096 245903 289098
rect 174537 289040 174542 289096
rect 174598 289040 245842 289096
rect 245898 289040 245903 289096
rect 174537 289038 245903 289040
rect 174537 289035 174603 289038
rect 245837 289035 245903 289038
rect 66805 288962 66871 288965
rect 66805 288960 68908 288962
rect 66805 288904 66810 288960
rect 66866 288904 68908 288960
rect 66805 288902 68908 288904
rect 66805 288899 66871 288902
rect 160870 288690 160876 288692
rect 156676 288630 160876 288690
rect 160870 288628 160876 288630
rect 160940 288628 160946 288692
rect 226517 288690 226583 288693
rect 271137 288690 271203 288693
rect 226517 288688 271203 288690
rect 226517 288632 226522 288688
rect 226578 288632 271142 288688
rect 271198 288632 271203 288688
rect 226517 288630 271203 288632
rect 226517 288627 226583 288630
rect 271137 288627 271203 288630
rect 201401 288554 201467 288557
rect 259545 288554 259611 288557
rect 201401 288552 259611 288554
rect 201401 288496 201406 288552
rect 201462 288496 259550 288552
rect 259606 288496 259611 288552
rect 201401 288494 259611 288496
rect 201401 288491 201467 288494
rect 259545 288491 259611 288494
rect 235165 288418 235231 288421
rect 235901 288418 235967 288421
rect 235165 288416 235967 288418
rect 235165 288360 235170 288416
rect 235226 288360 235906 288416
rect 235962 288360 235967 288416
rect 235165 288358 235967 288360
rect 235165 288355 235231 288358
rect 235901 288355 235967 288358
rect 240726 288356 240732 288420
rect 240796 288418 240802 288420
rect 240869 288418 240935 288421
rect 240796 288416 240935 288418
rect 240796 288360 240874 288416
rect 240930 288360 240935 288416
rect 240796 288358 240935 288360
rect 240796 288356 240802 288358
rect 240869 288355 240935 288358
rect 66621 287874 66687 287877
rect 66621 287872 68908 287874
rect 66621 287816 66626 287872
rect 66682 287816 68908 287872
rect 66621 287814 68908 287816
rect 66621 287811 66687 287814
rect 165153 287738 165219 287741
rect 184013 287738 184079 287741
rect 165153 287736 184079 287738
rect 165153 287680 165158 287736
rect 165214 287680 184018 287736
rect 184074 287680 184079 287736
rect 165153 287678 184079 287680
rect 165153 287675 165219 287678
rect 184013 287675 184079 287678
rect 233141 287738 233207 287741
rect 259729 287738 259795 287741
rect 583569 287738 583635 287741
rect 233141 287736 583635 287738
rect 233141 287680 233146 287736
rect 233202 287680 259734 287736
rect 259790 287680 583574 287736
rect 583630 287680 583635 287736
rect 233141 287678 583635 287680
rect 233141 287675 233207 287678
rect 259729 287675 259795 287678
rect 583569 287675 583635 287678
rect 158713 287602 158779 287605
rect 156676 287600 158779 287602
rect 156676 287544 158718 287600
rect 158774 287544 158779 287600
rect 156676 287542 158779 287544
rect 158713 287539 158779 287542
rect 180241 287602 180307 287605
rect 230749 287602 230815 287605
rect 180241 287600 230815 287602
rect 180241 287544 180246 287600
rect 180302 287544 230754 287600
rect 230810 287544 230815 287600
rect 180241 287542 230815 287544
rect 180241 287539 180307 287542
rect 230749 287539 230815 287542
rect 199326 287404 199332 287468
rect 199396 287466 199402 287468
rect 211797 287466 211863 287469
rect 199396 287464 211863 287466
rect 199396 287408 211802 287464
rect 211858 287408 211863 287464
rect 199396 287406 211863 287408
rect 199396 287404 199402 287406
rect 211797 287403 211863 287406
rect 185669 287330 185735 287333
rect 203149 287330 203215 287333
rect 185669 287328 203215 287330
rect 185669 287272 185674 287328
rect 185730 287272 203154 287328
rect 203210 287272 203215 287328
rect 185669 287270 203215 287272
rect 185669 287267 185735 287270
rect 203149 287267 203215 287270
rect 217409 287330 217475 287333
rect 221038 287330 221044 287332
rect 217409 287328 221044 287330
rect 217409 287272 217414 287328
rect 217470 287272 221044 287328
rect 217409 287270 221044 287272
rect 217409 287267 217475 287270
rect 221038 287268 221044 287270
rect 221108 287268 221114 287332
rect 223665 287330 223731 287333
rect 231894 287330 231900 287332
rect 223665 287328 231900 287330
rect 223665 287272 223670 287328
rect 223726 287272 231900 287328
rect 223665 287270 231900 287272
rect 223665 287267 223731 287270
rect 231894 287268 231900 287270
rect 231964 287268 231970 287332
rect 235165 287330 235231 287333
rect 260097 287330 260163 287333
rect 235165 287328 260163 287330
rect 235165 287272 235170 287328
rect 235226 287272 260102 287328
rect 260158 287272 260163 287328
rect 235165 287270 260163 287272
rect 235165 287267 235231 287270
rect 260097 287267 260163 287270
rect 220077 287194 220143 287197
rect 228214 287194 228220 287196
rect 220077 287192 228220 287194
rect 220077 287136 220082 287192
rect 220138 287136 228220 287192
rect 220077 287134 228220 287136
rect 220077 287131 220143 287134
rect 228214 287132 228220 287134
rect 228284 287132 228290 287196
rect 236637 287194 236703 287197
rect 238702 287194 238708 287196
rect 236637 287192 238708 287194
rect 236637 287136 236642 287192
rect 236698 287136 238708 287192
rect 236637 287134 238708 287136
rect 236637 287131 236703 287134
rect 238702 287132 238708 287134
rect 238772 287132 238778 287196
rect 240869 287194 240935 287197
rect 280981 287194 281047 287197
rect 240869 287192 281047 287194
rect 240869 287136 240874 287192
rect 240930 287136 280986 287192
rect 281042 287136 281047 287192
rect 240869 287134 281047 287136
rect 240869 287131 240935 287134
rect 280981 287131 281047 287134
rect 66345 286786 66411 286789
rect 66345 286784 68908 286786
rect 66345 286728 66350 286784
rect 66406 286728 68908 286784
rect 66345 286726 68908 286728
rect 66345 286723 66411 286726
rect 158713 286514 158779 286517
rect 156676 286512 158779 286514
rect 156676 286456 158718 286512
rect 158774 286456 158779 286512
rect 156676 286454 158779 286456
rect 158713 286451 158779 286454
rect 206093 286106 206159 286109
rect 244181 286106 244247 286109
rect 200070 286104 206159 286106
rect 200070 286048 206098 286104
rect 206154 286048 206159 286104
rect 200070 286046 206159 286048
rect 178861 285834 178927 285837
rect 200070 285834 200130 286046
rect 206093 286043 206159 286046
rect 238710 286104 244247 286106
rect 238710 286048 244186 286104
rect 244242 286048 244247 286104
rect 238710 286046 244247 286048
rect 205541 285970 205607 285973
rect 178861 285832 200130 285834
rect 178861 285776 178866 285832
rect 178922 285776 200130 285832
rect 178861 285774 200130 285776
rect 200254 285968 205607 285970
rect 200254 285912 205546 285968
rect 205602 285912 205607 285968
rect 200254 285910 205607 285912
rect 178861 285771 178927 285774
rect 53557 285700 53623 285701
rect 53557 285696 53604 285700
rect 53668 285698 53674 285700
rect 66805 285698 66871 285701
rect 162669 285698 162735 285701
rect 200254 285698 200314 285910
rect 205541 285907 205607 285910
rect 222929 285970 222995 285973
rect 234654 285970 234660 285972
rect 222929 285968 234660 285970
rect 222929 285912 222934 285968
rect 222990 285912 234660 285968
rect 222929 285910 234660 285912
rect 222929 285907 222995 285910
rect 234654 285908 234660 285910
rect 234724 285908 234730 285972
rect 238109 285970 238175 285973
rect 238710 285970 238770 286046
rect 244181 286043 244247 286046
rect 238109 285968 238770 285970
rect 238109 285912 238114 285968
rect 238170 285912 238770 285968
rect 238109 285910 238770 285912
rect 242893 285970 242959 285973
rect 244038 285970 244044 285972
rect 242893 285968 244044 285970
rect 242893 285912 242898 285968
rect 242954 285912 244044 285968
rect 242893 285910 244044 285912
rect 238109 285907 238175 285910
rect 242893 285907 242959 285910
rect 244038 285908 244044 285910
rect 244108 285908 244114 285972
rect 200389 285834 200455 285837
rect 202873 285834 202939 285837
rect 200389 285832 202939 285834
rect 200389 285776 200394 285832
rect 200450 285776 202878 285832
rect 202934 285776 202939 285832
rect 200389 285774 202939 285776
rect 200389 285771 200455 285774
rect 202873 285771 202939 285774
rect 214741 285834 214807 285837
rect 215385 285834 215451 285837
rect 214741 285832 215451 285834
rect 214741 285776 214746 285832
rect 214802 285776 215390 285832
rect 215446 285776 215451 285832
rect 214741 285774 215451 285776
rect 214741 285771 214807 285774
rect 215385 285771 215451 285774
rect 220169 285834 220235 285837
rect 220629 285834 220695 285837
rect 226926 285834 226932 285836
rect 220169 285832 226932 285834
rect 220169 285776 220174 285832
rect 220230 285776 220634 285832
rect 220690 285776 226932 285832
rect 220169 285774 226932 285776
rect 220169 285771 220235 285774
rect 220629 285771 220695 285774
rect 226926 285772 226932 285774
rect 226996 285772 227002 285836
rect 249006 285834 249012 285836
rect 238710 285774 249012 285834
rect 53557 285640 53562 285696
rect 53557 285636 53604 285640
rect 53668 285638 53714 285698
rect 66805 285696 68908 285698
rect 66805 285640 66810 285696
rect 66866 285640 68908 285696
rect 66805 285638 68908 285640
rect 162669 285696 200314 285698
rect 162669 285640 162674 285696
rect 162730 285640 200314 285696
rect 162669 285638 200314 285640
rect 53668 285636 53674 285638
rect 53557 285635 53623 285636
rect 66805 285635 66871 285638
rect 162669 285635 162735 285638
rect 200614 285636 200620 285700
rect 200684 285698 200690 285700
rect 200757 285698 200823 285701
rect 200684 285696 200823 285698
rect 200684 285640 200762 285696
rect 200818 285640 200823 285696
rect 200684 285638 200823 285640
rect 200684 285636 200690 285638
rect 200757 285635 200823 285638
rect 204897 285698 204963 285701
rect 207565 285698 207631 285701
rect 204897 285696 207631 285698
rect 204897 285640 204902 285696
rect 204958 285640 207570 285696
rect 207626 285640 207631 285696
rect 204897 285638 207631 285640
rect 204897 285635 204963 285638
rect 207565 285635 207631 285638
rect 209630 285636 209636 285700
rect 209700 285698 209706 285700
rect 214373 285698 214439 285701
rect 209700 285696 214439 285698
rect 209700 285640 214378 285696
rect 214434 285640 214439 285696
rect 209700 285638 214439 285640
rect 209700 285636 209706 285638
rect 214373 285635 214439 285638
rect 215334 285636 215340 285700
rect 215404 285698 215410 285700
rect 215845 285698 215911 285701
rect 215404 285696 215911 285698
rect 215404 285640 215850 285696
rect 215906 285640 215911 285696
rect 215404 285638 215911 285640
rect 215404 285636 215410 285638
rect 215845 285635 215911 285638
rect 225137 285698 225203 285701
rect 226190 285698 226196 285700
rect 225137 285696 226196 285698
rect 225137 285640 225142 285696
rect 225198 285640 226196 285696
rect 225137 285638 226196 285640
rect 225137 285635 225203 285638
rect 226190 285636 226196 285638
rect 226260 285636 226266 285700
rect 233969 285698 234035 285701
rect 236637 285698 236703 285701
rect 238710 285698 238770 285774
rect 249006 285772 249012 285774
rect 249076 285772 249082 285836
rect 233969 285696 238770 285698
rect 233969 285640 233974 285696
rect 234030 285640 236642 285696
rect 236698 285640 238770 285696
rect 233969 285638 238770 285640
rect 239949 285698 240015 285701
rect 268377 285698 268443 285701
rect 269021 285698 269087 285701
rect 239949 285696 269087 285698
rect 239949 285640 239954 285696
rect 240010 285640 268382 285696
rect 268438 285640 269026 285696
rect 269082 285640 269087 285696
rect 239949 285638 269087 285640
rect 233969 285635 234035 285638
rect 236637 285635 236703 285638
rect 239949 285635 240015 285638
rect 268377 285635 268443 285638
rect 269021 285635 269087 285638
rect 158713 285426 158779 285429
rect 156676 285424 158779 285426
rect 156676 285368 158718 285424
rect 158774 285368 158779 285424
rect 156676 285366 158779 285368
rect 158713 285363 158779 285366
rect 583520 285276 584960 285516
rect 158437 284882 158503 284885
rect 200297 284882 200363 284885
rect 158437 284880 200363 284882
rect 158437 284824 158442 284880
rect 158498 284824 200302 284880
rect 200358 284824 200363 284880
rect 158437 284822 200363 284824
rect 158437 284819 158503 284822
rect 200297 284819 200363 284822
rect 66713 284610 66779 284613
rect 198825 284610 198891 284613
rect 218605 284610 218671 284613
rect 66713 284608 68908 284610
rect 66713 284552 66718 284608
rect 66774 284552 68908 284608
rect 66713 284550 68908 284552
rect 198825 284608 218671 284610
rect 198825 284552 198830 284608
rect 198886 284552 218610 284608
rect 218666 284552 218671 284608
rect 198825 284550 218671 284552
rect 66713 284547 66779 284550
rect 198825 284547 198891 284550
rect 218605 284547 218671 284550
rect 242341 284610 242407 284613
rect 280889 284610 280955 284613
rect 242341 284608 280955 284610
rect 242341 284552 242346 284608
rect 242402 284552 280894 284608
rect 280950 284552 280955 284608
rect 242341 284550 280955 284552
rect 242341 284547 242407 284550
rect 280889 284547 280955 284550
rect 198774 284412 198780 284476
rect 198844 284474 198850 284476
rect 204253 284474 204319 284477
rect 198844 284472 204319 284474
rect 198844 284416 204258 284472
rect 204314 284416 204319 284472
rect 198844 284414 204319 284416
rect 198844 284412 198850 284414
rect 204253 284411 204319 284414
rect 212349 284474 212415 284477
rect 381537 284474 381603 284477
rect 212349 284472 381603 284474
rect 212349 284416 212354 284472
rect 212410 284416 381542 284472
rect 381598 284416 381603 284472
rect 212349 284414 381603 284416
rect 212349 284411 212415 284414
rect 381537 284411 381603 284414
rect 158713 284338 158779 284341
rect 156676 284336 158779 284338
rect 156676 284280 158718 284336
rect 158774 284280 158779 284336
rect 156676 284278 158779 284280
rect 158713 284275 158779 284278
rect 195421 284338 195487 284341
rect 203701 284338 203767 284341
rect 195421 284336 203767 284338
rect 195421 284280 195426 284336
rect 195482 284280 203706 284336
rect 203762 284280 203767 284336
rect 195421 284278 203767 284280
rect 195421 284275 195487 284278
rect 203701 284275 203767 284278
rect 208025 284338 208091 284341
rect 214741 284338 214807 284341
rect 583201 284338 583267 284341
rect 208025 284336 208226 284338
rect 208025 284280 208030 284336
rect 208086 284280 208226 284336
rect 208025 284278 208226 284280
rect 208025 284275 208091 284278
rect 208166 284204 208226 284278
rect 214741 284336 583267 284338
rect 214741 284280 214746 284336
rect 214802 284280 583206 284336
rect 583262 284280 583267 284336
rect 214741 284278 583267 284280
rect 214741 284275 214807 284278
rect 583201 284275 583267 284278
rect 208158 284140 208164 284204
rect 208228 284140 208234 284204
rect 191189 284066 191255 284069
rect 201401 284066 201467 284069
rect 191189 284064 201467 284066
rect 191189 284008 191194 284064
rect 191250 284008 201406 284064
rect 201462 284008 201467 284064
rect 191189 284006 201467 284008
rect 191189 284003 191255 284006
rect 201401 284003 201467 284006
rect 216029 284066 216095 284069
rect 216438 284066 216444 284068
rect 216029 284064 216444 284066
rect 216029 284008 216034 284064
rect 216090 284008 216444 284064
rect 216029 284006 216444 284008
rect 216029 284003 216095 284006
rect 216438 284004 216444 284006
rect 216508 284004 216514 284068
rect 201125 283930 201191 283933
rect 201350 283930 201356 283932
rect 201125 283928 201356 283930
rect 201125 283872 201130 283928
rect 201186 283872 201356 283928
rect 201125 283870 201356 283872
rect 201125 283867 201191 283870
rect 201350 283868 201356 283870
rect 201420 283868 201426 283932
rect 215518 283868 215524 283932
rect 215588 283930 215594 283932
rect 215937 283930 216003 283933
rect 215588 283928 216003 283930
rect 215588 283872 215942 283928
rect 215998 283872 216003 283928
rect 215588 283870 216003 283872
rect 215588 283868 215594 283870
rect 215937 283867 216003 283870
rect 219341 283930 219407 283933
rect 224677 283932 224743 283933
rect 220854 283930 220860 283932
rect 219341 283928 220860 283930
rect 219341 283872 219346 283928
rect 219402 283872 220860 283928
rect 219341 283870 220860 283872
rect 219341 283867 219407 283870
rect 220854 283868 220860 283870
rect 220924 283868 220930 283932
rect 224677 283930 224724 283932
rect 224632 283928 224724 283930
rect 224632 283872 224682 283928
rect 224632 283870 224724 283872
rect 224677 283868 224724 283870
rect 224788 283868 224794 283932
rect 227662 283868 227668 283932
rect 227732 283930 227738 283932
rect 227989 283930 228055 283933
rect 228766 283930 228772 283932
rect 227732 283928 228772 283930
rect 227732 283872 227994 283928
rect 228050 283872 228772 283928
rect 227732 283870 228772 283872
rect 227732 283868 227738 283870
rect 224677 283867 224743 283868
rect 227989 283867 228055 283870
rect 228766 283868 228772 283870
rect 228836 283868 228842 283932
rect 229461 283930 229527 283933
rect 231025 283932 231091 283933
rect 229686 283930 229692 283932
rect 229461 283928 229692 283930
rect 229461 283872 229466 283928
rect 229522 283872 229692 283928
rect 229461 283870 229692 283872
rect 229461 283867 229527 283870
rect 229686 283868 229692 283870
rect 229756 283868 229762 283932
rect 230974 283868 230980 283932
rect 231044 283930 231091 283932
rect 231044 283928 231136 283930
rect 231086 283872 231136 283928
rect 231044 283870 231136 283872
rect 231044 283868 231091 283870
rect 236494 283868 236500 283932
rect 236564 283930 236570 283932
rect 236729 283930 236795 283933
rect 236564 283928 236795 283930
rect 236564 283872 236734 283928
rect 236790 283872 236795 283928
rect 236564 283870 236795 283872
rect 236564 283868 236570 283870
rect 231025 283867 231091 283868
rect 236729 283867 236795 283870
rect 237966 283868 237972 283932
rect 238036 283930 238042 283932
rect 238201 283930 238267 283933
rect 238036 283928 238267 283930
rect 238036 283872 238206 283928
rect 238262 283872 238267 283928
rect 238036 283870 238267 283872
rect 238036 283868 238042 283870
rect 238201 283867 238267 283870
rect 245929 283794 245995 283797
rect 244076 283792 245995 283794
rect 66805 283522 66871 283525
rect 66805 283520 68908 283522
rect 66805 283464 66810 283520
rect 66866 283464 68908 283520
rect 66805 283462 68908 283464
rect 66805 283459 66871 283462
rect 158805 283250 158871 283253
rect 156676 283248 158871 283250
rect 156676 283192 158810 283248
rect 158866 283192 158871 283248
rect 156676 283190 158871 283192
rect 158805 283187 158871 283190
rect 173249 283250 173315 283253
rect 200254 283250 200314 283764
rect 244076 283736 245934 283792
rect 245990 283736 245995 283792
rect 244076 283734 245995 283736
rect 245929 283731 245995 283734
rect 244181 283522 244247 283525
rect 266261 283522 266327 283525
rect 244181 283520 266327 283522
rect 244181 283464 244186 283520
rect 244242 283464 266266 283520
rect 266322 283464 266327 283520
rect 244181 283462 266327 283464
rect 244181 283459 244247 283462
rect 266261 283459 266327 283462
rect 246941 283250 247007 283253
rect 173249 283248 200314 283250
rect 173249 283192 173254 283248
rect 173310 283192 200314 283248
rect 173249 283190 200314 283192
rect 244076 283248 247007 283250
rect 244076 283192 246946 283248
rect 247002 283192 247007 283248
rect 244076 283190 247007 283192
rect 173249 283187 173315 283190
rect 246941 283187 247007 283190
rect 197169 282978 197235 282981
rect 197169 282976 200284 282978
rect 197169 282920 197174 282976
rect 197230 282920 200284 282976
rect 197169 282918 200284 282920
rect 197169 282915 197235 282918
rect 67449 282434 67515 282437
rect 197353 282434 197419 282437
rect 245929 282434 245995 282437
rect 67449 282432 68908 282434
rect 67449 282376 67454 282432
rect 67510 282376 68908 282432
rect 67449 282374 68908 282376
rect 197353 282432 200284 282434
rect 197353 282376 197358 282432
rect 197414 282376 200284 282432
rect 197353 282374 200284 282376
rect 244076 282432 245995 282434
rect 244076 282376 245934 282432
rect 245990 282376 245995 282432
rect 244076 282374 245995 282376
rect 67449 282371 67515 282374
rect 197353 282371 197419 282374
rect 245929 282371 245995 282374
rect 159357 282298 159423 282301
rect 176561 282298 176627 282301
rect 185669 282298 185735 282301
rect 159357 282296 161490 282298
rect 159357 282240 159362 282296
rect 159418 282240 161490 282296
rect 159357 282238 161490 282240
rect 159357 282235 159423 282238
rect 158713 282162 158779 282165
rect 156676 282160 158779 282162
rect 156676 282104 158718 282160
rect 158774 282104 158779 282160
rect 156676 282102 158779 282104
rect 161430 282162 161490 282238
rect 176561 282296 185735 282298
rect 176561 282240 176566 282296
rect 176622 282240 185674 282296
rect 185730 282240 185735 282296
rect 176561 282238 185735 282240
rect 176561 282235 176627 282238
rect 185669 282235 185735 282238
rect 193949 282162 194015 282165
rect 161430 282160 194015 282162
rect 161430 282104 193954 282160
rect 194010 282104 194015 282160
rect 161430 282102 194015 282104
rect 158713 282099 158779 282102
rect 193949 282099 194015 282102
rect 197997 281618 198063 281621
rect 245745 281618 245811 281621
rect 197997 281616 200284 281618
rect 197997 281560 198002 281616
rect 198058 281560 200284 281616
rect 197997 281558 200284 281560
rect 244076 281616 245811 281618
rect 244076 281560 245750 281616
rect 245806 281560 245811 281616
rect 244076 281558 245811 281560
rect 197997 281555 198063 281558
rect 245745 281555 245811 281558
rect 65885 281346 65951 281349
rect 65885 281344 68908 281346
rect 65885 281288 65890 281344
rect 65946 281288 68908 281344
rect 65885 281286 68908 281288
rect 65885 281283 65951 281286
rect 158805 281074 158871 281077
rect 245653 281074 245719 281077
rect 156676 281072 158871 281074
rect 156676 281016 158810 281072
rect 158866 281016 158871 281072
rect 156676 281014 158871 281016
rect 244076 281072 245719 281074
rect 244076 281016 245658 281072
rect 245714 281016 245719 281072
rect 244076 281014 245719 281016
rect 158805 281011 158871 281014
rect 245653 281011 245719 281014
rect 197353 280802 197419 280805
rect 197353 280800 200284 280802
rect 197353 280744 197358 280800
rect 197414 280744 200284 280800
rect 197353 280742 200284 280744
rect 197353 280739 197419 280742
rect 198273 280530 198339 280533
rect 198273 280528 200314 280530
rect 198273 280472 198278 280528
rect 198334 280472 200314 280528
rect 198273 280470 200314 280472
rect 198273 280467 198339 280470
rect 67173 280258 67239 280261
rect 67766 280258 67772 280260
rect 67173 280256 67772 280258
rect -960 279972 480 280212
rect 67173 280200 67178 280256
rect 67234 280200 67772 280256
rect 67173 280198 67772 280200
rect 67173 280195 67239 280198
rect 67766 280196 67772 280198
rect 67836 280258 67842 280260
rect 67836 280198 68908 280258
rect 200254 280228 200314 280470
rect 245653 280258 245719 280261
rect 244076 280256 245719 280258
rect 244076 280200 245658 280256
rect 245714 280200 245719 280256
rect 244076 280198 245719 280200
rect 67836 280196 67842 280198
rect 245653 280195 245719 280198
rect 244774 280060 244780 280124
rect 244844 280122 244850 280124
rect 245653 280122 245719 280125
rect 244844 280120 245719 280122
rect 244844 280064 245658 280120
rect 245714 280064 245719 280120
rect 244844 280062 245719 280064
rect 244844 280060 244850 280062
rect 245653 280059 245719 280062
rect 255262 280060 255268 280124
rect 255332 280122 255338 280124
rect 255589 280122 255655 280125
rect 255332 280120 255655 280122
rect 255332 280064 255594 280120
rect 255650 280064 255655 280120
rect 255332 280062 255655 280064
rect 255332 280060 255338 280062
rect 255589 280059 255655 280062
rect 158713 279986 158779 279989
rect 156676 279984 158779 279986
rect 156676 279928 158718 279984
rect 158774 279928 158779 279984
rect 156676 279926 158779 279928
rect 158713 279923 158779 279926
rect 197353 279578 197419 279581
rect 197353 279576 200130 279578
rect 197353 279520 197358 279576
rect 197414 279520 200130 279576
rect 197353 279518 200130 279520
rect 197353 279515 197419 279518
rect 163589 279442 163655 279445
rect 198774 279442 198780 279444
rect 163589 279440 198780 279442
rect 163589 279384 163594 279440
rect 163650 279384 198780 279440
rect 163589 279382 198780 279384
rect 163589 279379 163655 279382
rect 198774 279380 198780 279382
rect 198844 279380 198850 279444
rect 200070 279442 200130 279518
rect 245929 279442 245995 279445
rect 200070 279382 200284 279442
rect 244076 279440 245995 279442
rect 244076 279384 245934 279440
rect 245990 279384 245995 279440
rect 244076 279382 245995 279384
rect 245929 279379 245995 279382
rect 194501 279306 194567 279309
rect 198774 279306 198780 279308
rect 194501 279304 198780 279306
rect 194501 279248 194506 279304
rect 194562 279248 198780 279304
rect 194501 279246 198780 279248
rect 194501 279243 194567 279246
rect 198774 279244 198780 279246
rect 198844 279244 198850 279308
rect 67173 279170 67239 279173
rect 67173 279168 68908 279170
rect 67173 279112 67178 279168
rect 67234 279112 68908 279168
rect 67173 279110 68908 279112
rect 67173 279107 67239 279110
rect 158713 278898 158779 278901
rect 245745 278898 245811 278901
rect 156676 278896 158779 278898
rect 156676 278840 158718 278896
rect 158774 278840 158779 278896
rect 156676 278838 158779 278840
rect 244076 278896 245811 278898
rect 244076 278840 245750 278896
rect 245806 278840 245811 278896
rect 244076 278838 245811 278840
rect 158713 278835 158779 278838
rect 245745 278835 245811 278838
rect 249977 278764 250043 278765
rect 249926 278762 249932 278764
rect 249886 278702 249932 278762
rect 249996 278760 250043 278764
rect 250038 278704 250043 278760
rect 249926 278700 249932 278702
rect 249996 278700 250043 278704
rect 249977 278699 250043 278700
rect 197353 278626 197419 278629
rect 197353 278624 200284 278626
rect 197353 278568 197358 278624
rect 197414 278568 200284 278624
rect 197353 278566 200284 278568
rect 197353 278563 197419 278566
rect 66805 278082 66871 278085
rect 180057 278082 180123 278085
rect 185577 278082 185643 278085
rect 66805 278080 68908 278082
rect 66805 278024 66810 278080
rect 66866 278024 68908 278080
rect 66805 278022 68908 278024
rect 180057 278080 185643 278082
rect 180057 278024 180062 278080
rect 180118 278024 185582 278080
rect 185638 278024 185643 278080
rect 180057 278022 185643 278024
rect 66805 278019 66871 278022
rect 180057 278019 180123 278022
rect 185577 278019 185643 278022
rect 198590 278020 198596 278084
rect 198660 278082 198666 278084
rect 244273 278082 244339 278085
rect 198660 278022 200284 278082
rect 244076 278080 244339 278082
rect 244076 278024 244278 278080
rect 244334 278024 244339 278080
rect 244076 278022 244339 278024
rect 198660 278020 198666 278022
rect 244273 278019 244339 278022
rect 157742 277810 157748 277812
rect 156676 277750 157748 277810
rect 157742 277748 157748 277750
rect 157812 277810 157818 277812
rect 159357 277810 159423 277813
rect 157812 277808 159423 277810
rect 157812 277752 159362 277808
rect 159418 277752 159423 277808
rect 157812 277750 159423 277752
rect 157812 277748 157818 277750
rect 159357 277747 159423 277750
rect 245745 277538 245811 277541
rect 244076 277536 245811 277538
rect 244076 277480 245750 277536
rect 245806 277480 245811 277536
rect 244076 277478 245811 277480
rect 245745 277475 245811 277478
rect 66805 277266 66871 277269
rect 197353 277266 197419 277269
rect 66805 277264 68908 277266
rect 66805 277208 66810 277264
rect 66866 277208 68908 277264
rect 66805 277206 68908 277208
rect 197353 277264 200284 277266
rect 197353 277208 197358 277264
rect 197414 277208 200284 277264
rect 197353 277206 200284 277208
rect 66805 277203 66871 277206
rect 197353 277203 197419 277206
rect 158713 276722 158779 276725
rect 156676 276720 158779 276722
rect 156676 276664 158718 276720
rect 158774 276664 158779 276720
rect 156676 276662 158779 276664
rect 158713 276659 158779 276662
rect 160686 276660 160692 276724
rect 160756 276722 160762 276724
rect 174537 276722 174603 276725
rect 160756 276720 174603 276722
rect 160756 276664 174542 276720
rect 174598 276664 174603 276720
rect 160756 276662 174603 276664
rect 160756 276660 160762 276662
rect 174537 276659 174603 276662
rect 197353 276722 197419 276725
rect 246113 276722 246179 276725
rect 197353 276720 200284 276722
rect 197353 276664 197358 276720
rect 197414 276664 200284 276720
rect 197353 276662 200284 276664
rect 244076 276720 246179 276722
rect 244076 276664 246118 276720
rect 246174 276664 246179 276720
rect 244076 276662 246179 276664
rect 197353 276659 197419 276662
rect 246113 276659 246179 276662
rect 66846 276116 66852 276180
rect 66916 276178 66922 276180
rect 66916 276118 68908 276178
rect 66916 276116 66922 276118
rect 197445 275906 197511 275909
rect 200021 275906 200087 275909
rect 245837 275906 245903 275909
rect 197445 275904 200284 275906
rect 197445 275848 197450 275904
rect 197506 275848 200026 275904
rect 200082 275848 200284 275904
rect 197445 275846 200284 275848
rect 244076 275904 245903 275906
rect 244076 275848 245842 275904
rect 245898 275848 245903 275904
rect 244076 275846 245903 275848
rect 197445 275843 197511 275846
rect 200021 275843 200087 275846
rect 245837 275843 245903 275846
rect 158805 275634 158871 275637
rect 156676 275632 158871 275634
rect 156676 275576 158810 275632
rect 158866 275576 158871 275632
rect 156676 275574 158871 275576
rect 158805 275571 158871 275574
rect 245694 275362 245700 275364
rect 244076 275302 245700 275362
rect 245694 275300 245700 275302
rect 245764 275300 245770 275364
rect 66621 275090 66687 275093
rect 197353 275090 197419 275093
rect 66621 275088 68908 275090
rect 66621 275032 66626 275088
rect 66682 275032 68908 275088
rect 66621 275030 68908 275032
rect 197353 275088 200284 275090
rect 197353 275032 197358 275088
rect 197414 275032 200284 275088
rect 197353 275030 200284 275032
rect 66621 275027 66687 275030
rect 197353 275027 197419 275030
rect 158713 274546 158779 274549
rect 156676 274544 158779 274546
rect 156676 274488 158718 274544
rect 158774 274488 158779 274544
rect 156676 274486 158779 274488
rect 158713 274483 158779 274486
rect 197353 274546 197419 274549
rect 245929 274546 245995 274549
rect 197353 274544 200284 274546
rect 197353 274488 197358 274544
rect 197414 274488 200284 274544
rect 197353 274486 200284 274488
rect 244076 274544 245995 274546
rect 244076 274488 245934 274544
rect 245990 274488 245995 274544
rect 244076 274486 245995 274488
rect 197353 274483 197419 274486
rect 245929 274483 245995 274486
rect 66989 274002 67055 274005
rect 66989 274000 68908 274002
rect 66989 273944 66994 274000
rect 67050 273944 68908 274000
rect 66989 273942 68908 273944
rect 66989 273939 67055 273942
rect 171869 273866 171935 273869
rect 183093 273866 183159 273869
rect 171869 273864 183159 273866
rect 171869 273808 171874 273864
rect 171930 273808 183098 273864
rect 183154 273808 183159 273864
rect 171869 273806 183159 273808
rect 171869 273803 171935 273806
rect 183093 273803 183159 273806
rect 197353 273730 197419 273733
rect 245929 273730 245995 273733
rect 197353 273728 200284 273730
rect 197353 273672 197358 273728
rect 197414 273672 200284 273728
rect 197353 273670 200284 273672
rect 244076 273728 245995 273730
rect 244076 273672 245934 273728
rect 245990 273672 245995 273728
rect 244076 273670 245995 273672
rect 197353 273667 197419 273670
rect 245929 273667 245995 273670
rect 158713 273458 158779 273461
rect 156676 273456 158779 273458
rect 156676 273400 158718 273456
rect 158774 273400 158779 273456
rect 156676 273398 158779 273400
rect 158713 273395 158779 273398
rect 246941 273186 247007 273189
rect 247125 273186 247191 273189
rect 244076 273184 247191 273186
rect 244076 273128 246946 273184
rect 247002 273128 247130 273184
rect 247186 273128 247191 273184
rect 244076 273126 247191 273128
rect 246941 273123 247007 273126
rect 247125 273123 247191 273126
rect 166901 273050 166967 273053
rect 156646 273048 166967 273050
rect 156646 272992 166906 273048
rect 166962 272992 166967 273048
rect 156646 272990 166967 272992
rect 66253 272914 66319 272917
rect 66253 272912 68908 272914
rect 66253 272856 66258 272912
rect 66314 272856 68908 272912
rect 66253 272854 68908 272856
rect 66253 272851 66319 272854
rect 156646 272340 156706 272990
rect 166901 272987 166967 272990
rect 197353 272914 197419 272917
rect 197353 272912 200284 272914
rect 197353 272856 197358 272912
rect 197414 272856 200284 272912
rect 197353 272854 200284 272856
rect 197353 272851 197419 272854
rect 166901 272506 166967 272509
rect 178534 272506 178540 272508
rect 166901 272504 178540 272506
rect 166901 272448 166906 272504
rect 166962 272448 178540 272504
rect 166901 272446 178540 272448
rect 166901 272443 166967 272446
rect 178534 272444 178540 272446
rect 178604 272444 178610 272508
rect 197445 272370 197511 272373
rect 245837 272370 245903 272373
rect 197445 272368 200284 272370
rect 197445 272312 197450 272368
rect 197506 272312 200284 272368
rect 197445 272310 200284 272312
rect 244076 272368 245903 272370
rect 244076 272312 245842 272368
rect 245898 272312 245903 272368
rect 244076 272310 245903 272312
rect 197445 272307 197511 272310
rect 245837 272307 245903 272310
rect 579797 272234 579863 272237
rect 583520 272234 584960 272324
rect 579797 272232 584960 272234
rect 579797 272176 579802 272232
rect 579858 272176 584960 272232
rect 579797 272174 584960 272176
rect 579797 272171 579863 272174
rect 583520 272084 584960 272174
rect 66069 271826 66135 271829
rect 66069 271824 68908 271826
rect 66069 271768 66074 271824
rect 66130 271768 68908 271824
rect 66069 271766 68908 271768
rect 66069 271763 66135 271766
rect 197353 271554 197419 271557
rect 247217 271554 247283 271557
rect 197353 271552 200284 271554
rect 197353 271496 197358 271552
rect 197414 271496 200284 271552
rect 197353 271494 200284 271496
rect 244076 271552 247283 271554
rect 244076 271496 247222 271552
rect 247278 271496 247283 271552
rect 244076 271494 247283 271496
rect 197353 271491 197419 271494
rect 247217 271491 247283 271494
rect 159357 271282 159423 271285
rect 156676 271280 159423 271282
rect 156676 271224 159362 271280
rect 159418 271224 159423 271280
rect 156676 271222 159423 271224
rect 159357 271219 159423 271222
rect 156781 271146 156847 271149
rect 199326 271146 199332 271148
rect 156781 271144 199332 271146
rect 156781 271088 156786 271144
rect 156842 271088 199332 271144
rect 156781 271086 199332 271088
rect 156781 271083 156847 271086
rect 199326 271084 199332 271086
rect 199396 271084 199402 271148
rect 198365 271010 198431 271013
rect 244549 271010 244615 271013
rect 198365 271008 200284 271010
rect 198365 270952 198370 271008
rect 198426 270952 200284 271008
rect 244076 271008 244615 271010
rect 244076 270980 244554 271008
rect 198365 270950 200284 270952
rect 244046 270952 244554 270980
rect 244610 270952 244615 271008
rect 244046 270950 244615 270952
rect 198365 270947 198431 270950
rect 67817 270738 67883 270741
rect 67817 270736 68908 270738
rect 67817 270680 67822 270736
rect 67878 270680 68908 270736
rect 67817 270678 68908 270680
rect 67817 270675 67883 270678
rect 244046 270602 244106 270950
rect 244549 270947 244615 270950
rect 285765 270602 285831 270605
rect 286041 270602 286107 270605
rect 244046 270600 286107 270602
rect 244046 270544 285770 270600
rect 285826 270544 286046 270600
rect 286102 270544 286107 270600
rect 244046 270542 286107 270544
rect 285765 270539 285831 270542
rect 286041 270539 286107 270542
rect 199469 270194 199535 270197
rect 245745 270194 245811 270197
rect 199469 270192 200284 270194
rect 67950 269588 67956 269652
rect 68020 269650 68026 269652
rect 68020 269590 68908 269650
rect 68020 269588 68026 269590
rect 156646 269378 156706 270164
rect 199469 270136 199474 270192
rect 199530 270136 200284 270192
rect 244076 270192 245811 270194
rect 244076 270164 245750 270192
rect 199469 270134 200284 270136
rect 244046 270136 245750 270164
rect 245806 270136 245811 270192
rect 244046 270134 245811 270136
rect 199469 270131 199535 270134
rect 244046 269922 244106 270134
rect 245745 270131 245811 270134
rect 244222 269922 244228 269924
rect 244046 269862 244228 269922
rect 244222 269860 244228 269862
rect 244292 269860 244298 269924
rect 245837 269650 245903 269653
rect 244076 269648 245903 269650
rect 244076 269592 245842 269648
rect 245898 269592 245903 269648
rect 244076 269590 245903 269592
rect 245837 269587 245903 269590
rect 160134 269378 160140 269380
rect 156646 269318 160140 269378
rect 160134 269316 160140 269318
rect 160204 269378 160210 269380
rect 162117 269378 162183 269381
rect 160204 269376 162183 269378
rect 160204 269320 162122 269376
rect 162178 269320 162183 269376
rect 160204 269318 162183 269320
rect 160204 269316 160210 269318
rect 162117 269315 162183 269318
rect 200070 269318 200284 269378
rect 169518 269180 169524 269244
rect 169588 269242 169594 269244
rect 169845 269242 169911 269245
rect 200070 269242 200130 269318
rect 169588 269240 200130 269242
rect 169588 269184 169850 269240
rect 169906 269184 200130 269240
rect 169588 269182 200130 269184
rect 169588 269180 169594 269182
rect 169845 269179 169911 269182
rect 158713 269106 158779 269109
rect 156676 269104 158779 269106
rect 156676 269048 158718 269104
rect 158774 269048 158779 269104
rect 156676 269046 158779 269048
rect 158713 269043 158779 269046
rect 243486 269044 243492 269108
rect 243556 269044 243562 269108
rect 197353 268834 197419 268837
rect 243494 268834 243554 269044
rect 251817 268834 251883 268837
rect 197353 268832 200284 268834
rect 197353 268776 197358 268832
rect 197414 268776 200284 268832
rect 243494 268832 251883 268834
rect 243494 268804 251822 268832
rect 197353 268774 200284 268776
rect 243524 268776 251822 268804
rect 251878 268776 251883 268832
rect 243524 268774 251883 268776
rect 197353 268771 197419 268774
rect 251817 268771 251883 268774
rect 66805 268562 66871 268565
rect 66805 268560 68908 268562
rect 66805 268504 66810 268560
rect 66866 268504 68908 268560
rect 66805 268502 68908 268504
rect 66805 268499 66871 268502
rect 53465 268426 53531 268429
rect 66846 268426 66852 268428
rect 53465 268424 66852 268426
rect 53465 268368 53470 268424
rect 53526 268368 66852 268424
rect 53465 268366 66852 268368
rect 53465 268363 53531 268366
rect 66846 268364 66852 268366
rect 66916 268364 66922 268428
rect 168649 268426 168715 268429
rect 175273 268426 175339 268429
rect 168649 268424 175339 268426
rect 168649 268368 168654 268424
rect 168710 268368 175278 268424
rect 175334 268368 175339 268424
rect 168649 268366 175339 268368
rect 168649 268363 168715 268366
rect 175273 268363 175339 268366
rect 258717 268426 258783 268429
rect 281758 268426 281764 268428
rect 258717 268424 281764 268426
rect 258717 268368 258722 268424
rect 258778 268368 281764 268424
rect 258717 268366 281764 268368
rect 258717 268363 258783 268366
rect 281758 268364 281764 268366
rect 281828 268364 281834 268428
rect 158713 268018 158779 268021
rect 156676 268016 158779 268018
rect 156676 267960 158718 268016
rect 158774 267960 158779 268016
rect 156676 267958 158779 267960
rect 158713 267955 158779 267958
rect 197445 268018 197511 268021
rect 246205 268018 246271 268021
rect 197445 268016 200284 268018
rect 197445 267960 197450 268016
rect 197506 267960 200284 268016
rect 197445 267958 200284 267960
rect 244076 268016 246271 268018
rect 244076 267960 246210 268016
rect 246266 267960 246271 268016
rect 244076 267958 246271 267960
rect 197445 267955 197511 267958
rect 246205 267955 246271 267958
rect 170489 267612 170555 267613
rect 170438 267548 170444 267612
rect 170508 267610 170555 267612
rect 170508 267608 170600 267610
rect 170550 267552 170600 267608
rect 170508 267550 170600 267552
rect 170508 267548 170555 267550
rect 170489 267547 170555 267548
rect 67398 267412 67404 267476
rect 67468 267474 67474 267476
rect 245929 267474 245995 267477
rect 67468 267414 68908 267474
rect 244076 267472 245995 267474
rect 244076 267416 245934 267472
rect 245990 267416 245995 267472
rect 244076 267414 245995 267416
rect 67468 267412 67474 267414
rect 245929 267411 245995 267414
rect 195329 267338 195395 267341
rect 195830 267338 195836 267340
rect 195329 267336 195836 267338
rect -960 267202 480 267292
rect 195329 267280 195334 267336
rect 195390 267280 195836 267336
rect 195329 267278 195836 267280
rect 195329 267275 195395 267278
rect 195830 267276 195836 267278
rect 195900 267338 195906 267340
rect 195900 267278 200130 267338
rect 195900 267276 195906 267278
rect 3325 267202 3391 267205
rect -960 267200 3391 267202
rect -960 267144 3330 267200
rect 3386 267144 3391 267200
rect -960 267142 3391 267144
rect 200070 267202 200130 267278
rect 200070 267142 200284 267202
rect -960 267052 480 267142
rect 3325 267139 3391 267142
rect 67541 266386 67607 266389
rect 156646 266386 156706 266900
rect 197353 266658 197419 266661
rect 197353 266656 200284 266658
rect 197353 266600 197358 266656
rect 197414 266600 200284 266656
rect 197353 266598 200284 266600
rect 244076 266598 248430 266658
rect 197353 266595 197419 266598
rect 170438 266522 170444 266524
rect 161430 266462 170444 266522
rect 161430 266386 161490 266462
rect 170438 266460 170444 266462
rect 170508 266460 170514 266524
rect 248370 266522 248430 266598
rect 258257 266522 258323 266525
rect 259361 266522 259427 266525
rect 248370 266520 259427 266522
rect 248370 266464 258262 266520
rect 258318 266464 259366 266520
rect 259422 266464 259427 266520
rect 248370 266462 259427 266464
rect 258257 266459 258323 266462
rect 259361 266459 259427 266462
rect 67541 266384 68908 266386
rect 67541 266328 67546 266384
rect 67602 266328 68908 266384
rect 67541 266326 68908 266328
rect 156646 266326 161490 266386
rect 164141 266386 164207 266389
rect 169702 266386 169708 266388
rect 164141 266384 169708 266386
rect 164141 266328 164146 266384
rect 164202 266328 169708 266384
rect 164141 266326 169708 266328
rect 67541 266323 67607 266326
rect 164141 266323 164207 266326
rect 169702 266324 169708 266326
rect 169772 266324 169778 266388
rect 245929 266386 245995 266389
rect 270033 266386 270099 266389
rect 270401 266386 270467 266389
rect 245929 266384 270467 266386
rect 245929 266328 245934 266384
rect 245990 266328 270038 266384
rect 270094 266328 270406 266384
rect 270462 266328 270467 266384
rect 245929 266326 270467 266328
rect 245929 266323 245995 266326
rect 270033 266323 270099 266326
rect 270401 266323 270467 266326
rect 246205 266250 246271 266253
rect 267825 266250 267891 266253
rect 269021 266250 269087 266253
rect 246205 266248 269087 266250
rect 246205 266192 246210 266248
rect 246266 266192 267830 266248
rect 267886 266192 269026 266248
rect 269082 266192 269087 266248
rect 246205 266190 269087 266192
rect 246205 266187 246271 266190
rect 267825 266187 267891 266190
rect 269021 266187 269087 266190
rect 159449 265842 159515 265845
rect 156676 265840 159515 265842
rect 156676 265784 159454 265840
rect 159510 265784 159515 265840
rect 156676 265782 159515 265784
rect 159449 265779 159515 265782
rect 199377 265842 199443 265845
rect 245929 265842 245995 265845
rect 199377 265840 200284 265842
rect 199377 265784 199382 265840
rect 199438 265784 200284 265840
rect 199377 265782 200284 265784
rect 244076 265840 245995 265842
rect 244076 265784 245934 265840
rect 245990 265784 245995 265840
rect 244076 265782 245995 265784
rect 199377 265779 199443 265782
rect 245929 265779 245995 265782
rect 168966 265508 168972 265572
rect 169036 265570 169042 265572
rect 198774 265570 198780 265572
rect 169036 265510 198780 265570
rect 169036 265508 169042 265510
rect 198774 265508 198780 265510
rect 198844 265508 198850 265572
rect 269021 265570 269087 265573
rect 583477 265570 583543 265573
rect 269021 265568 583543 265570
rect 269021 265512 269026 265568
rect 269082 265512 583482 265568
rect 583538 265512 583543 265568
rect 269021 265510 583543 265512
rect 269021 265507 269087 265510
rect 583477 265507 583543 265510
rect 66805 265298 66871 265301
rect 197445 265298 197511 265301
rect 246757 265298 246823 265301
rect 66805 265296 68908 265298
rect 66805 265240 66810 265296
rect 66866 265240 68908 265296
rect 66805 265238 68908 265240
rect 197445 265296 200284 265298
rect 197445 265240 197450 265296
rect 197506 265240 200284 265296
rect 197445 265238 200284 265240
rect 244076 265296 246823 265298
rect 244076 265240 246762 265296
rect 246818 265240 246823 265296
rect 244076 265238 246823 265240
rect 66805 265235 66871 265238
rect 197445 265235 197511 265238
rect 246757 265235 246823 265238
rect 157977 264754 158043 264757
rect 156676 264752 158043 264754
rect 156676 264696 157982 264752
rect 158038 264696 158043 264752
rect 156676 264694 158043 264696
rect 157977 264691 158043 264694
rect 197353 264482 197419 264485
rect 247125 264482 247191 264485
rect 197353 264480 200284 264482
rect 197353 264424 197358 264480
rect 197414 264424 200284 264480
rect 197353 264422 200284 264424
rect 244076 264480 247191 264482
rect 244076 264424 247130 264480
rect 247186 264424 247191 264480
rect 244076 264422 247191 264424
rect 197353 264419 197419 264422
rect 247125 264419 247191 264422
rect 66805 264210 66871 264213
rect 259361 264210 259427 264213
rect 583017 264210 583083 264213
rect 66805 264208 68908 264210
rect 66805 264152 66810 264208
rect 66866 264152 68908 264208
rect 66805 264150 68908 264152
rect 259361 264208 583083 264210
rect 259361 264152 259366 264208
rect 259422 264152 583022 264208
rect 583078 264152 583083 264208
rect 259361 264150 583083 264152
rect 66805 264147 66871 264150
rect 259361 264147 259427 264150
rect 583017 264147 583083 264150
rect 245837 263938 245903 263941
rect 244076 263936 245903 263938
rect 244076 263880 245842 263936
rect 245898 263880 245903 263936
rect 244076 263878 245903 263880
rect 245837 263875 245903 263878
rect 158713 263666 158779 263669
rect 156676 263664 158779 263666
rect 156676 263608 158718 263664
rect 158774 263608 158779 263664
rect 156676 263606 158779 263608
rect 158713 263603 158779 263606
rect 197353 263666 197419 263669
rect 197353 263664 200284 263666
rect 197353 263608 197358 263664
rect 197414 263608 200284 263664
rect 197353 263606 200284 263608
rect 197353 263603 197419 263606
rect 66805 263122 66871 263125
rect 198641 263122 198707 263125
rect 199326 263122 199332 263124
rect 66805 263120 68908 263122
rect 66805 263064 66810 263120
rect 66866 263064 68908 263120
rect 66805 263062 68908 263064
rect 198641 263120 199332 263122
rect 198641 263064 198646 263120
rect 198702 263064 199332 263120
rect 198641 263062 199332 263064
rect 66805 263059 66871 263062
rect 198641 263059 198707 263062
rect 199326 263060 199332 263062
rect 199396 263122 199402 263124
rect 245745 263122 245811 263125
rect 199396 263062 200284 263122
rect 244076 263120 245811 263122
rect 244076 263064 245750 263120
rect 245806 263064 245811 263120
rect 244076 263062 245811 263064
rect 199396 263060 199402 263062
rect 245745 263059 245811 263062
rect 160829 262578 160895 262581
rect 156676 262576 160895 262578
rect 156676 262520 160834 262576
rect 160890 262520 160895 262576
rect 156676 262518 160895 262520
rect 160829 262515 160895 262518
rect 198549 262306 198615 262309
rect 245929 262306 245995 262309
rect 198549 262304 200284 262306
rect 198549 262248 198554 262304
rect 198610 262248 200284 262304
rect 198549 262246 200284 262248
rect 244076 262304 245995 262306
rect 244076 262248 245934 262304
rect 245990 262248 245995 262304
rect 244076 262246 245995 262248
rect 198549 262243 198615 262246
rect 245929 262243 245995 262246
rect 66437 262034 66503 262037
rect 66437 262032 68908 262034
rect 66437 261976 66442 262032
rect 66498 261976 68908 262032
rect 66437 261974 68908 261976
rect 66437 261971 66503 261974
rect 158437 261490 158503 261493
rect 159357 261490 159423 261493
rect 156676 261488 159423 261490
rect 156676 261432 158442 261488
rect 158498 261432 159362 261488
rect 159418 261432 159423 261488
rect 156676 261430 159423 261432
rect 158437 261427 158503 261430
rect 159357 261427 159423 261430
rect 164049 261490 164115 261493
rect 197353 261490 197419 261493
rect 164049 261488 180810 261490
rect 164049 261432 164054 261488
rect 164110 261432 180810 261488
rect 164049 261430 180810 261432
rect 164049 261427 164115 261430
rect 66069 260946 66135 260949
rect 180750 260946 180810 261430
rect 197353 261488 200284 261490
rect 197353 261432 197358 261488
rect 197414 261432 200284 261488
rect 197353 261430 200284 261432
rect 197353 261427 197419 261430
rect 244046 261218 244106 261732
rect 249006 261428 249012 261492
rect 249076 261490 249082 261492
rect 580257 261490 580323 261493
rect 249076 261488 580323 261490
rect 249076 261432 580262 261488
rect 580318 261432 580323 261488
rect 249076 261430 580323 261432
rect 249076 261428 249082 261430
rect 580257 261427 580323 261430
rect 254025 261218 254091 261221
rect 244046 261216 254091 261218
rect 244046 261160 254030 261216
rect 254086 261160 254091 261216
rect 244046 261158 254091 261160
rect 254025 261155 254091 261158
rect 183553 260946 183619 260949
rect 246389 260946 246455 260949
rect 66069 260944 68908 260946
rect 66069 260888 66074 260944
rect 66130 260888 68908 260944
rect 66069 260886 68908 260888
rect 180750 260944 200284 260946
rect 180750 260888 183558 260944
rect 183614 260888 200284 260944
rect 180750 260886 200284 260888
rect 244076 260944 246455 260946
rect 244076 260888 246394 260944
rect 246450 260888 246455 260944
rect 244076 260886 246455 260888
rect 66069 260883 66135 260886
rect 183553 260883 183619 260886
rect 246389 260883 246455 260886
rect 66805 259858 66871 259861
rect 66805 259856 68908 259858
rect 66805 259800 66810 259856
rect 66866 259800 68908 259856
rect 66805 259798 68908 259800
rect 66805 259795 66871 259798
rect 156646 259586 156706 260372
rect 162158 260068 162164 260132
rect 162228 260130 162234 260132
rect 189073 260130 189139 260133
rect 162228 260128 189139 260130
rect 162228 260072 189078 260128
rect 189134 260072 189139 260128
rect 162228 260070 189139 260072
rect 162228 260068 162234 260070
rect 189073 260067 189139 260070
rect 197353 260130 197419 260133
rect 245837 260130 245903 260133
rect 197353 260128 200284 260130
rect 197353 260072 197358 260128
rect 197414 260072 200284 260128
rect 197353 260070 200284 260072
rect 244076 260128 245903 260130
rect 244076 260072 245842 260128
rect 245898 260072 245903 260128
rect 244076 260070 245903 260072
rect 197353 260067 197419 260070
rect 245837 260067 245903 260070
rect 159909 259586 159975 259589
rect 161974 259586 161980 259588
rect 156646 259584 161980 259586
rect 156646 259528 159914 259584
rect 159970 259528 161980 259584
rect 156646 259526 161980 259528
rect 159909 259523 159975 259526
rect 161974 259524 161980 259526
rect 162044 259524 162050 259588
rect 244406 259586 244412 259588
rect 244076 259526 244412 259586
rect 244406 259524 244412 259526
rect 244476 259586 244482 259588
rect 245929 259586 245995 259589
rect 244476 259584 245995 259586
rect 244476 259528 245934 259584
rect 245990 259528 245995 259584
rect 244476 259526 245995 259528
rect 244476 259524 244482 259526
rect 245929 259523 245995 259526
rect 195278 259450 195284 259452
rect 156646 259390 195284 259450
rect 156646 259284 156706 259390
rect 195278 259388 195284 259390
rect 195348 259388 195354 259452
rect 197353 259314 197419 259317
rect 197353 259312 200284 259314
rect 197353 259256 197358 259312
rect 197414 259256 200284 259312
rect 197353 259254 200284 259256
rect 197353 259251 197419 259254
rect 580165 258906 580231 258909
rect 583520 258906 584960 258996
rect 580165 258904 584960 258906
rect 580165 258848 580170 258904
rect 580226 258848 584960 258904
rect 580165 258846 584960 258848
rect 580165 258843 580231 258846
rect 197445 258770 197511 258773
rect 245929 258770 245995 258773
rect 197445 258768 200284 258770
rect 46841 257954 46907 257957
rect 65374 257954 65380 257956
rect 46841 257952 65380 257954
rect 46841 257896 46846 257952
rect 46902 257896 65380 257952
rect 46841 257894 65380 257896
rect 46841 257891 46907 257894
rect 65374 257892 65380 257894
rect 65444 257954 65450 257956
rect 68878 257954 68938 258740
rect 197445 258712 197450 258768
rect 197506 258712 200284 258768
rect 197445 258710 200284 258712
rect 244076 258768 245995 258770
rect 244076 258712 245934 258768
rect 245990 258712 245995 258768
rect 583520 258756 584960 258846
rect 244076 258710 245995 258712
rect 197445 258707 197511 258710
rect 245929 258707 245995 258710
rect 158713 258226 158779 258229
rect 245837 258226 245903 258229
rect 156676 258224 158779 258226
rect 156676 258168 158718 258224
rect 158774 258168 158779 258224
rect 156676 258166 158779 258168
rect 244076 258224 245903 258226
rect 244076 258168 245842 258224
rect 245898 258168 245903 258224
rect 244076 258166 245903 258168
rect 158713 258163 158779 258166
rect 245837 258163 245903 258166
rect 180241 257954 180307 257957
rect 65444 257894 68938 257954
rect 156830 257952 180307 257954
rect 156830 257896 180246 257952
rect 180302 257896 180307 257952
rect 156830 257894 180307 257896
rect 65444 257892 65450 257894
rect 156830 257818 156890 257894
rect 180241 257891 180307 257894
rect 197445 257954 197511 257957
rect 197445 257952 200284 257954
rect 197445 257896 197450 257952
rect 197506 257896 200284 257952
rect 197445 257894 200284 257896
rect 197445 257891 197511 257894
rect 156646 257758 156890 257818
rect 69430 257140 69490 257652
rect 69422 257076 69428 257140
rect 69492 257076 69498 257140
rect 156646 257108 156706 257758
rect 198089 257410 198155 257413
rect 246021 257410 246087 257413
rect 198089 257408 200284 257410
rect 198089 257352 198094 257408
rect 198150 257352 200284 257408
rect 198089 257350 200284 257352
rect 244076 257408 246087 257410
rect 244076 257352 246026 257408
rect 246082 257352 246087 257408
rect 244076 257350 246087 257352
rect 198089 257347 198155 257350
rect 246021 257347 246087 257350
rect 66805 256594 66871 256597
rect 197445 256594 197511 256597
rect 245929 256594 245995 256597
rect 66805 256592 68908 256594
rect 66805 256536 66810 256592
rect 66866 256536 68908 256592
rect 66805 256534 68908 256536
rect 197445 256592 200284 256594
rect 197445 256536 197450 256592
rect 197506 256536 200284 256592
rect 197445 256534 200284 256536
rect 244076 256592 245995 256594
rect 244076 256536 245934 256592
rect 245990 256536 245995 256592
rect 244076 256534 245995 256536
rect 66805 256531 66871 256534
rect 197445 256531 197511 256534
rect 245929 256531 245995 256534
rect 158805 256322 158871 256325
rect 156676 256320 158871 256322
rect 156676 256264 158810 256320
rect 158866 256264 158871 256320
rect 156676 256262 158871 256264
rect 158805 256259 158871 256262
rect 247718 256050 247724 256052
rect 244076 255990 247724 256050
rect 247718 255988 247724 255990
rect 247788 255988 247794 256052
rect 197353 255778 197419 255781
rect 197353 255776 200284 255778
rect 197353 255720 197358 255776
rect 197414 255720 200284 255776
rect 197353 255718 200284 255720
rect 197353 255715 197419 255718
rect 67265 255506 67331 255509
rect 67265 255504 68908 255506
rect 67265 255448 67270 255504
rect 67326 255448 68908 255504
rect 67265 255446 68908 255448
rect 67265 255443 67331 255446
rect 158713 255234 158779 255237
rect 156676 255232 158779 255234
rect 156676 255176 158718 255232
rect 158774 255176 158779 255232
rect 156676 255174 158779 255176
rect 158713 255171 158779 255174
rect 197353 255234 197419 255237
rect 244365 255234 244431 255237
rect 197353 255232 200284 255234
rect 197353 255176 197358 255232
rect 197414 255176 200284 255232
rect 197353 255174 200284 255176
rect 244076 255232 244431 255234
rect 244076 255176 244370 255232
rect 244426 255176 244431 255232
rect 244076 255174 244431 255176
rect 197353 255171 197419 255174
rect 244365 255171 244431 255174
rect 67950 254356 67956 254420
rect 68020 254418 68026 254420
rect 68020 254358 68908 254418
rect 68020 254356 68026 254358
rect 195094 254356 195100 254420
rect 195164 254418 195170 254420
rect 245929 254418 245995 254421
rect 195164 254358 200284 254418
rect 244076 254416 245995 254418
rect 244076 254360 245934 254416
rect 245990 254360 245995 254416
rect 244076 254358 245995 254360
rect 195164 254356 195170 254358
rect 245929 254355 245995 254358
rect -960 254146 480 254236
rect 3141 254146 3207 254149
rect 160001 254146 160067 254149
rect -960 254144 3207 254146
rect -960 254088 3146 254144
rect 3202 254088 3207 254144
rect -960 254086 3207 254088
rect 156676 254144 160067 254146
rect 156676 254088 160006 254144
rect 160062 254088 160067 254144
rect 156676 254086 160067 254088
rect -960 253996 480 254086
rect 3141 254083 3207 254086
rect 160001 254083 160067 254086
rect 244457 253874 244523 253877
rect 245469 253874 245535 253877
rect 244076 253872 245535 253874
rect 244076 253816 244462 253872
rect 244518 253816 245474 253872
rect 245530 253816 245535 253872
rect 244076 253814 245535 253816
rect 244457 253811 244523 253814
rect 245469 253811 245535 253814
rect 197353 253602 197419 253605
rect 197353 253600 200284 253602
rect 197353 253544 197358 253600
rect 197414 253544 200284 253600
rect 197353 253542 200284 253544
rect 197353 253539 197419 253542
rect 66989 253330 67055 253333
rect 66989 253328 68908 253330
rect 66989 253272 66994 253328
rect 67050 253272 68908 253328
rect 66989 253270 68908 253272
rect 66989 253267 67055 253270
rect 158713 253058 158779 253061
rect 156676 253056 158779 253058
rect 156676 253000 158718 253056
rect 158774 253000 158779 253056
rect 156676 252998 158779 253000
rect 158713 252995 158779 252998
rect 196617 253058 196683 253061
rect 244641 253058 244707 253061
rect 245469 253058 245535 253061
rect 196617 253056 200284 253058
rect 196617 253000 196622 253056
rect 196678 253000 200284 253056
rect 196617 252998 200284 253000
rect 244076 253056 245535 253058
rect 244076 253000 244646 253056
rect 244702 253000 245474 253056
rect 245530 253000 245535 253056
rect 244076 252998 245535 253000
rect 196617 252995 196683 252998
rect 244641 252995 244707 252998
rect 245469 252995 245535 252998
rect 176469 252650 176535 252653
rect 176469 252648 197370 252650
rect 176469 252592 176474 252648
rect 176530 252592 197370 252648
rect 176469 252590 197370 252592
rect 176469 252587 176535 252590
rect 190177 252514 190243 252517
rect 191189 252514 191255 252517
rect 190177 252512 191255 252514
rect 190177 252456 190182 252512
rect 190238 252456 191194 252512
rect 191250 252456 191255 252512
rect 190177 252454 191255 252456
rect 197310 252514 197370 252590
rect 197854 252588 197860 252652
rect 197924 252588 197930 252652
rect 197862 252514 197922 252588
rect 197310 252454 200314 252514
rect 190177 252451 190243 252454
rect 191189 252451 191255 252454
rect 66662 252180 66668 252244
rect 66732 252242 66738 252244
rect 66732 252182 68908 252242
rect 200254 252212 200314 252454
rect 248454 252242 248460 252244
rect 244076 252182 248460 252242
rect 66732 252180 66738 252182
rect 248454 252180 248460 252182
rect 248524 252180 248530 252244
rect 156646 251290 156706 251940
rect 162393 251834 162459 251837
rect 187601 251834 187667 251837
rect 197997 251834 198063 251837
rect 162393 251832 198063 251834
rect 162393 251776 162398 251832
rect 162454 251776 187606 251832
rect 187662 251776 198002 251832
rect 198058 251776 198063 251832
rect 162393 251774 198063 251776
rect 162393 251771 162459 251774
rect 187601 251771 187667 251774
rect 197997 251771 198063 251774
rect 197353 251698 197419 251701
rect 245929 251698 245995 251701
rect 197353 251696 200284 251698
rect 197353 251640 197358 251696
rect 197414 251640 200284 251696
rect 197353 251638 200284 251640
rect 244076 251696 245995 251698
rect 244076 251640 245934 251696
rect 245990 251640 245995 251696
rect 244076 251638 245995 251640
rect 197353 251635 197419 251638
rect 245929 251635 245995 251638
rect 168414 251290 168420 251292
rect 156646 251230 168420 251290
rect 168414 251228 168420 251230
rect 168484 251228 168490 251292
rect 66897 251154 66963 251157
rect 66897 251152 68908 251154
rect 66897 251096 66902 251152
rect 66958 251096 68908 251152
rect 66897 251094 68908 251096
rect 66897 251091 66963 251094
rect 160134 251092 160140 251156
rect 160204 251154 160210 251156
rect 161197 251154 161263 251157
rect 160204 251152 161263 251154
rect 160204 251096 161202 251152
rect 161258 251096 161263 251152
rect 160204 251094 161263 251096
rect 160204 251092 160210 251094
rect 161197 251091 161263 251094
rect 164969 251154 165035 251157
rect 192569 251154 192635 251157
rect 193029 251154 193095 251157
rect 164969 251152 193095 251154
rect 164969 251096 164974 251152
rect 165030 251096 192574 251152
rect 192630 251096 193034 251152
rect 193090 251096 193095 251152
rect 164969 251094 193095 251096
rect 164969 251091 165035 251094
rect 192569 251091 192635 251094
rect 193029 251091 193095 251094
rect 197905 250882 197971 250885
rect 244273 250882 244339 250885
rect 197905 250880 200284 250882
rect 156646 250202 156706 250852
rect 197905 250824 197910 250880
rect 197966 250824 200284 250880
rect 197905 250822 200284 250824
rect 244076 250880 244339 250882
rect 244076 250824 244278 250880
rect 244334 250824 244339 250880
rect 244076 250822 244339 250824
rect 197905 250819 197971 250822
rect 244273 250819 244339 250822
rect 180241 250474 180307 250477
rect 184381 250474 184447 250477
rect 180241 250472 184447 250474
rect 180241 250416 180246 250472
rect 180302 250416 184386 250472
rect 184442 250416 184447 250472
rect 180241 250414 184447 250416
rect 180241 250411 180307 250414
rect 184381 250411 184447 250414
rect 245745 250338 245811 250341
rect 244076 250336 245811 250338
rect 244076 250280 245750 250336
rect 245806 250280 245811 250336
rect 244076 250278 245811 250280
rect 245745 250275 245811 250278
rect 156646 250142 161490 250202
rect 66805 250066 66871 250069
rect 161430 250066 161490 250142
rect 174721 250066 174787 250069
rect 66805 250064 68908 250066
rect 66805 250008 66810 250064
rect 66866 250008 68908 250064
rect 66805 250006 68908 250008
rect 161430 250064 174787 250066
rect 161430 250008 174726 250064
rect 174782 250008 174787 250064
rect 161430 250006 174787 250008
rect 66805 250003 66871 250006
rect 174721 250003 174787 250006
rect 197353 250066 197419 250069
rect 197353 250064 200284 250066
rect 197353 250008 197358 250064
rect 197414 250008 200284 250064
rect 197353 250006 200284 250008
rect 197353 250003 197419 250006
rect 248454 249868 248460 249932
rect 248524 249930 248530 249932
rect 248597 249930 248663 249933
rect 248524 249928 248663 249930
rect 248524 249872 248602 249928
rect 248658 249872 248663 249928
rect 248524 249870 248663 249872
rect 248524 249868 248530 249870
rect 248597 249867 248663 249870
rect 158805 249794 158871 249797
rect 156676 249792 158871 249794
rect 156676 249736 158810 249792
rect 158866 249736 158871 249792
rect 156676 249734 158871 249736
rect 158805 249731 158871 249734
rect 173157 249794 173223 249797
rect 177297 249794 177363 249797
rect 173157 249792 177363 249794
rect 173157 249736 173162 249792
rect 173218 249736 177302 249792
rect 177358 249736 177363 249792
rect 173157 249734 177363 249736
rect 173157 249731 173223 249734
rect 177297 249731 177363 249734
rect 197353 249522 197419 249525
rect 245929 249522 245995 249525
rect 197353 249520 200284 249522
rect 197353 249464 197358 249520
rect 197414 249464 200284 249520
rect 197353 249462 200284 249464
rect 244076 249520 245995 249522
rect 244076 249464 245934 249520
rect 245990 249464 245995 249520
rect 244076 249462 245995 249464
rect 197353 249459 197419 249462
rect 245929 249459 245995 249462
rect 67766 248916 67772 248980
rect 67836 248978 67842 248980
rect 67836 248918 68908 248978
rect 67836 248916 67842 248918
rect 158713 248706 158779 248709
rect 156676 248704 158779 248706
rect 156676 248648 158718 248704
rect 158774 248648 158779 248704
rect 156676 248646 158779 248648
rect 158713 248643 158779 248646
rect 197445 248706 197511 248709
rect 245929 248706 245995 248709
rect 197445 248704 200284 248706
rect 197445 248648 197450 248704
rect 197506 248648 200284 248704
rect 197445 248646 200284 248648
rect 244076 248704 245995 248706
rect 244076 248648 245934 248704
rect 245990 248648 245995 248704
rect 244076 248646 245995 248648
rect 197445 248643 197511 248646
rect 245929 248643 245995 248646
rect 246941 248162 247007 248165
rect 244076 248160 247007 248162
rect 244076 248104 246946 248160
rect 247002 248104 247007 248160
rect 244076 248102 247007 248104
rect 246941 248099 247007 248102
rect 66897 247890 66963 247893
rect 197445 247890 197511 247893
rect 66897 247888 68908 247890
rect 66897 247832 66902 247888
rect 66958 247832 68908 247888
rect 66897 247830 68908 247832
rect 197445 247888 200284 247890
rect 197445 247832 197450 247888
rect 197506 247832 200284 247888
rect 197445 247830 200284 247832
rect 66897 247827 66963 247830
rect 197445 247827 197511 247830
rect 159398 247618 159404 247620
rect 156676 247558 159404 247618
rect 159398 247556 159404 247558
rect 159468 247556 159474 247620
rect 160870 247556 160876 247620
rect 160940 247618 160946 247620
rect 167821 247618 167887 247621
rect 160940 247616 167887 247618
rect 160940 247560 167826 247616
rect 167882 247560 167887 247616
rect 160940 247558 167887 247560
rect 160940 247556 160946 247558
rect 167821 247555 167887 247558
rect 174629 247346 174695 247349
rect 244457 247346 244523 247349
rect 174629 247344 200284 247346
rect 174629 247288 174634 247344
rect 174690 247288 200284 247344
rect 174629 247286 200284 247288
rect 244076 247344 244523 247346
rect 244076 247288 244462 247344
rect 244518 247288 244523 247344
rect 244076 247286 244523 247288
rect 174629 247283 174695 247286
rect 244457 247283 244523 247286
rect 160737 247210 160803 247213
rect 161381 247210 161447 247213
rect 181713 247210 181779 247213
rect 160737 247208 181779 247210
rect 160737 247152 160742 247208
rect 160798 247152 161386 247208
rect 161442 247152 181718 247208
rect 181774 247152 181779 247208
rect 160737 247150 181779 247152
rect 160737 247147 160803 247150
rect 161381 247147 161447 247150
rect 181713 247147 181779 247150
rect 66805 246802 66871 246805
rect 66805 246800 68908 246802
rect 66805 246744 66810 246800
rect 66866 246744 68908 246800
rect 66805 246742 68908 246744
rect 66805 246739 66871 246742
rect 245653 246530 245719 246533
rect 244076 246528 245719 246530
rect 156646 246258 156706 246500
rect 173157 246258 173223 246261
rect 199837 246258 199903 246261
rect 200254 246258 200314 246500
rect 244076 246472 245658 246528
rect 245714 246472 245719 246528
rect 244076 246470 245719 246472
rect 245653 246467 245719 246470
rect 156646 246256 173223 246258
rect 156646 246200 173162 246256
rect 173218 246200 173223 246256
rect 156646 246198 173223 246200
rect 173157 246195 173223 246198
rect 190410 246256 200314 246258
rect 190410 246200 199842 246256
rect 199898 246200 200314 246256
rect 190410 246198 200314 246200
rect 158110 245788 158116 245852
rect 158180 245850 158186 245852
rect 158621 245850 158687 245853
rect 182265 245850 182331 245853
rect 158180 245848 182331 245850
rect 158180 245792 158626 245848
rect 158682 245792 182270 245848
rect 182326 245792 182331 245848
rect 158180 245790 182331 245792
rect 158180 245788 158186 245790
rect 158621 245787 158687 245790
rect 182265 245787 182331 245790
rect 186221 245850 186287 245853
rect 186814 245850 186820 245852
rect 186221 245848 186820 245850
rect 186221 245792 186226 245848
rect 186282 245792 186820 245848
rect 186221 245790 186820 245792
rect 186221 245787 186287 245790
rect 186814 245788 186820 245790
rect 186884 245788 186890 245852
rect 67725 245714 67791 245717
rect 166441 245714 166507 245717
rect 190410 245714 190470 246198
rect 199837 246195 199903 246198
rect 197353 245986 197419 245989
rect 245745 245986 245811 245989
rect 197353 245984 200284 245986
rect 197353 245928 197358 245984
rect 197414 245928 200284 245984
rect 197353 245926 200284 245928
rect 244076 245984 245811 245986
rect 244076 245928 245750 245984
rect 245806 245928 245811 245984
rect 244076 245926 245811 245928
rect 197353 245923 197419 245926
rect 245745 245923 245811 245926
rect 67725 245712 68908 245714
rect 67725 245656 67730 245712
rect 67786 245656 68908 245712
rect 67725 245654 68908 245656
rect 166441 245712 190470 245714
rect 166441 245656 166446 245712
rect 166502 245656 190470 245712
rect 166441 245654 190470 245656
rect 245653 245714 245719 245717
rect 246113 245714 246179 245717
rect 245653 245712 246179 245714
rect 245653 245656 245658 245712
rect 245714 245656 246118 245712
rect 246174 245656 246179 245712
rect 245653 245654 246179 245656
rect 67725 245651 67791 245654
rect 166441 245651 166507 245654
rect 245653 245651 245719 245654
rect 246113 245651 246179 245654
rect 580165 245578 580231 245581
rect 583520 245578 584960 245668
rect 580165 245576 584960 245578
rect 580165 245520 580170 245576
rect 580226 245520 584960 245576
rect 580165 245518 584960 245520
rect 580165 245515 580231 245518
rect 583520 245428 584960 245518
rect 156646 244898 156706 245412
rect 197353 245170 197419 245173
rect 197353 245168 200284 245170
rect 197353 245112 197358 245168
rect 197414 245112 200284 245168
rect 197353 245110 200284 245112
rect 197353 245107 197419 245110
rect 156822 244972 156828 245036
rect 156892 245034 156898 245036
rect 168966 245034 168972 245036
rect 156892 244974 168972 245034
rect 156892 244972 156898 244974
rect 168966 244972 168972 244974
rect 169036 244972 169042 245036
rect 177389 245034 177455 245037
rect 185669 245034 185735 245037
rect 177389 245032 185735 245034
rect 177389 244976 177394 245032
rect 177450 244976 185674 245032
rect 185730 244976 185735 245032
rect 177389 244974 185735 244976
rect 177389 244971 177455 244974
rect 185669 244971 185735 244974
rect 244046 244901 244106 245140
rect 161289 244898 161355 244901
rect 181529 244898 181595 244901
rect 156646 244896 181595 244898
rect 156646 244840 161294 244896
rect 161350 244840 181534 244896
rect 181590 244840 181595 244896
rect 156646 244838 181595 244840
rect 161289 244835 161355 244838
rect 181529 244835 181595 244838
rect 243997 244896 244106 244901
rect 243997 244840 244002 244896
rect 244058 244840 244106 244896
rect 243997 244838 244106 244840
rect 243997 244835 244063 244838
rect 66345 244626 66411 244629
rect 245745 244626 245811 244629
rect 66345 244624 68908 244626
rect 66345 244568 66350 244624
rect 66406 244568 68908 244624
rect 66345 244566 68908 244568
rect 244076 244624 245811 244626
rect 244076 244568 245750 244624
rect 245806 244568 245811 244624
rect 244076 244566 245811 244568
rect 66345 244563 66411 244566
rect 245745 244563 245811 244566
rect 158713 244354 158779 244357
rect 156676 244352 158779 244354
rect 156676 244296 158718 244352
rect 158774 244296 158779 244352
rect 156676 244294 158779 244296
rect 158713 244291 158779 244294
rect 198457 244354 198523 244357
rect 198457 244352 200284 244354
rect 198457 244296 198462 244352
rect 198518 244296 200284 244352
rect 198457 244294 200284 244296
rect 198457 244291 198523 244294
rect 266353 244218 266419 244221
rect 244046 244216 266419 244218
rect 244046 244160 266358 244216
rect 266414 244160 266419 244216
rect 244046 244158 266419 244160
rect 197997 243810 198063 243813
rect 197997 243808 200284 243810
rect 197997 243752 198002 243808
rect 198058 243752 200284 243808
rect 244046 243780 244106 244158
rect 266353 244155 266419 244158
rect 197997 243750 200284 243752
rect 197997 243747 198063 243750
rect 176561 243674 176627 243677
rect 187141 243674 187207 243677
rect 176561 243672 187207 243674
rect 176561 243616 176566 243672
rect 176622 243616 187146 243672
rect 187202 243616 187207 243672
rect 176561 243614 187207 243616
rect 176561 243611 176627 243614
rect 187141 243611 187207 243614
rect 158161 243538 158227 243541
rect 191741 243538 191807 243541
rect 197445 243538 197511 243541
rect 158161 243536 197511 243538
rect 64638 242932 64644 242996
rect 64708 242994 64714 242996
rect 68878 242994 68938 243508
rect 158161 243480 158166 243536
rect 158222 243480 191746 243536
rect 191802 243480 197450 243536
rect 197506 243480 197511 243536
rect 158161 243478 197511 243480
rect 158161 243475 158227 243478
rect 191741 243475 191807 243478
rect 197445 243475 197511 243478
rect 158713 243266 158779 243269
rect 156676 243264 158779 243266
rect 156676 243208 158718 243264
rect 158774 243208 158779 243264
rect 156676 243206 158779 243208
rect 158713 243203 158779 243206
rect 64708 242934 68938 242994
rect 197353 242994 197419 242997
rect 245694 242994 245700 242996
rect 197353 242992 200284 242994
rect 197353 242936 197358 242992
rect 197414 242936 200284 242992
rect 197353 242934 200284 242936
rect 244076 242934 245700 242994
rect 64708 242932 64714 242934
rect 197353 242931 197419 242934
rect 245694 242932 245700 242934
rect 245764 242932 245770 242996
rect 67081 242858 67147 242861
rect 195329 242860 195395 242861
rect 67398 242858 67404 242860
rect 67081 242856 67404 242858
rect 67081 242800 67086 242856
rect 67142 242800 67404 242856
rect 67081 242798 67404 242800
rect 67081 242795 67147 242798
rect 67398 242796 67404 242798
rect 67468 242796 67474 242860
rect 195278 242858 195284 242860
rect 195238 242798 195284 242858
rect 195348 242856 195395 242860
rect 195390 242800 195395 242856
rect 195278 242796 195284 242798
rect 195348 242796 195395 242800
rect 195329 242795 195395 242796
rect 246389 242450 246455 242453
rect 244076 242448 246455 242450
rect 69430 241906 69490 242420
rect 244076 242392 246394 242448
rect 246450 242392 246455 242448
rect 244076 242390 246455 242392
rect 246389 242387 246455 242390
rect 157926 242178 157932 242180
rect 156676 242118 157932 242178
rect 157926 242116 157932 242118
rect 157996 242116 158002 242180
rect 197813 242178 197879 242181
rect 197813 242176 200284 242178
rect 197813 242120 197818 242176
rect 197874 242120 200284 242176
rect 197813 242118 200284 242120
rect 197813 242115 197879 242118
rect 80973 242044 81039 242045
rect 154665 242044 154731 242045
rect 80973 242042 81020 242044
rect 80928 242040 81020 242042
rect 80928 241984 80978 242040
rect 80928 241982 81020 241984
rect 80973 241980 81020 241982
rect 81084 241980 81090 242044
rect 154614 241980 154620 242044
rect 154684 242042 154731 242044
rect 154684 242040 154776 242042
rect 154726 241984 154776 242040
rect 154684 241982 154776 241984
rect 154684 241980 154731 241982
rect 80973 241979 81039 241980
rect 154665 241979 154731 241980
rect 69749 241906 69815 241909
rect 195278 241906 195284 241908
rect 69430 241904 69815 241906
rect 69430 241848 69754 241904
rect 69810 241848 69815 241904
rect 69430 241846 69815 241848
rect 69749 241843 69815 241846
rect 180750 241846 195284 241906
rect 67357 241770 67423 241773
rect 69657 241770 69723 241773
rect 67357 241768 69723 241770
rect 67357 241712 67362 241768
rect 67418 241712 69662 241768
rect 69718 241712 69723 241768
rect 67357 241710 69723 241712
rect 67357 241707 67423 241710
rect 69657 241707 69723 241710
rect 167821 241770 167887 241773
rect 180750 241770 180810 241846
rect 195278 241844 195284 241846
rect 195348 241844 195354 241908
rect 199929 241770 199995 241773
rect 167821 241768 180810 241770
rect 167821 241712 167826 241768
rect 167882 241712 180810 241768
rect 167821 241710 180810 241712
rect 195286 241768 199995 241770
rect 195286 241712 199934 241768
rect 199990 241712 199995 241768
rect 195286 241710 199995 241712
rect 167821 241707 167887 241710
rect 156689 241634 156755 241637
rect 170254 241634 170260 241636
rect 156689 241632 170260 241634
rect 156689 241576 156694 241632
rect 156750 241576 170260 241632
rect 156689 241574 170260 241576
rect 156689 241571 156755 241574
rect 170254 241572 170260 241574
rect 170324 241572 170330 241636
rect 180333 241634 180399 241637
rect 180609 241634 180675 241637
rect 195286 241634 195346 241710
rect 199929 241707 199995 241710
rect 180333 241632 195346 241634
rect 180333 241576 180338 241632
rect 180394 241576 180614 241632
rect 180670 241576 195346 241632
rect 180333 241574 195346 241576
rect 197077 241634 197143 241637
rect 197077 241632 200284 241634
rect 197077 241576 197082 241632
rect 197138 241576 200284 241632
rect 197077 241574 200284 241576
rect 180333 241571 180399 241574
rect 180609 241571 180675 241574
rect 197077 241571 197143 241574
rect 53649 241498 53715 241501
rect 83319 241498 83385 241501
rect 83549 241498 83615 241501
rect 53649 241496 83615 241498
rect 53649 241440 53654 241496
rect 53710 241440 83324 241496
rect 83380 241440 83554 241496
rect 83610 241440 83615 241496
rect 53649 241438 83615 241440
rect 53649 241435 53715 241438
rect 83319 241435 83385 241438
rect 83549 241435 83615 241438
rect 154159 241498 154225 241501
rect 156454 241498 156460 241500
rect 154159 241496 156460 241498
rect 154159 241440 154164 241496
rect 154220 241440 156460 241496
rect 154159 241438 156460 241440
rect 154159 241435 154225 241438
rect 156454 241436 156460 241438
rect 156524 241436 156530 241500
rect 146799 241362 146865 241365
rect 178769 241362 178835 241365
rect 146799 241360 178835 241362
rect 146799 241304 146804 241360
rect 146860 241304 178774 241360
rect 178830 241304 178835 241360
rect 146799 241302 178835 241304
rect 146799 241299 146865 241302
rect 178769 241299 178835 241302
rect 184749 241362 184815 241365
rect 186221 241362 186287 241365
rect 200021 241362 200087 241365
rect 243494 241364 243554 241604
rect 246297 241498 246363 241501
rect 299473 241498 299539 241501
rect 246297 241496 299539 241498
rect 246297 241440 246302 241496
rect 246358 241440 299478 241496
rect 299534 241440 299539 241496
rect 246297 241438 299539 241440
rect 246297 241435 246363 241438
rect 299473 241435 299539 241438
rect 184749 241360 200087 241362
rect 184749 241304 184754 241360
rect 184810 241304 186226 241360
rect 186282 241304 200026 241360
rect 200082 241304 200087 241360
rect 184749 241302 200087 241304
rect 184749 241299 184815 241302
rect 186221 241299 186287 241302
rect 200021 241299 200087 241302
rect 243486 241300 243492 241364
rect 243556 241300 243562 241364
rect 155125 241226 155191 241229
rect 158805 241226 158871 241229
rect 155125 241224 158871 241226
rect -960 241090 480 241180
rect 155125 241168 155130 241224
rect 155186 241168 158810 241224
rect 158866 241168 158871 241224
rect 155125 241166 158871 241168
rect 155125 241163 155191 241166
rect 158805 241163 158871 241166
rect 3509 241090 3575 241093
rect -960 241088 3575 241090
rect -960 241032 3514 241088
rect 3570 241032 3575 241088
rect -960 241030 3575 241032
rect -960 240940 480 241030
rect 3509 241027 3575 241030
rect 196985 240954 197051 240957
rect 196985 240952 200130 240954
rect 196985 240896 196990 240952
rect 197046 240896 200130 240952
rect 196985 240894 200130 240896
rect 196985 240891 197051 240894
rect 121361 240818 121427 240821
rect 151905 240818 151971 240821
rect 121361 240816 151971 240818
rect 121361 240760 121366 240816
rect 121422 240760 151910 240816
rect 151966 240760 151971 240816
rect 121361 240758 151971 240760
rect 121361 240755 121427 240758
rect 151905 240755 151971 240758
rect 157333 240818 157399 240821
rect 165153 240818 165219 240821
rect 157333 240816 165219 240818
rect 157333 240760 157338 240816
rect 157394 240760 165158 240816
rect 165214 240760 165219 240816
rect 157333 240758 165219 240760
rect 157333 240755 157399 240758
rect 165153 240755 165219 240758
rect 168373 240818 168439 240821
rect 197077 240818 197143 240821
rect 168373 240816 197143 240818
rect 168373 240760 168378 240816
rect 168434 240760 197082 240816
rect 197138 240760 197143 240816
rect 168373 240758 197143 240760
rect 200070 240818 200130 240894
rect 245653 240818 245719 240821
rect 200070 240758 200284 240818
rect 244076 240816 245719 240818
rect 244076 240760 245658 240816
rect 245714 240760 245719 240816
rect 244076 240758 245719 240760
rect 168373 240755 168439 240758
rect 197077 240755 197143 240758
rect 245653 240755 245719 240758
rect 121637 240274 121703 240277
rect 147213 240274 147279 240277
rect 245929 240274 245995 240277
rect 121637 240272 147279 240274
rect 121637 240216 121642 240272
rect 121698 240216 147218 240272
rect 147274 240216 147279 240272
rect 121637 240214 147279 240216
rect 244076 240272 245995 240274
rect 244076 240216 245934 240272
rect 245990 240216 245995 240272
rect 244076 240214 245995 240216
rect 121637 240211 121703 240214
rect 147213 240211 147279 240214
rect 245929 240211 245995 240214
rect 48129 240138 48195 240141
rect 77293 240138 77359 240141
rect 48129 240136 77359 240138
rect 48129 240080 48134 240136
rect 48190 240080 77298 240136
rect 77354 240080 77359 240136
rect 48129 240078 77359 240080
rect 48129 240075 48195 240078
rect 77293 240075 77359 240078
rect 155217 240138 155283 240141
rect 155769 240138 155835 240141
rect 155217 240136 155835 240138
rect 155217 240080 155222 240136
rect 155278 240080 155774 240136
rect 155830 240080 155835 240136
rect 155217 240078 155835 240080
rect 155217 240075 155283 240078
rect 155769 240075 155835 240078
rect 166809 240138 166875 240141
rect 168230 240138 168236 240140
rect 166809 240136 168236 240138
rect 166809 240080 166814 240136
rect 166870 240080 168236 240136
rect 166809 240078 168236 240080
rect 166809 240075 166875 240078
rect 168230 240076 168236 240078
rect 168300 240076 168306 240140
rect 199929 240138 199995 240141
rect 200573 240138 200639 240141
rect 202597 240140 202663 240141
rect 202597 240138 202644 240140
rect 199929 240136 200639 240138
rect 199929 240080 199934 240136
rect 199990 240080 200578 240136
rect 200634 240080 200639 240136
rect 199929 240078 200639 240080
rect 202552 240136 202644 240138
rect 202552 240080 202602 240136
rect 202552 240078 202644 240080
rect 199929 240075 199995 240078
rect 200573 240075 200639 240078
rect 202597 240076 202644 240078
rect 202708 240076 202714 240140
rect 202781 240138 202847 240141
rect 203190 240138 203196 240140
rect 202781 240136 203196 240138
rect 202781 240080 202786 240136
rect 202842 240080 203196 240136
rect 202781 240078 203196 240080
rect 202597 240075 202663 240076
rect 202781 240075 202847 240078
rect 203190 240076 203196 240078
rect 203260 240076 203266 240140
rect 207933 240138 207999 240141
rect 208209 240140 208275 240141
rect 208158 240138 208164 240140
rect 207933 240136 208164 240138
rect 208228 240138 208275 240140
rect 210693 240140 210759 240141
rect 213913 240140 213979 240141
rect 210693 240138 210740 240140
rect 208228 240136 208356 240138
rect 207933 240080 207938 240136
rect 207994 240080 208164 240136
rect 208270 240080 208356 240136
rect 207933 240078 208164 240080
rect 207933 240075 207999 240078
rect 208158 240076 208164 240078
rect 208228 240078 208356 240080
rect 210648 240136 210740 240138
rect 210648 240080 210698 240136
rect 210648 240078 210740 240080
rect 208228 240076 208275 240078
rect 208209 240075 208275 240076
rect 210693 240076 210740 240078
rect 210804 240076 210810 240140
rect 213862 240138 213868 240140
rect 213822 240078 213868 240138
rect 213932 240136 213979 240140
rect 213974 240080 213979 240136
rect 213862 240076 213868 240078
rect 213932 240076 213979 240080
rect 210693 240075 210759 240076
rect 213913 240075 213979 240076
rect 214189 240138 214255 240141
rect 217501 240140 217567 240141
rect 214414 240138 214420 240140
rect 214189 240136 214420 240138
rect 214189 240080 214194 240136
rect 214250 240080 214420 240136
rect 214189 240078 214420 240080
rect 214189 240075 214255 240078
rect 214414 240076 214420 240078
rect 214484 240076 214490 240140
rect 217501 240138 217548 240140
rect 217456 240136 217548 240138
rect 217612 240138 217618 240140
rect 217961 240138 218027 240141
rect 217612 240136 218027 240138
rect 217456 240080 217506 240136
rect 217612 240080 217966 240136
rect 218022 240080 218027 240136
rect 217456 240078 217548 240080
rect 217501 240076 217548 240078
rect 217612 240078 218027 240080
rect 217612 240076 217618 240078
rect 217501 240075 217567 240076
rect 217961 240075 218027 240078
rect 218421 240138 218487 240141
rect 218697 240138 218763 240141
rect 219198 240138 219204 240140
rect 218421 240136 219204 240138
rect 218421 240080 218426 240136
rect 218482 240080 218702 240136
rect 218758 240080 219204 240136
rect 218421 240078 219204 240080
rect 218421 240075 218487 240078
rect 218697 240075 218763 240078
rect 219198 240076 219204 240078
rect 219268 240076 219274 240140
rect 221038 240076 221044 240140
rect 221108 240138 221114 240140
rect 221365 240138 221431 240141
rect 221108 240136 221431 240138
rect 221108 240080 221370 240136
rect 221426 240080 221431 240136
rect 221108 240078 221431 240080
rect 221108 240076 221114 240078
rect 221365 240075 221431 240078
rect 230422 240076 230428 240140
rect 230492 240138 230498 240140
rect 230565 240138 230631 240141
rect 230492 240136 230631 240138
rect 230492 240080 230570 240136
rect 230626 240080 230631 240136
rect 230492 240078 230631 240080
rect 230492 240076 230498 240078
rect 230565 240075 230631 240078
rect 230749 240138 230815 240141
rect 230974 240138 230980 240140
rect 230749 240136 230980 240138
rect 230749 240080 230754 240136
rect 230810 240080 230980 240136
rect 230749 240078 230980 240080
rect 230749 240075 230815 240078
rect 230974 240076 230980 240078
rect 231044 240076 231050 240140
rect 231945 240138 232011 240141
rect 232078 240138 232084 240140
rect 231945 240136 232084 240138
rect 231945 240080 231950 240136
rect 232006 240080 232084 240136
rect 231945 240078 232084 240080
rect 231945 240075 232011 240078
rect 232078 240076 232084 240078
rect 232148 240076 232154 240140
rect 234470 240076 234476 240140
rect 234540 240138 234546 240140
rect 236453 240138 236519 240141
rect 234540 240136 236519 240138
rect 234540 240080 236458 240136
rect 236514 240080 236519 240136
rect 234540 240078 236519 240080
rect 234540 240076 234546 240078
rect 236453 240075 236519 240078
rect 237925 240138 237991 240141
rect 238702 240138 238708 240140
rect 237925 240136 238708 240138
rect 237925 240080 237930 240136
rect 237986 240080 238708 240136
rect 237925 240078 238708 240080
rect 237925 240075 237991 240078
rect 238702 240076 238708 240078
rect 238772 240076 238778 240140
rect 85113 240002 85179 240005
rect 207974 240002 207980 240004
rect 85113 240000 207980 240002
rect 85113 239944 85118 240000
rect 85174 239944 207980 240000
rect 85113 239942 207980 239944
rect 85113 239939 85179 239942
rect 207974 239940 207980 239942
rect 208044 240002 208050 240004
rect 208301 240002 208367 240005
rect 208044 240000 208367 240002
rect 208044 239944 208306 240000
rect 208362 239944 208367 240000
rect 208044 239942 208367 239944
rect 208044 239940 208050 239942
rect 208301 239939 208367 239942
rect 239213 240002 239279 240005
rect 259637 240002 259703 240005
rect 239213 240000 259703 240002
rect 239213 239944 239218 240000
rect 239274 239944 259642 240000
rect 259698 239944 259703 240000
rect 239213 239942 259703 239944
rect 239213 239939 239279 239942
rect 259637 239939 259703 239942
rect 80697 239594 80763 239597
rect 87597 239594 87663 239597
rect 80697 239592 87663 239594
rect 80697 239536 80702 239592
rect 80758 239536 87602 239592
rect 87658 239536 87663 239592
rect 80697 239534 87663 239536
rect 80697 239531 80763 239534
rect 87597 239531 87663 239534
rect 113633 239594 113699 239597
rect 205541 239594 205607 239597
rect 113633 239592 205607 239594
rect 113633 239536 113638 239592
rect 113694 239536 205546 239592
rect 205602 239536 205607 239592
rect 113633 239534 205607 239536
rect 113633 239531 113699 239534
rect 205541 239531 205607 239534
rect 207657 239594 207723 239597
rect 248454 239594 248460 239596
rect 207657 239592 248460 239594
rect 207657 239536 207662 239592
rect 207718 239536 248460 239592
rect 207657 239534 248460 239536
rect 207657 239531 207723 239534
rect 248454 239532 248460 239534
rect 248524 239532 248530 239596
rect 71681 239458 71747 239461
rect 86217 239458 86283 239461
rect 71681 239456 86283 239458
rect 71681 239400 71686 239456
rect 71742 239400 86222 239456
rect 86278 239400 86283 239456
rect 71681 239398 86283 239400
rect 71681 239395 71747 239398
rect 86217 239395 86283 239398
rect 122281 239458 122347 239461
rect 213821 239458 213887 239461
rect 122281 239456 213887 239458
rect 122281 239400 122286 239456
rect 122342 239400 213826 239456
rect 213882 239400 213887 239456
rect 122281 239398 213887 239400
rect 122281 239395 122347 239398
rect 213821 239395 213887 239398
rect 241237 239458 241303 239461
rect 262857 239458 262923 239461
rect 241237 239456 262923 239458
rect 241237 239400 241242 239456
rect 241298 239400 262862 239456
rect 262918 239400 262923 239456
rect 241237 239398 262923 239400
rect 241237 239395 241303 239398
rect 262857 239395 262923 239398
rect 39941 238642 40007 238645
rect 71773 238642 71839 238645
rect 39941 238640 71839 238642
rect 39941 238584 39946 238640
rect 40002 238584 71778 238640
rect 71834 238584 71839 238640
rect 39941 238582 71839 238584
rect 39941 238579 40007 238582
rect 71773 238579 71839 238582
rect 205817 238642 205883 238645
rect 206870 238642 206876 238644
rect 205817 238640 206876 238642
rect 205817 238584 205822 238640
rect 205878 238584 206876 238640
rect 205817 238582 206876 238584
rect 205817 238579 205883 238582
rect 206870 238580 206876 238582
rect 206940 238580 206946 238644
rect 212574 238580 212580 238644
rect 212644 238642 212650 238644
rect 213637 238642 213703 238645
rect 212644 238640 213703 238642
rect 212644 238584 213642 238640
rect 213698 238584 213703 238640
rect 212644 238582 213703 238584
rect 212644 238580 212650 238582
rect 213637 238579 213703 238582
rect 222326 238580 222332 238644
rect 222396 238642 222402 238644
rect 223481 238642 223547 238645
rect 222396 238640 223547 238642
rect 222396 238584 223486 238640
rect 223542 238584 223547 238640
rect 222396 238582 223547 238584
rect 222396 238580 222402 238582
rect 223481 238579 223547 238582
rect 235901 238642 235967 238645
rect 243854 238642 243860 238644
rect 235901 238640 243860 238642
rect 235901 238584 235906 238640
rect 235962 238584 243860 238640
rect 235901 238582 243860 238584
rect 235901 238579 235967 238582
rect 243854 238580 243860 238582
rect 243924 238580 243930 238644
rect 69105 238506 69171 238509
rect 180333 238506 180399 238509
rect 69105 238504 180399 238506
rect 69105 238448 69110 238504
rect 69166 238448 180338 238504
rect 180394 238448 180399 238504
rect 69105 238446 180399 238448
rect 69105 238443 69171 238446
rect 180333 238443 180399 238446
rect 196934 238444 196940 238508
rect 197004 238506 197010 238508
rect 204253 238506 204319 238509
rect 197004 238504 204319 238506
rect 197004 238448 204258 238504
rect 204314 238448 204319 238504
rect 197004 238446 204319 238448
rect 197004 238444 197010 238446
rect 204253 238443 204319 238446
rect 219525 238506 219591 238509
rect 224902 238506 224908 238508
rect 219525 238504 224908 238506
rect 219525 238448 219530 238504
rect 219586 238448 224908 238504
rect 219525 238446 224908 238448
rect 219525 238443 219591 238446
rect 224902 238444 224908 238446
rect 224972 238444 224978 238508
rect 226190 238444 226196 238508
rect 226260 238506 226266 238508
rect 232589 238506 232655 238509
rect 226260 238504 232655 238506
rect 226260 238448 232594 238504
rect 232650 238448 232655 238504
rect 226260 238446 232655 238448
rect 226260 238444 226266 238446
rect 232589 238443 232655 238446
rect 243537 238506 243603 238509
rect 260189 238506 260255 238509
rect 243537 238504 260255 238506
rect 243537 238448 243542 238504
rect 243598 238448 260194 238504
rect 260250 238448 260255 238504
rect 243537 238446 260255 238448
rect 243537 238443 243603 238446
rect 260189 238443 260255 238446
rect 114553 238370 114619 238373
rect 220997 238370 221063 238373
rect 114553 238368 221063 238370
rect 114553 238312 114558 238368
rect 114614 238312 221002 238368
rect 221058 238312 221063 238368
rect 114553 238310 221063 238312
rect 114553 238307 114619 238310
rect 220997 238307 221063 238310
rect 226701 238370 226767 238373
rect 285857 238370 285923 238373
rect 226701 238368 285923 238370
rect 226701 238312 226706 238368
rect 226762 238312 285862 238368
rect 285918 238312 285923 238368
rect 226701 238310 285923 238312
rect 226701 238307 226767 238310
rect 285857 238307 285923 238310
rect 96613 238234 96679 238237
rect 214189 238234 214255 238237
rect 96613 238232 214255 238234
rect 96613 238176 96618 238232
rect 96674 238176 214194 238232
rect 214250 238176 214255 238232
rect 96613 238174 214255 238176
rect 96613 238171 96679 238174
rect 214189 238171 214255 238174
rect 213821 238098 213887 238101
rect 226701 238098 226767 238101
rect 213821 238096 226767 238098
rect 213821 238040 213826 238096
rect 213882 238040 226706 238096
rect 226762 238040 226767 238096
rect 213821 238038 226767 238040
rect 213821 238035 213887 238038
rect 226701 238035 226767 238038
rect 71773 237418 71839 237421
rect 72417 237418 72483 237421
rect 71773 237416 72483 237418
rect 71773 237360 71778 237416
rect 71834 237360 72422 237416
rect 72478 237360 72483 237416
rect 71773 237358 72483 237360
rect 71773 237355 71839 237358
rect 72417 237355 72483 237358
rect 204253 237418 204319 237421
rect 205357 237418 205423 237421
rect 204253 237416 205423 237418
rect 204253 237360 204258 237416
rect 204314 237360 205362 237416
rect 205418 237360 205423 237416
rect 204253 237358 205423 237360
rect 204253 237355 204319 237358
rect 205357 237355 205423 237358
rect 78489 237284 78555 237285
rect 78438 237282 78444 237284
rect 78398 237222 78444 237282
rect 78508 237280 78555 237284
rect 78550 237224 78555 237280
rect 78438 237220 78444 237222
rect 78508 237220 78555 237224
rect 83958 237220 83964 237284
rect 84028 237282 84034 237284
rect 89713 237282 89779 237285
rect 84028 237280 89779 237282
rect 84028 237224 89718 237280
rect 89774 237224 89779 237280
rect 84028 237222 89779 237224
rect 84028 237220 84034 237222
rect 78489 237219 78555 237220
rect 89713 237219 89779 237222
rect 138013 237282 138079 237285
rect 142981 237282 143047 237285
rect 138013 237280 143047 237282
rect 138013 237224 138018 237280
rect 138074 237224 142986 237280
rect 143042 237224 143047 237280
rect 138013 237222 143047 237224
rect 138013 237219 138079 237222
rect 142981 237219 143047 237222
rect 152089 237282 152155 237285
rect 160829 237282 160895 237285
rect 152089 237280 160895 237282
rect 152089 237224 152094 237280
rect 152150 237224 160834 237280
rect 160890 237224 160895 237280
rect 152089 237222 160895 237224
rect 152089 237219 152155 237222
rect 160829 237219 160895 237222
rect 164141 237282 164207 237285
rect 207013 237282 207079 237285
rect 164141 237280 207079 237282
rect 164141 237224 164146 237280
rect 164202 237224 207018 237280
rect 207074 237224 207079 237280
rect 164141 237222 207079 237224
rect 164141 237219 164207 237222
rect 207013 237219 207079 237222
rect 208393 237282 208459 237285
rect 209221 237282 209287 237285
rect 317505 237282 317571 237285
rect 208393 237280 317571 237282
rect 208393 237224 208398 237280
rect 208454 237224 209226 237280
rect 209282 237224 317510 237280
rect 317566 237224 317571 237280
rect 208393 237222 317571 237224
rect 208393 237219 208459 237222
rect 209221 237219 209287 237222
rect 317505 237219 317571 237222
rect 143533 237146 143599 237149
rect 173249 237146 173315 237149
rect 143533 237144 173315 237146
rect 143533 237088 143538 237144
rect 143594 237088 173254 237144
rect 173310 237088 173315 237144
rect 143533 237086 173315 237088
rect 143533 237083 143599 237086
rect 173249 237083 173315 237086
rect 185577 237146 185643 237149
rect 210325 237146 210391 237149
rect 185577 237144 210391 237146
rect 185577 237088 185582 237144
rect 185638 237088 210330 237144
rect 210386 237088 210391 237144
rect 185577 237086 210391 237088
rect 185577 237083 185643 237086
rect 210325 237083 210391 237086
rect 231209 237146 231275 237149
rect 309869 237146 309935 237149
rect 231209 237144 309935 237146
rect 231209 237088 231214 237144
rect 231270 237088 309874 237144
rect 309930 237088 309935 237144
rect 231209 237086 309935 237088
rect 231209 237083 231275 237086
rect 309869 237083 309935 237086
rect 147673 237010 147739 237013
rect 158069 237010 158135 237013
rect 147673 237008 158135 237010
rect 147673 236952 147678 237008
rect 147734 236952 158074 237008
rect 158130 236952 158135 237008
rect 147673 236950 158135 236952
rect 147673 236947 147739 236950
rect 158069 236947 158135 236950
rect 191281 237010 191347 237013
rect 242709 237010 242775 237013
rect 191281 237008 242775 237010
rect 191281 236952 191286 237008
rect 191342 236952 242714 237008
rect 242770 236952 242775 237008
rect 191281 236950 242775 236952
rect 191281 236947 191347 236950
rect 242709 236947 242775 236950
rect 73470 236676 73476 236740
rect 73540 236738 73546 236740
rect 103421 236738 103487 236741
rect 73540 236736 103487 236738
rect 73540 236680 103426 236736
rect 103482 236680 103487 236736
rect 73540 236678 103487 236680
rect 73540 236676 73546 236678
rect 103421 236675 103487 236678
rect 107653 236738 107719 236741
rect 146845 236738 146911 236741
rect 107653 236736 146911 236738
rect 107653 236680 107658 236736
rect 107714 236680 146850 236736
rect 146906 236680 146911 236736
rect 107653 236678 146911 236680
rect 107653 236675 107719 236678
rect 146845 236675 146911 236678
rect 67265 236602 67331 236605
rect 142797 236602 142863 236605
rect 67265 236600 142863 236602
rect 67265 236544 67270 236600
rect 67326 236544 142802 236600
rect 142858 236544 142863 236600
rect 67265 236542 142863 236544
rect 67265 236539 67331 236542
rect 142797 236539 142863 236542
rect 89713 236058 89779 236061
rect 90357 236058 90423 236061
rect 89713 236056 90423 236058
rect 89713 236000 89718 236056
rect 89774 236000 90362 236056
rect 90418 236000 90423 236056
rect 89713 235998 90423 236000
rect 89713 235995 89779 235998
rect 90357 235995 90423 235998
rect 159265 236058 159331 236061
rect 159541 236058 159607 236061
rect 191741 236058 191807 236061
rect 159265 236056 191807 236058
rect 159265 236000 159270 236056
rect 159326 236000 159546 236056
rect 159602 236000 191746 236056
rect 191802 236000 191807 236056
rect 159265 235998 191807 236000
rect 159265 235995 159331 235998
rect 159541 235995 159607 235998
rect 191741 235995 191807 235998
rect 52177 235922 52243 235925
rect 93945 235922 94011 235925
rect 95141 235922 95207 235925
rect 52177 235920 95207 235922
rect 52177 235864 52182 235920
rect 52238 235864 93950 235920
rect 94006 235864 95146 235920
rect 95202 235864 95207 235920
rect 52177 235862 95207 235864
rect 52177 235859 52243 235862
rect 93945 235859 94011 235862
rect 95141 235859 95207 235862
rect 114645 235922 114711 235925
rect 154062 235922 154068 235924
rect 114645 235920 154068 235922
rect 114645 235864 114650 235920
rect 114706 235864 154068 235920
rect 114645 235862 154068 235864
rect 114645 235859 114711 235862
rect 154062 235860 154068 235862
rect 154132 235922 154138 235924
rect 208393 235922 208459 235925
rect 154132 235920 208459 235922
rect 154132 235864 208398 235920
rect 208454 235864 208459 235920
rect 154132 235862 208459 235864
rect 154132 235860 154138 235862
rect 208393 235859 208459 235862
rect 212717 235922 212783 235925
rect 239397 235922 239463 235925
rect 212717 235920 239463 235922
rect 212717 235864 212722 235920
rect 212778 235864 239402 235920
rect 239458 235864 239463 235920
rect 212717 235862 239463 235864
rect 212717 235859 212783 235862
rect 239397 235859 239463 235862
rect 240685 235922 240751 235925
rect 342345 235922 342411 235925
rect 240685 235920 342411 235922
rect 240685 235864 240690 235920
rect 240746 235864 342350 235920
rect 342406 235864 342411 235920
rect 240685 235862 342411 235864
rect 240685 235859 240751 235862
rect 342345 235859 342411 235862
rect 142981 235786 143047 235789
rect 162393 235786 162459 235789
rect 142981 235784 162459 235786
rect 142981 235728 142986 235784
rect 143042 235728 162398 235784
rect 162454 235728 162459 235784
rect 142981 235726 162459 235728
rect 142981 235723 143047 235726
rect 162393 235723 162459 235726
rect 172053 235786 172119 235789
rect 208853 235786 208919 235789
rect 172053 235784 208919 235786
rect 172053 235728 172058 235784
rect 172114 235728 208858 235784
rect 208914 235728 208919 235784
rect 172053 235726 208919 235728
rect 172053 235723 172119 235726
rect 208853 235723 208919 235726
rect 216581 235786 216647 235789
rect 263593 235786 263659 235789
rect 298737 235786 298803 235789
rect 216581 235784 298803 235786
rect 216581 235728 216586 235784
rect 216642 235728 263598 235784
rect 263654 235728 298742 235784
rect 298798 235728 298803 235784
rect 216581 235726 298803 235728
rect 216581 235723 216647 235726
rect 263593 235723 263659 235726
rect 298737 235723 298803 235726
rect 184054 235588 184060 235652
rect 184124 235650 184130 235652
rect 204437 235650 204503 235653
rect 184124 235648 204503 235650
rect 184124 235592 204442 235648
rect 204498 235592 204503 235648
rect 184124 235590 204503 235592
rect 184124 235588 184130 235590
rect 204437 235587 204503 235590
rect 228357 235650 228423 235653
rect 230197 235650 230263 235653
rect 228357 235648 230263 235650
rect 228357 235592 228362 235648
rect 228418 235592 230202 235648
rect 230258 235592 230263 235648
rect 228357 235590 230263 235592
rect 228357 235587 228423 235590
rect 230197 235587 230263 235590
rect 239213 235652 239279 235653
rect 239213 235648 239260 235652
rect 239324 235650 239330 235652
rect 247217 235650 247283 235653
rect 239324 235648 247283 235650
rect 239213 235592 239218 235648
rect 239324 235592 247222 235648
rect 247278 235592 247283 235648
rect 239213 235588 239260 235592
rect 239324 235590 247283 235592
rect 239324 235588 239330 235590
rect 239213 235587 239279 235588
rect 247217 235587 247283 235590
rect 95141 235242 95207 235245
rect 143349 235242 143415 235245
rect 95141 235240 143415 235242
rect 95141 235184 95146 235240
rect 95202 235184 143354 235240
rect 143410 235184 143415 235240
rect 95141 235182 143415 235184
rect 95141 235179 95207 235182
rect 143349 235179 143415 235182
rect 150433 235242 150499 235245
rect 158110 235242 158116 235244
rect 150433 235240 158116 235242
rect 150433 235184 150438 235240
rect 150494 235184 158116 235240
rect 150433 235182 158116 235184
rect 150433 235179 150499 235182
rect 158110 235180 158116 235182
rect 158180 235180 158186 235244
rect 164049 234698 164115 234701
rect 166993 234698 167059 234701
rect 164049 234696 167059 234698
rect 164049 234640 164054 234696
rect 164110 234640 166998 234696
rect 167054 234640 167059 234696
rect 164049 234638 167059 234640
rect 164049 234635 164115 234638
rect 166993 234635 167059 234638
rect 211889 234698 211955 234701
rect 212717 234698 212783 234701
rect 211889 234696 212783 234698
rect 211889 234640 211894 234696
rect 211950 234640 212722 234696
rect 212778 234640 212783 234696
rect 211889 234638 212783 234640
rect 211889 234635 211955 234638
rect 212717 234635 212783 234638
rect 65977 234562 66043 234565
rect 209773 234562 209839 234565
rect 210969 234562 211035 234565
rect 65977 234560 211035 234562
rect 65977 234504 65982 234560
rect 66038 234504 209778 234560
rect 209834 234504 210974 234560
rect 211030 234504 211035 234560
rect 65977 234502 211035 234504
rect 65977 234499 66043 234502
rect 209773 234499 209839 234502
rect 210969 234499 211035 234502
rect 215293 234562 215359 234565
rect 216029 234562 216095 234565
rect 574737 234562 574803 234565
rect 215293 234560 574803 234562
rect 215293 234504 215298 234560
rect 215354 234504 216034 234560
rect 216090 234504 574742 234560
rect 574798 234504 574803 234560
rect 215293 234502 574803 234504
rect 215293 234499 215359 234502
rect 216029 234499 216095 234502
rect 574737 234499 574803 234502
rect 146201 234426 146267 234429
rect 178033 234426 178099 234429
rect 146201 234424 178099 234426
rect 146201 234368 146206 234424
rect 146262 234368 178038 234424
rect 178094 234368 178099 234424
rect 146201 234366 178099 234368
rect 146201 234363 146267 234366
rect 178033 234363 178099 234366
rect 183093 234426 183159 234429
rect 228173 234426 228239 234429
rect 183093 234424 228239 234426
rect 183093 234368 183098 234424
rect 183154 234368 228178 234424
rect 228234 234368 228239 234424
rect 183093 234366 228239 234368
rect 183093 234363 183159 234366
rect 228173 234363 228239 234366
rect 232957 234426 233023 234429
rect 272609 234426 272675 234429
rect 232957 234424 272675 234426
rect 232957 234368 232962 234424
rect 233018 234368 272614 234424
rect 272670 234368 272675 234424
rect 232957 234366 272675 234368
rect 232957 234363 233023 234366
rect 272609 234363 272675 234366
rect 194317 234290 194383 234293
rect 202965 234290 203031 234293
rect 204161 234290 204227 234293
rect 194317 234288 204227 234290
rect 194317 234232 194322 234288
rect 194378 234232 202970 234288
rect 203026 234232 204166 234288
rect 204222 234232 204227 234288
rect 194317 234230 204227 234232
rect 194317 234227 194383 234230
rect 202965 234227 203031 234230
rect 204161 234227 204227 234230
rect 221457 234290 221523 234293
rect 255497 234290 255563 234293
rect 221457 234288 255563 234290
rect 221457 234232 221462 234288
rect 221518 234232 255502 234288
rect 255558 234232 255563 234288
rect 221457 234230 255563 234232
rect 221457 234227 221523 234230
rect 255497 234227 255563 234230
rect 178033 234154 178099 234157
rect 178677 234154 178743 234157
rect 178033 234152 178743 234154
rect 178033 234096 178038 234152
rect 178094 234096 178682 234152
rect 178738 234096 178743 234152
rect 178033 234094 178743 234096
rect 178033 234091 178099 234094
rect 178677 234091 178743 234094
rect 132585 233882 132651 233885
rect 158621 233882 158687 233885
rect 159214 233882 159220 233884
rect 132585 233880 159220 233882
rect 132585 233824 132590 233880
rect 132646 233824 158626 233880
rect 158682 233824 159220 233880
rect 132585 233822 159220 233824
rect 132585 233819 132651 233822
rect 158621 233819 158687 233822
rect 159214 233820 159220 233822
rect 159284 233820 159290 233884
rect 244457 233202 244523 233205
rect 180750 233200 244523 233202
rect 180750 233144 244462 233200
rect 244518 233144 244523 233200
rect 180750 233142 244523 233144
rect 117405 233066 117471 233069
rect 173801 233066 173867 233069
rect 117405 233064 173867 233066
rect 117405 233008 117410 233064
rect 117466 233008 173806 233064
rect 173862 233008 173867 233064
rect 117405 233006 173867 233008
rect 117405 233003 117471 233006
rect 173801 233003 173867 233006
rect 129825 232930 129891 232933
rect 164233 232930 164299 232933
rect 180750 232930 180810 233142
rect 244457 233139 244523 233142
rect 223297 233066 223363 233069
rect 262949 233066 263015 233069
rect 223297 233064 263015 233066
rect 223297 233008 223302 233064
rect 223358 233008 262954 233064
rect 263010 233008 263015 233064
rect 223297 233006 263015 233008
rect 223297 233003 223363 233006
rect 262949 233003 263015 233006
rect 129825 232928 180810 232930
rect 129825 232872 129830 232928
rect 129886 232872 164238 232928
rect 164294 232872 180810 232928
rect 129825 232870 180810 232872
rect 583477 232930 583543 232933
rect 583477 232928 583586 232930
rect 583477 232872 583482 232928
rect 583538 232872 583586 232928
rect 129825 232867 129891 232870
rect 164233 232867 164299 232870
rect 583477 232867 583586 232872
rect 57605 232794 57671 232797
rect 167821 232794 167887 232797
rect 57605 232792 167887 232794
rect 57605 232736 57610 232792
rect 57666 232736 167826 232792
rect 167882 232736 167887 232792
rect 57605 232734 167887 232736
rect 57605 232731 57671 232734
rect 167821 232731 167887 232734
rect 173801 232658 173867 232661
rect 195329 232658 195395 232661
rect 173801 232656 195395 232658
rect 173801 232600 173806 232656
rect 173862 232600 195334 232656
rect 195390 232600 195395 232656
rect 173801 232598 195395 232600
rect 173801 232595 173867 232598
rect 195329 232595 195395 232598
rect 199929 232658 199995 232661
rect 208485 232658 208551 232661
rect 199929 232656 208551 232658
rect 199929 232600 199934 232656
rect 199990 232600 208490 232656
rect 208546 232600 208551 232656
rect 199929 232598 208551 232600
rect 199929 232595 199995 232598
rect 208485 232595 208551 232598
rect 175181 232522 175247 232525
rect 226149 232522 226215 232525
rect 583526 232522 583586 232867
rect 175181 232520 226215 232522
rect 175181 232464 175186 232520
rect 175242 232464 226154 232520
rect 226210 232464 226215 232520
rect 175181 232462 226215 232464
rect 175181 232459 175247 232462
rect 226149 232459 226215 232462
rect 583342 232476 583586 232522
rect 583342 232462 584960 232476
rect 583342 232386 583402 232462
rect 583520 232386 584960 232462
rect 583342 232326 584960 232386
rect 583520 232236 584960 232326
rect 146845 231842 146911 231845
rect 156638 231842 156644 231844
rect 146845 231840 156644 231842
rect 146845 231784 146850 231840
rect 146906 231784 156644 231840
rect 146845 231782 156644 231784
rect 146845 231779 146911 231782
rect 156638 231780 156644 231782
rect 156708 231780 156714 231844
rect 64689 231706 64755 231709
rect 215293 231706 215359 231709
rect 64689 231704 215359 231706
rect 64689 231648 64694 231704
rect 64750 231648 215298 231704
rect 215354 231648 215359 231704
rect 64689 231646 215359 231648
rect 64689 231643 64755 231646
rect 215293 231643 215359 231646
rect 191741 231570 191807 231573
rect 208393 231570 208459 231573
rect 191741 231568 208459 231570
rect 191741 231512 191746 231568
rect 191802 231512 208398 231568
rect 208454 231512 208459 231568
rect 191741 231510 208459 231512
rect 191741 231507 191807 231510
rect 208393 231507 208459 231510
rect 59077 231434 59143 231437
rect 245694 231434 245700 231436
rect 59077 231432 245700 231434
rect 59077 231376 59082 231432
rect 59138 231376 245700 231432
rect 59077 231374 245700 231376
rect 59077 231371 59143 231374
rect 245694 231372 245700 231374
rect 245764 231372 245770 231436
rect 210969 231162 211035 231165
rect 582925 231162 582991 231165
rect 210969 231160 582991 231162
rect 210969 231104 210974 231160
rect 211030 231104 582930 231160
rect 582986 231104 582991 231160
rect 210969 231102 582991 231104
rect 210969 231099 211035 231102
rect 582925 231099 582991 231102
rect 83457 230482 83523 230485
rect 239765 230482 239831 230485
rect 83457 230480 239831 230482
rect 83457 230424 83462 230480
rect 83518 230424 239770 230480
rect 239826 230424 239831 230480
rect 83457 230422 239831 230424
rect 83457 230419 83523 230422
rect 239765 230419 239831 230422
rect 63217 230346 63283 230349
rect 198549 230346 198615 230349
rect 203517 230346 203583 230349
rect 63217 230344 203583 230346
rect 63217 230288 63222 230344
rect 63278 230288 198554 230344
rect 198610 230288 203522 230344
rect 203578 230288 203583 230344
rect 63217 230286 203583 230288
rect 63217 230283 63283 230286
rect 198549 230283 198615 230286
rect 203517 230283 203583 230286
rect 57697 230210 57763 230213
rect 163589 230210 163655 230213
rect 57697 230208 163655 230210
rect 57697 230152 57702 230208
rect 57758 230152 163594 230208
rect 163650 230152 163655 230208
rect 57697 230150 163655 230152
rect 57697 230147 57763 230150
rect 163589 230147 163655 230150
rect 195278 229740 195284 229804
rect 195348 229802 195354 229804
rect 268469 229802 268535 229805
rect 195348 229800 268535 229802
rect 195348 229744 268474 229800
rect 268530 229744 268535 229800
rect 195348 229742 268535 229744
rect 195348 229740 195354 229742
rect 268469 229739 268535 229742
rect 67633 228986 67699 228989
rect 231209 228986 231275 228989
rect 67633 228984 231275 228986
rect 67633 228928 67638 228984
rect 67694 228928 231214 228984
rect 231270 228928 231275 228984
rect 67633 228926 231275 228928
rect 67633 228923 67699 228926
rect 231209 228923 231275 228926
rect 70894 228788 70900 228852
rect 70964 228850 70970 228852
rect 102777 228850 102843 228853
rect 232957 228850 233023 228853
rect 70964 228848 233023 228850
rect 70964 228792 102782 228848
rect 102838 228792 232962 228848
rect 233018 228792 233023 228848
rect 70964 228790 233023 228792
rect 70964 228788 70970 228790
rect 102777 228787 102843 228790
rect 232957 228787 233023 228790
rect 135161 228714 135227 228717
rect 173014 228714 173020 228716
rect 135161 228712 173020 228714
rect 135161 228656 135166 228712
rect 135222 228656 173020 228712
rect 135161 228654 173020 228656
rect 135161 228651 135227 228654
rect 173014 228652 173020 228654
rect 173084 228652 173090 228716
rect 177941 228714 178007 228717
rect 212165 228714 212231 228717
rect 177941 228712 212231 228714
rect 177941 228656 177946 228712
rect 178002 228656 212170 228712
rect 212226 228656 212231 228712
rect 177941 228654 212231 228656
rect 177941 228651 178007 228654
rect 212165 228651 212231 228654
rect 212165 228306 212231 228309
rect 574737 228306 574803 228309
rect 212165 228304 574803 228306
rect 212165 228248 212170 228304
rect 212226 228248 574742 228304
rect 574798 228248 574803 228304
rect 212165 228246 574803 228248
rect 212165 228243 212231 228246
rect 574737 228243 574803 228246
rect -960 227884 480 228124
rect 177297 227762 177363 227765
rect 177941 227762 178007 227765
rect 177297 227760 178007 227762
rect 177297 227704 177302 227760
rect 177358 227704 177946 227760
rect 178002 227704 178007 227760
rect 177297 227702 178007 227704
rect 177297 227699 177363 227702
rect 177941 227699 178007 227702
rect 82670 227564 82676 227628
rect 82740 227626 82746 227628
rect 245929 227626 245995 227629
rect 82740 227624 245995 227626
rect 82740 227568 245934 227624
rect 245990 227568 245995 227624
rect 82740 227566 245995 227568
rect 82740 227564 82746 227566
rect 245929 227563 245995 227566
rect 144913 227490 144979 227493
rect 236821 227490 236887 227493
rect 144913 227488 236887 227490
rect 144913 227432 144918 227488
rect 144974 227432 236826 227488
rect 236882 227432 236887 227488
rect 144913 227430 236887 227432
rect 144913 227427 144979 227430
rect 236821 227427 236887 227430
rect 63125 226946 63191 226949
rect 146937 226946 147003 226949
rect 63125 226944 147003 226946
rect 63125 226888 63130 226944
rect 63186 226888 146942 226944
rect 146998 226888 147003 226944
rect 63125 226886 147003 226888
rect 63125 226883 63191 226886
rect 146937 226883 147003 226886
rect 236821 226946 236887 226949
rect 302141 226946 302207 226949
rect 236821 226944 302207 226946
rect 236821 226888 236826 226944
rect 236882 226888 302146 226944
rect 302202 226888 302207 226944
rect 236821 226886 302207 226888
rect 236821 226883 236887 226886
rect 302141 226883 302207 226886
rect 184749 226268 184815 226269
rect 184749 226264 184796 226268
rect 184860 226266 184866 226268
rect 184749 226208 184754 226264
rect 184749 226204 184796 226208
rect 184860 226206 184906 226266
rect 184860 226204 184866 226206
rect 184749 226203 184815 226204
rect 137277 226130 137343 226133
rect 171777 226130 171843 226133
rect 242934 226130 242940 226132
rect 137277 226128 242940 226130
rect 137277 226072 137282 226128
rect 137338 226072 171782 226128
rect 171838 226072 242940 226128
rect 137277 226070 242940 226072
rect 137277 226067 137343 226070
rect 171777 226067 171843 226070
rect 242934 226068 242940 226070
rect 243004 226068 243010 226132
rect 52269 225994 52335 225997
rect 227621 225994 227687 225997
rect 52269 225992 227687 225994
rect 52269 225936 52274 225992
rect 52330 225936 227626 225992
rect 227682 225936 227687 225992
rect 52269 225934 227687 225936
rect 52269 225931 52335 225934
rect 227621 225931 227687 225934
rect 69606 225660 69612 225724
rect 69676 225722 69682 225724
rect 195237 225722 195303 225725
rect 69676 225720 195303 225722
rect 69676 225664 195242 225720
rect 195298 225664 195303 225720
rect 69676 225662 195303 225664
rect 69676 225660 69682 225662
rect 195237 225659 195303 225662
rect 195329 225586 195395 225589
rect 583753 225586 583819 225589
rect 195329 225584 583819 225586
rect 195329 225528 195334 225584
rect 195390 225528 583758 225584
rect 583814 225528 583819 225584
rect 195329 225526 583819 225528
rect 195329 225523 195395 225526
rect 583753 225523 583819 225526
rect 58985 224906 59051 224909
rect 270033 224906 270099 224909
rect 270401 224906 270467 224909
rect 58985 224904 270467 224906
rect 58985 224848 58990 224904
rect 59046 224848 270038 224904
rect 270094 224848 270406 224904
rect 270462 224848 270467 224904
rect 58985 224846 270467 224848
rect 58985 224843 59051 224846
rect 270033 224843 270099 224846
rect 270401 224843 270467 224846
rect 66161 224770 66227 224773
rect 234981 224770 235047 224773
rect 66161 224768 235047 224770
rect 66161 224712 66166 224768
rect 66222 224712 234986 224768
rect 235042 224712 235047 224768
rect 66161 224710 235047 224712
rect 66161 224707 66227 224710
rect 234981 224707 235047 224710
rect 100937 224634 101003 224637
rect 102041 224634 102107 224637
rect 160870 224634 160876 224636
rect 100937 224632 160876 224634
rect 100937 224576 100942 224632
rect 100998 224576 102046 224632
rect 102102 224576 160876 224632
rect 100937 224574 160876 224576
rect 100937 224571 101003 224574
rect 102041 224571 102107 224574
rect 160870 224572 160876 224574
rect 160940 224572 160946 224636
rect 270401 224226 270467 224229
rect 279509 224226 279575 224229
rect 270401 224224 279575 224226
rect 270401 224168 270406 224224
rect 270462 224168 279514 224224
rect 279570 224168 279575 224224
rect 270401 224166 279575 224168
rect 270401 224163 270467 224166
rect 279509 224163 279575 224166
rect 147489 223546 147555 223549
rect 218697 223546 218763 223549
rect 233233 223548 233299 223549
rect 147489 223544 219450 223546
rect 147489 223488 147494 223544
rect 147550 223488 218702 223544
rect 218758 223488 219450 223544
rect 147489 223486 219450 223488
rect 147489 223483 147555 223486
rect 218697 223483 218763 223486
rect 166809 223410 166875 223413
rect 166809 223408 200130 223410
rect 166809 223352 166814 223408
rect 166870 223352 200130 223408
rect 166809 223350 200130 223352
rect 166809 223347 166875 223350
rect 32397 222866 32463 222869
rect 169845 222866 169911 222869
rect 32397 222864 169911 222866
rect 32397 222808 32402 222864
rect 32458 222808 169850 222864
rect 169906 222808 169911 222864
rect 32397 222806 169911 222808
rect 200070 222866 200130 223350
rect 219390 223002 219450 223486
rect 233182 223484 233188 223548
rect 233252 223546 233299 223548
rect 233252 223544 233344 223546
rect 233294 223488 233344 223544
rect 233252 223486 233344 223488
rect 233252 223484 233299 223486
rect 233233 223483 233299 223484
rect 285673 223002 285739 223005
rect 219390 223000 285739 223002
rect 219390 222944 285678 223000
rect 285734 222944 285739 223000
rect 219390 222942 285739 222944
rect 285673 222939 285739 222942
rect 204989 222866 205055 222869
rect 583661 222866 583727 222869
rect 200070 222864 583727 222866
rect 200070 222808 204994 222864
rect 205050 222808 583666 222864
rect 583722 222808 583727 222864
rect 200070 222806 583727 222808
rect 32397 222803 32463 222806
rect 169845 222803 169911 222806
rect 204989 222803 205055 222806
rect 583661 222803 583727 222806
rect 215109 222324 215175 222325
rect 215109 222320 215156 222324
rect 215220 222322 215226 222324
rect 215109 222264 215114 222320
rect 215109 222260 215156 222264
rect 215220 222262 215266 222322
rect 215220 222260 215226 222262
rect 215109 222259 215175 222260
rect 139393 222186 139459 222189
rect 231853 222186 231919 222189
rect 139393 222184 231919 222186
rect 139393 222128 139398 222184
rect 139454 222128 231858 222184
rect 231914 222128 231919 222184
rect 139393 222126 231919 222128
rect 139393 222123 139459 222126
rect 231853 222123 231919 222126
rect 111057 222050 111123 222053
rect 201493 222050 201559 222053
rect 202229 222050 202295 222053
rect 111057 222048 202295 222050
rect 111057 221992 111062 222048
rect 111118 221992 201498 222048
rect 201554 221992 202234 222048
rect 202290 221992 202295 222048
rect 111057 221990 202295 221992
rect 111057 221987 111123 221990
rect 201493 221987 201559 221990
rect 202229 221987 202295 221990
rect 159357 221914 159423 221917
rect 228357 221914 228423 221917
rect 159357 221912 228423 221914
rect 159357 221856 159362 221912
rect 159418 221856 228362 221912
rect 228418 221856 228423 221912
rect 159357 221854 228423 221856
rect 159357 221851 159423 221854
rect 228357 221851 228423 221854
rect 43437 221506 43503 221509
rect 159541 221506 159607 221509
rect 43437 221504 159607 221506
rect 43437 221448 43442 221504
rect 43498 221448 159546 221504
rect 159602 221448 159607 221504
rect 43437 221446 159607 221448
rect 43437 221443 43503 221446
rect 159541 221443 159607 221446
rect 61837 220826 61903 220829
rect 195094 220826 195100 220828
rect 61837 220824 195100 220826
rect 61837 220768 61842 220824
rect 61898 220768 195100 220824
rect 61837 220766 195100 220768
rect 61837 220763 61903 220766
rect 195094 220764 195100 220766
rect 195164 220764 195170 220828
rect 143441 220690 143507 220693
rect 160737 220690 160803 220693
rect 143441 220688 160803 220690
rect 143441 220632 143446 220688
rect 143502 220632 160742 220688
rect 160798 220632 160803 220688
rect 143441 220630 160803 220632
rect 143441 220627 143507 220630
rect 160737 220627 160803 220630
rect 75678 220084 75684 220148
rect 75748 220146 75754 220148
rect 309869 220146 309935 220149
rect 75748 220144 309935 220146
rect 75748 220088 309874 220144
rect 309930 220088 309935 220144
rect 75748 220086 309935 220088
rect 75748 220084 75754 220086
rect 309869 220083 309935 220086
rect 227713 219602 227779 219605
rect 228214 219602 228220 219604
rect 227713 219600 228220 219602
rect 227713 219544 227718 219600
rect 227774 219544 228220 219600
rect 227713 219542 228220 219544
rect 227713 219539 227779 219542
rect 228214 219540 228220 219542
rect 228284 219602 228290 219604
rect 231117 219602 231183 219605
rect 228284 219600 231183 219602
rect 228284 219544 231122 219600
rect 231178 219544 231183 219600
rect 228284 219542 231183 219544
rect 228284 219540 228290 219542
rect 231117 219539 231183 219542
rect 209773 219466 209839 219469
rect 211061 219466 211127 219469
rect 291193 219466 291259 219469
rect 209773 219464 291259 219466
rect 209773 219408 209778 219464
rect 209834 219408 211066 219464
rect 211122 219408 291198 219464
rect 291254 219408 291259 219464
rect 209773 219406 291259 219408
rect 209773 219403 209839 219406
rect 211061 219403 211127 219406
rect 291193 219403 291259 219406
rect 93853 219330 93919 219333
rect 95141 219330 95207 219333
rect 380893 219330 380959 219333
rect 93853 219328 380959 219330
rect 93853 219272 93858 219328
rect 93914 219272 95146 219328
rect 95202 219272 380898 219328
rect 380954 219272 380959 219328
rect 93853 219270 380959 219272
rect 93853 219267 93919 219270
rect 95141 219267 95207 219270
rect 380893 219267 380959 219270
rect 64505 219194 64571 219197
rect 180149 219194 180215 219197
rect 64505 219192 180215 219194
rect 64505 219136 64510 219192
rect 64566 219136 180154 219192
rect 180210 219136 180215 219192
rect 64505 219134 180215 219136
rect 64505 219131 64571 219134
rect 180149 219131 180215 219134
rect 185669 219194 185735 219197
rect 266353 219194 266419 219197
rect 185669 219192 266419 219194
rect 185669 219136 185674 219192
rect 185730 219136 266358 219192
rect 266414 219136 266419 219192
rect 185669 219134 266419 219136
rect 185669 219131 185735 219134
rect 266353 219131 266419 219134
rect 150341 219058 150407 219061
rect 172094 219058 172100 219060
rect 150341 219056 172100 219058
rect 150341 219000 150346 219056
rect 150402 219000 172100 219056
rect 150341 218998 172100 219000
rect 150341 218995 150407 218998
rect 172094 218996 172100 218998
rect 172164 218996 172170 219060
rect 583201 219058 583267 219061
rect 583520 219058 584960 219148
rect 583201 219056 584960 219058
rect 583201 219000 583206 219056
rect 583262 219000 584960 219056
rect 583201 218998 584960 219000
rect 583201 218995 583267 218998
rect 583520 218908 584960 218998
rect 69749 217970 69815 217973
rect 251357 217970 251423 217973
rect 69749 217968 251423 217970
rect 69749 217912 69754 217968
rect 69810 217912 251362 217968
rect 251418 217912 251423 217968
rect 69749 217910 251423 217912
rect 69749 217907 69815 217910
rect 251357 217907 251423 217910
rect 53557 217834 53623 217837
rect 176469 217834 176535 217837
rect 53557 217832 180810 217834
rect 53557 217776 53562 217832
rect 53618 217776 176474 217832
rect 176530 217776 180810 217832
rect 53557 217774 180810 217776
rect 53557 217771 53623 217774
rect 176469 217771 176535 217774
rect 112989 217698 113055 217701
rect 177982 217698 177988 217700
rect 112989 217696 177988 217698
rect 112989 217640 112994 217696
rect 113050 217640 177988 217696
rect 112989 217638 177988 217640
rect 112989 217635 113055 217638
rect 177982 217636 177988 217638
rect 178052 217636 178058 217700
rect 180750 217426 180810 217774
rect 204897 217426 204963 217429
rect 180750 217424 204963 217426
rect 180750 217368 204902 217424
rect 204958 217368 204963 217424
rect 180750 217366 204963 217368
rect 204897 217363 204963 217366
rect 177982 217228 177988 217292
rect 178052 217290 178058 217292
rect 298134 217290 298140 217292
rect 178052 217230 298140 217290
rect 178052 217228 178058 217230
rect 298134 217228 298140 217230
rect 298204 217228 298210 217292
rect 91001 216474 91067 216477
rect 187693 216474 187759 216477
rect 91001 216472 187759 216474
rect 91001 216416 91006 216472
rect 91062 216416 187698 216472
rect 187754 216416 187759 216472
rect 91001 216414 187759 216416
rect 91001 216411 91067 216414
rect 187693 216411 187759 216414
rect 146937 216338 147003 216341
rect 268377 216338 268443 216341
rect 269021 216338 269087 216341
rect 146937 216336 269087 216338
rect 146937 216280 146942 216336
rect 146998 216280 268382 216336
rect 268438 216280 269026 216336
rect 269082 216280 269087 216336
rect 146937 216278 269087 216280
rect 146937 216275 147003 216278
rect 268377 216275 268443 216278
rect 269021 216275 269087 216278
rect 175273 216066 175339 216069
rect 176510 216066 176516 216068
rect 175273 216064 176516 216066
rect 175273 216008 175278 216064
rect 175334 216008 176516 216064
rect 175273 216006 176516 216008
rect 175273 216003 175339 216006
rect 176510 216004 176516 216006
rect 176580 216004 176586 216068
rect 187693 216066 187759 216069
rect 188797 216066 188863 216069
rect 298093 216066 298159 216069
rect 187693 216064 298159 216066
rect 187693 216008 187698 216064
rect 187754 216008 188802 216064
rect 188858 216008 298098 216064
rect 298154 216008 298159 216064
rect 187693 216006 298159 216008
rect 187693 216003 187759 216006
rect 188797 216003 188863 216006
rect 298093 216003 298159 216006
rect 56501 215930 56567 215933
rect 195145 215930 195211 215933
rect 56501 215928 195211 215930
rect 56501 215872 56506 215928
rect 56562 215872 195150 215928
rect 195206 215872 195211 215928
rect 56501 215870 195211 215872
rect 56501 215867 56567 215870
rect 195145 215867 195211 215870
rect 211337 215930 211403 215933
rect 241421 215930 241487 215933
rect 241646 215930 241652 215932
rect 211337 215928 241652 215930
rect 211337 215872 211342 215928
rect 211398 215872 241426 215928
rect 241482 215872 241652 215928
rect 211337 215870 241652 215872
rect 211337 215867 211403 215870
rect 241421 215867 241487 215870
rect 241646 215868 241652 215870
rect 241716 215868 241722 215932
rect 269021 215930 269087 215933
rect 285029 215930 285095 215933
rect 269021 215928 285095 215930
rect 269021 215872 269026 215928
rect 269082 215872 285034 215928
rect 285090 215872 285095 215928
rect 269021 215870 285095 215872
rect 269021 215867 269087 215870
rect 285029 215867 285095 215870
rect 136449 215250 136515 215253
rect 188838 215250 188844 215252
rect 136449 215248 188844 215250
rect 136449 215192 136454 215248
rect 136510 215192 188844 215248
rect 136449 215190 188844 215192
rect 136449 215187 136515 215190
rect 188838 215188 188844 215190
rect 188908 215250 188914 215252
rect 259453 215250 259519 215253
rect 260741 215250 260807 215253
rect 188908 215190 190470 215250
rect 188908 215188 188914 215190
rect -960 214978 480 215068
rect 3417 214978 3483 214981
rect -960 214976 3483 214978
rect -960 214920 3422 214976
rect 3478 214920 3483 214976
rect -960 214918 3483 214920
rect -960 214828 480 214918
rect 3417 214915 3483 214918
rect 190410 214706 190470 215190
rect 219390 215248 260807 215250
rect 219390 215192 259458 215248
rect 259514 215192 260746 215248
rect 260802 215192 260807 215248
rect 219390 215190 260807 215192
rect 213269 215114 213335 215117
rect 219390 215114 219450 215190
rect 259453 215187 259519 215190
rect 260741 215187 260807 215190
rect 249885 215116 249951 215117
rect 249885 215114 249932 215116
rect 213269 215112 219450 215114
rect 213269 215056 213274 215112
rect 213330 215056 219450 215112
rect 213269 215054 219450 215056
rect 249840 215112 249932 215114
rect 249840 215056 249890 215112
rect 249840 215054 249932 215056
rect 213269 215051 213335 215054
rect 249885 215052 249932 215054
rect 249996 215052 250002 215116
rect 249885 215051 249951 215052
rect 302734 214706 302740 214708
rect 190410 214646 302740 214706
rect 302734 214644 302740 214646
rect 302804 214644 302810 214708
rect 77293 214570 77359 214573
rect 215201 214570 215267 214573
rect 215518 214570 215524 214572
rect 77293 214568 215524 214570
rect 77293 214512 77298 214568
rect 77354 214512 215206 214568
rect 215262 214512 215524 214568
rect 77293 214510 215524 214512
rect 77293 214507 77359 214510
rect 215201 214507 215267 214510
rect 215518 214508 215524 214510
rect 215588 214508 215594 214572
rect 183277 213892 183343 213893
rect 183277 213888 183324 213892
rect 183388 213890 183394 213892
rect 240133 213890 240199 213893
rect 240869 213890 240935 213893
rect 183277 213832 183282 213888
rect 183277 213828 183324 213832
rect 183388 213830 183434 213890
rect 219390 213888 240935 213890
rect 219390 213832 240138 213888
rect 240194 213832 240874 213888
rect 240930 213832 240935 213888
rect 219390 213830 240935 213832
rect 183388 213828 183394 213830
rect 183277 213827 183343 213828
rect 195145 213754 195211 213757
rect 219390 213754 219450 213830
rect 240133 213827 240199 213830
rect 240869 213827 240935 213830
rect 195145 213752 219450 213754
rect 195145 213696 195150 213752
rect 195206 213696 219450 213752
rect 195145 213694 219450 213696
rect 195145 213691 195211 213694
rect 50797 213618 50863 213621
rect 209773 213618 209839 213621
rect 50797 213616 209839 213618
rect 50797 213560 50802 213616
rect 50858 213560 209778 213616
rect 209834 213560 209839 213616
rect 50797 213558 209839 213560
rect 50797 213555 50863 213558
rect 209773 213555 209839 213558
rect 66662 213148 66668 213212
rect 66732 213210 66738 213212
rect 583477 213210 583543 213213
rect 66732 213208 583543 213210
rect 66732 213152 583482 213208
rect 583538 213152 583543 213208
rect 66732 213150 583543 213152
rect 66732 213148 66738 213150
rect 583477 213147 583543 213150
rect 87137 212530 87203 212533
rect 189073 212530 189139 212533
rect 87137 212528 189139 212530
rect 87137 212472 87142 212528
rect 87198 212472 189078 212528
rect 189134 212472 189139 212528
rect 87137 212470 189139 212472
rect 87137 212467 87203 212470
rect 189073 212467 189139 212470
rect 237373 212530 237439 212533
rect 237966 212530 237972 212532
rect 237373 212528 237972 212530
rect 237373 212472 237378 212528
rect 237434 212472 237972 212528
rect 237373 212470 237972 212472
rect 237373 212467 237439 212470
rect 237966 212468 237972 212470
rect 238036 212468 238042 212532
rect 100661 212394 100727 212397
rect 100661 212392 161490 212394
rect 100661 212336 100666 212392
rect 100722 212336 161490 212392
rect 100661 212334 161490 212336
rect 100661 212331 100727 212334
rect 161430 211850 161490 212334
rect 198457 211986 198523 211989
rect 207657 211986 207723 211989
rect 198457 211984 207723 211986
rect 198457 211928 198462 211984
rect 198518 211928 207662 211984
rect 207718 211928 207723 211984
rect 198457 211926 207723 211928
rect 198457 211923 198523 211926
rect 207657 211923 207723 211926
rect 208301 211986 208367 211989
rect 279417 211986 279483 211989
rect 208301 211984 279483 211986
rect 208301 211928 208306 211984
rect 208362 211928 279422 211984
rect 279478 211928 279483 211984
rect 208301 211926 279483 211928
rect 208301 211923 208367 211926
rect 279417 211923 279483 211926
rect 174670 211850 174676 211852
rect 161430 211790 174676 211850
rect 174670 211788 174676 211790
rect 174740 211850 174746 211852
rect 303613 211850 303679 211853
rect 174740 211848 303679 211850
rect 174740 211792 303618 211848
rect 303674 211792 303679 211848
rect 174740 211790 303679 211792
rect 174740 211788 174746 211790
rect 303613 211787 303679 211790
rect 209681 211308 209747 211309
rect 209630 211306 209636 211308
rect 209590 211246 209636 211306
rect 209700 211304 209747 211308
rect 209742 211248 209747 211304
rect 209630 211244 209636 211246
rect 209700 211244 209747 211248
rect 209681 211243 209747 211244
rect 97993 211170 98059 211173
rect 99281 211170 99347 211173
rect 97993 211168 99347 211170
rect 97993 211112 97998 211168
rect 98054 211112 99286 211168
rect 99342 211112 99347 211168
rect 97993 211110 99347 211112
rect 97993 211107 98059 211110
rect 99281 211107 99347 211110
rect 128353 211034 128419 211037
rect 231945 211034 232011 211037
rect 128353 211032 232011 211034
rect 128353 210976 128358 211032
rect 128414 210976 231950 211032
rect 232006 210976 232011 211032
rect 128353 210974 232011 210976
rect 128353 210971 128419 210974
rect 231945 210971 232011 210974
rect 75821 210898 75887 210901
rect 162158 210898 162164 210900
rect 75821 210896 162164 210898
rect 75821 210840 75826 210896
rect 75882 210840 162164 210896
rect 75821 210838 162164 210840
rect 75821 210835 75887 210838
rect 162158 210836 162164 210838
rect 162228 210836 162234 210900
rect 99281 210762 99347 210765
rect 163446 210762 163452 210764
rect 99281 210760 163452 210762
rect 99281 210704 99286 210760
rect 99342 210704 163452 210760
rect 99281 210702 163452 210704
rect 99281 210699 99347 210702
rect 163446 210700 163452 210702
rect 163516 210700 163522 210764
rect 191649 210354 191715 210357
rect 220261 210354 220327 210357
rect 191649 210352 220327 210354
rect 191649 210296 191654 210352
rect 191710 210296 220266 210352
rect 220322 210296 220327 210352
rect 191649 210294 220327 210296
rect 191649 210291 191715 210294
rect 220261 210291 220327 210294
rect 161197 209810 161263 209813
rect 335353 209810 335419 209813
rect 161197 209808 335419 209810
rect 161197 209752 161202 209808
rect 161258 209752 335358 209808
rect 335414 209752 335419 209808
rect 161197 209750 335419 209752
rect 161197 209747 161263 209750
rect 335353 209747 335419 209750
rect 82813 209674 82879 209677
rect 207749 209674 207815 209677
rect 82813 209672 207815 209674
rect 82813 209616 82818 209672
rect 82874 209616 207754 209672
rect 207810 209616 207815 209672
rect 82813 209614 207815 209616
rect 82813 209611 82879 209614
rect 207749 209611 207815 209614
rect 93761 209538 93827 209541
rect 179270 209538 179276 209540
rect 93761 209536 179276 209538
rect 93761 209480 93766 209536
rect 93822 209480 179276 209536
rect 93761 209478 179276 209480
rect 93761 209475 93827 209478
rect 179270 209476 179276 209478
rect 179340 209476 179346 209540
rect 118693 209402 118759 209405
rect 187785 209402 187851 209405
rect 118693 209400 187851 209402
rect 118693 209344 118698 209400
rect 118754 209344 187790 209400
rect 187846 209344 187851 209400
rect 118693 209342 187851 209344
rect 118693 209339 118759 209342
rect 187785 209339 187851 209342
rect 203609 209130 203675 209133
rect 289905 209130 289971 209133
rect 203609 209128 289971 209130
rect 203609 209072 203614 209128
rect 203670 209072 289910 209128
rect 289966 209072 289971 209128
rect 203609 209070 289971 209072
rect 203609 209067 203675 209070
rect 289905 209067 289971 209070
rect 179270 208932 179276 208996
rect 179340 208994 179346 208996
rect 340965 208994 341031 208997
rect 179340 208992 341031 208994
rect 179340 208936 340970 208992
rect 341026 208936 341031 208992
rect 179340 208934 341031 208936
rect 179340 208932 179346 208934
rect 340965 208931 341031 208934
rect 187785 208450 187851 208453
rect 188613 208450 188679 208453
rect 187785 208448 188679 208450
rect 187785 208392 187790 208448
rect 187846 208392 188618 208448
rect 188674 208392 188679 208448
rect 187785 208390 188679 208392
rect 187785 208387 187851 208390
rect 188613 208387 188679 208390
rect 86769 208314 86835 208317
rect 192702 208314 192708 208316
rect 86769 208312 192708 208314
rect 86769 208256 86774 208312
rect 86830 208256 192708 208312
rect 86769 208254 192708 208256
rect 86769 208251 86835 208254
rect 192702 208252 192708 208254
rect 192772 208252 192778 208316
rect 214557 207770 214623 207773
rect 283097 207770 283163 207773
rect 214557 207768 283163 207770
rect 214557 207712 214562 207768
rect 214618 207712 283102 207768
rect 283158 207712 283163 207768
rect 214557 207710 283163 207712
rect 214557 207707 214623 207710
rect 283097 207707 283163 207710
rect 117129 207634 117195 207637
rect 293166 207634 293172 207636
rect 117129 207632 293172 207634
rect 117129 207576 117134 207632
rect 117190 207576 293172 207632
rect 117129 207574 293172 207576
rect 117129 207571 117195 207574
rect 293166 207572 293172 207574
rect 293236 207634 293242 207636
rect 375465 207634 375531 207637
rect 293236 207632 375531 207634
rect 293236 207576 375470 207632
rect 375526 207576 375531 207632
rect 293236 207574 375531 207576
rect 293236 207572 293242 207574
rect 375465 207571 375531 207574
rect 192702 207164 192708 207228
rect 192772 207226 192778 207228
rect 195329 207226 195395 207229
rect 192772 207224 195395 207226
rect 192772 207168 195334 207224
rect 195390 207168 195395 207224
rect 192772 207166 195395 207168
rect 192772 207164 192778 207166
rect 195329 207163 195395 207166
rect 146937 207090 147003 207093
rect 205817 207090 205883 207093
rect 206461 207090 206527 207093
rect 146937 207088 206527 207090
rect 146937 207032 146942 207088
rect 146998 207032 205822 207088
rect 205878 207032 206466 207088
rect 206522 207032 206527 207088
rect 146937 207030 206527 207032
rect 146937 207027 147003 207030
rect 205817 207027 205883 207030
rect 206461 207027 206527 207030
rect 96521 206954 96587 206957
rect 96521 206952 180810 206954
rect 96521 206896 96526 206952
rect 96582 206896 180810 206952
rect 96521 206894 180810 206896
rect 96521 206891 96587 206894
rect 87597 206818 87663 206821
rect 146937 206818 147003 206821
rect 87597 206816 147003 206818
rect 87597 206760 87602 206816
rect 87658 206760 146942 206816
rect 146998 206760 147003 206816
rect 87597 206758 147003 206760
rect 87597 206755 87663 206758
rect 146937 206755 147003 206758
rect 180750 206410 180810 206894
rect 191598 206410 191604 206412
rect 180750 206350 191604 206410
rect 191598 206348 191604 206350
rect 191668 206410 191674 206412
rect 342897 206410 342963 206413
rect 191668 206408 342963 206410
rect 191668 206352 342902 206408
rect 342958 206352 342963 206408
rect 191668 206350 342963 206352
rect 191668 206348 191674 206350
rect 342897 206347 342963 206350
rect 81341 206274 81407 206277
rect 305729 206274 305795 206277
rect 583569 206274 583635 206277
rect 81341 206272 305795 206274
rect 81341 206216 81346 206272
rect 81402 206216 305734 206272
rect 305790 206216 305795 206272
rect 81341 206214 305795 206216
rect 81341 206211 81407 206214
rect 305729 206211 305795 206214
rect 583526 206272 583635 206274
rect 583526 206216 583574 206272
rect 583630 206216 583635 206272
rect 583526 206211 583635 206216
rect 583526 205866 583586 206211
rect 583342 205820 583586 205866
rect 583342 205806 584960 205820
rect 583342 205730 583402 205806
rect 583520 205730 584960 205806
rect 583342 205670 584960 205730
rect 131021 205594 131087 205597
rect 197118 205594 197124 205596
rect 131021 205592 197124 205594
rect 131021 205536 131026 205592
rect 131082 205536 197124 205592
rect 131021 205534 197124 205536
rect 131021 205531 131087 205534
rect 197118 205532 197124 205534
rect 197188 205594 197194 205596
rect 197188 205534 200130 205594
rect 583520 205580 584960 205670
rect 197188 205532 197194 205534
rect 200070 205050 200130 205534
rect 296713 205050 296779 205053
rect 200070 205048 296779 205050
rect 200070 204992 296718 205048
rect 296774 204992 296779 205048
rect 200070 204990 296779 204992
rect 296713 204987 296779 204990
rect 67081 204914 67147 204917
rect 583569 204914 583635 204917
rect 67081 204912 583635 204914
rect 67081 204856 67086 204912
rect 67142 204856 583574 204912
rect 583630 204856 583635 204912
rect 67081 204854 583635 204856
rect 67081 204851 67147 204854
rect 583569 204851 583635 204854
rect 54937 204234 55003 204237
rect 218053 204234 218119 204237
rect 54937 204232 218119 204234
rect 54937 204176 54942 204232
rect 54998 204176 218058 204232
rect 218114 204176 218119 204232
rect 54937 204174 218119 204176
rect 54937 204171 55003 204174
rect 218053 204171 218119 204174
rect 151721 204098 151787 204101
rect 240777 204098 240843 204101
rect 151721 204096 240843 204098
rect 151721 204040 151726 204096
rect 151782 204040 240782 204096
rect 240838 204040 240843 204096
rect 151721 204038 240843 204040
rect 151721 204035 151787 204038
rect 240777 204035 240843 204038
rect 102041 203554 102107 203557
rect 180057 203554 180123 203557
rect 102041 203552 180123 203554
rect 102041 203496 102046 203552
rect 102102 203496 180062 203552
rect 180118 203496 180123 203552
rect 102041 203494 180123 203496
rect 102041 203491 102107 203494
rect 180057 203491 180123 203494
rect 188337 203554 188403 203557
rect 256693 203554 256759 203557
rect 188337 203552 256759 203554
rect 188337 203496 188342 203552
rect 188398 203496 256698 203552
rect 256754 203496 256759 203552
rect 188337 203494 256759 203496
rect 188337 203491 188403 203494
rect 256693 203491 256759 203494
rect 121361 202874 121427 202877
rect 169201 202874 169267 202877
rect 121361 202872 169267 202874
rect 121361 202816 121366 202872
rect 121422 202816 169206 202872
rect 169262 202816 169267 202872
rect 121361 202814 169267 202816
rect 121361 202811 121427 202814
rect 169201 202811 169267 202814
rect 129641 202738 129707 202741
rect 162117 202738 162183 202741
rect 129641 202736 162183 202738
rect 129641 202680 129646 202736
rect 129702 202680 162122 202736
rect 162178 202680 162183 202736
rect 129641 202678 162183 202680
rect 129641 202675 129707 202678
rect 162117 202675 162183 202678
rect 169385 202330 169451 202333
rect 199326 202330 199332 202332
rect 169385 202328 199332 202330
rect 169385 202272 169390 202328
rect 169446 202272 199332 202328
rect 169385 202270 199332 202272
rect 169385 202267 169451 202270
rect 199326 202268 199332 202270
rect 199396 202330 199402 202332
rect 281625 202330 281691 202333
rect 199396 202328 281691 202330
rect 199396 202272 281630 202328
rect 281686 202272 281691 202328
rect 199396 202270 281691 202272
rect 199396 202268 199402 202270
rect 281625 202267 281691 202270
rect 166257 202194 166323 202197
rect 313273 202194 313339 202197
rect 166257 202192 313339 202194
rect 166257 202136 166262 202192
rect 166318 202136 313278 202192
rect 313334 202136 313339 202192
rect 166257 202134 313339 202136
rect 166257 202131 166323 202134
rect 313273 202131 313339 202134
rect -960 201922 480 202012
rect 3417 201922 3483 201925
rect -960 201920 3483 201922
rect -960 201864 3422 201920
rect 3478 201864 3483 201920
rect -960 201862 3483 201864
rect -960 201772 480 201862
rect 3417 201859 3483 201862
rect 67950 201316 67956 201380
rect 68020 201378 68026 201380
rect 213269 201378 213335 201381
rect 68020 201376 213335 201378
rect 68020 201320 213274 201376
rect 213330 201320 213335 201376
rect 68020 201318 213335 201320
rect 68020 201316 68026 201318
rect 213269 201315 213335 201318
rect 136541 201242 136607 201245
rect 166349 201242 166415 201245
rect 136541 201240 166415 201242
rect 136541 201184 136546 201240
rect 136602 201184 166354 201240
rect 166410 201184 166415 201240
rect 136541 201182 166415 201184
rect 136541 201179 136607 201182
rect 166349 201179 166415 201182
rect 192569 200834 192635 200837
rect 273989 200834 274055 200837
rect 192569 200832 274055 200834
rect 192569 200776 192574 200832
rect 192630 200776 273994 200832
rect 274050 200776 274055 200832
rect 192569 200774 274055 200776
rect 192569 200771 192635 200774
rect 273989 200771 274055 200774
rect 155861 200698 155927 200701
rect 300117 200698 300183 200701
rect 155861 200696 300183 200698
rect 155861 200640 155866 200696
rect 155922 200640 300122 200696
rect 300178 200640 300183 200696
rect 155861 200638 300183 200640
rect 155861 200635 155927 200638
rect 300117 200635 300183 200638
rect 180241 199610 180307 199613
rect 224902 199610 224908 199612
rect 180241 199608 224908 199610
rect 180241 199552 180246 199608
rect 180302 199552 224908 199608
rect 180241 199550 224908 199552
rect 180241 199547 180307 199550
rect 224902 199548 224908 199550
rect 224972 199548 224978 199612
rect 158621 199474 158687 199477
rect 182817 199474 182883 199477
rect 158621 199472 182883 199474
rect 158621 199416 158626 199472
rect 158682 199416 182822 199472
rect 182878 199416 182883 199472
rect 158621 199414 182883 199416
rect 158621 199411 158687 199414
rect 182817 199411 182883 199414
rect 197077 199474 197143 199477
rect 317505 199474 317571 199477
rect 197077 199472 317571 199474
rect 197077 199416 197082 199472
rect 197138 199416 317510 199472
rect 317566 199416 317571 199472
rect 197077 199414 317571 199416
rect 197077 199411 197143 199414
rect 317505 199411 317571 199414
rect 92381 199338 92447 199341
rect 246246 199338 246252 199340
rect 92381 199336 246252 199338
rect 92381 199280 92386 199336
rect 92442 199280 246252 199336
rect 92381 199278 246252 199280
rect 92381 199275 92447 199278
rect 246246 199276 246252 199278
rect 246316 199276 246322 199340
rect 79869 198658 79935 198661
rect 284293 198658 284359 198661
rect 79869 198656 284359 198658
rect 79869 198600 79874 198656
rect 79930 198600 284298 198656
rect 284354 198600 284359 198656
rect 79869 198598 284359 198600
rect 79869 198595 79935 198598
rect 284293 198595 284359 198598
rect 178677 197978 178743 197981
rect 248454 197978 248460 197980
rect 178677 197976 248460 197978
rect 178677 197920 178682 197976
rect 178738 197920 248460 197976
rect 178677 197918 248460 197920
rect 178677 197915 178743 197918
rect 248454 197916 248460 197918
rect 248524 197916 248530 197980
rect 86861 197298 86927 197301
rect 211654 197298 211660 197300
rect 86861 197296 211660 197298
rect 86861 197240 86866 197296
rect 86922 197240 211660 197296
rect 86861 197238 211660 197240
rect 86861 197235 86927 197238
rect 211654 197236 211660 197238
rect 211724 197298 211730 197300
rect 212390 197298 212396 197300
rect 211724 197238 212396 197298
rect 211724 197236 211730 197238
rect 212390 197236 212396 197238
rect 212460 197236 212466 197300
rect 190453 197162 190519 197165
rect 246021 197162 246087 197165
rect 190453 197160 246087 197162
rect 190453 197104 190458 197160
rect 190514 197104 246026 197160
rect 246082 197104 246087 197160
rect 190453 197102 246087 197104
rect 190453 197099 190519 197102
rect 246021 197099 246087 197102
rect 173014 196692 173020 196756
rect 173084 196754 173090 196756
rect 188429 196754 188495 196757
rect 173084 196752 188495 196754
rect 173084 196696 188434 196752
rect 188490 196696 188495 196752
rect 173084 196694 188495 196696
rect 173084 196692 173090 196694
rect 188429 196691 188495 196694
rect 122741 196618 122807 196621
rect 197997 196618 198063 196621
rect 122741 196616 198063 196618
rect 122741 196560 122746 196616
rect 122802 196560 198002 196616
rect 198058 196560 198063 196616
rect 122741 196558 198063 196560
rect 122741 196555 122807 196558
rect 197997 196555 198063 196558
rect 212390 196556 212396 196620
rect 212460 196618 212466 196620
rect 258574 196618 258580 196620
rect 212460 196558 258580 196618
rect 212460 196556 212466 196558
rect 258574 196556 258580 196558
rect 258644 196556 258650 196620
rect 174721 195938 174787 195941
rect 267825 195938 267891 195941
rect 268377 195938 268443 195941
rect 174721 195936 268443 195938
rect 174721 195880 174726 195936
rect 174782 195880 267830 195936
rect 267886 195880 268382 195936
rect 268438 195880 268443 195936
rect 174721 195878 268443 195880
rect 174721 195875 174787 195878
rect 267825 195875 267891 195878
rect 268377 195875 268443 195878
rect 188613 195394 188679 195397
rect 291469 195394 291535 195397
rect 188613 195392 291535 195394
rect 188613 195336 188618 195392
rect 188674 195336 291474 195392
rect 291530 195336 291535 195392
rect 188613 195334 291535 195336
rect 188613 195331 188679 195334
rect 291469 195331 291535 195334
rect 72417 195258 72483 195261
rect 351913 195258 351979 195261
rect 72417 195256 351979 195258
rect 72417 195200 72422 195256
rect 72478 195200 351918 195256
rect 351974 195200 351979 195256
rect 72417 195198 351979 195200
rect 72417 195195 72483 195198
rect 351913 195195 351979 195198
rect 60457 194578 60523 194581
rect 233509 194578 233575 194581
rect 60457 194576 233575 194578
rect 60457 194520 60462 194576
rect 60518 194520 233514 194576
rect 233570 194520 233575 194576
rect 60457 194518 233575 194520
rect 60457 194515 60523 194518
rect 233509 194515 233575 194518
rect 88977 193898 89043 193901
rect 322933 193898 322999 193901
rect 88977 193896 322999 193898
rect 88977 193840 88982 193896
rect 89038 193840 322938 193896
rect 322994 193840 322999 193896
rect 88977 193838 322999 193840
rect 88977 193835 89043 193838
rect 322933 193835 322999 193838
rect 93117 193218 93183 193221
rect 211797 193218 211863 193221
rect 93117 193216 211863 193218
rect 93117 193160 93122 193216
rect 93178 193160 211802 193216
rect 211858 193160 211863 193216
rect 93117 193158 211863 193160
rect 93117 193155 93183 193158
rect 211797 193155 211863 193158
rect 200757 192674 200823 192677
rect 244181 192674 244247 192677
rect 200757 192672 244247 192674
rect 200757 192616 200762 192672
rect 200818 192616 244186 192672
rect 244242 192616 244247 192672
rect 200757 192614 244247 192616
rect 200757 192611 200823 192614
rect 244181 192611 244247 192614
rect 79961 192538 80027 192541
rect 220721 192538 220787 192541
rect 220854 192538 220860 192540
rect 79961 192536 220860 192538
rect 79961 192480 79966 192536
rect 80022 192480 220726 192536
rect 220782 192480 220860 192536
rect 79961 192478 220860 192480
rect 79961 192475 80027 192478
rect 220721 192475 220787 192478
rect 220854 192476 220860 192478
rect 220924 192476 220930 192540
rect 223389 192538 223455 192541
rect 279325 192538 279391 192541
rect 223389 192536 279391 192538
rect 223389 192480 223394 192536
rect 223450 192480 279330 192536
rect 279386 192480 279391 192536
rect 223389 192478 279391 192480
rect 223389 192475 223455 192478
rect 279325 192475 279391 192478
rect 582649 192538 582715 192541
rect 583520 192538 584960 192628
rect 582649 192536 584960 192538
rect 582649 192480 582654 192536
rect 582710 192480 584960 192536
rect 582649 192478 584960 192480
rect 582649 192475 582715 192478
rect 583520 192388 584960 192478
rect 195513 191178 195579 191181
rect 236085 191178 236151 191181
rect 195513 191176 236151 191178
rect 195513 191120 195518 191176
rect 195574 191120 236090 191176
rect 236146 191120 236151 191176
rect 195513 191118 236151 191120
rect 195513 191115 195579 191118
rect 236085 191115 236151 191118
rect 104801 191042 104867 191045
rect 316677 191042 316743 191045
rect 104801 191040 316743 191042
rect 104801 190984 104806 191040
rect 104862 190984 316682 191040
rect 316738 190984 316743 191040
rect 104801 190982 316743 190984
rect 104801 190979 104867 190982
rect 316677 190979 316743 190982
rect 64781 190362 64847 190365
rect 266261 190362 266327 190365
rect 64781 190360 266327 190362
rect 64781 190304 64786 190360
rect 64842 190304 266266 190360
rect 266322 190304 266327 190360
rect 64781 190302 266327 190304
rect 64781 190299 64847 190302
rect 266261 190299 266327 190302
rect 266261 189818 266327 189821
rect 302509 189818 302575 189821
rect 266261 189816 302575 189818
rect 266261 189760 266266 189816
rect 266322 189760 302514 189816
rect 302570 189760 302575 189816
rect 266261 189758 302575 189760
rect 266261 189755 266327 189758
rect 302509 189755 302575 189758
rect 107561 189682 107627 189685
rect 287646 189682 287652 189684
rect 107561 189680 287652 189682
rect 107561 189624 107566 189680
rect 107622 189624 287652 189680
rect 107561 189622 287652 189624
rect 107561 189619 107627 189622
rect 287646 189620 287652 189622
rect 287716 189682 287722 189684
rect 288382 189682 288388 189684
rect 287716 189622 288388 189682
rect 287716 189620 287722 189622
rect 288382 189620 288388 189622
rect 288452 189620 288458 189684
rect 242934 189076 242940 189140
rect 243004 189138 243010 189140
rect 243905 189138 243971 189141
rect 243004 189136 243971 189138
rect 243004 189080 243910 189136
rect 243966 189080 243971 189136
rect 243004 189078 243971 189080
rect 243004 189076 243010 189078
rect 243905 189075 243971 189078
rect -960 188866 480 188956
rect 3509 188866 3575 188869
rect -960 188864 3575 188866
rect -960 188808 3514 188864
rect 3570 188808 3575 188864
rect -960 188806 3575 188808
rect -960 188716 480 188806
rect 3509 188803 3575 188806
rect 206369 188594 206435 188597
rect 237414 188594 237420 188596
rect 206369 188592 237420 188594
rect 206369 188536 206374 188592
rect 206430 188536 237420 188592
rect 206369 188534 237420 188536
rect 206369 188531 206435 188534
rect 237414 188532 237420 188534
rect 237484 188532 237490 188596
rect 216438 188396 216444 188460
rect 216508 188458 216514 188460
rect 284518 188458 284524 188460
rect 216508 188398 284524 188458
rect 216508 188396 216514 188398
rect 284518 188396 284524 188398
rect 284588 188396 284594 188460
rect 77150 188260 77156 188324
rect 77220 188322 77226 188324
rect 324313 188322 324379 188325
rect 77220 188320 324379 188322
rect 77220 188264 324318 188320
rect 324374 188264 324379 188320
rect 77220 188262 324379 188264
rect 77220 188260 77226 188262
rect 324313 188259 324379 188262
rect 61929 187642 61995 187645
rect 195421 187642 195487 187645
rect 61929 187640 195487 187642
rect 61929 187584 61934 187640
rect 61990 187584 195426 187640
rect 195482 187584 195487 187640
rect 61929 187582 195487 187584
rect 61929 187579 61995 187582
rect 195421 187579 195487 187582
rect 186129 187098 186195 187101
rect 301037 187098 301103 187101
rect 186129 187096 301103 187098
rect 186129 187040 186134 187096
rect 186190 187040 301042 187096
rect 301098 187040 301103 187096
rect 186129 187038 301103 187040
rect 186129 187035 186195 187038
rect 301037 187035 301103 187038
rect 99281 186962 99347 186965
rect 240225 186962 240291 186965
rect 99281 186960 240291 186962
rect 99281 186904 99286 186960
rect 99342 186904 240230 186960
rect 240286 186904 240291 186960
rect 99281 186902 240291 186904
rect 99281 186899 99347 186902
rect 240225 186899 240291 186902
rect 95141 186282 95207 186285
rect 230197 186282 230263 186285
rect 95141 186280 230263 186282
rect 95141 186224 95146 186280
rect 95202 186224 230202 186280
rect 230258 186224 230263 186280
rect 95141 186222 230263 186224
rect 95141 186219 95207 186222
rect 230197 186219 230263 186222
rect 220721 185874 220787 185877
rect 233366 185874 233372 185876
rect 220721 185872 233372 185874
rect 220721 185816 220726 185872
rect 220782 185816 233372 185872
rect 220721 185814 233372 185816
rect 220721 185811 220787 185814
rect 233366 185812 233372 185814
rect 233436 185812 233442 185876
rect 231117 185738 231183 185741
rect 232078 185738 232084 185740
rect 231117 185736 232084 185738
rect 231117 185680 231122 185736
rect 231178 185680 232084 185736
rect 231117 185678 232084 185680
rect 231117 185675 231183 185678
rect 232078 185676 232084 185678
rect 232148 185676 232154 185740
rect 142061 185602 142127 185605
rect 332593 185602 332659 185605
rect 338849 185602 338915 185605
rect 142061 185600 338915 185602
rect 142061 185544 142066 185600
rect 142122 185544 332598 185600
rect 332654 185544 338854 185600
rect 338910 185544 338915 185600
rect 142061 185542 338915 185544
rect 142061 185539 142127 185542
rect 332593 185539 332659 185542
rect 338849 185539 338915 185542
rect 233049 185058 233115 185061
rect 299606 185058 299612 185060
rect 233049 185056 299612 185058
rect 233049 185000 233054 185056
rect 233110 185000 299612 185056
rect 233049 184998 299612 185000
rect 233049 184995 233115 184998
rect 299606 184996 299612 184998
rect 299676 184996 299682 185060
rect 217409 184514 217475 184517
rect 230657 184514 230723 184517
rect 217409 184512 230723 184514
rect 217409 184456 217414 184512
rect 217470 184456 230662 184512
rect 230718 184456 230723 184512
rect 217409 184454 230723 184456
rect 217409 184451 217475 184454
rect 230657 184451 230723 184454
rect 166901 184378 166967 184381
rect 280153 184378 280219 184381
rect 166901 184376 280219 184378
rect 166901 184320 166906 184376
rect 166962 184320 280158 184376
rect 280214 184320 280219 184376
rect 166901 184318 280219 184320
rect 166901 184315 166967 184318
rect 280153 184315 280219 184318
rect 154481 184242 154547 184245
rect 316033 184242 316099 184245
rect 371233 184242 371299 184245
rect 154481 184240 371299 184242
rect 154481 184184 154486 184240
rect 154542 184184 316038 184240
rect 316094 184184 371238 184240
rect 371294 184184 371299 184240
rect 154481 184182 371299 184184
rect 154481 184179 154547 184182
rect 316033 184179 316099 184182
rect 371233 184179 371299 184182
rect 103421 183698 103487 183701
rect 192477 183698 192543 183701
rect 103421 183696 192543 183698
rect 103421 183640 103426 183696
rect 103482 183640 192482 183696
rect 192538 183640 192543 183696
rect 103421 183638 192543 183640
rect 103421 183635 103487 183638
rect 192477 183635 192543 183638
rect 195421 183154 195487 183157
rect 240317 183154 240383 183157
rect 195421 183152 240383 183154
rect 195421 183096 195426 183152
rect 195482 183096 240322 183152
rect 240378 183096 240383 183152
rect 195421 183094 240383 183096
rect 195421 183091 195487 183094
rect 240317 183091 240383 183094
rect 269849 183154 269915 183157
rect 280470 183154 280476 183156
rect 269849 183152 280476 183154
rect 269849 183096 269854 183152
rect 269910 183096 280476 183152
rect 269849 183094 280476 183096
rect 269849 183091 269915 183094
rect 280470 183092 280476 183094
rect 280540 183092 280546 183156
rect 186998 182956 187004 183020
rect 187068 183018 187074 183020
rect 196709 183018 196775 183021
rect 187068 183016 196775 183018
rect 187068 182960 196714 183016
rect 196770 182960 196775 183016
rect 187068 182958 196775 182960
rect 187068 182956 187074 182958
rect 196709 182955 196775 182958
rect 220077 183018 220143 183021
rect 279233 183018 279299 183021
rect 220077 183016 279299 183018
rect 220077 182960 220082 183016
rect 220138 182960 279238 183016
rect 279294 182960 279299 183016
rect 220077 182958 279299 182960
rect 220077 182955 220143 182958
rect 279233 182955 279299 182958
rect 279509 183018 279575 183021
rect 288566 183018 288572 183020
rect 279509 183016 288572 183018
rect 279509 182960 279514 183016
rect 279570 182960 288572 183016
rect 279509 182958 288572 182960
rect 279509 182955 279575 182958
rect 288566 182956 288572 182958
rect 288636 182956 288642 183020
rect 159909 182882 159975 182885
rect 360285 182882 360351 182885
rect 159909 182880 360351 182882
rect 159909 182824 159914 182880
rect 159970 182824 360290 182880
rect 360346 182824 360351 182880
rect 159909 182822 360351 182824
rect 159909 182819 159975 182822
rect 360285 182819 360351 182822
rect 115841 182338 115907 182341
rect 180149 182338 180215 182341
rect 115841 182336 180215 182338
rect 115841 182280 115846 182336
rect 115902 182280 180154 182336
rect 180210 182280 180215 182336
rect 115841 182278 180215 182280
rect 115841 182275 115907 182278
rect 180149 182275 180215 182278
rect 99465 182202 99531 182205
rect 167637 182202 167703 182205
rect 99465 182200 167703 182202
rect 99465 182144 99470 182200
rect 99526 182144 167642 182200
rect 167698 182144 167703 182200
rect 99465 182142 167703 182144
rect 99465 182139 99531 182142
rect 167637 182139 167703 182142
rect 280889 182066 280955 182069
rect 283005 182066 283071 182069
rect 280889 182064 283071 182066
rect 280889 182008 280894 182064
rect 280950 182008 283010 182064
rect 283066 182008 283071 182064
rect 280889 182006 283071 182008
rect 280889 182003 280955 182006
rect 283005 182003 283071 182006
rect 222837 181658 222903 181661
rect 234705 181658 234771 181661
rect 222837 181656 234771 181658
rect 222837 181600 222842 181656
rect 222898 181600 234710 181656
rect 234766 181600 234771 181656
rect 222837 181598 234771 181600
rect 222837 181595 222903 181598
rect 234705 181595 234771 181598
rect 204161 181522 204227 181525
rect 280286 181522 280292 181524
rect 204161 181520 280292 181522
rect 204161 181464 204166 181520
rect 204222 181464 280292 181520
rect 204161 181462 280292 181464
rect 204161 181459 204227 181462
rect 280286 181460 280292 181462
rect 280356 181460 280362 181524
rect 210417 181386 210483 181389
rect 294137 181386 294203 181389
rect 210417 181384 294203 181386
rect 210417 181328 210422 181384
rect 210478 181328 294142 181384
rect 294198 181328 294203 181384
rect 210417 181326 294203 181328
rect 210417 181323 210483 181326
rect 294137 181323 294203 181326
rect 224902 181188 224908 181252
rect 224972 181250 224978 181252
rect 229001 181250 229067 181253
rect 224972 181248 229067 181250
rect 224972 181192 229006 181248
rect 229062 181192 229067 181248
rect 224972 181190 229067 181192
rect 224972 181188 224978 181190
rect 229001 181187 229067 181190
rect 98453 180978 98519 180981
rect 184565 180978 184631 180981
rect 98453 180976 184631 180978
rect 98453 180920 98458 180976
rect 98514 180920 184570 180976
rect 184626 180920 184631 180976
rect 98453 180918 184631 180920
rect 98453 180915 98519 180918
rect 184565 180915 184631 180918
rect 100753 180842 100819 180845
rect 188521 180842 188587 180845
rect 100753 180840 188587 180842
rect 100753 180784 100758 180840
rect 100814 180784 188526 180840
rect 188582 180784 188587 180840
rect 100753 180782 188587 180784
rect 100753 180779 100819 180782
rect 188521 180779 188587 180782
rect 183461 180706 183527 180709
rect 226241 180706 226307 180709
rect 183461 180704 226307 180706
rect 183461 180648 183466 180704
rect 183522 180648 226246 180704
rect 226302 180648 226307 180704
rect 183461 180646 226307 180648
rect 183461 180643 183527 180646
rect 226241 180643 226307 180646
rect 226926 180236 226932 180300
rect 226996 180298 227002 180300
rect 234797 180298 234863 180301
rect 226996 180296 234863 180298
rect 226996 180240 234802 180296
rect 234858 180240 234863 180296
rect 226996 180238 234863 180240
rect 226996 180236 227002 180238
rect 234797 180235 234863 180238
rect 273989 180298 274055 180301
rect 287094 180298 287100 180300
rect 273989 180296 287100 180298
rect 273989 180240 273994 180296
rect 274050 180240 287100 180296
rect 273989 180238 287100 180240
rect 273989 180235 274055 180238
rect 287094 180236 287100 180238
rect 287164 180236 287170 180300
rect 224718 180100 224724 180164
rect 224788 180162 224794 180164
rect 235993 180162 236059 180165
rect 224788 180160 236059 180162
rect 224788 180104 235998 180160
rect 236054 180104 236059 180160
rect 224788 180102 236059 180104
rect 224788 180100 224794 180102
rect 235993 180099 236059 180102
rect 237966 180100 237972 180164
rect 238036 180162 238042 180164
rect 242249 180162 242315 180165
rect 238036 180160 242315 180162
rect 238036 180104 242254 180160
rect 242310 180104 242315 180160
rect 238036 180102 242315 180104
rect 238036 180100 238042 180102
rect 242249 180099 242315 180102
rect 268469 180162 268535 180165
rect 290590 180162 290596 180164
rect 268469 180160 290596 180162
rect 268469 180104 268474 180160
rect 268530 180104 290596 180160
rect 268469 180102 290596 180104
rect 268469 180099 268535 180102
rect 290590 180100 290596 180102
rect 290660 180100 290666 180164
rect 184381 180026 184447 180029
rect 273253 180026 273319 180029
rect 184381 180024 273319 180026
rect 184381 179968 184386 180024
rect 184442 179968 273258 180024
rect 273314 179968 273319 180024
rect 184381 179966 273319 179968
rect 184381 179963 184447 179966
rect 273253 179963 273319 179966
rect 114369 179618 114435 179621
rect 166441 179618 166507 179621
rect 114369 179616 166507 179618
rect 114369 179560 114374 179616
rect 114430 179560 166446 179616
rect 166502 179560 166507 179616
rect 114369 179558 166507 179560
rect 114369 179555 114435 179558
rect 166441 179555 166507 179558
rect 97349 179482 97415 179485
rect 166257 179482 166323 179485
rect 97349 179480 166323 179482
rect 97349 179424 97354 179480
rect 97410 179424 166262 179480
rect 166318 179424 166323 179480
rect 97349 179422 166323 179424
rect 97349 179419 97415 179422
rect 166257 179419 166323 179422
rect 580257 179210 580323 179213
rect 583520 179210 584960 179300
rect 580257 179208 584960 179210
rect 580257 179152 580262 179208
rect 580318 179152 584960 179208
rect 580257 179150 584960 179152
rect 580257 179147 580323 179150
rect 583520 179060 584960 179150
rect 226977 178938 227043 178941
rect 229185 178938 229251 178941
rect 226977 178936 229251 178938
rect 226977 178880 226982 178936
rect 227038 178880 229190 178936
rect 229246 178880 229251 178936
rect 226977 178878 229251 178880
rect 226977 178875 227043 178878
rect 229185 178875 229251 178878
rect 276013 178938 276079 178941
rect 281901 178938 281967 178941
rect 276013 178936 281967 178938
rect 276013 178880 276018 178936
rect 276074 178880 281906 178936
rect 281962 178880 281967 178936
rect 276013 178878 281967 178880
rect 276013 178875 276079 178878
rect 281901 178875 281967 178878
rect 194501 178802 194567 178805
rect 241646 178802 241652 178804
rect 194501 178800 241652 178802
rect 194501 178744 194506 178800
rect 194562 178744 241652 178800
rect 194501 178742 241652 178744
rect 194501 178739 194567 178742
rect 241646 178740 241652 178742
rect 241716 178740 241722 178804
rect 271137 178802 271203 178805
rect 284334 178802 284340 178804
rect 271137 178800 284340 178802
rect 271137 178744 271142 178800
rect 271198 178744 284340 178800
rect 271137 178742 284340 178744
rect 271137 178739 271203 178742
rect 284334 178740 284340 178742
rect 284404 178740 284410 178804
rect 213821 178666 213887 178669
rect 227713 178666 227779 178669
rect 213821 178664 227779 178666
rect 213821 178608 213826 178664
rect 213882 178608 227718 178664
rect 227774 178608 227779 178664
rect 213821 178606 227779 178608
rect 213821 178603 213887 178606
rect 227713 178603 227779 178606
rect 228766 178604 228772 178668
rect 228836 178666 228842 178668
rect 278998 178666 279004 178668
rect 228836 178606 279004 178666
rect 228836 178604 228842 178606
rect 278998 178604 279004 178606
rect 279068 178604 279074 178668
rect 164877 178394 164943 178397
rect 110646 178392 164943 178394
rect 110646 178336 164882 178392
rect 164938 178336 164943 178392
rect 110646 178334 164943 178336
rect 110646 177988 110706 178334
rect 164877 178331 164943 178334
rect 116894 178196 116900 178260
rect 116964 178258 116970 178260
rect 171777 178258 171843 178261
rect 116964 178256 171843 178258
rect 116964 178200 171782 178256
rect 171838 178200 171843 178256
rect 116964 178198 171843 178200
rect 116964 178196 116970 178198
rect 171777 178195 171843 178198
rect 207749 178122 207815 178125
rect 110830 178120 207815 178122
rect 110830 178064 207754 178120
rect 207810 178064 207815 178120
rect 110830 178062 207815 178064
rect 110638 177924 110644 177988
rect 110708 177924 110714 177988
rect 109534 177788 109540 177852
rect 109604 177850 109610 177852
rect 110830 177850 110890 178062
rect 207749 178059 207815 178062
rect 109604 177790 110890 177850
rect 109604 177788 109610 177790
rect 98310 177516 98316 177580
rect 98380 177578 98386 177580
rect 98453 177578 98519 177581
rect 100753 177580 100819 177581
rect 100702 177578 100708 177580
rect 98380 177576 98519 177578
rect 98380 177520 98458 177576
rect 98514 177520 98519 177576
rect 98380 177518 98519 177520
rect 100662 177518 100708 177578
rect 100772 177576 100819 177580
rect 100814 177520 100819 177576
rect 98380 177516 98386 177518
rect 98453 177515 98519 177518
rect 100702 177516 100708 177518
rect 100772 177516 100819 177520
rect 105670 177516 105676 177580
rect 105740 177578 105746 177580
rect 105905 177578 105971 177581
rect 105740 177576 105971 177578
rect 105740 177520 105910 177576
rect 105966 177520 105971 177576
rect 105740 177518 105971 177520
rect 105740 177516 105746 177518
rect 100753 177515 100819 177516
rect 105905 177515 105971 177518
rect 106958 177516 106964 177580
rect 107028 177578 107034 177580
rect 107561 177578 107627 177581
rect 107028 177576 107627 177578
rect 107028 177520 107566 177576
rect 107622 177520 107627 177576
rect 107028 177518 107627 177520
rect 107028 177516 107034 177518
rect 107561 177515 107627 177518
rect 113214 177516 113220 177580
rect 113284 177578 113290 177580
rect 114185 177578 114251 177581
rect 115841 177580 115907 177581
rect 115790 177578 115796 177580
rect 113284 177576 114251 177578
rect 113284 177520 114190 177576
rect 114246 177520 114251 177576
rect 113284 177518 114251 177520
rect 115750 177518 115796 177578
rect 115860 177576 115907 177580
rect 115902 177520 115907 177576
rect 113284 177516 113290 177518
rect 114185 177515 114251 177518
rect 115790 177516 115796 177518
rect 115860 177516 115907 177520
rect 118366 177516 118372 177580
rect 118436 177578 118442 177580
rect 118601 177578 118667 177581
rect 121913 177580 121979 177581
rect 121862 177578 121868 177580
rect 118436 177576 118667 177578
rect 118436 177520 118606 177576
rect 118662 177520 118667 177576
rect 118436 177518 118667 177520
rect 121822 177518 121868 177578
rect 121932 177576 121979 177580
rect 121974 177520 121979 177576
rect 118436 177516 118442 177518
rect 115841 177515 115907 177516
rect 118601 177515 118667 177518
rect 121862 177516 121868 177518
rect 121932 177516 121979 177520
rect 124438 177516 124444 177580
rect 124508 177578 124514 177580
rect 125501 177578 125567 177581
rect 124508 177576 125567 177578
rect 124508 177520 125506 177576
rect 125562 177520 125567 177576
rect 124508 177518 125567 177520
rect 124508 177516 124514 177518
rect 121913 177515 121979 177516
rect 125501 177515 125567 177518
rect 127014 177516 127020 177580
rect 127084 177578 127090 177580
rect 127985 177578 128051 177581
rect 132401 177580 132467 177581
rect 132350 177578 132356 177580
rect 127084 177576 128051 177578
rect 127084 177520 127990 177576
rect 128046 177520 128051 177576
rect 127084 177518 128051 177520
rect 132310 177518 132356 177578
rect 132420 177576 132467 177580
rect 132462 177520 132467 177576
rect 127084 177516 127090 177518
rect 127985 177515 128051 177518
rect 132350 177516 132356 177518
rect 132420 177516 132467 177520
rect 133086 177516 133092 177580
rect 133156 177578 133162 177580
rect 133781 177578 133847 177581
rect 133156 177576 133847 177578
rect 133156 177520 133786 177576
rect 133842 177520 133847 177576
rect 133156 177518 133847 177520
rect 133156 177516 133162 177518
rect 132401 177515 132467 177516
rect 133781 177515 133847 177518
rect 189717 177442 189783 177445
rect 226517 177442 226583 177445
rect 189717 177440 226583 177442
rect 189717 177384 189722 177440
rect 189778 177384 226522 177440
rect 226578 177384 226583 177440
rect 189717 177382 226583 177384
rect 189717 177379 189783 177382
rect 226517 177379 226583 177382
rect 227713 177442 227779 177445
rect 240409 177442 240475 177445
rect 227713 177440 240475 177442
rect 227713 177384 227718 177440
rect 227774 177384 240414 177440
rect 240470 177384 240475 177440
rect 227713 177382 240475 177384
rect 227713 177379 227779 177382
rect 240409 177379 240475 177382
rect 276749 177442 276815 177445
rect 283782 177442 283788 177444
rect 276749 177440 283788 177442
rect 276749 177384 276754 177440
rect 276810 177384 283788 177440
rect 276749 177382 283788 177384
rect 276749 177379 276815 177382
rect 283782 177380 283788 177382
rect 283852 177380 283858 177444
rect 192661 177306 192727 177309
rect 240542 177306 240548 177308
rect 192661 177304 240548 177306
rect 192661 177248 192666 177304
rect 192722 177248 240548 177304
rect 192661 177246 240548 177248
rect 192661 177243 192727 177246
rect 240542 177244 240548 177246
rect 240612 177244 240618 177308
rect 255814 177244 255820 177308
rect 255884 177306 255890 177308
rect 264973 177306 265039 177309
rect 255884 177304 265039 177306
rect 255884 177248 264978 177304
rect 265034 177248 265039 177304
rect 255884 177246 265039 177248
rect 255884 177244 255890 177246
rect 264973 177243 265039 177246
rect 273253 177306 273319 177309
rect 279366 177306 279372 177308
rect 273253 177304 279372 177306
rect 273253 177248 273258 177304
rect 273314 177248 279372 177304
rect 273253 177246 279372 177248
rect 273253 177243 273319 177246
rect 279366 177244 279372 177246
rect 279436 177244 279442 177308
rect 112110 177108 112116 177172
rect 112180 177170 112186 177172
rect 113081 177170 113147 177173
rect 114369 177172 114435 177173
rect 114318 177170 114324 177172
rect 112180 177168 113147 177170
rect 112180 177112 113086 177168
rect 113142 177112 113147 177168
rect 112180 177110 113147 177112
rect 114278 177110 114324 177170
rect 114388 177168 114435 177172
rect 114430 177112 114435 177168
rect 112180 177108 112186 177110
rect 113081 177107 113147 177110
rect 114318 177108 114324 177110
rect 114388 177108 114435 177112
rect 119470 177108 119476 177172
rect 119540 177170 119546 177172
rect 119889 177170 119955 177173
rect 119540 177168 119955 177170
rect 119540 177112 119894 177168
rect 119950 177112 119955 177168
rect 119540 177110 119955 177112
rect 119540 177108 119546 177110
rect 114369 177107 114435 177108
rect 119889 177107 119955 177110
rect 134374 177108 134380 177172
rect 134444 177170 134450 177172
rect 134793 177170 134859 177173
rect 134444 177168 134859 177170
rect 134444 177112 134798 177168
rect 134854 177112 134859 177168
rect 134444 177110 134859 177112
rect 134444 177108 134450 177110
rect 134793 177107 134859 177110
rect 104566 176972 104572 177036
rect 104636 177034 104642 177036
rect 195421 177034 195487 177037
rect 104636 177032 195487 177034
rect 104636 176976 195426 177032
rect 195482 176976 195487 177032
rect 104636 176974 195487 176976
rect 104636 176972 104642 176974
rect 195421 176971 195487 176974
rect 229134 176972 229140 177036
rect 229204 177034 229210 177036
rect 229369 177034 229435 177037
rect 229204 177032 229435 177034
rect 229204 176976 229374 177032
rect 229430 176976 229435 177032
rect 229204 176974 229435 176976
rect 229204 176972 229210 176974
rect 229369 176971 229435 176974
rect 97022 176836 97028 176900
rect 97092 176898 97098 176900
rect 97349 176898 97415 176901
rect 97092 176896 97415 176898
rect 97092 176840 97354 176896
rect 97410 176840 97415 176896
rect 97092 176838 97415 176840
rect 97092 176836 97098 176838
rect 97349 176835 97415 176838
rect 101990 176836 101996 176900
rect 102060 176898 102066 176900
rect 169017 176898 169083 176901
rect 102060 176896 169083 176898
rect 102060 176840 169022 176896
rect 169078 176840 169083 176896
rect 102060 176838 169083 176840
rect 102060 176836 102066 176838
rect 169017 176835 169083 176838
rect 224861 176898 224927 176901
rect 230606 176898 230612 176900
rect 224861 176896 230612 176898
rect 224861 176840 224866 176896
rect 224922 176840 230612 176896
rect 224861 176838 230612 176840
rect 224861 176835 224927 176838
rect 230606 176836 230612 176838
rect 230676 176836 230682 176900
rect 285029 176898 285095 176901
rect 285806 176898 285812 176900
rect 285029 176896 285812 176898
rect 285029 176840 285034 176896
rect 285090 176840 285812 176896
rect 285029 176838 285812 176840
rect 285029 176835 285095 176838
rect 285806 176836 285812 176838
rect 285876 176836 285882 176900
rect 99465 176762 99531 176765
rect 103421 176762 103487 176765
rect 99422 176760 99531 176762
rect 99422 176704 99470 176760
rect 99526 176704 99531 176760
rect 99422 176699 99531 176704
rect 103286 176760 103487 176762
rect 103286 176704 103426 176760
rect 103482 176704 103487 176760
rect 103286 176702 103487 176704
rect 99422 176492 99482 176699
rect 103286 176492 103346 176702
rect 103421 176699 103487 176702
rect 123150 176700 123156 176764
rect 123220 176762 123226 176764
rect 123293 176762 123359 176765
rect 123220 176760 123359 176762
rect 123220 176704 123298 176760
rect 123354 176704 123359 176760
rect 123220 176702 123359 176704
rect 123220 176700 123226 176702
rect 123293 176699 123359 176702
rect 125726 176700 125732 176764
rect 125796 176762 125802 176764
rect 126789 176762 126855 176765
rect 129457 176764 129523 176765
rect 148225 176764 148291 176765
rect 129406 176762 129412 176764
rect 125796 176760 126855 176762
rect 125796 176704 126794 176760
rect 126850 176704 126855 176760
rect 125796 176702 126855 176704
rect 129366 176702 129412 176762
rect 129476 176760 129523 176764
rect 148174 176762 148180 176764
rect 129518 176704 129523 176760
rect 125796 176700 125802 176702
rect 126789 176699 126855 176702
rect 129406 176700 129412 176702
rect 129476 176700 129523 176704
rect 148134 176702 148180 176762
rect 148244 176760 148291 176764
rect 148286 176704 148291 176760
rect 148174 176700 148180 176702
rect 148244 176700 148291 176704
rect 158846 176700 158852 176764
rect 158916 176762 158922 176764
rect 158989 176762 159055 176765
rect 158916 176760 159055 176762
rect 158916 176704 158994 176760
rect 159050 176704 159055 176760
rect 158916 176702 159055 176704
rect 158916 176700 158922 176702
rect 129457 176699 129523 176700
rect 148225 176699 148291 176700
rect 158989 176699 159055 176702
rect 226333 176762 226399 176765
rect 290089 176762 290155 176765
rect 226333 176760 290155 176762
rect 226333 176704 226338 176760
rect 226394 176704 290094 176760
rect 290150 176704 290155 176760
rect 226333 176702 290155 176704
rect 226333 176699 226399 176702
rect 290089 176699 290155 176702
rect 128169 176492 128235 176493
rect 99414 176428 99420 176492
rect 99484 176428 99490 176492
rect 103278 176428 103284 176492
rect 103348 176428 103354 176492
rect 128118 176490 128124 176492
rect 128078 176430 128124 176490
rect 128188 176488 128235 176492
rect 128230 176432 128235 176488
rect 128118 176428 128124 176430
rect 128188 176428 128235 176432
rect 128169 176427 128235 176428
rect 231301 176082 231367 176085
rect 248689 176082 248755 176085
rect 231301 176080 248755 176082
rect -960 175796 480 176036
rect 231301 176024 231306 176080
rect 231362 176024 248694 176080
rect 248750 176024 248755 176080
rect 231301 176022 248755 176024
rect 231301 176019 231367 176022
rect 248689 176019 248755 176022
rect 171869 175946 171935 175949
rect 244406 175946 244412 175948
rect 171869 175944 244412 175946
rect 171869 175888 171874 175944
rect 171930 175888 244412 175944
rect 171869 175886 244412 175888
rect 171869 175883 171935 175886
rect 244406 175884 244412 175886
rect 244476 175884 244482 175948
rect 229369 175810 229435 175813
rect 236177 175810 236243 175813
rect 229369 175808 236243 175810
rect 229369 175752 229374 175808
rect 229430 175752 236182 175808
rect 236238 175752 236243 175808
rect 229369 175750 236243 175752
rect 229369 175747 229435 175750
rect 236177 175747 236243 175750
rect 130745 175676 130811 175677
rect 135713 175676 135779 175677
rect 130694 175674 130700 175676
rect 130654 175614 130700 175674
rect 130764 175672 130811 175676
rect 135662 175674 135668 175676
rect 130806 175616 130811 175672
rect 130694 175612 130700 175614
rect 130764 175612 130811 175616
rect 135622 175614 135668 175674
rect 135732 175672 135779 175676
rect 135774 175616 135779 175672
rect 135662 175612 135668 175614
rect 135732 175612 135779 175616
rect 130745 175611 130811 175612
rect 135713 175611 135779 175612
rect 213913 175674 213979 175677
rect 230657 175674 230723 175677
rect 213913 175672 217028 175674
rect 213913 175616 213918 175672
rect 213974 175616 217028 175672
rect 213913 175614 217028 175616
rect 228988 175672 230723 175674
rect 228988 175616 230662 175672
rect 230718 175616 230723 175672
rect 228988 175614 230723 175616
rect 213913 175611 213979 175614
rect 230657 175611 230723 175614
rect 264973 175674 265039 175677
rect 264973 175672 268180 175674
rect 264973 175616 264978 175672
rect 265034 175616 268180 175672
rect 264973 175614 268180 175616
rect 264973 175611 265039 175614
rect 120758 175476 120764 175540
rect 120828 175538 120834 175540
rect 166533 175538 166599 175541
rect 281717 175538 281783 175541
rect 120828 175536 166599 175538
rect 120828 175480 166538 175536
rect 166594 175480 166599 175536
rect 120828 175478 166599 175480
rect 279956 175536 281783 175538
rect 279956 175480 281722 175536
rect 281778 175480 281783 175536
rect 279956 175478 281783 175480
rect 120828 175476 120834 175478
rect 166533 175475 166599 175478
rect 281717 175475 281783 175478
rect 108062 175340 108068 175404
rect 108132 175402 108138 175404
rect 170489 175402 170555 175405
rect 108132 175400 170555 175402
rect 108132 175344 170494 175400
rect 170550 175344 170555 175400
rect 108132 175342 170555 175344
rect 108132 175340 108138 175342
rect 170489 175339 170555 175342
rect 168281 175266 168347 175269
rect 214557 175266 214623 175269
rect 231301 175266 231367 175269
rect 168281 175264 214623 175266
rect 168281 175208 168286 175264
rect 168342 175208 214562 175264
rect 214618 175208 214623 175264
rect 168281 175206 214623 175208
rect 228988 175264 231367 175266
rect 228988 175208 231306 175264
rect 231362 175208 231367 175264
rect 228988 175206 231367 175208
rect 168281 175203 168347 175206
rect 214557 175203 214623 175206
rect 231301 175203 231367 175206
rect 236085 175266 236151 175269
rect 236678 175266 236684 175268
rect 236085 175264 236684 175266
rect 236085 175208 236090 175264
rect 236146 175208 236684 175264
rect 236085 175206 236684 175208
rect 236085 175203 236151 175206
rect 236678 175204 236684 175206
rect 236748 175204 236754 175268
rect 240225 175266 240291 175269
rect 241278 175266 241284 175268
rect 240225 175264 241284 175266
rect 240225 175208 240230 175264
rect 240286 175208 241284 175264
rect 240225 175206 241284 175208
rect 240225 175203 240291 175206
rect 241278 175204 241284 175206
rect 241348 175204 241354 175268
rect 265617 175266 265683 175269
rect 265617 175264 268180 175266
rect 265617 175208 265622 175264
rect 265678 175208 268180 175264
rect 265617 175206 268180 175208
rect 265617 175203 265683 175206
rect 279366 175204 279372 175268
rect 279436 175204 279442 175268
rect 235441 175130 235507 175133
rect 236494 175130 236500 175132
rect 235441 175128 236500 175130
rect 235441 175072 235446 175128
rect 235502 175072 236500 175128
rect 235441 175070 236500 175072
rect 235441 175067 235507 175070
rect 236494 175068 236500 175070
rect 236564 175068 236570 175132
rect 213913 174994 213979 174997
rect 213913 174992 217028 174994
rect 213913 174936 213918 174992
rect 213974 174936 217028 174992
rect 213913 174934 217028 174936
rect 213913 174931 213979 174934
rect 264973 174858 265039 174861
rect 264973 174856 268180 174858
rect 264973 174800 264978 174856
rect 265034 174800 268180 174856
rect 264973 174798 268180 174800
rect 264973 174795 265039 174798
rect 232221 174722 232287 174725
rect 228988 174720 232287 174722
rect 228988 174664 232226 174720
rect 232282 174664 232287 174720
rect 279374 174692 279434 175204
rect 228988 174662 232287 174664
rect 232221 174659 232287 174662
rect 258030 174390 268180 174450
rect 214005 174314 214071 174317
rect 240358 174314 240364 174316
rect 214005 174312 217028 174314
rect 214005 174256 214010 174312
rect 214066 174256 217028 174312
rect 214005 174254 217028 174256
rect 228988 174254 240364 174314
rect 214005 174251 214071 174254
rect 240358 174252 240364 174254
rect 240428 174252 240434 174316
rect 257337 174314 257403 174317
rect 258030 174314 258090 174390
rect 257337 174312 258090 174314
rect 257337 174256 257342 174312
rect 257398 174256 258090 174312
rect 257337 174254 258090 174256
rect 257337 174251 257403 174254
rect 265065 174042 265131 174045
rect 282177 174042 282243 174045
rect 265065 174040 268180 174042
rect 265065 173984 265070 174040
rect 265126 173984 268180 174040
rect 265065 173982 268180 173984
rect 279956 174040 282243 174042
rect 279956 173984 282182 174040
rect 282238 173984 282243 174040
rect 279956 173982 282243 173984
rect 265065 173979 265131 173982
rect 282177 173979 282243 173982
rect 242341 173906 242407 173909
rect 247718 173906 247724 173908
rect 242341 173904 247724 173906
rect 242341 173848 242346 173904
rect 242402 173848 247724 173904
rect 242341 173846 247724 173848
rect 242341 173843 242407 173846
rect 247718 173844 247724 173846
rect 247788 173844 247794 173908
rect 229093 173770 229159 173773
rect 228988 173768 229159 173770
rect 228988 173712 229098 173768
rect 229154 173712 229159 173768
rect 228988 173710 229159 173712
rect 229093 173707 229159 173710
rect 279366 173708 279372 173772
rect 279436 173708 279442 173772
rect 214925 173634 214991 173637
rect 264237 173634 264303 173637
rect 214925 173632 217028 173634
rect 214925 173576 214930 173632
rect 214986 173576 217028 173632
rect 214925 173574 217028 173576
rect 264237 173632 268180 173634
rect 264237 173576 264242 173632
rect 264298 173576 268180 173632
rect 264237 173574 268180 173576
rect 214925 173571 214991 173574
rect 264237 173571 264303 173574
rect 260833 173362 260899 173365
rect 228988 173360 260899 173362
rect 228988 173304 260838 173360
rect 260894 173304 260899 173360
rect 228988 173302 260899 173304
rect 260833 173299 260899 173302
rect 279374 173196 279434 173708
rect 213913 172954 213979 172957
rect 213913 172952 217028 172954
rect 213913 172896 213918 172952
rect 213974 172896 217028 172952
rect 213913 172894 217028 172896
rect 213913 172891 213979 172894
rect 244222 172818 244228 172820
rect 228988 172758 244228 172818
rect 244222 172756 244228 172758
rect 244292 172756 244298 172820
rect 257613 172818 257679 172821
rect 268150 172818 268210 173060
rect 257613 172816 268210 172818
rect 257613 172760 257618 172816
rect 257674 172760 268210 172816
rect 257613 172758 268210 172760
rect 257613 172755 257679 172758
rect 264973 172682 265039 172685
rect 264973 172680 268180 172682
rect 264973 172624 264978 172680
rect 265034 172624 268180 172680
rect 264973 172622 268180 172624
rect 264973 172619 265039 172622
rect 282453 172546 282519 172549
rect 279956 172544 282519 172546
rect 279956 172488 282458 172544
rect 282514 172488 282519 172544
rect 279956 172486 282519 172488
rect 282453 172483 282519 172486
rect 230749 172410 230815 172413
rect 228988 172408 230815 172410
rect 228988 172352 230754 172408
rect 230810 172352 230815 172408
rect 228988 172350 230815 172352
rect 230749 172347 230815 172350
rect 280102 172348 280108 172412
rect 280172 172410 280178 172412
rect 280470 172410 280476 172412
rect 280172 172350 280476 172410
rect 280172 172348 280178 172350
rect 280470 172348 280476 172350
rect 280540 172348 280546 172412
rect 213913 172274 213979 172277
rect 265065 172274 265131 172277
rect 279325 172274 279391 172277
rect 213913 172272 217028 172274
rect 213913 172216 213918 172272
rect 213974 172216 217028 172272
rect 213913 172214 217028 172216
rect 265065 172272 268180 172274
rect 265065 172216 265070 172272
rect 265126 172216 268180 172272
rect 265065 172214 268180 172216
rect 279325 172272 279434 172274
rect 279325 172216 279330 172272
rect 279386 172216 279434 172272
rect 213913 172211 213979 172214
rect 265065 172211 265131 172214
rect 279325 172211 279434 172216
rect 231393 171866 231459 171869
rect 228988 171864 231459 171866
rect 228988 171808 231398 171864
rect 231454 171808 231459 171864
rect 228988 171806 231459 171808
rect 231393 171803 231459 171806
rect 164724 171594 165354 171600
rect 167913 171594 167979 171597
rect 164724 171592 167979 171594
rect 164724 171540 167918 171592
rect 165294 171536 167918 171540
rect 167974 171536 167979 171592
rect 165294 171534 167979 171536
rect 167913 171531 167979 171534
rect 214005 171594 214071 171597
rect 250713 171594 250779 171597
rect 268150 171594 268210 171836
rect 279374 171700 279434 172211
rect 214005 171592 217028 171594
rect 214005 171536 214010 171592
rect 214066 171536 217028 171592
rect 214005 171534 217028 171536
rect 250713 171592 268210 171594
rect 250713 171536 250718 171592
rect 250774 171536 268210 171592
rect 250713 171534 268210 171536
rect 214005 171531 214071 171534
rect 250713 171531 250779 171534
rect 231301 171458 231367 171461
rect 228988 171456 231367 171458
rect 228988 171400 231306 171456
rect 231362 171400 231367 171456
rect 228988 171398 231367 171400
rect 231301 171395 231367 171398
rect 264973 171458 265039 171461
rect 264973 171456 268180 171458
rect 264973 171400 264978 171456
rect 265034 171400 268180 171456
rect 264973 171398 268180 171400
rect 264973 171395 265039 171398
rect 233366 171186 233372 171188
rect 230798 171126 233372 171186
rect 213913 171050 213979 171053
rect 213913 171048 217028 171050
rect 213913 170992 213918 171048
rect 213974 170992 217028 171048
rect 213913 170990 217028 170992
rect 213913 170987 213979 170990
rect 230798 170914 230858 171126
rect 233366 171124 233372 171126
rect 233436 171124 233442 171188
rect 265065 171050 265131 171053
rect 265065 171048 268180 171050
rect 265065 170992 265070 171048
rect 265126 170992 268180 171048
rect 265065 170990 268180 170992
rect 265065 170987 265131 170990
rect 282269 170914 282335 170917
rect 228988 170854 230858 170914
rect 279956 170912 282335 170914
rect 279956 170856 282274 170912
rect 282330 170856 282335 170912
rect 279956 170854 282335 170856
rect 282269 170851 282335 170854
rect 279550 170580 279556 170644
rect 279620 170580 279626 170644
rect 231853 170506 231919 170509
rect 228988 170504 231919 170506
rect 228988 170448 231858 170504
rect 231914 170448 231919 170504
rect 228988 170446 231919 170448
rect 231853 170443 231919 170446
rect 265157 170506 265223 170509
rect 265157 170504 268180 170506
rect 265157 170448 265162 170504
rect 265218 170448 268180 170504
rect 265157 170446 268180 170448
rect 265157 170443 265223 170446
rect 185577 170370 185643 170373
rect 214005 170370 214071 170373
rect 240961 170370 241027 170373
rect 249793 170370 249859 170373
rect 185577 170368 200130 170370
rect 185577 170312 185582 170368
rect 185638 170312 200130 170368
rect 185577 170310 200130 170312
rect 185577 170307 185643 170310
rect 200070 170234 200130 170310
rect 214005 170368 217028 170370
rect 214005 170312 214010 170368
rect 214066 170312 217028 170368
rect 214005 170310 217028 170312
rect 240961 170368 249859 170370
rect 240961 170312 240966 170368
rect 241022 170312 249798 170368
rect 249854 170312 249859 170368
rect 240961 170310 249859 170312
rect 214005 170307 214071 170310
rect 240961 170307 241027 170310
rect 249793 170307 249859 170310
rect 214097 170234 214163 170237
rect 200070 170232 214163 170234
rect 200070 170176 214102 170232
rect 214158 170176 214163 170232
rect 279558 170204 279618 170580
rect 200070 170174 214163 170176
rect 214097 170171 214163 170174
rect 264973 170098 265039 170101
rect 264973 170096 268180 170098
rect 264973 170040 264978 170096
rect 265034 170040 268180 170096
rect 264973 170038 268180 170040
rect 264973 170035 265039 170038
rect 230565 169962 230631 169965
rect 228988 169960 230631 169962
rect 228988 169904 230570 169960
rect 230626 169904 230631 169960
rect 228988 169902 230631 169904
rect 230565 169899 230631 169902
rect 213913 169690 213979 169693
rect 264973 169690 265039 169693
rect 213913 169688 217028 169690
rect 213913 169632 213918 169688
rect 213974 169632 217028 169688
rect 213913 169630 217028 169632
rect 264973 169688 268180 169690
rect 264973 169632 264978 169688
rect 265034 169632 268180 169688
rect 264973 169630 268180 169632
rect 213913 169627 213979 169630
rect 264973 169627 265039 169630
rect 230606 169554 230612 169556
rect 228988 169494 230612 169554
rect 230606 169492 230612 169494
rect 230676 169492 230682 169556
rect 282821 169418 282887 169421
rect 279956 169416 282887 169418
rect 279956 169360 282826 169416
rect 282882 169360 282887 169416
rect 279956 169358 282887 169360
rect 282821 169355 282887 169358
rect 265249 169282 265315 169285
rect 265249 169280 268180 169282
rect 265249 169224 265254 169280
rect 265310 169224 268180 169280
rect 265249 169222 268180 169224
rect 265249 169219 265315 169222
rect 214005 169010 214071 169013
rect 230565 169010 230631 169013
rect 214005 169008 217028 169010
rect 214005 168952 214010 169008
rect 214066 168952 217028 169008
rect 214005 168950 217028 168952
rect 228988 169008 230631 169010
rect 228988 168952 230570 169008
rect 230626 168952 230631 169008
rect 228988 168950 230631 168952
rect 214005 168947 214071 168950
rect 230565 168947 230631 168950
rect 265065 168874 265131 168877
rect 265065 168872 268180 168874
rect 265065 168816 265070 168872
rect 265126 168816 268180 168872
rect 265065 168814 268180 168816
rect 265065 168811 265131 168814
rect 280245 168738 280311 168741
rect 279956 168736 280311 168738
rect 279956 168680 280250 168736
rect 280306 168680 280311 168736
rect 279956 168678 280311 168680
rect 280245 168675 280311 168678
rect 231117 168602 231183 168605
rect 228988 168600 231183 168602
rect 228988 168544 231122 168600
rect 231178 168544 231183 168600
rect 228988 168542 231183 168544
rect 231117 168539 231183 168542
rect 253473 168466 253539 168469
rect 253473 168464 268180 168466
rect 253473 168408 253478 168464
rect 253534 168408 268180 168464
rect 253473 168406 268180 168408
rect 253473 168403 253539 168406
rect 213913 168330 213979 168333
rect 213913 168328 217028 168330
rect 213913 168272 213918 168328
rect 213974 168272 217028 168328
rect 213913 168270 217028 168272
rect 213913 168267 213979 168270
rect 231393 168058 231459 168061
rect 228988 168056 231459 168058
rect 228988 168000 231398 168056
rect 231454 168000 231459 168056
rect 228988 167998 231459 168000
rect 231393 167995 231459 167998
rect 265065 167922 265131 167925
rect 282269 167922 282335 167925
rect 265065 167920 268180 167922
rect 265065 167864 265070 167920
rect 265126 167864 268180 167920
rect 265065 167862 268180 167864
rect 279956 167920 282335 167922
rect 279956 167864 282274 167920
rect 282330 167864 282335 167920
rect 279956 167862 282335 167864
rect 265065 167859 265131 167862
rect 282269 167859 282335 167862
rect 214005 167650 214071 167653
rect 231894 167650 231900 167652
rect 214005 167648 217028 167650
rect 214005 167592 214010 167648
rect 214066 167592 217028 167648
rect 214005 167590 217028 167592
rect 228988 167590 231900 167650
rect 214005 167587 214071 167590
rect 231894 167588 231900 167590
rect 231964 167588 231970 167652
rect 254853 167650 254919 167653
rect 265157 167650 265223 167653
rect 254853 167648 265223 167650
rect 254853 167592 254858 167648
rect 254914 167592 265162 167648
rect 265218 167592 265223 167648
rect 254853 167590 265223 167592
rect 254853 167587 254919 167590
rect 265157 167587 265223 167590
rect 264973 167514 265039 167517
rect 264973 167512 268180 167514
rect 264973 167456 264978 167512
rect 265034 167456 268180 167512
rect 264973 167454 268180 167456
rect 264973 167451 265039 167454
rect 230974 167180 230980 167244
rect 231044 167242 231050 167244
rect 231044 167182 234630 167242
rect 231044 167180 231050 167182
rect 231393 167106 231459 167109
rect 228988 167104 231459 167106
rect 228988 167048 231398 167104
rect 231454 167048 231459 167104
rect 228988 167046 231459 167048
rect 234570 167106 234630 167182
rect 236177 167106 236243 167109
rect 234570 167104 236243 167106
rect 234570 167048 236182 167104
rect 236238 167048 236243 167104
rect 234570 167046 236243 167048
rect 231393 167043 231459 167046
rect 236177 167043 236243 167046
rect 260097 167106 260163 167109
rect 287094 167106 287100 167108
rect 260097 167104 268180 167106
rect 260097 167048 260102 167104
rect 260158 167048 268180 167104
rect 260097 167046 268180 167048
rect 279956 167046 287100 167106
rect 260097 167043 260163 167046
rect 287094 167044 287100 167046
rect 287164 167044 287170 167108
rect 213913 166970 213979 166973
rect 213913 166968 217028 166970
rect 213913 166912 213918 166968
rect 213974 166912 217028 166968
rect 213913 166910 217028 166912
rect 213913 166907 213979 166910
rect 231761 166698 231827 166701
rect 228988 166696 231827 166698
rect 228988 166640 231766 166696
rect 231822 166640 231827 166696
rect 228988 166638 231827 166640
rect 231761 166635 231827 166638
rect 265065 166698 265131 166701
rect 265065 166696 268180 166698
rect 265065 166640 265070 166696
rect 265126 166640 268180 166696
rect 265065 166638 268180 166640
rect 265065 166635 265131 166638
rect 214097 166426 214163 166429
rect 235349 166426 235415 166429
rect 244457 166426 244523 166429
rect 265249 166426 265315 166429
rect 280981 166426 281047 166429
rect 214097 166424 217028 166426
rect 214097 166368 214102 166424
rect 214158 166368 217028 166424
rect 214097 166366 217028 166368
rect 235349 166424 244523 166426
rect 235349 166368 235354 166424
rect 235410 166368 244462 166424
rect 244518 166368 244523 166424
rect 235349 166366 244523 166368
rect 214097 166363 214163 166366
rect 235349 166363 235415 166366
rect 244457 166363 244523 166366
rect 258030 166424 265315 166426
rect 258030 166368 265254 166424
rect 265310 166368 265315 166424
rect 258030 166366 265315 166368
rect 279956 166424 281047 166426
rect 279956 166368 280986 166424
rect 281042 166368 281047 166424
rect 279956 166366 281047 166368
rect 239673 166290 239739 166293
rect 258030 166290 258090 166366
rect 265249 166363 265315 166366
rect 280981 166363 281047 166366
rect 239673 166288 258090 166290
rect 239673 166232 239678 166288
rect 239734 166232 258090 166288
rect 239673 166230 258090 166232
rect 264973 166290 265039 166293
rect 264973 166288 268180 166290
rect 264973 166232 264978 166288
rect 265034 166232 268180 166288
rect 264973 166230 268180 166232
rect 239673 166227 239739 166230
rect 264973 166227 265039 166230
rect 229461 166154 229527 166157
rect 228988 166152 229527 166154
rect 228988 166096 229466 166152
rect 229522 166096 229527 166152
rect 228988 166094 229527 166096
rect 229461 166091 229527 166094
rect 265157 165882 265223 165885
rect 580165 165882 580231 165885
rect 583520 165882 584960 165972
rect 265157 165880 268180 165882
rect 265157 165824 265162 165880
rect 265218 165824 268180 165880
rect 265157 165822 268180 165824
rect 580165 165880 584960 165882
rect 580165 165824 580170 165880
rect 580226 165824 584960 165880
rect 580165 165822 584960 165824
rect 265157 165819 265223 165822
rect 580165 165819 580231 165822
rect 214005 165746 214071 165749
rect 238845 165746 238911 165749
rect 214005 165744 217028 165746
rect 214005 165688 214010 165744
rect 214066 165688 217028 165744
rect 214005 165686 217028 165688
rect 228988 165744 238911 165746
rect 228988 165688 238850 165744
rect 238906 165688 238911 165744
rect 583520 165732 584960 165822
rect 228988 165686 238911 165688
rect 214005 165683 214071 165686
rect 238845 165683 238911 165686
rect 282821 165610 282887 165613
rect 279956 165608 282887 165610
rect 279956 165552 282826 165608
rect 282882 165552 282887 165608
rect 279956 165550 282887 165552
rect 282821 165547 282887 165550
rect 265065 165338 265131 165341
rect 265065 165336 268180 165338
rect 265065 165280 265070 165336
rect 265126 165280 268180 165336
rect 265065 165278 268180 165280
rect 265065 165275 265131 165278
rect 231485 165202 231551 165205
rect 228988 165200 231551 165202
rect 228988 165144 231490 165200
rect 231546 165144 231551 165200
rect 228988 165142 231551 165144
rect 231485 165139 231551 165142
rect 213913 165066 213979 165069
rect 265157 165066 265223 165069
rect 213913 165064 217028 165066
rect 213913 165008 213918 165064
rect 213974 165008 217028 165064
rect 213913 165006 217028 165008
rect 258030 165064 265223 165066
rect 258030 165008 265162 165064
rect 265218 165008 265223 165064
rect 258030 165006 265223 165008
rect 213913 165003 213979 165006
rect 232589 164930 232655 164933
rect 258030 164930 258090 165006
rect 265157 165003 265223 165006
rect 232589 164928 258090 164930
rect 232589 164872 232594 164928
rect 232650 164872 258090 164928
rect 232589 164870 258090 164872
rect 264973 164930 265039 164933
rect 281901 164930 281967 164933
rect 264973 164928 268180 164930
rect 264973 164872 264978 164928
rect 265034 164872 268180 164928
rect 264973 164870 268180 164872
rect 279956 164928 281967 164930
rect 279956 164872 281906 164928
rect 281962 164872 281967 164928
rect 279956 164870 281967 164872
rect 232589 164867 232655 164870
rect 264973 164867 265039 164870
rect 281901 164867 281967 164870
rect 232037 164794 232103 164797
rect 228988 164792 232103 164794
rect 228988 164736 232042 164792
rect 232098 164736 232103 164792
rect 228988 164734 232103 164736
rect 232037 164731 232103 164734
rect 265249 164522 265315 164525
rect 265249 164520 268180 164522
rect 265249 164464 265254 164520
rect 265310 164464 268180 164520
rect 265249 164462 268180 164464
rect 265249 164459 265315 164462
rect 214005 164386 214071 164389
rect 233417 164386 233483 164389
rect 214005 164384 217028 164386
rect 214005 164328 214010 164384
rect 214066 164328 217028 164384
rect 214005 164326 217028 164328
rect 228988 164384 233483 164386
rect 228988 164328 233422 164384
rect 233478 164328 233483 164384
rect 228988 164326 233483 164328
rect 214005 164323 214071 164326
rect 233417 164323 233483 164326
rect 264973 164114 265039 164117
rect 282821 164114 282887 164117
rect 264973 164112 268180 164114
rect 264973 164056 264978 164112
rect 265034 164056 268180 164112
rect 264973 164054 268180 164056
rect 279956 164112 282887 164114
rect 279956 164056 282826 164112
rect 282882 164056 282887 164112
rect 279956 164054 282887 164056
rect 264973 164051 265039 164054
rect 282821 164051 282887 164054
rect 231025 163842 231091 163845
rect 228988 163840 231091 163842
rect 228988 163784 231030 163840
rect 231086 163784 231091 163840
rect 228988 163782 231091 163784
rect 231025 163779 231091 163782
rect 213913 163706 213979 163709
rect 265065 163706 265131 163709
rect 213913 163704 217028 163706
rect 213913 163648 213918 163704
rect 213974 163648 217028 163704
rect 213913 163646 217028 163648
rect 265065 163704 268180 163706
rect 265065 163648 265070 163704
rect 265126 163648 268180 163704
rect 265065 163646 268180 163648
rect 213913 163643 213979 163646
rect 265065 163643 265131 163646
rect 240317 163434 240383 163437
rect 228988 163432 240383 163434
rect 228988 163376 240322 163432
rect 240378 163376 240383 163432
rect 228988 163374 240383 163376
rect 240317 163371 240383 163374
rect 265157 163298 265223 163301
rect 281625 163298 281691 163301
rect 265157 163296 268180 163298
rect 265157 163240 265162 163296
rect 265218 163240 268180 163296
rect 265157 163238 268180 163240
rect 279956 163296 281691 163298
rect 279956 163240 281630 163296
rect 281686 163240 281691 163296
rect 279956 163238 281691 163240
rect 265157 163235 265223 163238
rect 281625 163235 281691 163238
rect 214005 163026 214071 163029
rect 214005 163024 217028 163026
rect -960 162890 480 162980
rect 214005 162968 214010 163024
rect 214066 162968 217028 163024
rect 214005 162966 217028 162968
rect 214005 162963 214071 162966
rect 3233 162890 3299 162893
rect 231669 162890 231735 162893
rect -960 162888 3299 162890
rect -960 162832 3238 162888
rect 3294 162832 3299 162888
rect -960 162830 3299 162832
rect 228988 162888 231735 162890
rect 228988 162832 231674 162888
rect 231730 162832 231735 162888
rect 228988 162830 231735 162832
rect -960 162740 480 162830
rect 3233 162827 3299 162830
rect 231669 162827 231735 162830
rect 242249 162890 242315 162893
rect 242249 162888 268180 162890
rect 242249 162832 242254 162888
rect 242310 162832 268180 162888
rect 242249 162830 268180 162832
rect 242249 162827 242315 162830
rect 260373 162754 260439 162757
rect 265249 162754 265315 162757
rect 260373 162752 265315 162754
rect 260373 162696 260378 162752
rect 260434 162696 265254 162752
rect 265310 162696 265315 162752
rect 260373 162694 265315 162696
rect 260373 162691 260439 162694
rect 265249 162691 265315 162694
rect 280153 162618 280219 162621
rect 279956 162616 280219 162618
rect 279956 162560 280158 162616
rect 280214 162560 280219 162616
rect 279956 162558 280219 162560
rect 280153 162555 280219 162558
rect 253933 162482 253999 162485
rect 228988 162480 253999 162482
rect 228988 162424 253938 162480
rect 253994 162424 253999 162480
rect 228988 162422 253999 162424
rect 253933 162419 253999 162422
rect 213913 162346 213979 162349
rect 264973 162346 265039 162349
rect 213913 162344 217028 162346
rect 213913 162288 213918 162344
rect 213974 162288 217028 162344
rect 213913 162286 217028 162288
rect 264973 162344 268180 162346
rect 264973 162288 264978 162344
rect 265034 162288 268180 162344
rect 264973 162286 268180 162288
rect 213913 162283 213979 162286
rect 264973 162283 265039 162286
rect 230933 161938 230999 161941
rect 228988 161936 230999 161938
rect 228988 161880 230938 161936
rect 230994 161880 230999 161936
rect 228988 161878 230999 161880
rect 230933 161875 230999 161878
rect 265065 161938 265131 161941
rect 265065 161936 268180 161938
rect 265065 161880 265070 161936
rect 265126 161880 268180 161936
rect 265065 161878 268180 161880
rect 265065 161875 265131 161878
rect 214005 161802 214071 161805
rect 282821 161802 282887 161805
rect 214005 161800 217028 161802
rect 214005 161744 214010 161800
rect 214066 161744 217028 161800
rect 214005 161742 217028 161744
rect 279956 161800 282887 161802
rect 279956 161744 282826 161800
rect 282882 161744 282887 161800
rect 279956 161742 282887 161744
rect 214005 161739 214071 161742
rect 282821 161739 282887 161742
rect 237414 161530 237420 161532
rect 228988 161470 237420 161530
rect 237414 161468 237420 161470
rect 237484 161468 237490 161532
rect 253197 161530 253263 161533
rect 253197 161528 268180 161530
rect 253197 161472 253202 161528
rect 253258 161472 268180 161528
rect 253197 161470 268180 161472
rect 253197 161467 253263 161470
rect 213913 161122 213979 161125
rect 265065 161122 265131 161125
rect 282821 161122 282887 161125
rect 213913 161120 217028 161122
rect 213913 161064 213918 161120
rect 213974 161064 217028 161120
rect 213913 161062 217028 161064
rect 265065 161120 268180 161122
rect 265065 161064 265070 161120
rect 265126 161064 268180 161120
rect 265065 161062 268180 161064
rect 279956 161120 282887 161122
rect 279956 161064 282826 161120
rect 282882 161064 282887 161120
rect 279956 161062 282887 161064
rect 213913 161059 213979 161062
rect 265065 161059 265131 161062
rect 282821 161059 282887 161062
rect 248505 160986 248571 160989
rect 228988 160984 248571 160986
rect 228988 160928 248510 160984
rect 248566 160928 248571 160984
rect 228988 160926 248571 160928
rect 248505 160923 248571 160926
rect 195421 160714 195487 160717
rect 214097 160714 214163 160717
rect 195421 160712 214163 160714
rect 195421 160656 195426 160712
rect 195482 160656 214102 160712
rect 214158 160656 214163 160712
rect 195421 160654 214163 160656
rect 195421 160651 195487 160654
rect 214097 160651 214163 160654
rect 231209 160578 231275 160581
rect 228988 160576 231275 160578
rect 228988 160520 231214 160576
rect 231270 160520 231275 160576
rect 228988 160518 231275 160520
rect 231209 160515 231275 160518
rect 214005 160442 214071 160445
rect 250437 160442 250503 160445
rect 268150 160442 268210 160684
rect 214005 160440 217028 160442
rect 214005 160384 214010 160440
rect 214066 160384 217028 160440
rect 214005 160382 217028 160384
rect 250437 160440 268210 160442
rect 250437 160384 250442 160440
rect 250498 160384 268210 160440
rect 250437 160382 268210 160384
rect 214005 160379 214071 160382
rect 250437 160379 250503 160382
rect 264973 160306 265039 160309
rect 281717 160306 281783 160309
rect 264973 160304 268180 160306
rect 264973 160248 264978 160304
rect 265034 160248 268180 160304
rect 264973 160246 268180 160248
rect 279956 160304 281783 160306
rect 279956 160248 281722 160304
rect 281778 160248 281783 160304
rect 279956 160246 281783 160248
rect 264973 160243 265039 160246
rect 281717 160243 281783 160246
rect 231761 160034 231827 160037
rect 228988 160032 231827 160034
rect 228988 159976 231766 160032
rect 231822 159976 231827 160032
rect 228988 159974 231827 159976
rect 231761 159971 231827 159974
rect 213913 159762 213979 159765
rect 265065 159762 265131 159765
rect 213913 159760 217028 159762
rect 213913 159704 213918 159760
rect 213974 159704 217028 159760
rect 213913 159702 217028 159704
rect 265065 159760 268180 159762
rect 265065 159704 265070 159760
rect 265126 159704 268180 159760
rect 265065 159702 268180 159704
rect 213913 159699 213979 159702
rect 265065 159699 265131 159702
rect 230974 159626 230980 159628
rect 228988 159566 230980 159626
rect 230974 159564 230980 159566
rect 231044 159564 231050 159628
rect 281901 159490 281967 159493
rect 279956 159488 281967 159490
rect 279956 159432 281906 159488
rect 281962 159432 281967 159488
rect 279956 159430 281967 159432
rect 281901 159427 281967 159430
rect 214097 159082 214163 159085
rect 231393 159082 231459 159085
rect 214097 159080 217028 159082
rect 214097 159024 214102 159080
rect 214158 159024 217028 159080
rect 214097 159022 217028 159024
rect 228988 159080 231459 159082
rect 228988 159024 231398 159080
rect 231454 159024 231459 159080
rect 228988 159022 231459 159024
rect 214097 159019 214163 159022
rect 231393 159019 231459 159022
rect 232497 159082 232563 159085
rect 268150 159082 268210 159324
rect 232497 159080 268210 159082
rect 232497 159024 232502 159080
rect 232558 159024 268210 159080
rect 232497 159022 268210 159024
rect 232497 159019 232563 159022
rect 264973 158946 265039 158949
rect 264973 158944 268180 158946
rect 264973 158888 264978 158944
rect 265034 158888 268180 158944
rect 264973 158886 268180 158888
rect 264973 158883 265039 158886
rect 282361 158810 282427 158813
rect 279956 158808 282427 158810
rect 279956 158752 282366 158808
rect 282422 158752 282427 158808
rect 279956 158750 282427 158752
rect 282361 158747 282427 158750
rect 231669 158674 231735 158677
rect 228988 158672 231735 158674
rect 228988 158616 231674 158672
rect 231730 158616 231735 158672
rect 228988 158614 231735 158616
rect 231669 158611 231735 158614
rect 265065 158538 265131 158541
rect 265065 158536 268180 158538
rect 265065 158480 265070 158536
rect 265126 158480 268180 158536
rect 265065 158478 268180 158480
rect 265065 158475 265131 158478
rect 213913 158402 213979 158405
rect 213913 158400 217028 158402
rect 213913 158344 213918 158400
rect 213974 158344 217028 158400
rect 213913 158342 217028 158344
rect 213913 158339 213979 158342
rect 231209 158130 231275 158133
rect 228988 158128 231275 158130
rect 228988 158072 231214 158128
rect 231270 158072 231275 158128
rect 228988 158070 231275 158072
rect 231209 158067 231275 158070
rect 231577 158130 231643 158133
rect 251265 158130 251331 158133
rect 231577 158128 251331 158130
rect 231577 158072 231582 158128
rect 231638 158072 251270 158128
rect 251326 158072 251331 158128
rect 231577 158070 251331 158072
rect 231577 158067 231643 158070
rect 251265 158067 251331 158070
rect 264973 158130 265039 158133
rect 264973 158128 268180 158130
rect 264973 158072 264978 158128
rect 265034 158072 268180 158128
rect 264973 158070 268180 158072
rect 264973 158067 265039 158070
rect 231669 157994 231735 157997
rect 260189 157994 260255 157997
rect 282821 157994 282887 157997
rect 231669 157992 260255 157994
rect 231669 157936 231674 157992
rect 231730 157936 260194 157992
rect 260250 157936 260255 157992
rect 231669 157934 260255 157936
rect 279956 157992 282887 157994
rect 279956 157936 282826 157992
rect 282882 157936 282887 157992
rect 279956 157934 282887 157936
rect 231669 157931 231735 157934
rect 260189 157931 260255 157934
rect 282821 157931 282887 157934
rect 214005 157722 214071 157725
rect 230841 157722 230907 157725
rect 214005 157720 217028 157722
rect 214005 157664 214010 157720
rect 214066 157664 217028 157720
rect 214005 157662 217028 157664
rect 228988 157720 230907 157722
rect 228988 157664 230846 157720
rect 230902 157664 230907 157720
rect 228988 157662 230907 157664
rect 214005 157659 214071 157662
rect 230841 157659 230907 157662
rect 265341 157722 265407 157725
rect 265341 157720 268180 157722
rect 265341 157664 265346 157720
rect 265402 157664 268180 157720
rect 265341 157662 268180 157664
rect 265341 157659 265407 157662
rect 264329 157450 264395 157453
rect 265157 157450 265223 157453
rect 264329 157448 265223 157450
rect 264329 157392 264334 157448
rect 264390 157392 265162 157448
rect 265218 157392 265223 157448
rect 264329 157390 265223 157392
rect 264329 157387 264395 157390
rect 265157 157387 265223 157390
rect 281758 157314 281764 157316
rect 279956 157254 281764 157314
rect 281758 157252 281764 157254
rect 281828 157252 281834 157316
rect 213913 157178 213979 157181
rect 231669 157178 231735 157181
rect 213913 157176 217028 157178
rect 213913 157120 213918 157176
rect 213974 157120 217028 157176
rect 213913 157118 217028 157120
rect 228988 157176 231735 157178
rect 228988 157120 231674 157176
rect 231730 157120 231735 157176
rect 228988 157118 231735 157120
rect 213913 157115 213979 157118
rect 231669 157115 231735 157118
rect 265065 157178 265131 157181
rect 265065 157176 268180 157178
rect 265065 157120 265070 157176
rect 265126 157120 268180 157176
rect 265065 157118 268180 157120
rect 265065 157115 265131 157118
rect 231761 156770 231827 156773
rect 228988 156768 231827 156770
rect 228988 156712 231766 156768
rect 231822 156712 231827 156768
rect 228988 156710 231827 156712
rect 231761 156707 231827 156710
rect 230381 156634 230447 156637
rect 239254 156634 239260 156636
rect 230381 156632 239260 156634
rect 230381 156576 230386 156632
rect 230442 156576 239260 156632
rect 230381 156574 239260 156576
rect 230381 156571 230447 156574
rect 239254 156572 239260 156574
rect 239324 156572 239330 156636
rect 214005 156498 214071 156501
rect 251909 156498 251975 156501
rect 268150 156498 268210 156740
rect 281574 156498 281580 156500
rect 214005 156496 217028 156498
rect 214005 156440 214010 156496
rect 214066 156440 217028 156496
rect 214005 156438 217028 156440
rect 251909 156496 268210 156498
rect 251909 156440 251914 156496
rect 251970 156440 268210 156496
rect 251909 156438 268210 156440
rect 279956 156438 281580 156498
rect 214005 156435 214071 156438
rect 251909 156435 251975 156438
rect 281574 156436 281580 156438
rect 281644 156436 281650 156500
rect 264973 156362 265039 156365
rect 264973 156360 268180 156362
rect 264973 156304 264978 156360
rect 265034 156304 268180 156360
rect 264973 156302 268180 156304
rect 264973 156299 265039 156302
rect 231761 156226 231827 156229
rect 228988 156224 231827 156226
rect 228988 156168 231766 156224
rect 231822 156168 231827 156224
rect 228988 156166 231827 156168
rect 231761 156163 231827 156166
rect 265157 155954 265223 155957
rect 279325 155954 279391 155957
rect 265157 155952 268180 155954
rect 265157 155896 265162 155952
rect 265218 155896 268180 155952
rect 265157 155894 268180 155896
rect 279325 155952 279434 155954
rect 279325 155896 279330 155952
rect 279386 155896 279434 155952
rect 265157 155891 265223 155894
rect 279325 155891 279434 155896
rect 213913 155818 213979 155821
rect 229185 155818 229251 155821
rect 213913 155816 217028 155818
rect 213913 155760 213918 155816
rect 213974 155760 217028 155816
rect 213913 155758 217028 155760
rect 228988 155816 229251 155818
rect 228988 155760 229190 155816
rect 229246 155760 229251 155816
rect 228988 155758 229251 155760
rect 213913 155755 213979 155758
rect 229185 155755 229251 155758
rect 279374 155652 279434 155891
rect 231485 155274 231551 155277
rect 228988 155272 231551 155274
rect 228988 155216 231490 155272
rect 231546 155216 231551 155272
rect 228988 155214 231551 155216
rect 231485 155211 231551 155214
rect 260281 155274 260347 155277
rect 268150 155274 268210 155516
rect 260281 155272 268210 155274
rect 260281 155216 260286 155272
rect 260342 155216 268210 155272
rect 260281 155214 268210 155216
rect 260281 155211 260347 155214
rect 214005 155138 214071 155141
rect 214005 155136 217028 155138
rect 214005 155080 214010 155136
rect 214066 155080 217028 155136
rect 214005 155078 217028 155080
rect 258030 155078 268180 155138
rect 214005 155075 214071 155078
rect 233969 155002 234035 155005
rect 258030 155002 258090 155078
rect 281625 155002 281691 155005
rect 233969 155000 258090 155002
rect 233969 154944 233974 155000
rect 234030 154944 258090 155000
rect 233969 154942 258090 154944
rect 279956 155000 281691 155002
rect 279956 154944 281630 155000
rect 281686 154944 281691 155000
rect 279956 154942 281691 154944
rect 233969 154939 234035 154942
rect 281625 154939 281691 154942
rect 234654 154866 234660 154868
rect 228988 154806 234660 154866
rect 234654 154804 234660 154806
rect 234724 154804 234730 154868
rect 264973 154594 265039 154597
rect 264973 154592 268180 154594
rect 264973 154536 264978 154592
rect 265034 154536 268180 154592
rect 264973 154534 268180 154536
rect 264973 154531 265039 154534
rect 214005 154458 214071 154461
rect 214005 154456 217028 154458
rect 214005 154400 214010 154456
rect 214066 154400 217028 154456
rect 214005 154398 217028 154400
rect 214005 154395 214071 154398
rect 231669 154322 231735 154325
rect 228988 154320 231735 154322
rect 228988 154264 231674 154320
rect 231730 154264 231735 154320
rect 228988 154262 231735 154264
rect 231669 154259 231735 154262
rect 265709 154186 265775 154189
rect 281625 154186 281691 154189
rect 265709 154184 268180 154186
rect 265709 154128 265714 154184
rect 265770 154128 268180 154184
rect 265709 154126 268180 154128
rect 279956 154184 281691 154186
rect 279956 154128 281630 154184
rect 281686 154128 281691 154184
rect 279956 154126 281691 154128
rect 265709 154123 265775 154126
rect 281625 154123 281691 154126
rect 231761 153914 231827 153917
rect 228988 153912 231827 153914
rect 228988 153856 231766 153912
rect 231822 153856 231827 153912
rect 228988 153854 231827 153856
rect 231761 153851 231827 153854
rect 213913 153778 213979 153781
rect 234245 153778 234311 153781
rect 247033 153778 247099 153781
rect 213913 153776 217028 153778
rect 213913 153720 213918 153776
rect 213974 153720 217028 153776
rect 213913 153718 217028 153720
rect 234245 153776 247099 153778
rect 234245 153720 234250 153776
rect 234306 153720 247038 153776
rect 247094 153720 247099 153776
rect 234245 153718 247099 153720
rect 213913 153715 213979 153718
rect 234245 153715 234311 153718
rect 247033 153715 247099 153718
rect 265065 153778 265131 153781
rect 282177 153778 282243 153781
rect 289813 153778 289879 153781
rect 265065 153776 268180 153778
rect 265065 153720 265070 153776
rect 265126 153720 268180 153776
rect 265065 153718 268180 153720
rect 282177 153776 289879 153778
rect 282177 153720 282182 153776
rect 282238 153720 289818 153776
rect 289874 153720 289879 153776
rect 282177 153718 289879 153720
rect 265065 153715 265131 153718
rect 282177 153715 282243 153718
rect 289813 153715 289879 153718
rect 283097 153506 283163 153509
rect 279956 153504 283163 153506
rect 279956 153448 283102 153504
rect 283158 153448 283163 153504
rect 279956 153446 283163 153448
rect 283097 153443 283163 153446
rect 231485 153370 231551 153373
rect 228988 153368 231551 153370
rect 228988 153312 231490 153368
rect 231546 153312 231551 153368
rect 228988 153310 231551 153312
rect 231485 153307 231551 153310
rect 264973 153370 265039 153373
rect 264973 153368 268180 153370
rect 264973 153312 264978 153368
rect 265034 153312 268180 153368
rect 264973 153310 268180 153312
rect 264973 153307 265039 153310
rect 214005 153098 214071 153101
rect 230565 153098 230631 153101
rect 233182 153098 233188 153100
rect 214005 153096 217028 153098
rect 214005 153040 214010 153096
rect 214066 153040 217028 153096
rect 214005 153038 217028 153040
rect 230565 153096 233188 153098
rect 230565 153040 230570 153096
rect 230626 153040 233188 153096
rect 230565 153038 233188 153040
rect 214005 153035 214071 153038
rect 230565 153035 230631 153038
rect 233182 153036 233188 153038
rect 233252 153036 233258 153100
rect 231485 152962 231551 152965
rect 228988 152960 231551 152962
rect 228988 152904 231490 152960
rect 231546 152904 231551 152960
rect 228988 152902 231551 152904
rect 231485 152899 231551 152902
rect 264973 152962 265039 152965
rect 264973 152960 268180 152962
rect 264973 152904 264978 152960
rect 265034 152904 268180 152960
rect 264973 152902 268180 152904
rect 264973 152899 265039 152902
rect 281625 152690 281691 152693
rect 279956 152688 281691 152690
rect 279956 152632 281630 152688
rect 281686 152632 281691 152688
rect 279956 152630 281691 152632
rect 281625 152627 281691 152630
rect 583385 152690 583451 152693
rect 583520 152690 584960 152780
rect 583385 152688 584960 152690
rect 583385 152632 583390 152688
rect 583446 152632 584960 152688
rect 583385 152630 584960 152632
rect 583385 152627 583451 152630
rect 214557 152554 214623 152557
rect 240542 152554 240548 152556
rect 214557 152552 217028 152554
rect 214557 152496 214562 152552
rect 214618 152496 217028 152552
rect 214557 152494 217028 152496
rect 228988 152494 240548 152554
rect 214557 152491 214623 152494
rect 240542 152492 240548 152494
rect 240612 152492 240618 152556
rect 265249 152554 265315 152557
rect 265249 152552 268180 152554
rect 265249 152496 265254 152552
rect 265310 152496 268180 152552
rect 583520 152540 584960 152630
rect 265249 152494 268180 152496
rect 265249 152491 265315 152494
rect 172094 152356 172100 152420
rect 172164 152418 172170 152420
rect 193949 152418 194015 152421
rect 172164 152416 194015 152418
rect 172164 152360 193954 152416
rect 194010 152360 194015 152416
rect 172164 152358 194015 152360
rect 172164 152356 172170 152358
rect 193949 152355 194015 152358
rect 231577 152010 231643 152013
rect 228988 152008 231643 152010
rect 228988 151952 231582 152008
rect 231638 151952 231643 152008
rect 228988 151950 231643 151952
rect 231577 151947 231643 151950
rect 258717 152010 258783 152013
rect 258717 152008 268180 152010
rect 258717 151952 258722 152008
rect 258778 151952 268180 152008
rect 258717 151950 268180 151952
rect 258717 151947 258783 151950
rect 213177 151874 213243 151877
rect 281717 151874 281783 151877
rect 213177 151872 217028 151874
rect 213177 151816 213182 151872
rect 213238 151816 217028 151872
rect 213177 151814 217028 151816
rect 279956 151872 281783 151874
rect 279956 151816 281722 151872
rect 281778 151816 281783 151872
rect 279956 151814 281783 151816
rect 213177 151811 213243 151814
rect 281717 151811 281783 151814
rect 230565 151602 230631 151605
rect 228988 151600 230631 151602
rect 228988 151544 230570 151600
rect 230626 151544 230631 151600
rect 228988 151542 230631 151544
rect 230565 151539 230631 151542
rect 265065 151602 265131 151605
rect 265065 151600 268180 151602
rect 265065 151544 265070 151600
rect 265126 151544 268180 151600
rect 265065 151542 268180 151544
rect 265065 151539 265131 151542
rect 214005 151194 214071 151197
rect 264973 151194 265039 151197
rect 281625 151194 281691 151197
rect 214005 151192 217028 151194
rect 214005 151136 214010 151192
rect 214066 151136 217028 151192
rect 214005 151134 217028 151136
rect 264973 151192 268180 151194
rect 264973 151136 264978 151192
rect 265034 151136 268180 151192
rect 264973 151134 268180 151136
rect 279956 151192 281691 151194
rect 279956 151136 281630 151192
rect 281686 151136 281691 151192
rect 279956 151134 281691 151136
rect 214005 151131 214071 151134
rect 264973 151131 265039 151134
rect 281625 151131 281691 151134
rect 231485 151058 231551 151061
rect 228988 151056 231551 151058
rect 228988 151000 231490 151056
rect 231546 151000 231551 151056
rect 228988 150998 231551 151000
rect 231485 150995 231551 150998
rect 231761 151058 231827 151061
rect 244406 151058 244412 151060
rect 231761 151056 244412 151058
rect 231761 151000 231766 151056
rect 231822 151000 244412 151056
rect 231761 150998 244412 151000
rect 231761 150995 231827 150998
rect 244406 150996 244412 150998
rect 244476 150996 244482 151060
rect 265249 150786 265315 150789
rect 265249 150784 268180 150786
rect 265249 150728 265254 150784
rect 265310 150728 268180 150784
rect 265249 150726 268180 150728
rect 265249 150723 265315 150726
rect 231669 150650 231735 150653
rect 228988 150648 231735 150650
rect 228988 150592 231674 150648
rect 231730 150592 231735 150648
rect 228988 150590 231735 150592
rect 231669 150587 231735 150590
rect 213913 150514 213979 150517
rect 246297 150514 246363 150517
rect 249742 150514 249748 150516
rect 213913 150512 217028 150514
rect 213913 150456 213918 150512
rect 213974 150456 217028 150512
rect 213913 150454 217028 150456
rect 246297 150512 249748 150514
rect 246297 150456 246302 150512
rect 246358 150456 249748 150512
rect 246297 150454 249748 150456
rect 213913 150451 213979 150454
rect 246297 150451 246363 150454
rect 249742 150452 249748 150454
rect 249812 150452 249818 150516
rect 281625 150378 281691 150381
rect 279956 150376 281691 150378
rect 247718 150106 247724 150108
rect 228988 150046 247724 150106
rect 247718 150044 247724 150046
rect 247788 150044 247794 150108
rect 268150 150106 268210 150348
rect 279956 150320 281630 150376
rect 281686 150320 281691 150376
rect 279956 150318 281691 150320
rect 281625 150315 281691 150318
rect 258030 150046 268210 150106
rect -960 149834 480 149924
rect 3509 149834 3575 149837
rect -960 149832 3575 149834
rect -960 149776 3514 149832
rect 3570 149776 3575 149832
rect -960 149774 3575 149776
rect -960 149684 480 149774
rect 3509 149771 3575 149774
rect 203609 149290 203675 149293
rect 216998 149290 217058 149804
rect 229134 149698 229140 149700
rect 228988 149638 229140 149698
rect 229134 149636 229140 149638
rect 229204 149636 229210 149700
rect 257521 149698 257587 149701
rect 258030 149698 258090 150046
rect 264973 149970 265039 149973
rect 264973 149968 268180 149970
rect 264973 149912 264978 149968
rect 265034 149912 268180 149968
rect 264973 149910 268180 149912
rect 264973 149907 265039 149910
rect 281717 149698 281783 149701
rect 257521 149696 258090 149698
rect 257521 149640 257526 149696
rect 257582 149640 258090 149696
rect 257521 149638 258090 149640
rect 279956 149696 281783 149698
rect 279956 149640 281722 149696
rect 281778 149640 281783 149696
rect 279956 149638 281783 149640
rect 257521 149635 257587 149638
rect 281717 149635 281783 149638
rect 265065 149562 265131 149565
rect 265065 149560 268180 149562
rect 265065 149504 265070 149560
rect 265126 149504 268180 149560
rect 265065 149502 268180 149504
rect 265065 149499 265131 149502
rect 203609 149288 217058 149290
rect 203609 149232 203614 149288
rect 203670 149232 217058 149288
rect 203609 149230 217058 149232
rect 203609 149227 203675 149230
rect 214097 149154 214163 149157
rect 242934 149154 242940 149156
rect 214097 149152 217028 149154
rect 214097 149096 214102 149152
rect 214158 149096 217028 149152
rect 214097 149094 217028 149096
rect 228988 149094 242940 149154
rect 214097 149091 214163 149094
rect 242934 149092 242940 149094
rect 243004 149092 243010 149156
rect 267089 149018 267155 149021
rect 267089 149016 268180 149018
rect 267089 148960 267094 149016
rect 267150 148960 268180 149016
rect 267089 148958 268180 148960
rect 267089 148955 267155 148958
rect 281809 148882 281875 148885
rect 279956 148880 281875 148882
rect 279956 148824 281814 148880
rect 281870 148824 281875 148880
rect 279956 148822 281875 148824
rect 281809 148819 281875 148822
rect 231485 148746 231551 148749
rect 228988 148744 231551 148746
rect 228988 148688 231490 148744
rect 231546 148688 231551 148744
rect 228988 148686 231551 148688
rect 231485 148683 231551 148686
rect 265801 148610 265867 148613
rect 265801 148608 268180 148610
rect 265801 148552 265806 148608
rect 265862 148552 268180 148608
rect 265801 148550 268180 148552
rect 265801 148547 265867 148550
rect 213913 148474 213979 148477
rect 250621 148474 250687 148477
rect 265065 148474 265131 148477
rect 213913 148472 217028 148474
rect 213913 148416 213918 148472
rect 213974 148416 217028 148472
rect 213913 148414 217028 148416
rect 250621 148472 265131 148474
rect 250621 148416 250626 148472
rect 250682 148416 265070 148472
rect 265126 148416 265131 148472
rect 250621 148414 265131 148416
rect 213913 148411 213979 148414
rect 250621 148411 250687 148414
rect 265065 148411 265131 148414
rect 231577 148338 231643 148341
rect 251173 148338 251239 148341
rect 231577 148336 251239 148338
rect 231577 148280 231582 148336
rect 231638 148280 251178 148336
rect 251234 148280 251239 148336
rect 231577 148278 251239 148280
rect 231577 148275 231643 148278
rect 251173 148275 251239 148278
rect 279325 148338 279391 148341
rect 280061 148338 280127 148341
rect 279325 148336 280127 148338
rect 279325 148280 279330 148336
rect 279386 148280 280066 148336
rect 280122 148280 280127 148336
rect 279325 148278 280127 148280
rect 279325 148275 279391 148278
rect 280061 148275 280127 148278
rect 231761 148202 231827 148205
rect 228988 148200 231827 148202
rect 228988 148144 231766 148200
rect 231822 148144 231827 148200
rect 228988 148142 231827 148144
rect 231761 148139 231827 148142
rect 265157 148202 265223 148205
rect 265157 148200 268180 148202
rect 265157 148144 265162 148200
rect 265218 148144 268180 148200
rect 265157 148142 268180 148144
rect 265157 148139 265223 148142
rect 229134 148004 229140 148068
rect 229204 148066 229210 148068
rect 230381 148066 230447 148069
rect 281625 148066 281691 148069
rect 229204 148064 230447 148066
rect 229204 148008 230386 148064
rect 230442 148008 230447 148064
rect 229204 148006 230447 148008
rect 279956 148064 281691 148066
rect 279956 148008 281630 148064
rect 281686 148008 281691 148064
rect 279956 148006 281691 148008
rect 229204 148004 229210 148006
rect 230381 148003 230447 148006
rect 281625 148003 281691 148006
rect 213913 147930 213979 147933
rect 229737 147930 229803 147933
rect 230422 147930 230428 147932
rect 213913 147928 217028 147930
rect 213913 147872 213918 147928
rect 213974 147872 217028 147928
rect 213913 147870 217028 147872
rect 229737 147928 230428 147930
rect 229737 147872 229742 147928
rect 229798 147872 230428 147928
rect 229737 147870 230428 147872
rect 213913 147867 213979 147870
rect 229737 147867 229803 147870
rect 230422 147868 230428 147870
rect 230492 147868 230498 147932
rect 248597 147794 248663 147797
rect 228988 147792 248663 147794
rect 228988 147736 248602 147792
rect 248658 147736 248663 147792
rect 228988 147734 248663 147736
rect 248597 147731 248663 147734
rect 264973 147794 265039 147797
rect 264973 147792 268180 147794
rect 264973 147736 264978 147792
rect 265034 147736 268180 147792
rect 264973 147734 268180 147736
rect 264973 147731 265039 147734
rect 264973 147386 265039 147389
rect 282821 147386 282887 147389
rect 264973 147384 268180 147386
rect 264973 147328 264978 147384
rect 265034 147328 268180 147384
rect 264973 147326 268180 147328
rect 279956 147384 282887 147386
rect 279956 147328 282826 147384
rect 282882 147328 282887 147384
rect 279956 147326 282887 147328
rect 264973 147323 265039 147326
rect 282821 147323 282887 147326
rect 214005 147250 214071 147253
rect 232078 147250 232084 147252
rect 214005 147248 217028 147250
rect 214005 147192 214010 147248
rect 214066 147192 217028 147248
rect 214005 147190 217028 147192
rect 228988 147190 232084 147250
rect 214005 147187 214071 147190
rect 232078 147188 232084 147190
rect 232148 147188 232154 147252
rect 231761 147114 231827 147117
rect 249926 147114 249932 147116
rect 231761 147112 249932 147114
rect 231761 147056 231766 147112
rect 231822 147056 249932 147112
rect 231761 147054 249932 147056
rect 231761 147051 231827 147054
rect 249926 147052 249932 147054
rect 249996 147052 250002 147116
rect 231710 146916 231716 146980
rect 231780 146978 231786 146980
rect 244549 146978 244615 146981
rect 231780 146976 244615 146978
rect 231780 146920 244554 146976
rect 244610 146920 244615 146976
rect 231780 146918 244615 146920
rect 231780 146916 231786 146918
rect 244549 146915 244615 146918
rect 245193 146978 245259 146981
rect 265249 146978 265315 146981
rect 245193 146976 265315 146978
rect 245193 146920 245198 146976
rect 245254 146920 265254 146976
rect 265310 146920 265315 146976
rect 245193 146918 265315 146920
rect 245193 146915 245259 146918
rect 265249 146915 265315 146918
rect 265433 146978 265499 146981
rect 265433 146976 268180 146978
rect 265433 146920 265438 146976
rect 265494 146920 268180 146976
rect 265433 146918 268180 146920
rect 265433 146915 265499 146918
rect 229093 146842 229159 146845
rect 228988 146840 229159 146842
rect 228988 146784 229098 146840
rect 229154 146784 229159 146840
rect 228988 146782 229159 146784
rect 229093 146779 229159 146782
rect 213913 146570 213979 146573
rect 283782 146570 283788 146572
rect 213913 146568 217028 146570
rect 213913 146512 213918 146568
rect 213974 146512 217028 146568
rect 213913 146510 217028 146512
rect 279956 146510 283788 146570
rect 213913 146507 213979 146510
rect 283782 146508 283788 146510
rect 283852 146508 283858 146572
rect 265065 146434 265131 146437
rect 265065 146432 268180 146434
rect 265065 146376 265070 146432
rect 265126 146376 268180 146432
rect 265065 146374 268180 146376
rect 265065 146371 265131 146374
rect 230013 146298 230079 146301
rect 228988 146296 230079 146298
rect 228988 146240 230018 146296
rect 230074 146240 230079 146296
rect 228988 146238 230079 146240
rect 230013 146235 230079 146238
rect 265065 146026 265131 146029
rect 265065 146024 268180 146026
rect 265065 145968 265070 146024
rect 265126 145968 268180 146024
rect 265065 145966 268180 145968
rect 265065 145963 265131 145966
rect 215937 145890 216003 145893
rect 231710 145890 231716 145892
rect 215937 145888 217028 145890
rect 215937 145832 215942 145888
rect 215998 145832 217028 145888
rect 215937 145830 217028 145832
rect 228988 145830 231716 145890
rect 215937 145827 216003 145830
rect 231710 145828 231716 145830
rect 231780 145828 231786 145892
rect 280889 145890 280955 145893
rect 279956 145888 280955 145890
rect 279956 145832 280894 145888
rect 280950 145832 280955 145888
rect 279956 145830 280955 145832
rect 280889 145827 280955 145830
rect 229829 145618 229895 145621
rect 265157 145618 265223 145621
rect 229829 145616 265223 145618
rect 229829 145560 229834 145616
rect 229890 145560 265162 145616
rect 265218 145560 265223 145616
rect 229829 145558 265223 145560
rect 229829 145555 229895 145558
rect 265157 145555 265223 145558
rect 267690 145558 268180 145618
rect 234061 145482 234127 145485
rect 267690 145482 267750 145558
rect 234061 145480 267750 145482
rect 234061 145424 234066 145480
rect 234122 145424 267750 145480
rect 234061 145422 267750 145424
rect 234061 145419 234127 145422
rect 236678 145346 236684 145348
rect 228988 145286 236684 145346
rect 236678 145284 236684 145286
rect 236748 145284 236754 145348
rect 213913 145210 213979 145213
rect 264973 145210 265039 145213
rect 213913 145208 217028 145210
rect 213913 145152 213918 145208
rect 213974 145152 217028 145208
rect 213913 145150 217028 145152
rect 264973 145208 268180 145210
rect 264973 145152 264978 145208
rect 265034 145152 268180 145208
rect 264973 145150 268180 145152
rect 213913 145147 213979 145150
rect 264973 145147 265039 145150
rect 282361 145074 282427 145077
rect 279956 145072 282427 145074
rect 279956 145016 282366 145072
rect 282422 145016 282427 145072
rect 279956 145014 282427 145016
rect 282361 145011 282427 145014
rect 231669 144938 231735 144941
rect 228988 144936 231735 144938
rect 228988 144880 231674 144936
rect 231730 144880 231735 144936
rect 228988 144878 231735 144880
rect 231669 144875 231735 144878
rect 264605 144802 264671 144805
rect 279417 144802 279483 144805
rect 264605 144800 268180 144802
rect 264605 144744 264610 144800
rect 264666 144744 268180 144800
rect 264605 144742 268180 144744
rect 279374 144800 279483 144802
rect 279374 144744 279422 144800
rect 279478 144744 279483 144800
rect 264605 144739 264671 144742
rect 279374 144739 279483 144744
rect 214005 144530 214071 144533
rect 214005 144528 217028 144530
rect 214005 144472 214010 144528
rect 214066 144472 217028 144528
rect 214005 144470 217028 144472
rect 214005 144467 214071 144470
rect 231577 144394 231643 144397
rect 228988 144392 231643 144394
rect 228988 144336 231582 144392
rect 231638 144336 231643 144392
rect 228988 144334 231643 144336
rect 231577 144331 231643 144334
rect 230422 144060 230428 144124
rect 230492 144122 230498 144124
rect 248454 144122 248460 144124
rect 230492 144062 248460 144122
rect 230492 144060 230498 144062
rect 248454 144060 248460 144062
rect 248524 144060 248530 144124
rect 242157 143986 242223 143989
rect 228988 143984 242223 143986
rect 228988 143928 242162 143984
rect 242218 143928 242223 143984
rect 228988 143926 242223 143928
rect 242157 143923 242223 143926
rect 242341 143986 242407 143989
rect 268150 143986 268210 144364
rect 279374 144228 279434 144739
rect 242341 143984 268210 143986
rect 242341 143928 242346 143984
rect 242402 143928 268210 143984
rect 242341 143926 268210 143928
rect 242341 143923 242407 143926
rect 213913 143850 213979 143853
rect 264973 143850 265039 143853
rect 213913 143848 217028 143850
rect 213913 143792 213918 143848
rect 213974 143792 217028 143848
rect 213913 143790 217028 143792
rect 264973 143848 268180 143850
rect 264973 143792 264978 143848
rect 265034 143792 268180 143848
rect 264973 143790 268180 143792
rect 213913 143787 213979 143790
rect 264973 143787 265039 143790
rect 288566 143578 288572 143580
rect 279956 143518 288572 143578
rect 288566 143516 288572 143518
rect 288636 143516 288642 143580
rect 231761 143442 231827 143445
rect 228988 143440 231827 143442
rect 228988 143384 231766 143440
rect 231822 143384 231827 143440
rect 228988 143382 231827 143384
rect 231761 143379 231827 143382
rect 264973 143442 265039 143445
rect 264973 143440 268180 143442
rect 264973 143384 264978 143440
rect 265034 143384 268180 143440
rect 264973 143382 268180 143384
rect 264973 143379 265039 143382
rect 213913 143306 213979 143309
rect 213913 143304 217028 143306
rect 213913 143248 213918 143304
rect 213974 143248 217028 143304
rect 213913 143246 217028 143248
rect 213913 143243 213979 143246
rect 231669 143034 231735 143037
rect 228988 143032 231735 143034
rect 228988 142976 231674 143032
rect 231730 142976 231735 143032
rect 228988 142974 231735 142976
rect 231669 142971 231735 142974
rect 258030 142974 268180 143034
rect 254761 142898 254827 142901
rect 258030 142898 258090 142974
rect 254761 142896 258090 142898
rect 254761 142840 254766 142896
rect 254822 142840 258090 142896
rect 254761 142838 258090 142840
rect 254761 142835 254827 142838
rect 170254 142700 170260 142764
rect 170324 142762 170330 142764
rect 191097 142762 191163 142765
rect 170324 142760 191163 142762
rect 170324 142704 191102 142760
rect 191158 142704 191163 142760
rect 170324 142702 191163 142704
rect 170324 142700 170330 142702
rect 191097 142699 191163 142702
rect 242433 142762 242499 142765
rect 265433 142762 265499 142765
rect 282821 142762 282887 142765
rect 242433 142760 265499 142762
rect 242433 142704 242438 142760
rect 242494 142704 265438 142760
rect 265494 142704 265499 142760
rect 242433 142702 265499 142704
rect 279956 142760 282887 142762
rect 279956 142704 282826 142760
rect 282882 142704 282887 142760
rect 279956 142702 282887 142704
rect 242433 142699 242499 142702
rect 265433 142699 265499 142702
rect 282821 142699 282887 142702
rect 216029 142626 216095 142629
rect 265157 142626 265223 142629
rect 216029 142624 217028 142626
rect 216029 142568 216034 142624
rect 216090 142568 217028 142624
rect 216029 142566 217028 142568
rect 265157 142624 268180 142626
rect 265157 142568 265162 142624
rect 265218 142568 268180 142624
rect 265157 142566 268180 142568
rect 216029 142563 216095 142566
rect 265157 142563 265223 142566
rect 237966 142490 237972 142492
rect 228988 142430 237972 142490
rect 237966 142428 237972 142430
rect 238036 142428 238042 142492
rect 265617 142218 265683 142221
rect 265617 142216 268180 142218
rect 265617 142160 265622 142216
rect 265678 142160 268180 142216
rect 265617 142158 268180 142160
rect 265617 142155 265683 142158
rect 231117 142082 231183 142085
rect 282821 142082 282887 142085
rect 228988 142080 231183 142082
rect 228988 142024 231122 142080
rect 231178 142024 231183 142080
rect 228988 142022 231183 142024
rect 279956 142080 282887 142082
rect 279956 142024 282826 142080
rect 282882 142024 282887 142080
rect 279956 142022 282887 142024
rect 231117 142019 231183 142022
rect 282821 142019 282887 142022
rect 213913 141946 213979 141949
rect 213913 141944 217028 141946
rect 213913 141888 213918 141944
rect 213974 141888 217028 141944
rect 213913 141886 217028 141888
rect 213913 141883 213979 141886
rect 258030 141750 268180 141810
rect 230422 141674 230428 141676
rect 228988 141614 230428 141674
rect 230422 141612 230428 141614
rect 230492 141612 230498 141676
rect 232446 141612 232452 141676
rect 232516 141674 232522 141676
rect 258030 141674 258090 141750
rect 232516 141614 258090 141674
rect 232516 141612 232522 141614
rect 230974 141476 230980 141540
rect 231044 141538 231050 141540
rect 250713 141538 250779 141541
rect 231044 141536 250779 141538
rect 231044 141480 250718 141536
rect 250774 141480 250779 141536
rect 231044 141478 250779 141480
rect 231044 141476 231050 141478
rect 250713 141475 250779 141478
rect 231710 141340 231716 141404
rect 231780 141402 231786 141404
rect 257337 141402 257403 141405
rect 231780 141400 257403 141402
rect 231780 141344 257342 141400
rect 257398 141344 257403 141400
rect 231780 141342 257403 141344
rect 231780 141340 231786 141342
rect 257337 141339 257403 141342
rect 214097 141266 214163 141269
rect 265065 141266 265131 141269
rect 282085 141266 282151 141269
rect 214097 141264 217028 141266
rect 214097 141208 214102 141264
rect 214158 141208 217028 141264
rect 214097 141206 217028 141208
rect 265065 141264 268180 141266
rect 265065 141208 265070 141264
rect 265126 141208 268180 141264
rect 265065 141206 268180 141208
rect 279956 141264 282151 141266
rect 279956 141208 282090 141264
rect 282146 141208 282151 141264
rect 279956 141206 282151 141208
rect 214097 141203 214163 141206
rect 265065 141203 265131 141206
rect 282085 141203 282151 141206
rect 229134 141130 229140 141132
rect 228988 141070 229140 141130
rect 229134 141068 229140 141070
rect 229204 141068 229210 141132
rect 264421 140858 264487 140861
rect 264421 140856 268180 140858
rect 264421 140800 264426 140856
rect 264482 140800 268180 140856
rect 264421 140798 268180 140800
rect 264421 140795 264487 140798
rect 231761 140722 231827 140725
rect 228988 140720 231827 140722
rect 228988 140664 231766 140720
rect 231822 140664 231827 140720
rect 228988 140662 231827 140664
rect 231761 140659 231827 140662
rect 233877 140722 233943 140725
rect 246665 140722 246731 140725
rect 233877 140720 246731 140722
rect 233877 140664 233882 140720
rect 233938 140664 246670 140720
rect 246726 140664 246731 140720
rect 233877 140662 246731 140664
rect 233877 140659 233943 140662
rect 246665 140659 246731 140662
rect 213913 140586 213979 140589
rect 213913 140584 217028 140586
rect 213913 140528 213918 140584
rect 213974 140528 217028 140584
rect 213913 140526 217028 140528
rect 213913 140523 213979 140526
rect 266854 140388 266860 140452
rect 266924 140450 266930 140452
rect 284518 140450 284524 140452
rect 266924 140390 268180 140450
rect 279956 140390 284524 140450
rect 266924 140388 266930 140390
rect 284518 140388 284524 140390
rect 284588 140388 284594 140452
rect 241513 140178 241579 140181
rect 228988 140176 241579 140178
rect 228988 140120 241518 140176
rect 241574 140120 241579 140176
rect 228988 140118 241579 140120
rect 241513 140115 241579 140118
rect 244774 139980 244780 140044
rect 244844 140042 244850 140044
rect 265157 140042 265223 140045
rect 244844 140040 265223 140042
rect 244844 139984 265162 140040
rect 265218 139984 265223 140040
rect 244844 139982 265223 139984
rect 244844 139980 244850 139982
rect 265157 139979 265223 139982
rect 265341 140042 265407 140045
rect 265341 140040 268180 140042
rect 265341 139984 265346 140040
rect 265402 139984 268180 140040
rect 265341 139982 268180 139984
rect 265341 139979 265407 139982
rect 214005 139906 214071 139909
rect 214005 139904 217028 139906
rect 214005 139848 214010 139904
rect 214066 139848 217028 139904
rect 214005 139846 217028 139848
rect 214005 139843 214071 139846
rect 230749 139770 230815 139773
rect 282821 139770 282887 139773
rect 228988 139768 230815 139770
rect 228988 139712 230754 139768
rect 230810 139712 230815 139768
rect 228988 139710 230815 139712
rect 279956 139768 282887 139770
rect 279956 139712 282826 139768
rect 282882 139712 282887 139768
rect 279956 139710 282887 139712
rect 230749 139707 230815 139710
rect 282821 139707 282887 139710
rect 258030 139574 268180 139634
rect 246389 139498 246455 139501
rect 258030 139498 258090 139574
rect 246389 139496 258090 139498
rect 246389 139440 246394 139496
rect 246450 139440 258090 139496
rect 246389 139438 258090 139440
rect 246389 139435 246455 139438
rect 583293 139362 583359 139365
rect 583520 139362 584960 139452
rect 583293 139360 584960 139362
rect 583293 139304 583298 139360
rect 583354 139304 584960 139360
rect 583293 139302 584960 139304
rect 583293 139299 583359 139302
rect 214833 139226 214899 139229
rect 229737 139226 229803 139229
rect 214833 139224 217028 139226
rect 214833 139168 214838 139224
rect 214894 139168 217028 139224
rect 214833 139166 217028 139168
rect 228988 139224 229803 139226
rect 228988 139168 229742 139224
rect 229798 139168 229803 139224
rect 228988 139166 229803 139168
rect 214833 139163 214899 139166
rect 229737 139163 229803 139166
rect 264973 139226 265039 139229
rect 264973 139224 268180 139226
rect 264973 139168 264978 139224
rect 265034 139168 268180 139224
rect 583520 139212 584960 139302
rect 264973 139166 268180 139168
rect 264973 139163 265039 139166
rect 282821 138954 282887 138957
rect 279956 138952 282887 138954
rect 279956 138896 282826 138952
rect 282882 138896 282887 138952
rect 279956 138894 282887 138896
rect 282821 138891 282887 138894
rect 241646 138818 241652 138820
rect 228988 138758 241652 138818
rect 241646 138756 241652 138758
rect 241716 138756 241722 138820
rect 213913 138682 213979 138685
rect 213913 138680 217028 138682
rect 213913 138624 213918 138680
rect 213974 138624 217028 138680
rect 213913 138622 217028 138624
rect 213913 138619 213979 138622
rect 237966 138620 237972 138684
rect 238036 138682 238042 138684
rect 265065 138682 265131 138685
rect 238036 138680 265131 138682
rect 238036 138624 265070 138680
rect 265126 138624 265131 138680
rect 238036 138622 265131 138624
rect 238036 138620 238042 138622
rect 265065 138619 265131 138622
rect 267774 138620 267780 138684
rect 267844 138682 267850 138684
rect 267844 138622 268180 138682
rect 267844 138620 267850 138622
rect 231485 138274 231551 138277
rect 228988 138272 231551 138274
rect 228988 138216 231490 138272
rect 231546 138216 231551 138272
rect 228988 138214 231551 138216
rect 231485 138211 231551 138214
rect 266997 138274 267063 138277
rect 282821 138274 282887 138277
rect 266997 138272 268180 138274
rect 266997 138216 267002 138272
rect 267058 138216 268180 138272
rect 266997 138214 268180 138216
rect 279956 138272 282887 138274
rect 279956 138216 282826 138272
rect 282882 138216 282887 138272
rect 279956 138214 282887 138216
rect 266997 138211 267063 138214
rect 282821 138211 282887 138214
rect 214005 138002 214071 138005
rect 214005 138000 217028 138002
rect 214005 137944 214010 138000
rect 214066 137944 217028 138000
rect 214005 137942 217028 137944
rect 214005 137939 214071 137942
rect 229921 137866 229987 137869
rect 228988 137864 229987 137866
rect 228988 137808 229926 137864
rect 229982 137808 229987 137864
rect 228988 137806 229987 137808
rect 229921 137803 229987 137806
rect 264973 137866 265039 137869
rect 264973 137864 268180 137866
rect 264973 137808 264978 137864
rect 265034 137808 268180 137864
rect 264973 137806 268180 137808
rect 264973 137803 265039 137806
rect 282821 137458 282887 137461
rect 279956 137456 282887 137458
rect 214741 137322 214807 137325
rect 229686 137322 229692 137324
rect 214741 137320 217028 137322
rect 214741 137264 214746 137320
rect 214802 137264 217028 137320
rect 214741 137262 217028 137264
rect 228988 137262 229692 137322
rect 214741 137259 214807 137262
rect 229686 137260 229692 137262
rect 229756 137260 229762 137324
rect 239397 137186 239463 137189
rect 268150 137186 268210 137428
rect 279956 137400 282826 137456
rect 282882 137400 282887 137456
rect 279956 137398 282887 137400
rect 282821 137395 282887 137398
rect 239397 137184 268210 137186
rect 239397 137128 239402 137184
rect 239458 137128 268210 137184
rect 239397 137126 268210 137128
rect 239397 137123 239463 137126
rect 258030 136990 268180 137050
rect 231577 136914 231643 136917
rect 228988 136912 231643 136914
rect -960 136778 480 136868
rect 228988 136856 231582 136912
rect 231638 136856 231643 136912
rect 228988 136854 231643 136856
rect 231577 136851 231643 136854
rect 242157 136914 242223 136917
rect 258030 136914 258090 136990
rect 242157 136912 258090 136914
rect 242157 136856 242162 136912
rect 242218 136856 258090 136912
rect 242157 136854 258090 136856
rect 242157 136851 242223 136854
rect 3509 136778 3575 136781
rect -960 136776 3575 136778
rect -960 136720 3514 136776
rect 3570 136720 3575 136776
rect -960 136718 3575 136720
rect -960 136628 480 136718
rect 3509 136715 3575 136718
rect 213361 136642 213427 136645
rect 265065 136642 265131 136645
rect 282821 136642 282887 136645
rect 213361 136640 217028 136642
rect 213361 136584 213366 136640
rect 213422 136584 217028 136640
rect 213361 136582 217028 136584
rect 265065 136640 268180 136642
rect 265065 136584 265070 136640
rect 265126 136584 268180 136640
rect 265065 136582 268180 136584
rect 279956 136640 282887 136642
rect 279956 136584 282826 136640
rect 282882 136584 282887 136640
rect 279956 136582 282887 136584
rect 213361 136579 213427 136582
rect 265065 136579 265131 136582
rect 282821 136579 282887 136582
rect 245653 136370 245719 136373
rect 282821 136370 282887 136373
rect 228988 136368 245719 136370
rect 228988 136312 245658 136368
rect 245714 136312 245719 136368
rect 228988 136310 245719 136312
rect 245653 136307 245719 136310
rect 279926 136368 282887 136370
rect 279926 136312 282826 136368
rect 282882 136312 282887 136368
rect 279926 136310 282887 136312
rect 213913 135962 213979 135965
rect 230565 135962 230631 135965
rect 213913 135960 217028 135962
rect 213913 135904 213918 135960
rect 213974 135904 217028 135960
rect 213913 135902 217028 135904
rect 228988 135960 230631 135962
rect 228988 135904 230570 135960
rect 230626 135904 230631 135960
rect 228988 135902 230631 135904
rect 213913 135899 213979 135902
rect 230565 135899 230631 135902
rect 249149 135962 249215 135965
rect 262765 135962 262831 135965
rect 249149 135960 262831 135962
rect 249149 135904 249154 135960
rect 249210 135904 262770 135960
rect 262826 135904 262831 135960
rect 249149 135902 262831 135904
rect 249149 135899 249215 135902
rect 262765 135899 262831 135902
rect 229737 135826 229803 135829
rect 268150 135826 268210 136204
rect 279926 135932 279986 136310
rect 282821 136307 282887 136310
rect 229737 135824 268210 135826
rect 229737 135768 229742 135824
rect 229798 135768 268210 135824
rect 229737 135766 268210 135768
rect 229737 135763 229803 135766
rect 264973 135690 265039 135693
rect 264973 135688 268180 135690
rect 264973 135632 264978 135688
rect 265034 135632 268180 135688
rect 264973 135630 268180 135632
rect 264973 135627 265039 135630
rect 231485 135418 231551 135421
rect 228988 135416 231551 135418
rect 228988 135360 231490 135416
rect 231546 135360 231551 135416
rect 228988 135358 231551 135360
rect 231485 135355 231551 135358
rect 262765 135418 262831 135421
rect 262765 135416 268210 135418
rect 262765 135360 262770 135416
rect 262826 135360 268210 135416
rect 262765 135358 268210 135360
rect 262765 135355 262831 135358
rect 213913 135282 213979 135285
rect 213913 135280 217028 135282
rect 213913 135224 213918 135280
rect 213974 135224 217028 135280
rect 268150 135252 268210 135358
rect 213913 135222 217028 135224
rect 213913 135219 213979 135222
rect 279366 135220 279372 135284
rect 279436 135220 279442 135284
rect 279374 135116 279434 135220
rect 231710 135010 231716 135012
rect 228988 134950 231716 135010
rect 231710 134948 231716 134950
rect 231780 134948 231786 135012
rect 213913 134602 213979 134605
rect 268150 134602 268210 134844
rect 213913 134600 217028 134602
rect 213913 134544 213918 134600
rect 213974 134544 217028 134600
rect 213913 134542 217028 134544
rect 258030 134542 268210 134602
rect 213913 134539 213979 134542
rect 231025 134466 231091 134469
rect 228988 134464 231091 134466
rect 228988 134408 231030 134464
rect 231086 134408 231091 134464
rect 228988 134406 231091 134408
rect 231025 134403 231091 134406
rect 233734 134132 233740 134196
rect 233804 134194 233810 134196
rect 258030 134194 258090 134542
rect 267089 134466 267155 134469
rect 282453 134466 282519 134469
rect 267089 134464 268180 134466
rect 267089 134408 267094 134464
rect 267150 134408 268180 134464
rect 267089 134406 268180 134408
rect 279956 134464 282519 134466
rect 279956 134408 282458 134464
rect 282514 134408 282519 134464
rect 279956 134406 282519 134408
rect 267089 134403 267155 134406
rect 282453 134403 282519 134406
rect 233804 134134 258090 134194
rect 233804 134132 233810 134134
rect 231577 134058 231643 134061
rect 228988 134056 231643 134058
rect 228988 134000 231582 134056
rect 231638 134000 231643 134056
rect 228988 133998 231643 134000
rect 231577 133995 231643 133998
rect 264973 134058 265039 134061
rect 264973 134056 268180 134058
rect 264973 134000 264978 134056
rect 265034 134000 268180 134056
rect 264973 133998 268180 134000
rect 264973 133995 265039 133998
rect 213269 133922 213335 133925
rect 213269 133920 217028 133922
rect 213269 133864 213274 133920
rect 213330 133864 217028 133920
rect 213269 133862 217028 133864
rect 213269 133859 213335 133862
rect 282821 133650 282887 133653
rect 279956 133648 282887 133650
rect 230841 133514 230907 133517
rect 228988 133512 230907 133514
rect 228988 133456 230846 133512
rect 230902 133456 230907 133512
rect 228988 133454 230907 133456
rect 230841 133451 230907 133454
rect 214005 133378 214071 133381
rect 214005 133376 217028 133378
rect 214005 133320 214010 133376
rect 214066 133320 217028 133376
rect 214005 133318 217028 133320
rect 214005 133315 214071 133318
rect 268150 133242 268210 133620
rect 279956 133592 282826 133648
rect 282882 133592 282887 133648
rect 279956 133590 282887 133592
rect 282821 133587 282887 133590
rect 258030 133182 268210 133242
rect 231761 133106 231827 133109
rect 228988 133104 231827 133106
rect 228988 133048 231766 133104
rect 231822 133048 231827 133104
rect 228988 133046 231827 133048
rect 231761 133043 231827 133046
rect 229921 132834 229987 132837
rect 258030 132834 258090 133182
rect 264094 133044 264100 133108
rect 264164 133106 264170 133108
rect 264164 133046 268180 133106
rect 264164 133044 264170 133046
rect 282729 132834 282795 132837
rect 229921 132832 258090 132834
rect 229921 132776 229926 132832
rect 229982 132776 258090 132832
rect 229921 132774 258090 132776
rect 279956 132832 282795 132834
rect 279956 132776 282734 132832
rect 282790 132776 282795 132832
rect 279956 132774 282795 132776
rect 229921 132771 229987 132774
rect 282729 132771 282795 132774
rect 213913 132698 213979 132701
rect 264973 132698 265039 132701
rect 213913 132696 217028 132698
rect 213913 132640 213918 132696
rect 213974 132640 217028 132696
rect 213913 132638 217028 132640
rect 264973 132696 268180 132698
rect 264973 132640 264978 132696
rect 265034 132640 268180 132696
rect 264973 132638 268180 132640
rect 213913 132635 213979 132638
rect 264973 132635 265039 132638
rect 231669 132562 231735 132565
rect 228988 132560 231735 132562
rect 228988 132504 231674 132560
rect 231730 132504 231735 132560
rect 228988 132502 231735 132504
rect 231669 132499 231735 132502
rect 264973 132290 265039 132293
rect 264973 132288 268180 132290
rect 264973 132232 264978 132288
rect 265034 132232 268180 132288
rect 264973 132230 268180 132232
rect 264973 132227 265039 132230
rect 230974 132154 230980 132156
rect 228988 132094 230980 132154
rect 230974 132092 230980 132094
rect 231044 132092 231050 132156
rect 282177 132154 282243 132157
rect 279956 132152 282243 132154
rect 279956 132096 282182 132152
rect 282238 132096 282243 132152
rect 279956 132094 282243 132096
rect 282177 132091 282243 132094
rect 213913 132018 213979 132021
rect 213913 132016 217028 132018
rect 213913 131960 213918 132016
rect 213974 131960 217028 132016
rect 213913 131958 217028 131960
rect 213913 131955 213979 131958
rect 231301 131610 231367 131613
rect 228988 131608 231367 131610
rect 228988 131552 231306 131608
rect 231362 131552 231367 131608
rect 228988 131550 231367 131552
rect 231301 131547 231367 131550
rect 253289 131610 253355 131613
rect 268150 131610 268210 131852
rect 253289 131608 268210 131610
rect 253289 131552 253294 131608
rect 253350 131552 268210 131608
rect 253289 131550 268210 131552
rect 253289 131547 253355 131550
rect 262806 131412 262812 131476
rect 262876 131474 262882 131476
rect 262876 131414 268180 131474
rect 262876 131412 262882 131414
rect 214005 131338 214071 131341
rect 282821 131338 282887 131341
rect 214005 131336 217028 131338
rect 214005 131280 214010 131336
rect 214066 131280 217028 131336
rect 214005 131278 217028 131280
rect 279956 131336 282887 131338
rect 279956 131280 282826 131336
rect 282882 131280 282887 131336
rect 279956 131278 282887 131280
rect 214005 131275 214071 131278
rect 282821 131275 282887 131278
rect 231669 131202 231735 131205
rect 228988 131200 231735 131202
rect 228988 131144 231674 131200
rect 231730 131144 231735 131200
rect 228988 131142 231735 131144
rect 231669 131139 231735 131142
rect 254853 131066 254919 131069
rect 238710 131064 254919 131066
rect 238710 131008 254858 131064
rect 254914 131008 254919 131064
rect 238710 131006 254919 131008
rect 213913 130658 213979 130661
rect 238710 130658 238770 131006
rect 254853 131003 254919 131006
rect 264973 131066 265039 131069
rect 264973 131064 268180 131066
rect 264973 131008 264978 131064
rect 265034 131008 268180 131064
rect 264973 131006 268180 131008
rect 264973 131003 265039 131006
rect 282821 130658 282887 130661
rect 213913 130656 217028 130658
rect 213913 130600 213918 130656
rect 213974 130600 217028 130656
rect 213913 130598 217028 130600
rect 228988 130598 238770 130658
rect 279956 130656 282887 130658
rect 279956 130600 282826 130656
rect 282882 130600 282887 130656
rect 279956 130598 282887 130600
rect 213913 130595 213979 130598
rect 282821 130595 282887 130598
rect 265065 130522 265131 130525
rect 265065 130520 268180 130522
rect 265065 130464 265070 130520
rect 265126 130464 268180 130520
rect 265065 130462 268180 130464
rect 265065 130459 265131 130462
rect 231209 130250 231275 130253
rect 228988 130248 231275 130250
rect 228988 130192 231214 130248
rect 231270 130192 231275 130248
rect 228988 130190 231275 130192
rect 231209 130187 231275 130190
rect 258030 130054 268180 130114
rect 214649 129978 214715 129981
rect 214649 129976 217028 129978
rect 214649 129920 214654 129976
rect 214710 129920 217028 129976
rect 214649 129918 217028 129920
rect 214649 129915 214715 129918
rect 250294 129916 250300 129980
rect 250364 129978 250370 129980
rect 258030 129978 258090 130054
rect 250364 129918 258090 129978
rect 250364 129916 250370 129918
rect 230565 129842 230631 129845
rect 282729 129842 282795 129845
rect 228988 129840 230631 129842
rect 228988 129784 230570 129840
rect 230626 129784 230631 129840
rect 228988 129782 230631 129784
rect 279956 129840 282795 129842
rect 279956 129784 282734 129840
rect 282790 129784 282795 129840
rect 279956 129782 282795 129784
rect 230565 129779 230631 129782
rect 282729 129779 282795 129782
rect 265157 129706 265223 129709
rect 265157 129704 268180 129706
rect 265157 129648 265162 129704
rect 265218 129648 268180 129704
rect 265157 129646 268180 129648
rect 265157 129643 265223 129646
rect 66161 129298 66227 129301
rect 68142 129298 68816 129304
rect 66161 129296 68816 129298
rect 66161 129240 66166 129296
rect 66222 129244 68816 129296
rect 214557 129298 214623 129301
rect 231761 129298 231827 129301
rect 214557 129296 217028 129298
rect 66222 129240 68202 129244
rect 66161 129238 68202 129240
rect 214557 129240 214562 129296
rect 214618 129240 217028 129296
rect 214557 129238 217028 129240
rect 228988 129296 231827 129298
rect 228988 129240 231766 129296
rect 231822 129240 231827 129296
rect 228988 129238 231827 129240
rect 66161 129235 66227 129238
rect 214557 129235 214623 129238
rect 231761 129235 231827 129238
rect 264973 129298 265039 129301
rect 264973 129296 268180 129298
rect 264973 129240 264978 129296
rect 265034 129240 268180 129296
rect 264973 129238 268180 129240
rect 264973 129235 265039 129238
rect 231158 128964 231164 129028
rect 231228 129026 231234 129028
rect 250437 129026 250503 129029
rect 281809 129026 281875 129029
rect 231228 129024 250503 129026
rect 231228 128968 250442 129024
rect 250498 128968 250503 129024
rect 231228 128966 250503 128968
rect 279956 129024 281875 129026
rect 279956 128968 281814 129024
rect 281870 128968 281875 129024
rect 279956 128966 281875 128968
rect 231228 128964 231234 128966
rect 250437 128963 250503 128966
rect 281809 128963 281875 128966
rect 231669 128890 231735 128893
rect 228988 128888 231735 128890
rect 228988 128832 231674 128888
rect 231730 128832 231735 128888
rect 228988 128830 231735 128832
rect 231669 128827 231735 128830
rect 258030 128830 268180 128890
rect 213913 128754 213979 128757
rect 236637 128754 236703 128757
rect 258030 128754 258090 128830
rect 213913 128752 217028 128754
rect 213913 128696 213918 128752
rect 213974 128696 217028 128752
rect 213913 128694 217028 128696
rect 236637 128752 258090 128754
rect 236637 128696 236642 128752
rect 236698 128696 258090 128752
rect 236637 128694 258090 128696
rect 213913 128691 213979 128694
rect 236637 128691 236703 128694
rect 267590 128420 267596 128484
rect 267660 128482 267666 128484
rect 267660 128422 268180 128482
rect 267660 128420 267666 128422
rect 231117 128346 231183 128349
rect 282821 128346 282887 128349
rect 228988 128344 231183 128346
rect 228988 128288 231122 128344
rect 231178 128288 231183 128344
rect 228988 128286 231183 128288
rect 279956 128344 282887 128346
rect 279956 128288 282826 128344
rect 282882 128288 282887 128344
rect 279956 128286 282887 128288
rect 231117 128283 231183 128286
rect 282821 128283 282887 128286
rect 67633 128074 67699 128077
rect 68142 128074 68816 128080
rect 67633 128072 68816 128074
rect 67633 128016 67638 128072
rect 67694 128020 68816 128072
rect 214005 128074 214071 128077
rect 214005 128072 217028 128074
rect 67694 128016 68202 128020
rect 67633 128014 68202 128016
rect 214005 128016 214010 128072
rect 214066 128016 217028 128072
rect 214005 128014 217028 128016
rect 67633 128011 67699 128014
rect 214005 128011 214071 128014
rect 231761 127938 231827 127941
rect 228988 127936 231827 127938
rect 228988 127880 231766 127936
rect 231822 127880 231827 127936
rect 228988 127878 231827 127880
rect 231761 127875 231827 127878
rect 265801 127938 265867 127941
rect 265801 127936 268180 127938
rect 265801 127880 265806 127936
rect 265862 127880 268180 127936
rect 265801 127878 268180 127880
rect 265801 127875 265867 127878
rect 231117 127802 231183 127805
rect 243905 127802 243971 127805
rect 231117 127800 243971 127802
rect 231117 127744 231122 127800
rect 231178 127744 243910 127800
rect 243966 127744 243971 127800
rect 231117 127742 243971 127744
rect 231117 127739 231183 127742
rect 243905 127739 243971 127742
rect 231301 127666 231367 127669
rect 249333 127666 249399 127669
rect 231301 127664 249399 127666
rect 231301 127608 231306 127664
rect 231362 127608 249338 127664
rect 249394 127608 249399 127664
rect 231301 127606 249399 127608
rect 231301 127603 231367 127606
rect 249333 127603 249399 127606
rect 264973 127530 265039 127533
rect 282729 127530 282795 127533
rect 264973 127528 268180 127530
rect 264973 127472 264978 127528
rect 265034 127472 268180 127528
rect 264973 127470 268180 127472
rect 279956 127528 282795 127530
rect 279956 127472 282734 127528
rect 282790 127472 282795 127528
rect 279956 127470 282795 127472
rect 264973 127467 265039 127470
rect 282729 127467 282795 127470
rect 213913 127394 213979 127397
rect 230749 127394 230815 127397
rect 213913 127392 217028 127394
rect 213913 127336 213918 127392
rect 213974 127336 217028 127392
rect 213913 127334 217028 127336
rect 228988 127392 230815 127394
rect 228988 127336 230754 127392
rect 230810 127336 230815 127392
rect 228988 127334 230815 127336
rect 213913 127331 213979 127334
rect 230749 127331 230815 127334
rect 242014 127060 242020 127124
rect 242084 127122 242090 127124
rect 242084 127062 268180 127122
rect 242084 127060 242090 127062
rect 231761 126986 231827 126989
rect 228988 126984 231827 126986
rect 228988 126928 231766 126984
rect 231822 126928 231827 126984
rect 228988 126926 231827 126928
rect 231761 126923 231827 126926
rect 280286 126850 280292 126852
rect 279956 126790 280292 126850
rect 280286 126788 280292 126790
rect 280356 126788 280362 126852
rect 214005 126714 214071 126717
rect 214005 126712 217028 126714
rect 214005 126656 214010 126712
rect 214066 126656 217028 126712
rect 214005 126654 217028 126656
rect 214005 126651 214071 126654
rect 265065 126578 265131 126581
rect 258030 126576 265131 126578
rect 258030 126520 265070 126576
rect 265126 126520 265131 126576
rect 258030 126518 265131 126520
rect 230565 126442 230631 126445
rect 228988 126440 230631 126442
rect 228988 126384 230570 126440
rect 230626 126384 230631 126440
rect 228988 126382 230631 126384
rect 230565 126379 230631 126382
rect 67449 126306 67515 126309
rect 68142 126306 68816 126312
rect 67449 126304 68816 126306
rect 67449 126248 67454 126304
rect 67510 126252 68816 126304
rect 67510 126248 68202 126252
rect 67449 126246 68202 126248
rect 67449 126243 67515 126246
rect 244958 126244 244964 126308
rect 245028 126306 245034 126308
rect 258030 126306 258090 126518
rect 265065 126515 265131 126518
rect 268150 126442 268210 126684
rect 245028 126246 258090 126306
rect 262814 126382 268210 126442
rect 245028 126244 245034 126246
rect 213913 126034 213979 126037
rect 230841 126034 230907 126037
rect 213913 126032 217028 126034
rect 213913 125976 213918 126032
rect 213974 125976 217028 126032
rect 213913 125974 217028 125976
rect 228988 126032 230907 126034
rect 228988 125976 230846 126032
rect 230902 125976 230907 126032
rect 228988 125974 230907 125976
rect 213913 125971 213979 125974
rect 230841 125971 230907 125974
rect 230974 125972 230980 126036
rect 231044 126034 231050 126036
rect 262814 126034 262874 126382
rect 265893 126306 265959 126309
rect 265893 126304 268180 126306
rect 265893 126248 265898 126304
rect 265954 126248 268180 126304
rect 265893 126246 268180 126248
rect 265893 126243 265959 126246
rect 282361 126034 282427 126037
rect 231044 125974 262874 126034
rect 279956 126032 282427 126034
rect 279956 125976 282366 126032
rect 282422 125976 282427 126032
rect 279956 125974 282427 125976
rect 231044 125972 231050 125974
rect 282361 125971 282427 125974
rect 583109 126034 583175 126037
rect 583520 126034 584960 126124
rect 583109 126032 584960 126034
rect 583109 125976 583114 126032
rect 583170 125976 584960 126032
rect 583109 125974 584960 125976
rect 583109 125971 583175 125974
rect 264973 125898 265039 125901
rect 264973 125896 268180 125898
rect 264973 125840 264978 125896
rect 265034 125840 268180 125896
rect 583520 125884 584960 125974
rect 264973 125838 268180 125840
rect 264973 125835 265039 125838
rect 232589 125490 232655 125493
rect 228988 125488 232655 125490
rect 228988 125432 232594 125488
rect 232650 125432 232655 125488
rect 228988 125430 232655 125432
rect 232589 125427 232655 125430
rect 214005 125354 214071 125357
rect 214005 125352 217028 125354
rect 214005 125296 214010 125352
rect 214066 125296 217028 125352
rect 214005 125294 217028 125296
rect 214005 125291 214071 125294
rect 65977 125218 66043 125221
rect 68142 125218 68816 125224
rect 65977 125216 68816 125218
rect 65977 125160 65982 125216
rect 66038 125164 68816 125216
rect 66038 125160 68202 125164
rect 65977 125158 68202 125160
rect 65977 125155 66043 125158
rect 231761 125082 231827 125085
rect 228988 125080 231827 125082
rect 228988 125024 231766 125080
rect 231822 125024 231827 125080
rect 228988 125022 231827 125024
rect 231761 125019 231827 125022
rect 262765 125082 262831 125085
rect 268150 125082 268210 125324
rect 282821 125218 282887 125221
rect 279956 125216 282887 125218
rect 279956 125160 282826 125216
rect 282882 125160 282887 125216
rect 279956 125158 282887 125160
rect 282821 125155 282887 125158
rect 262765 125080 268210 125082
rect 262765 125024 262770 125080
rect 262826 125024 268210 125080
rect 262765 125022 268210 125024
rect 262765 125019 262831 125022
rect 258030 124886 268180 124946
rect 239673 124810 239739 124813
rect 258030 124810 258090 124886
rect 239673 124808 258090 124810
rect 239673 124752 239678 124808
rect 239734 124752 258090 124808
rect 239673 124750 258090 124752
rect 239673 124747 239739 124750
rect 213913 124674 213979 124677
rect 232773 124674 232839 124677
rect 262765 124674 262831 124677
rect 213913 124672 217028 124674
rect 213913 124616 213918 124672
rect 213974 124616 217028 124672
rect 213913 124614 217028 124616
rect 232773 124672 262831 124674
rect 232773 124616 232778 124672
rect 232834 124616 262770 124672
rect 262826 124616 262831 124672
rect 232773 124614 262831 124616
rect 213913 124611 213979 124614
rect 232773 124611 232839 124614
rect 262765 124611 262831 124614
rect 231485 124538 231551 124541
rect 228988 124536 231551 124538
rect 228988 124480 231490 124536
rect 231546 124480 231551 124536
rect 228988 124478 231551 124480
rect 231485 124475 231551 124478
rect 264973 124538 265039 124541
rect 282729 124538 282795 124541
rect 264973 124536 268180 124538
rect 264973 124480 264978 124536
rect 265034 124480 268180 124536
rect 264973 124478 268180 124480
rect 279956 124536 282795 124538
rect 279956 124480 282734 124536
rect 282790 124480 282795 124536
rect 279956 124478 282795 124480
rect 264973 124475 265039 124478
rect 282729 124475 282795 124478
rect 213913 124130 213979 124133
rect 231761 124130 231827 124133
rect 213913 124128 217028 124130
rect 213913 124072 213918 124128
rect 213974 124072 217028 124128
rect 213913 124070 217028 124072
rect 228988 124128 231827 124130
rect 228988 124072 231766 124128
rect 231822 124072 231827 124128
rect 228988 124070 231827 124072
rect 213913 124067 213979 124070
rect 231761 124067 231827 124070
rect 267181 124130 267247 124133
rect 267181 124128 268180 124130
rect 267181 124072 267186 124128
rect 267242 124072 268180 124128
rect 267181 124070 268180 124072
rect 267181 124067 267247 124070
rect -960 123572 480 123812
rect 264973 123722 265039 123725
rect 282821 123722 282887 123725
rect 264973 123720 268180 123722
rect 264973 123664 264978 123720
rect 265034 123664 268180 123720
rect 264973 123662 268180 123664
rect 279956 123720 282887 123722
rect 279956 123664 282826 123720
rect 282882 123664 282887 123720
rect 279956 123662 282887 123664
rect 264973 123659 265039 123662
rect 282821 123659 282887 123662
rect 66069 123586 66135 123589
rect 68142 123586 68816 123592
rect 231669 123586 231735 123589
rect 66069 123584 68816 123586
rect 66069 123528 66074 123584
rect 66130 123532 68816 123584
rect 228988 123584 231735 123586
rect 66130 123528 68202 123532
rect 66069 123526 68202 123528
rect 228988 123528 231674 123584
rect 231730 123528 231735 123584
rect 228988 123526 231735 123528
rect 66069 123523 66135 123526
rect 231669 123523 231735 123526
rect 216121 123450 216187 123453
rect 216121 123448 217028 123450
rect 216121 123392 216126 123448
rect 216182 123392 217028 123448
rect 216121 123390 217028 123392
rect 216121 123387 216187 123390
rect 230013 123314 230079 123317
rect 230013 123312 268180 123314
rect 230013 123256 230018 123312
rect 230074 123256 268180 123312
rect 230013 123254 268180 123256
rect 230013 123251 230079 123254
rect 230933 123178 230999 123181
rect 228988 123176 230999 123178
rect 228988 123120 230938 123176
rect 230994 123120 230999 123176
rect 228988 123118 230999 123120
rect 230933 123115 230999 123118
rect 282085 123042 282151 123045
rect 279956 123040 282151 123042
rect 279956 122984 282090 123040
rect 282146 122984 282151 123040
rect 279956 122982 282151 122984
rect 282085 122979 282151 122982
rect 265617 122906 265683 122909
rect 265617 122904 268180 122906
rect 265617 122848 265622 122904
rect 265678 122848 268180 122904
rect 265617 122846 268180 122848
rect 265617 122843 265683 122846
rect 214005 122770 214071 122773
rect 264329 122770 264395 122773
rect 214005 122768 217028 122770
rect 214005 122712 214010 122768
rect 214066 122712 217028 122768
rect 214005 122710 217028 122712
rect 238710 122768 264395 122770
rect 238710 122712 264334 122768
rect 264390 122712 264395 122768
rect 238710 122710 264395 122712
rect 214005 122707 214071 122710
rect 64965 122634 65031 122637
rect 68142 122634 68816 122640
rect 238710 122634 238770 122710
rect 264329 122707 264395 122710
rect 64965 122632 68816 122634
rect 64965 122576 64970 122632
rect 65026 122580 68816 122632
rect 65026 122576 68202 122580
rect 64965 122574 68202 122576
rect 228988 122574 238770 122634
rect 64965 122571 65031 122574
rect 231761 122226 231827 122229
rect 228988 122224 231827 122226
rect 228988 122168 231766 122224
rect 231822 122168 231827 122224
rect 228988 122166 231827 122168
rect 231761 122163 231827 122166
rect 213913 122090 213979 122093
rect 240777 122090 240843 122093
rect 268150 122090 268210 122332
rect 282821 122226 282887 122229
rect 279956 122224 282887 122226
rect 279956 122168 282826 122224
rect 282882 122168 282887 122224
rect 279956 122166 282887 122168
rect 282821 122163 282887 122166
rect 213913 122088 217028 122090
rect 213913 122032 213918 122088
rect 213974 122032 217028 122088
rect 213913 122030 217028 122032
rect 240777 122088 268210 122090
rect 240777 122032 240782 122088
rect 240838 122032 268210 122088
rect 240777 122030 268210 122032
rect 213913 122027 213979 122030
rect 240777 122027 240843 122030
rect 264973 121954 265039 121957
rect 264973 121952 268180 121954
rect 264973 121896 264978 121952
rect 265034 121896 268180 121952
rect 264973 121894 268180 121896
rect 264973 121891 265039 121894
rect 231117 121682 231183 121685
rect 228988 121680 231183 121682
rect 228988 121624 231122 121680
rect 231178 121624 231183 121680
rect 228988 121622 231183 121624
rect 231117 121619 231183 121622
rect 64781 121546 64847 121549
rect 64965 121546 65031 121549
rect 64781 121544 65031 121546
rect 64781 121488 64786 121544
rect 64842 121488 64970 121544
rect 65026 121488 65031 121544
rect 64781 121486 65031 121488
rect 64781 121483 64847 121486
rect 64965 121483 65031 121486
rect 265065 121546 265131 121549
rect 265065 121544 268180 121546
rect 265065 121488 265070 121544
rect 265126 121488 268180 121544
rect 265065 121486 268180 121488
rect 265065 121483 265131 121486
rect 214005 121410 214071 121413
rect 262857 121410 262923 121413
rect 282821 121410 282887 121413
rect 214005 121408 217028 121410
rect 214005 121352 214010 121408
rect 214066 121352 217028 121408
rect 214005 121350 217028 121352
rect 238710 121408 262923 121410
rect 238710 121352 262862 121408
rect 262918 121352 262923 121408
rect 238710 121350 262923 121352
rect 279956 121408 282887 121410
rect 279956 121352 282826 121408
rect 282882 121352 282887 121408
rect 279956 121350 282887 121352
rect 214005 121347 214071 121350
rect 238710 121274 238770 121350
rect 262857 121347 262923 121350
rect 282821 121347 282887 121350
rect 228988 121214 238770 121274
rect 264973 121138 265039 121141
rect 264973 121136 268180 121138
rect 264973 121080 264978 121136
rect 265034 121080 268180 121136
rect 264973 121078 268180 121080
rect 264973 121075 265039 121078
rect 67357 120866 67423 120869
rect 68142 120866 68816 120872
rect 67357 120864 68816 120866
rect 67357 120808 67362 120864
rect 67418 120812 68816 120864
rect 67418 120808 68202 120812
rect 67357 120806 68202 120808
rect 67357 120803 67423 120806
rect 213913 120730 213979 120733
rect 230749 120730 230815 120733
rect 213913 120728 217028 120730
rect 213913 120672 213918 120728
rect 213974 120672 217028 120728
rect 213913 120670 217028 120672
rect 228988 120728 230815 120730
rect 228988 120672 230754 120728
rect 230810 120672 230815 120728
rect 228988 120670 230815 120672
rect 213913 120667 213979 120670
rect 230749 120667 230815 120670
rect 265065 120730 265131 120733
rect 282085 120730 282151 120733
rect 265065 120728 268180 120730
rect 265065 120672 265070 120728
rect 265126 120672 268180 120728
rect 265065 120670 268180 120672
rect 279956 120728 282151 120730
rect 279956 120672 282090 120728
rect 282146 120672 282151 120728
rect 279956 120670 282151 120672
rect 265065 120667 265131 120670
rect 282085 120667 282151 120670
rect 230565 120322 230631 120325
rect 228988 120320 230631 120322
rect 228988 120264 230570 120320
rect 230626 120264 230631 120320
rect 228988 120262 230631 120264
rect 230565 120259 230631 120262
rect 258030 120262 268180 120322
rect 251817 120186 251883 120189
rect 258030 120186 258090 120262
rect 251817 120184 258090 120186
rect 251817 120128 251822 120184
rect 251878 120128 258090 120184
rect 251817 120126 258090 120128
rect 251817 120123 251883 120126
rect 214097 120050 214163 120053
rect 231761 120050 231827 120053
rect 257429 120050 257495 120053
rect 214097 120048 217028 120050
rect 214097 119992 214102 120048
rect 214158 119992 217028 120048
rect 214097 119990 217028 119992
rect 231761 120048 257495 120050
rect 231761 119992 231766 120048
rect 231822 119992 257434 120048
rect 257490 119992 257495 120048
rect 231761 119990 257495 119992
rect 214097 119987 214163 119990
rect 231761 119987 231827 119990
rect 257429 119987 257495 119990
rect 282821 119914 282887 119917
rect 279956 119912 282887 119914
rect 279956 119856 282826 119912
rect 282882 119856 282887 119912
rect 279956 119854 282887 119856
rect 282821 119851 282887 119854
rect 231158 119778 231164 119780
rect 228988 119718 231164 119778
rect 231158 119716 231164 119718
rect 231228 119716 231234 119780
rect 264973 119778 265039 119781
rect 264973 119776 268180 119778
rect 264973 119720 264978 119776
rect 265034 119720 268180 119776
rect 264973 119718 268180 119720
rect 264973 119715 265039 119718
rect 193949 119506 194015 119509
rect 213177 119506 213243 119509
rect 193949 119504 213243 119506
rect 193949 119448 193954 119504
rect 194010 119448 213182 119504
rect 213238 119448 213243 119504
rect 193949 119446 213243 119448
rect 193949 119443 194015 119446
rect 213177 119443 213243 119446
rect 213913 119506 213979 119509
rect 213913 119504 217028 119506
rect 213913 119448 213918 119504
rect 213974 119448 217028 119504
rect 213913 119446 217028 119448
rect 213913 119443 213979 119446
rect 166206 119308 166212 119372
rect 166276 119370 166282 119372
rect 210509 119370 210575 119373
rect 231761 119370 231827 119373
rect 166276 119368 210575 119370
rect 166276 119312 210514 119368
rect 210570 119312 210575 119368
rect 166276 119310 210575 119312
rect 228988 119368 231827 119370
rect 228988 119312 231766 119368
rect 231822 119312 231827 119368
rect 228988 119310 231827 119312
rect 166276 119308 166282 119310
rect 210509 119307 210575 119310
rect 231761 119307 231827 119310
rect 264237 119370 264303 119373
rect 264237 119368 268180 119370
rect 264237 119312 264242 119368
rect 264298 119312 268180 119368
rect 264237 119310 268180 119312
rect 264237 119307 264303 119310
rect 231209 119234 231275 119237
rect 247861 119234 247927 119237
rect 281533 119234 281599 119237
rect 231209 119232 247927 119234
rect 231209 119176 231214 119232
rect 231270 119176 247866 119232
rect 247922 119176 247927 119232
rect 231209 119174 247927 119176
rect 279956 119232 281599 119234
rect 279956 119176 281538 119232
rect 281594 119176 281599 119232
rect 279956 119174 281599 119176
rect 231209 119171 231275 119174
rect 247861 119171 247927 119174
rect 281533 119171 281599 119174
rect 231485 118962 231551 118965
rect 228988 118960 231551 118962
rect 228988 118904 231490 118960
rect 231546 118904 231551 118960
rect 228988 118902 231551 118904
rect 231485 118899 231551 118902
rect 262857 118962 262923 118965
rect 262857 118960 268180 118962
rect 262857 118904 262862 118960
rect 262918 118904 268180 118960
rect 262857 118902 268180 118904
rect 262857 118899 262923 118902
rect 214005 118826 214071 118829
rect 214005 118824 217028 118826
rect 214005 118768 214010 118824
rect 214066 118768 217028 118824
rect 214005 118766 217028 118768
rect 214005 118763 214071 118766
rect 264973 118554 265039 118557
rect 264973 118552 268180 118554
rect 264973 118496 264978 118552
rect 265034 118496 268180 118552
rect 264973 118494 268180 118496
rect 264973 118491 265039 118494
rect 232497 118418 232563 118421
rect 282821 118418 282887 118421
rect 228988 118416 232563 118418
rect 228988 118360 232502 118416
rect 232558 118360 232563 118416
rect 228988 118358 232563 118360
rect 279956 118416 282887 118418
rect 279956 118360 282826 118416
rect 282882 118360 282887 118416
rect 279956 118358 282887 118360
rect 232497 118355 232563 118358
rect 282821 118355 282887 118358
rect 214005 118146 214071 118149
rect 214005 118144 217028 118146
rect 214005 118088 214010 118144
rect 214066 118088 217028 118144
rect 214005 118086 217028 118088
rect 214005 118083 214071 118086
rect 231393 118010 231459 118013
rect 228988 118008 231459 118010
rect 228988 117952 231398 118008
rect 231454 117952 231459 118008
rect 228988 117950 231459 117952
rect 231393 117947 231459 117950
rect 234153 117874 234219 117877
rect 268150 117874 268210 118116
rect 282729 118010 282795 118013
rect 302325 118010 302391 118013
rect 282729 118008 302391 118010
rect 282729 117952 282734 118008
rect 282790 117952 302330 118008
rect 302386 117952 302391 118008
rect 282729 117950 302391 117952
rect 282729 117947 282795 117950
rect 302325 117947 302391 117950
rect 234153 117872 268210 117874
rect 234153 117816 234158 117872
rect 234214 117816 268210 117872
rect 234153 117814 268210 117816
rect 234153 117811 234219 117814
rect 213913 117466 213979 117469
rect 231761 117466 231827 117469
rect 213913 117464 217028 117466
rect 213913 117408 213918 117464
rect 213974 117408 217028 117464
rect 213913 117406 217028 117408
rect 228988 117464 231827 117466
rect 228988 117408 231766 117464
rect 231822 117408 231827 117464
rect 228988 117406 231827 117408
rect 213913 117403 213979 117406
rect 231761 117403 231827 117406
rect 238017 117466 238083 117469
rect 268150 117466 268210 117708
rect 282821 117602 282887 117605
rect 279956 117600 282887 117602
rect 279956 117544 282826 117600
rect 282882 117544 282887 117600
rect 279956 117542 282887 117544
rect 282821 117539 282887 117542
rect 238017 117464 268210 117466
rect 238017 117408 238022 117464
rect 238078 117408 268210 117464
rect 238017 117406 268210 117408
rect 238017 117403 238083 117406
rect 290641 117332 290707 117333
rect 290590 117330 290596 117332
rect 290550 117270 290596 117330
rect 290660 117328 290707 117332
rect 290702 117272 290707 117328
rect 290590 117268 290596 117270
rect 290660 117268 290707 117272
rect 290641 117267 290707 117268
rect 231301 117194 231367 117197
rect 230246 117192 231367 117194
rect 230246 117136 231306 117192
rect 231362 117136 231367 117192
rect 230246 117134 231367 117136
rect 230246 117058 230306 117134
rect 231301 117131 231367 117134
rect 265065 117194 265131 117197
rect 265065 117192 268180 117194
rect 265065 117136 265070 117192
rect 265126 117136 268180 117192
rect 265065 117134 268180 117136
rect 265065 117131 265131 117134
rect 228988 116998 230306 117058
rect 282821 116922 282887 116925
rect 279956 116920 282887 116922
rect 279956 116864 282826 116920
rect 282882 116864 282887 116920
rect 279956 116862 282887 116864
rect 282821 116859 282887 116862
rect 214005 116786 214071 116789
rect 264973 116786 265039 116789
rect 214005 116784 217028 116786
rect 214005 116728 214010 116784
rect 214066 116728 217028 116784
rect 214005 116726 217028 116728
rect 264973 116784 268180 116786
rect 264973 116728 264978 116784
rect 265034 116728 268180 116784
rect 264973 116726 268180 116728
rect 214005 116723 214071 116726
rect 264973 116723 265039 116726
rect 230933 116514 230999 116517
rect 228988 116512 230999 116514
rect 228988 116456 230938 116512
rect 230994 116456 230999 116512
rect 228988 116454 230999 116456
rect 230933 116451 230999 116454
rect 231117 116514 231183 116517
rect 239581 116514 239647 116517
rect 231117 116512 239647 116514
rect 231117 116456 231122 116512
rect 231178 116456 239586 116512
rect 239642 116456 239647 116512
rect 231117 116454 239647 116456
rect 231117 116451 231183 116454
rect 239581 116451 239647 116454
rect 213913 116106 213979 116109
rect 230749 116106 230815 116109
rect 213913 116104 217028 116106
rect 213913 116048 213918 116104
rect 213974 116048 217028 116104
rect 213913 116046 217028 116048
rect 228988 116104 230815 116106
rect 228988 116048 230754 116104
rect 230810 116048 230815 116104
rect 228988 116046 230815 116048
rect 213913 116043 213979 116046
rect 230749 116043 230815 116046
rect 243537 116106 243603 116109
rect 268150 116106 268210 116348
rect 282729 116106 282795 116109
rect 243537 116104 268210 116106
rect 243537 116048 243542 116104
rect 243598 116048 268210 116104
rect 243537 116046 268210 116048
rect 279956 116104 282795 116106
rect 279956 116048 282734 116104
rect 282790 116048 282795 116104
rect 279956 116046 282795 116048
rect 243537 116043 243603 116046
rect 282729 116043 282795 116046
rect 235257 115970 235323 115973
rect 235257 115968 268180 115970
rect 235257 115912 235262 115968
rect 235318 115912 268180 115968
rect 235257 115910 268180 115912
rect 235257 115907 235323 115910
rect 231761 115562 231827 115565
rect 228988 115560 231827 115562
rect 228988 115504 231766 115560
rect 231822 115504 231827 115560
rect 228988 115502 231827 115504
rect 231761 115499 231827 115502
rect 214005 115426 214071 115429
rect 214005 115424 217028 115426
rect 214005 115368 214010 115424
rect 214066 115368 217028 115424
rect 214005 115366 217028 115368
rect 214005 115363 214071 115366
rect 268150 115290 268210 115532
rect 282821 115426 282887 115429
rect 279956 115424 282887 115426
rect 279956 115368 282826 115424
rect 282882 115368 282887 115424
rect 279956 115366 282887 115368
rect 282821 115363 282887 115366
rect 258030 115230 268210 115290
rect 231209 115154 231275 115157
rect 228988 115152 231275 115154
rect 228988 115096 231214 115152
rect 231270 115096 231275 115152
rect 228988 115094 231275 115096
rect 231209 115091 231275 115094
rect 213913 114882 213979 114885
rect 213913 114880 217028 114882
rect 213913 114824 213918 114880
rect 213974 114824 217028 114880
rect 213913 114822 217028 114824
rect 213913 114819 213979 114822
rect 229686 114820 229692 114884
rect 229756 114882 229762 114884
rect 258030 114882 258090 115230
rect 265065 115154 265131 115157
rect 265065 115152 268180 115154
rect 265065 115096 265070 115152
rect 265126 115096 268180 115152
rect 265065 115094 268180 115096
rect 265065 115091 265131 115094
rect 229756 114822 258090 114882
rect 229756 114820 229762 114822
rect 231025 114610 231091 114613
rect 228988 114608 231091 114610
rect 228988 114552 231030 114608
rect 231086 114552 231091 114608
rect 228988 114550 231091 114552
rect 231025 114547 231091 114550
rect 264973 114610 265039 114613
rect 282637 114610 282703 114613
rect 264973 114608 268180 114610
rect 264973 114552 264978 114608
rect 265034 114552 268180 114608
rect 264973 114550 268180 114552
rect 279956 114608 282703 114610
rect 279956 114552 282642 114608
rect 282698 114552 282703 114608
rect 279956 114550 282703 114552
rect 264973 114547 265039 114550
rect 282637 114547 282703 114550
rect 260281 114474 260347 114477
rect 238710 114472 260347 114474
rect 238710 114416 260286 114472
rect 260342 114416 260347 114472
rect 238710 114414 260347 114416
rect 213913 114202 213979 114205
rect 238710 114202 238770 114414
rect 260281 114411 260347 114414
rect 213913 114200 217028 114202
rect 213913 114144 213918 114200
rect 213974 114144 217028 114200
rect 213913 114142 217028 114144
rect 228988 114142 238770 114202
rect 213913 114139 213979 114142
rect 268150 113930 268210 114172
rect 258030 113870 268210 113930
rect 231577 113658 231643 113661
rect 228988 113656 231643 113658
rect 228988 113600 231582 113656
rect 231638 113600 231643 113656
rect 228988 113598 231643 113600
rect 231577 113595 231643 113598
rect 232681 113522 232747 113525
rect 258030 113522 258090 113870
rect 265065 113794 265131 113797
rect 282821 113794 282887 113797
rect 265065 113792 268180 113794
rect 265065 113736 265070 113792
rect 265126 113736 268180 113792
rect 265065 113734 268180 113736
rect 279956 113792 282887 113794
rect 279956 113736 282826 113792
rect 282882 113736 282887 113792
rect 279956 113734 282887 113736
rect 265065 113731 265131 113734
rect 282821 113731 282887 113734
rect 232681 113520 258090 113522
rect 202229 113386 202295 113389
rect 216998 113386 217058 113492
rect 232681 113464 232686 113520
rect 232742 113464 258090 113520
rect 232681 113462 258090 113464
rect 232681 113459 232747 113462
rect 202229 113384 217058 113386
rect 202229 113328 202234 113384
rect 202290 113328 217058 113384
rect 202229 113326 217058 113328
rect 264973 113386 265039 113389
rect 264973 113384 268180 113386
rect 264973 113328 264978 113384
rect 265034 113328 268180 113384
rect 264973 113326 268180 113328
rect 202229 113323 202295 113326
rect 264973 113323 265039 113326
rect 230565 113250 230631 113253
rect 228988 113248 230631 113250
rect 228988 113192 230570 113248
rect 230626 113192 230631 113248
rect 228988 113190 230631 113192
rect 230565 113187 230631 113190
rect 282821 113114 282887 113117
rect 279956 113112 282887 113114
rect 279956 113056 282826 113112
rect 282882 113056 282887 113112
rect 279956 113054 282887 113056
rect 282821 113051 282887 113054
rect 214005 112842 214071 112845
rect 214005 112840 217028 112842
rect 214005 112784 214010 112840
rect 214066 112784 217028 112840
rect 214005 112782 217028 112784
rect 214005 112779 214071 112782
rect 231761 112706 231827 112709
rect 268150 112706 268210 112948
rect 582833 112842 582899 112845
rect 583520 112842 584960 112932
rect 582833 112840 584960 112842
rect 582833 112784 582838 112840
rect 582894 112784 584960 112840
rect 582833 112782 584960 112784
rect 582833 112779 582899 112782
rect 228988 112704 231827 112706
rect 228988 112648 231766 112704
rect 231822 112648 231827 112704
rect 228988 112646 231827 112648
rect 231761 112643 231827 112646
rect 262814 112646 268210 112706
rect 583520 112692 584960 112782
rect 232497 112434 232563 112437
rect 260465 112434 260531 112437
rect 232497 112432 260531 112434
rect 232497 112376 232502 112432
rect 232558 112376 260470 112432
rect 260526 112376 260531 112432
rect 232497 112374 260531 112376
rect 232497 112371 232563 112374
rect 260465 112371 260531 112374
rect 231669 112298 231735 112301
rect 228988 112296 231735 112298
rect 228988 112240 231674 112296
rect 231730 112240 231735 112296
rect 228988 112238 231735 112240
rect 231669 112235 231735 112238
rect 213913 112162 213979 112165
rect 253197 112162 253263 112165
rect 262814 112162 262874 112646
rect 264973 112570 265039 112573
rect 264973 112568 268180 112570
rect 264973 112512 264978 112568
rect 265034 112512 268180 112568
rect 264973 112510 268180 112512
rect 264973 112507 265039 112510
rect 282177 112298 282243 112301
rect 279956 112296 282243 112298
rect 279956 112240 282182 112296
rect 282238 112240 282243 112296
rect 279956 112238 282243 112240
rect 282177 112235 282243 112238
rect 213913 112160 217028 112162
rect 213913 112104 213918 112160
rect 213974 112104 217028 112160
rect 213913 112102 217028 112104
rect 253197 112160 262874 112162
rect 253197 112104 253202 112160
rect 253258 112104 262874 112160
rect 253197 112102 262874 112104
rect 213913 112099 213979 112102
rect 253197 112099 253263 112102
rect 265985 112026 266051 112029
rect 265985 112024 268180 112026
rect 265985 111968 265990 112024
rect 266046 111968 268180 112024
rect 265985 111966 268180 111968
rect 265985 111963 266051 111966
rect 164724 111754 165354 111760
rect 167821 111754 167887 111757
rect 249057 111754 249123 111757
rect 164724 111752 167887 111754
rect 164724 111700 167826 111752
rect 165294 111696 167826 111700
rect 167882 111696 167887 111752
rect 165294 111694 167887 111696
rect 228988 111752 249123 111754
rect 228988 111696 249062 111752
rect 249118 111696 249123 111752
rect 228988 111694 249123 111696
rect 167821 111691 167887 111694
rect 249057 111691 249123 111694
rect 264973 111618 265039 111621
rect 282085 111618 282151 111621
rect 264973 111616 268180 111618
rect 264973 111560 264978 111616
rect 265034 111560 268180 111616
rect 264973 111558 268180 111560
rect 279956 111616 282151 111618
rect 279956 111560 282090 111616
rect 282146 111560 282151 111616
rect 279956 111558 282151 111560
rect 264973 111555 265039 111558
rect 282085 111555 282151 111558
rect 214005 111482 214071 111485
rect 214005 111480 217028 111482
rect 214005 111424 214010 111480
rect 214066 111424 217028 111480
rect 214005 111422 217028 111424
rect 214005 111419 214071 111422
rect 231393 111346 231459 111349
rect 228988 111344 231459 111346
rect 228988 111288 231398 111344
rect 231454 111288 231459 111344
rect 228988 111286 231459 111288
rect 231393 111283 231459 111286
rect 267733 111210 267799 111213
rect 267733 111208 268180 111210
rect 267733 111152 267738 111208
rect 267794 111152 268180 111208
rect 267733 111150 268180 111152
rect 267733 111147 267799 111150
rect 213913 110802 213979 110805
rect 230565 110802 230631 110805
rect 282821 110802 282887 110805
rect 213913 110800 217028 110802
rect -960 110666 480 110756
rect 213913 110744 213918 110800
rect 213974 110744 217028 110800
rect 213913 110742 217028 110744
rect 228988 110800 230631 110802
rect 228988 110744 230570 110800
rect 230626 110744 230631 110800
rect 228988 110742 230631 110744
rect 213913 110739 213979 110742
rect 230565 110739 230631 110742
rect 258030 110742 268180 110802
rect 279956 110800 282887 110802
rect 279956 110744 282826 110800
rect 282882 110744 282887 110800
rect 279956 110742 282887 110744
rect 3141 110666 3207 110669
rect -960 110664 3207 110666
rect -960 110608 3146 110664
rect 3202 110608 3207 110664
rect -960 110606 3207 110608
rect -960 110516 480 110606
rect 3141 110603 3207 110606
rect 249333 110666 249399 110669
rect 258030 110666 258090 110742
rect 282821 110739 282887 110742
rect 249333 110664 258090 110666
rect 249333 110608 249338 110664
rect 249394 110608 258090 110664
rect 249333 110606 258090 110608
rect 249333 110603 249399 110606
rect 258717 110394 258783 110397
rect 228988 110392 258783 110394
rect 228988 110336 258722 110392
rect 258778 110336 258783 110392
rect 228988 110334 258783 110336
rect 258717 110331 258783 110334
rect 265065 110394 265131 110397
rect 265065 110392 268180 110394
rect 265065 110336 265070 110392
rect 265126 110336 268180 110392
rect 265065 110334 268180 110336
rect 265065 110331 265131 110334
rect 214005 110258 214071 110261
rect 214005 110256 217028 110258
rect 214005 110200 214010 110256
rect 214066 110200 217028 110256
rect 214005 110198 217028 110200
rect 214005 110195 214071 110198
rect 164724 110122 165354 110128
rect 168189 110122 168255 110125
rect 164724 110120 168255 110122
rect 164724 110068 168194 110120
rect 165294 110064 168194 110068
rect 168250 110064 168255 110120
rect 165294 110062 168255 110064
rect 168189 110059 168255 110062
rect 264329 109986 264395 109989
rect 281717 109986 281783 109989
rect 264329 109984 268180 109986
rect 264329 109928 264334 109984
rect 264390 109928 268180 109984
rect 264329 109926 268180 109928
rect 279956 109984 281783 109986
rect 279956 109928 281722 109984
rect 281778 109928 281783 109984
rect 279956 109926 281783 109928
rect 264329 109923 264395 109926
rect 281717 109923 281783 109926
rect 230749 109850 230815 109853
rect 228988 109848 230815 109850
rect 228988 109792 230754 109848
rect 230810 109792 230815 109848
rect 228988 109790 230815 109792
rect 230749 109787 230815 109790
rect 213913 109578 213979 109581
rect 213913 109576 217028 109578
rect 213913 109520 213918 109576
rect 213974 109520 217028 109576
rect 213913 109518 217028 109520
rect 258030 109518 268180 109578
rect 213913 109515 213979 109518
rect 231761 109442 231827 109445
rect 228988 109440 231827 109442
rect 228988 109384 231766 109440
rect 231822 109384 231827 109440
rect 228988 109382 231827 109384
rect 231761 109379 231827 109382
rect 245101 109442 245167 109445
rect 258030 109442 258090 109518
rect 245101 109440 258090 109442
rect 245101 109384 245106 109440
rect 245162 109384 258090 109440
rect 245101 109382 258090 109384
rect 245101 109379 245167 109382
rect 282637 109306 282703 109309
rect 279956 109304 282703 109306
rect 279956 109248 282642 109304
rect 282698 109248 282703 109304
rect 279956 109246 282703 109248
rect 282637 109243 282703 109246
rect 259361 109170 259427 109173
rect 263542 109170 263548 109172
rect 259361 109168 263548 109170
rect 259361 109112 259366 109168
rect 259422 109112 263548 109168
rect 259361 109110 263548 109112
rect 259361 109107 259427 109110
rect 263542 109108 263548 109110
rect 263612 109108 263618 109172
rect 264973 109034 265039 109037
rect 264973 109032 268180 109034
rect 264973 108976 264978 109032
rect 265034 108976 268180 109032
rect 264973 108974 268180 108976
rect 264973 108971 265039 108974
rect 214005 108898 214071 108901
rect 245193 108898 245259 108901
rect 214005 108896 217028 108898
rect 214005 108840 214010 108896
rect 214066 108840 217028 108896
rect 214005 108838 217028 108840
rect 228988 108896 245259 108898
rect 228988 108840 245198 108896
rect 245254 108840 245259 108896
rect 228988 108838 245259 108840
rect 214005 108835 214071 108838
rect 245193 108835 245259 108838
rect 164724 108762 165354 108768
rect 167913 108762 167979 108765
rect 164724 108760 167979 108762
rect 164724 108708 167918 108760
rect 165294 108704 167918 108708
rect 167974 108704 167979 108760
rect 165294 108702 167979 108704
rect 167913 108699 167979 108702
rect 265341 108626 265407 108629
rect 265341 108624 268180 108626
rect 265341 108568 265346 108624
rect 265402 108568 268180 108624
rect 265341 108566 268180 108568
rect 265341 108563 265407 108566
rect 231761 108490 231827 108493
rect 281717 108490 281783 108493
rect 228988 108488 231827 108490
rect 228988 108432 231766 108488
rect 231822 108432 231827 108488
rect 228988 108430 231827 108432
rect 279956 108488 281783 108490
rect 279956 108432 281722 108488
rect 281778 108432 281783 108488
rect 279956 108430 281783 108432
rect 231761 108427 231827 108430
rect 281717 108427 281783 108430
rect 213913 108218 213979 108221
rect 213913 108216 217028 108218
rect 213913 108160 213918 108216
rect 213974 108160 217028 108216
rect 213913 108158 217028 108160
rect 213913 108155 213979 108158
rect 231485 107946 231551 107949
rect 228988 107944 231551 107946
rect 228988 107888 231490 107944
rect 231546 107888 231551 107944
rect 228988 107886 231551 107888
rect 231485 107883 231551 107886
rect 250529 107946 250595 107949
rect 268150 107946 268210 108188
rect 250529 107944 268210 107946
rect 250529 107888 250534 107944
rect 250590 107888 268210 107944
rect 250529 107886 268210 107888
rect 250529 107883 250595 107886
rect 262121 107810 262187 107813
rect 282821 107810 282887 107813
rect 262121 107808 268180 107810
rect 262121 107752 262126 107808
rect 262182 107752 268180 107808
rect 262121 107750 268180 107752
rect 279956 107808 282887 107810
rect 279956 107752 282826 107808
rect 282882 107752 282887 107808
rect 279956 107750 282887 107752
rect 262121 107747 262187 107750
rect 282821 107747 282887 107750
rect 214005 107538 214071 107541
rect 250621 107538 250687 107541
rect 214005 107536 217028 107538
rect 214005 107480 214010 107536
rect 214066 107480 217028 107536
rect 214005 107478 217028 107480
rect 228988 107536 250687 107538
rect 228988 107480 250626 107536
rect 250682 107480 250687 107536
rect 228988 107478 250687 107480
rect 214005 107475 214071 107478
rect 250621 107475 250687 107478
rect 264973 107402 265039 107405
rect 264973 107400 268180 107402
rect 264973 107344 264978 107400
rect 265034 107344 268180 107400
rect 264973 107342 268180 107344
rect 264973 107339 265039 107342
rect 231761 107130 231827 107133
rect 228988 107128 231827 107130
rect 228988 107072 231766 107128
rect 231822 107072 231827 107128
rect 228988 107070 231827 107072
rect 231761 107067 231827 107070
rect 282821 106994 282887 106997
rect 279956 106992 282887 106994
rect 213913 106858 213979 106861
rect 213913 106856 217028 106858
rect 213913 106800 213918 106856
rect 213974 106800 217028 106856
rect 213913 106798 217028 106800
rect 213913 106795 213979 106798
rect 231485 106586 231551 106589
rect 228988 106584 231551 106586
rect 228988 106528 231490 106584
rect 231546 106528 231551 106584
rect 228988 106526 231551 106528
rect 231485 106523 231551 106526
rect 256049 106586 256115 106589
rect 268150 106586 268210 106964
rect 279956 106936 282826 106992
rect 282882 106936 282887 106992
rect 279956 106934 282887 106936
rect 282821 106931 282887 106934
rect 256049 106584 268210 106586
rect 256049 106528 256054 106584
rect 256110 106528 268210 106584
rect 256049 106526 268210 106528
rect 256049 106523 256115 106526
rect 264881 106450 264947 106453
rect 264881 106448 268180 106450
rect 264881 106392 264886 106448
rect 264942 106392 268180 106448
rect 264881 106390 268180 106392
rect 264881 106387 264947 106390
rect 214005 106178 214071 106181
rect 229829 106178 229895 106181
rect 282821 106178 282887 106181
rect 214005 106176 217028 106178
rect 214005 106120 214010 106176
rect 214066 106120 217028 106176
rect 214005 106118 217028 106120
rect 228988 106176 229895 106178
rect 228988 106120 229834 106176
rect 229890 106120 229895 106176
rect 228988 106118 229895 106120
rect 279956 106176 282887 106178
rect 279956 106120 282826 106176
rect 282882 106120 282887 106176
rect 279956 106118 282887 106120
rect 214005 106115 214071 106118
rect 229829 106115 229895 106118
rect 282821 106115 282887 106118
rect 260281 105770 260347 105773
rect 268150 105770 268210 106012
rect 260281 105768 268210 105770
rect 260281 105712 260286 105768
rect 260342 105712 268210 105768
rect 260281 105710 268210 105712
rect 260281 105707 260347 105710
rect 231761 105634 231827 105637
rect 228988 105632 231827 105634
rect 209221 105226 209287 105229
rect 216998 105226 217058 105604
rect 228988 105576 231766 105632
rect 231822 105576 231827 105632
rect 228988 105574 231827 105576
rect 231761 105571 231827 105574
rect 238109 105498 238175 105501
rect 244958 105498 244964 105500
rect 238109 105496 244964 105498
rect 238109 105440 238114 105496
rect 238170 105440 244964 105496
rect 238109 105438 244964 105440
rect 238109 105435 238175 105438
rect 244958 105436 244964 105438
rect 245028 105436 245034 105500
rect 233969 105362 234035 105365
rect 268150 105362 268210 105604
rect 282821 105498 282887 105501
rect 279956 105496 282887 105498
rect 279956 105440 282826 105496
rect 282882 105440 282887 105496
rect 279956 105438 282887 105440
rect 282821 105435 282887 105438
rect 233969 105360 268210 105362
rect 233969 105304 233974 105360
rect 234030 105304 268210 105360
rect 233969 105302 268210 105304
rect 233969 105299 234035 105302
rect 230933 105226 230999 105229
rect 209221 105224 217058 105226
rect 209221 105168 209226 105224
rect 209282 105168 217058 105224
rect 209221 105166 217058 105168
rect 228988 105224 230999 105226
rect 228988 105168 230938 105224
rect 230994 105168 230999 105224
rect 228988 105166 230999 105168
rect 209221 105163 209287 105166
rect 230933 105163 230999 105166
rect 264973 105226 265039 105229
rect 264973 105224 268180 105226
rect 264973 105168 264978 105224
rect 265034 105168 268180 105224
rect 264973 105166 268180 105168
rect 264973 105163 265039 105166
rect 213913 104954 213979 104957
rect 213913 104952 217028 104954
rect 213913 104896 213918 104952
rect 213974 104896 217028 104952
rect 213913 104894 217028 104896
rect 213913 104891 213979 104894
rect 242433 104682 242499 104685
rect 228988 104680 242499 104682
rect 228988 104624 242438 104680
rect 242494 104624 242499 104680
rect 228988 104622 242499 104624
rect 242433 104619 242499 104622
rect 268150 104546 268210 104788
rect 282821 104682 282887 104685
rect 279956 104680 282887 104682
rect 279956 104624 282826 104680
rect 282882 104624 282887 104680
rect 279956 104622 282887 104624
rect 282821 104619 282887 104622
rect 258030 104486 268210 104546
rect 213913 104274 213979 104277
rect 230933 104274 230999 104277
rect 213913 104272 217028 104274
rect 213913 104216 213918 104272
rect 213974 104216 217028 104272
rect 213913 104214 217028 104216
rect 228988 104272 230999 104274
rect 228988 104216 230938 104272
rect 230994 104216 230999 104272
rect 228988 104214 230999 104216
rect 213913 104211 213979 104214
rect 230933 104211 230999 104214
rect 238201 104002 238267 104005
rect 258030 104002 258090 104486
rect 264973 104410 265039 104413
rect 264973 104408 268180 104410
rect 264973 104352 264978 104408
rect 265034 104352 268180 104408
rect 264973 104350 268180 104352
rect 264973 104347 265039 104350
rect 281533 104002 281599 104005
rect 238201 104000 258090 104002
rect 238201 103944 238206 104000
rect 238262 103944 258090 104000
rect 238201 103942 258090 103944
rect 279956 104000 281599 104002
rect 279956 103944 281538 104000
rect 281594 103944 281599 104000
rect 279956 103942 281599 103944
rect 238201 103939 238267 103942
rect 281533 103939 281599 103942
rect 260046 103804 260052 103868
rect 260116 103866 260122 103868
rect 260116 103806 268180 103866
rect 260116 103804 260122 103806
rect 231301 103730 231367 103733
rect 228988 103728 231367 103730
rect 228988 103672 231306 103728
rect 231362 103672 231367 103728
rect 228988 103670 231367 103672
rect 231301 103667 231367 103670
rect 168230 103532 168236 103596
rect 168300 103594 168306 103596
rect 168300 103534 217028 103594
rect 168300 103532 168306 103534
rect 265065 103458 265131 103461
rect 265065 103456 268180 103458
rect 265065 103400 265070 103456
rect 265126 103400 268180 103456
rect 265065 103398 268180 103400
rect 265065 103395 265131 103398
rect 234061 103322 234127 103325
rect 228988 103320 234127 103322
rect 228988 103264 234066 103320
rect 234122 103264 234127 103320
rect 228988 103262 234127 103264
rect 234061 103259 234127 103262
rect 282085 103186 282151 103189
rect 279956 103184 282151 103186
rect 279956 103128 282090 103184
rect 282146 103128 282151 103184
rect 279956 103126 282151 103128
rect 282085 103123 282151 103126
rect 263542 102988 263548 103052
rect 263612 103050 263618 103052
rect 263612 102990 268180 103050
rect 263612 102988 263618 102990
rect 213913 102914 213979 102917
rect 213913 102912 217028 102914
rect 213913 102856 213918 102912
rect 213974 102856 217028 102912
rect 213913 102854 217028 102856
rect 213913 102851 213979 102854
rect 231761 102778 231827 102781
rect 228988 102776 231827 102778
rect 228988 102720 231766 102776
rect 231822 102720 231827 102776
rect 228988 102718 231827 102720
rect 231761 102715 231827 102718
rect 264973 102642 265039 102645
rect 264973 102640 268180 102642
rect 264973 102584 264978 102640
rect 265034 102584 268180 102640
rect 264973 102582 268180 102584
rect 264973 102579 265039 102582
rect 65885 102370 65951 102373
rect 68142 102370 68816 102376
rect 231485 102370 231551 102373
rect 285806 102370 285812 102372
rect 65885 102368 68816 102370
rect 65885 102312 65890 102368
rect 65946 102316 68816 102368
rect 228988 102368 231551 102370
rect 65946 102312 68202 102316
rect 65885 102310 68202 102312
rect 228988 102312 231490 102368
rect 231546 102312 231551 102368
rect 228988 102310 231551 102312
rect 279956 102310 285812 102370
rect 65885 102307 65951 102310
rect 231485 102307 231551 102310
rect 285806 102308 285812 102310
rect 285876 102308 285882 102372
rect 214005 102234 214071 102237
rect 246481 102234 246547 102237
rect 214005 102232 217028 102234
rect 214005 102176 214010 102232
rect 214066 102176 217028 102232
rect 214005 102174 217028 102176
rect 246481 102232 268180 102234
rect 246481 102176 246486 102232
rect 246542 102176 268180 102232
rect 246481 102174 268180 102176
rect 214005 102171 214071 102174
rect 246481 102171 246547 102174
rect 230657 101826 230723 101829
rect 228988 101824 230723 101826
rect 228988 101768 230662 101824
rect 230718 101768 230723 101824
rect 228988 101766 230723 101768
rect 230657 101763 230723 101766
rect 264973 101826 265039 101829
rect 264973 101824 268180 101826
rect 264973 101768 264978 101824
rect 265034 101768 268180 101824
rect 264973 101766 268180 101768
rect 264973 101763 265039 101766
rect 282269 101690 282335 101693
rect 279956 101688 282335 101690
rect 279956 101632 282274 101688
rect 282330 101632 282335 101688
rect 279956 101630 282335 101632
rect 282269 101627 282335 101630
rect 214005 101554 214071 101557
rect 231301 101554 231367 101557
rect 250713 101554 250779 101557
rect 214005 101552 217028 101554
rect 214005 101496 214010 101552
rect 214066 101496 217028 101552
rect 214005 101494 217028 101496
rect 231301 101552 250779 101554
rect 231301 101496 231306 101552
rect 231362 101496 250718 101552
rect 250774 101496 250779 101552
rect 231301 101494 250779 101496
rect 214005 101491 214071 101494
rect 231301 101491 231367 101494
rect 250713 101491 250779 101494
rect 230565 101418 230631 101421
rect 228988 101416 230631 101418
rect 228988 101360 230570 101416
rect 230626 101360 230631 101416
rect 228988 101358 230631 101360
rect 230565 101355 230631 101358
rect 265065 101282 265131 101285
rect 265065 101280 268180 101282
rect 265065 101224 265070 101280
rect 265126 101224 268180 101280
rect 265065 101222 268180 101224
rect 265065 101219 265131 101222
rect 213913 101010 213979 101013
rect 213913 101008 217028 101010
rect 213913 100952 213918 101008
rect 213974 100952 217028 101008
rect 213913 100950 217028 100952
rect 213913 100947 213979 100950
rect 231669 100874 231735 100877
rect 228988 100872 231735 100874
rect 228988 100816 231674 100872
rect 231730 100816 231735 100872
rect 228988 100814 231735 100816
rect 231669 100811 231735 100814
rect 253381 100874 253447 100877
rect 281533 100874 281599 100877
rect 253381 100872 268180 100874
rect 253381 100816 253386 100872
rect 253442 100816 268180 100872
rect 253381 100814 268180 100816
rect 279956 100872 281599 100874
rect 279956 100816 281538 100872
rect 281594 100816 281599 100872
rect 279956 100814 281599 100816
rect 253381 100811 253447 100814
rect 281533 100811 281599 100814
rect 67725 100738 67791 100741
rect 68142 100738 68816 100744
rect 67725 100736 68816 100738
rect 67725 100680 67730 100736
rect 67786 100684 68816 100736
rect 231669 100738 231735 100741
rect 244774 100738 244780 100740
rect 231669 100736 244780 100738
rect 67786 100680 68202 100684
rect 67725 100678 68202 100680
rect 231669 100680 231674 100736
rect 231730 100680 244780 100736
rect 231669 100678 244780 100680
rect 67725 100675 67791 100678
rect 231669 100675 231735 100678
rect 244774 100676 244780 100678
rect 244844 100676 244850 100740
rect 279325 100602 279391 100605
rect 279325 100600 279434 100602
rect 279325 100544 279330 100600
rect 279386 100544 279434 100600
rect 279325 100539 279434 100544
rect 230657 100466 230723 100469
rect 228988 100464 230723 100466
rect 228988 100408 230662 100464
rect 230718 100408 230723 100464
rect 228988 100406 230723 100408
rect 230657 100403 230723 100406
rect 267641 100466 267707 100469
rect 267641 100464 268180 100466
rect 267641 100408 267646 100464
rect 267702 100408 268180 100464
rect 267641 100406 268180 100408
rect 267641 100403 267707 100406
rect 214097 100330 214163 100333
rect 214097 100328 217028 100330
rect 214097 100272 214102 100328
rect 214158 100272 217028 100328
rect 214097 100270 217028 100272
rect 214097 100267 214163 100270
rect 279374 100164 279434 100539
rect 196709 100058 196775 100061
rect 214005 100058 214071 100061
rect 196709 100056 214071 100058
rect 196709 100000 196714 100056
rect 196770 100000 214010 100056
rect 214066 100000 214071 100056
rect 196709 99998 214071 100000
rect 196709 99995 196775 99998
rect 214005 99995 214071 99998
rect 231669 99922 231735 99925
rect 228988 99920 231735 99922
rect 228988 99864 231674 99920
rect 231730 99864 231735 99920
rect 228988 99862 231735 99864
rect 231669 99859 231735 99862
rect 249057 99786 249123 99789
rect 268150 99786 268210 100028
rect 249057 99784 268210 99786
rect 249057 99728 249062 99784
rect 249118 99728 268210 99784
rect 249057 99726 268210 99728
rect 249057 99723 249123 99726
rect 213913 99650 213979 99653
rect 251909 99650 251975 99653
rect 213913 99648 217028 99650
rect 213913 99592 213918 99648
rect 213974 99592 217028 99648
rect 213913 99590 217028 99592
rect 251909 99648 268180 99650
rect 251909 99592 251914 99648
rect 251970 99592 268180 99648
rect 251909 99590 268180 99592
rect 213913 99587 213979 99590
rect 251909 99587 251975 99590
rect 231761 99514 231827 99517
rect 228988 99512 231827 99514
rect 228988 99456 231766 99512
rect 231822 99456 231827 99512
rect 228988 99454 231827 99456
rect 231761 99451 231827 99454
rect 583017 99514 583083 99517
rect 583520 99514 584960 99604
rect 583017 99512 584960 99514
rect 583017 99456 583022 99512
rect 583078 99456 584960 99512
rect 583017 99454 584960 99456
rect 583017 99451 583083 99454
rect 281625 99378 281691 99381
rect 279956 99376 281691 99378
rect 279956 99320 281630 99376
rect 281686 99320 281691 99376
rect 583520 99364 584960 99454
rect 279956 99318 281691 99320
rect 281625 99315 281691 99318
rect 265065 99242 265131 99245
rect 265065 99240 268180 99242
rect 265065 99184 265070 99240
rect 265126 99184 268180 99240
rect 265065 99182 268180 99184
rect 265065 99179 265131 99182
rect 231117 98970 231183 98973
rect 228988 98968 231183 98970
rect 200849 98426 200915 98429
rect 216998 98426 217058 98940
rect 228988 98912 231122 98968
rect 231178 98912 231183 98968
rect 228988 98910 231183 98912
rect 231117 98907 231183 98910
rect 265801 98834 265867 98837
rect 258030 98832 265867 98834
rect 258030 98776 265806 98832
rect 265862 98776 265867 98832
rect 258030 98774 265867 98776
rect 254761 98698 254827 98701
rect 258030 98698 258090 98774
rect 265801 98771 265867 98774
rect 254761 98696 258090 98698
rect 254761 98640 254766 98696
rect 254822 98640 258090 98696
rect 254761 98638 258090 98640
rect 264973 98698 265039 98701
rect 264973 98696 268180 98698
rect 264973 98640 264978 98696
rect 265034 98640 268180 98696
rect 264973 98638 268180 98640
rect 254761 98635 254827 98638
rect 264973 98635 265039 98638
rect 232446 98562 232452 98564
rect 228988 98502 232452 98562
rect 232446 98500 232452 98502
rect 232516 98500 232522 98564
rect 200849 98424 217058 98426
rect 200849 98368 200854 98424
rect 200910 98368 217058 98424
rect 200849 98366 217058 98368
rect 200849 98363 200915 98366
rect 213913 98290 213979 98293
rect 265985 98290 266051 98293
rect 213913 98288 217028 98290
rect 213913 98232 213918 98288
rect 213974 98232 217028 98288
rect 213913 98230 217028 98232
rect 265985 98288 268180 98290
rect 265985 98232 265990 98288
rect 266046 98232 268180 98288
rect 265985 98230 268180 98232
rect 213913 98227 213979 98230
rect 265985 98227 266051 98230
rect 279374 98157 279434 98532
rect 279325 98152 279434 98157
rect 279325 98096 279330 98152
rect 279386 98096 279434 98152
rect 279325 98094 279434 98096
rect 279325 98091 279391 98094
rect 237966 98018 237972 98020
rect 228988 97958 237972 98018
rect 237966 97956 237972 97958
rect 238036 97956 238042 98020
rect 229093 97884 229159 97885
rect 229093 97880 229140 97884
rect 229204 97882 229210 97884
rect 265065 97882 265131 97885
rect 281993 97882 282059 97885
rect 229093 97824 229098 97880
rect 229093 97820 229140 97824
rect 229204 97822 229250 97882
rect 265065 97880 268180 97882
rect 265065 97824 265070 97880
rect 265126 97824 268180 97880
rect 265065 97822 268180 97824
rect 279956 97880 282059 97882
rect 279956 97824 281998 97880
rect 282054 97824 282059 97880
rect 279956 97822 282059 97824
rect 229204 97820 229210 97822
rect 229093 97819 229159 97820
rect 265065 97819 265131 97822
rect 281993 97819 282059 97822
rect -960 97610 480 97700
rect 3509 97610 3575 97613
rect -960 97608 3575 97610
rect -960 97552 3514 97608
rect 3570 97552 3575 97608
rect -960 97550 3575 97552
rect -960 97460 480 97550
rect 3509 97547 3575 97550
rect 213913 97610 213979 97613
rect 230749 97610 230815 97613
rect 213913 97608 217028 97610
rect 213913 97552 213918 97608
rect 213974 97552 217028 97608
rect 213913 97550 217028 97552
rect 228988 97608 230815 97610
rect 228988 97552 230754 97608
rect 230810 97552 230815 97608
rect 228988 97550 230815 97552
rect 213913 97547 213979 97550
rect 230749 97547 230815 97550
rect 265709 97474 265775 97477
rect 265709 97472 268180 97474
rect 265709 97416 265714 97472
rect 265770 97416 268180 97472
rect 265709 97414 268180 97416
rect 265709 97411 265775 97414
rect 229185 97204 229251 97205
rect 229134 97202 229140 97204
rect 229094 97142 229140 97202
rect 229204 97200 229251 97204
rect 229246 97144 229251 97200
rect 229134 97140 229140 97142
rect 229204 97140 229251 97144
rect 229185 97139 229251 97140
rect 231117 97066 231183 97069
rect 284334 97066 284340 97068
rect 228988 97064 231778 97066
rect 228988 97008 231122 97064
rect 231178 97008 231778 97064
rect 228988 97006 231778 97008
rect 231117 97003 231183 97006
rect 214649 96930 214715 96933
rect 214649 96928 217028 96930
rect 214649 96872 214654 96928
rect 214710 96872 217028 96928
rect 214649 96870 217028 96872
rect 214649 96867 214715 96870
rect 230565 96658 230631 96661
rect 228988 96656 230631 96658
rect 228988 96600 230570 96656
rect 230626 96600 230631 96656
rect 228988 96598 230631 96600
rect 230565 96595 230631 96598
rect 231718 96522 231778 97006
rect 268518 96796 268578 97036
rect 279956 97006 284340 97066
rect 284334 97004 284340 97006
rect 284404 97004 284410 97068
rect 268510 96732 268516 96796
rect 268580 96732 268586 96796
rect 264973 96658 265039 96661
rect 264973 96656 268180 96658
rect 264973 96600 264978 96656
rect 265034 96600 268180 96656
rect 264973 96598 268180 96600
rect 264973 96595 265039 96598
rect 255313 96522 255379 96525
rect 255865 96522 255931 96525
rect 231718 96520 255931 96522
rect 231718 96464 255318 96520
rect 255374 96464 255870 96520
rect 255926 96464 255931 96520
rect 231718 96462 255931 96464
rect 255313 96459 255379 96462
rect 255865 96459 255931 96462
rect 213913 96386 213979 96389
rect 213913 96384 217028 96386
rect 213913 96328 213918 96384
rect 213974 96328 217028 96384
rect 213913 96326 217028 96328
rect 213913 96323 213979 96326
rect 230473 96250 230539 96253
rect 228988 96248 230539 96250
rect 228988 96192 230478 96248
rect 230534 96192 230539 96248
rect 228988 96190 230539 96192
rect 230473 96187 230539 96190
rect 264973 96250 265039 96253
rect 264973 96248 268180 96250
rect 264973 96192 264978 96248
rect 265034 96192 268180 96248
rect 264973 96190 268180 96192
rect 264973 96187 265039 96190
rect 228357 95842 228423 95845
rect 263542 95842 263548 95844
rect 228357 95840 263548 95842
rect 228357 95784 228362 95840
rect 228418 95784 263548 95840
rect 228357 95782 263548 95784
rect 228357 95779 228423 95782
rect 263542 95780 263548 95782
rect 263612 95780 263618 95844
rect 278773 95842 278839 95845
rect 279374 95842 279434 96356
rect 278773 95840 279434 95842
rect 278773 95784 278778 95840
rect 278834 95784 279434 95840
rect 278773 95782 279434 95784
rect 278773 95779 278839 95782
rect 223614 95508 223620 95572
rect 223684 95570 223690 95572
rect 228950 95570 228956 95572
rect 223684 95510 228956 95570
rect 223684 95508 223690 95510
rect 228950 95508 228956 95510
rect 229020 95508 229026 95572
rect 223430 95372 223436 95436
rect 223500 95434 223506 95436
rect 228766 95434 228772 95436
rect 223500 95374 228772 95434
rect 223500 95372 223506 95374
rect 228766 95372 228772 95374
rect 228836 95372 228842 95436
rect 201350 95100 201356 95164
rect 201420 95162 201426 95164
rect 278773 95162 278839 95165
rect 201420 95160 278839 95162
rect 201420 95104 278778 95160
rect 278834 95104 278839 95160
rect 201420 95102 278839 95104
rect 201420 95100 201426 95102
rect 278773 95099 278839 95102
rect 65885 95026 65951 95029
rect 165521 95026 165587 95029
rect 65885 95024 165587 95026
rect 65885 94968 65890 95024
rect 65946 94968 165526 95024
rect 165582 94968 165587 95024
rect 65885 94966 165587 94968
rect 65885 94963 65951 94966
rect 165521 94963 165587 94966
rect 268510 94964 268516 95028
rect 268580 95026 268586 95028
rect 270585 95026 270651 95029
rect 268580 95024 270651 95026
rect 268580 94968 270590 95024
rect 270646 94968 270651 95024
rect 268580 94966 270651 94968
rect 268580 94964 268586 94966
rect 270585 94963 270651 94966
rect 107745 94756 107811 94757
rect 117129 94756 117195 94757
rect 107696 94692 107702 94756
rect 107766 94754 107811 94756
rect 107766 94752 107858 94754
rect 107806 94696 107858 94752
rect 107766 94694 107858 94696
rect 107766 94692 107811 94694
rect 117080 94692 117086 94756
rect 117150 94754 117195 94756
rect 117150 94752 117242 94754
rect 117190 94696 117242 94752
rect 117150 94694 117242 94696
rect 117150 94692 117195 94694
rect 151486 94692 151492 94756
rect 151556 94754 151562 94756
rect 151760 94754 151766 94756
rect 151556 94694 151766 94754
rect 151556 94692 151562 94694
rect 151760 94692 151766 94694
rect 151830 94692 151836 94756
rect 107745 94691 107811 94692
rect 117129 94691 117195 94692
rect 171961 94482 172027 94485
rect 212441 94482 212507 94485
rect 171961 94480 212507 94482
rect 171961 94424 171966 94480
rect 172022 94424 212446 94480
rect 212502 94424 212507 94480
rect 171961 94422 212507 94424
rect 171961 94419 172027 94422
rect 212441 94419 212507 94422
rect 225597 94482 225663 94485
rect 241053 94482 241119 94485
rect 225597 94480 241119 94482
rect 225597 94424 225602 94480
rect 225658 94424 241058 94480
rect 241114 94424 241119 94480
rect 225597 94422 241119 94424
rect 225597 94419 225663 94422
rect 241053 94419 241119 94422
rect 165429 94210 165495 94213
rect 172145 94210 172211 94213
rect 165429 94208 172211 94210
rect 165429 94152 165434 94208
rect 165490 94152 172150 94208
rect 172206 94152 172211 94208
rect 165429 94150 172211 94152
rect 165429 94147 165495 94150
rect 172145 94147 172211 94150
rect 99598 94012 99604 94076
rect 99668 94074 99674 94076
rect 176193 94074 176259 94077
rect 99668 94072 176259 94074
rect 99668 94016 176198 94072
rect 176254 94016 176259 94072
rect 99668 94014 176259 94016
rect 99668 94012 99674 94014
rect 176193 94011 176259 94014
rect 219382 94012 219388 94076
rect 219452 94012 219458 94076
rect 219390 93941 219450 94012
rect 91318 93876 91324 93940
rect 91388 93938 91394 93940
rect 167821 93938 167887 93941
rect 219341 93938 219450 93941
rect 91388 93936 167887 93938
rect 91388 93880 167826 93936
rect 167882 93880 167887 93936
rect 91388 93878 167887 93880
rect 219296 93936 219450 93938
rect 219296 93880 219346 93936
rect 219402 93880 219450 93936
rect 219296 93878 219450 93880
rect 226977 93938 227043 93941
rect 229921 93938 229987 93941
rect 226977 93936 229987 93938
rect 226977 93880 226982 93936
rect 227038 93880 229926 93936
rect 229982 93880 229987 93936
rect 226977 93878 229987 93880
rect 91388 93876 91394 93878
rect 167821 93875 167887 93878
rect 219341 93875 219407 93878
rect 226977 93875 227043 93878
rect 229921 93875 229987 93878
rect 114318 93740 114324 93804
rect 114388 93802 114394 93804
rect 213361 93802 213427 93805
rect 114388 93800 213427 93802
rect 114388 93744 213366 93800
rect 213422 93744 213427 93800
rect 114388 93742 213427 93744
rect 114388 93740 114394 93742
rect 213361 93739 213427 93742
rect 129406 93604 129412 93668
rect 129476 93666 129482 93668
rect 184381 93666 184447 93669
rect 129476 93664 184447 93666
rect 129476 93608 184386 93664
rect 184442 93608 184447 93664
rect 129476 93606 184447 93608
rect 129476 93604 129482 93606
rect 184381 93603 184447 93606
rect 95049 93532 95115 93533
rect 115841 93532 115907 93533
rect 94998 93530 95004 93532
rect 94958 93470 95004 93530
rect 95068 93528 95115 93532
rect 115790 93530 115796 93532
rect 95110 93472 95115 93528
rect 94998 93468 95004 93470
rect 95068 93468 95115 93472
rect 115750 93470 115796 93530
rect 115860 93528 115907 93532
rect 115902 93472 115907 93528
rect 115790 93468 115796 93470
rect 115860 93468 115907 93472
rect 95049 93467 95115 93468
rect 115841 93467 115907 93468
rect 103329 93260 103395 93261
rect 110321 93260 110387 93261
rect 103278 93258 103284 93260
rect 103238 93198 103284 93258
rect 103348 93256 103395 93260
rect 110270 93258 110276 93260
rect 103390 93200 103395 93256
rect 103278 93196 103284 93198
rect 103348 93196 103395 93200
rect 110230 93198 110276 93258
rect 110340 93256 110387 93260
rect 110382 93200 110387 93256
rect 110270 93196 110276 93198
rect 110340 93196 110387 93200
rect 103329 93195 103395 93196
rect 110321 93195 110387 93196
rect 222929 93258 222995 93261
rect 260046 93258 260052 93260
rect 222929 93256 260052 93258
rect 222929 93200 222934 93256
rect 222990 93200 260052 93256
rect 222929 93198 260052 93200
rect 222929 93195 222995 93198
rect 260046 93196 260052 93198
rect 260116 93196 260122 93260
rect 267590 93196 267596 93260
rect 267660 93258 267666 93260
rect 270493 93258 270559 93261
rect 267660 93256 270559 93258
rect 267660 93200 270498 93256
rect 270554 93200 270559 93256
rect 267660 93198 270559 93200
rect 267660 93196 267666 93198
rect 270493 93195 270559 93198
rect 181529 93122 181595 93125
rect 285673 93122 285739 93125
rect 181529 93120 285739 93122
rect 181529 93064 181534 93120
rect 181590 93064 285678 93120
rect 285734 93064 285739 93120
rect 181529 93062 285739 93064
rect 181529 93059 181595 93062
rect 285673 93059 285739 93062
rect 162209 92578 162275 92581
rect 165521 92578 165587 92581
rect 162209 92576 165587 92578
rect 162209 92520 162214 92576
rect 162270 92520 165526 92576
rect 165582 92520 165587 92576
rect 162209 92518 165587 92520
rect 162209 92515 162275 92518
rect 165521 92515 165587 92518
rect 267774 92516 267780 92580
rect 267844 92578 267850 92580
rect 269113 92578 269179 92581
rect 267844 92576 269179 92578
rect 267844 92520 269118 92576
rect 269174 92520 269179 92576
rect 267844 92518 269179 92520
rect 267844 92516 267850 92518
rect 269113 92515 269179 92518
rect 86769 92444 86835 92445
rect 86718 92442 86724 92444
rect 86678 92382 86724 92442
rect 86788 92440 86835 92444
rect 86830 92384 86835 92440
rect 86718 92380 86724 92382
rect 86788 92380 86835 92384
rect 88926 92380 88932 92444
rect 88996 92442 89002 92444
rect 89069 92442 89135 92445
rect 102041 92444 102107 92445
rect 112345 92444 112411 92445
rect 132401 92444 132467 92445
rect 101990 92442 101996 92444
rect 88996 92440 89135 92442
rect 88996 92384 89074 92440
rect 89130 92384 89135 92440
rect 88996 92382 89135 92384
rect 101950 92382 101996 92442
rect 102060 92440 102107 92444
rect 112294 92442 112300 92444
rect 102102 92384 102107 92440
rect 88996 92380 89002 92382
rect 86769 92379 86835 92380
rect 89069 92379 89135 92382
rect 101990 92380 101996 92382
rect 102060 92380 102107 92384
rect 112254 92382 112300 92442
rect 112364 92440 112411 92444
rect 132350 92442 132356 92444
rect 112406 92384 112411 92440
rect 112294 92380 112300 92382
rect 112364 92380 112411 92384
rect 132310 92382 132356 92442
rect 132420 92440 132467 92444
rect 132462 92384 132467 92440
rect 132350 92380 132356 92382
rect 132420 92380 132467 92384
rect 134374 92380 134380 92444
rect 134444 92442 134450 92444
rect 134701 92442 134767 92445
rect 136081 92444 136147 92445
rect 136030 92442 136036 92444
rect 134444 92440 134767 92442
rect 134444 92384 134706 92440
rect 134762 92384 134767 92440
rect 134444 92382 134767 92384
rect 135990 92382 136036 92442
rect 136100 92440 136147 92444
rect 136142 92384 136147 92440
rect 134444 92380 134450 92382
rect 102041 92379 102107 92380
rect 112345 92379 112411 92380
rect 132401 92379 132467 92380
rect 134701 92379 134767 92382
rect 136030 92380 136036 92382
rect 136100 92380 136147 92384
rect 136081 92379 136147 92380
rect 85798 92244 85804 92308
rect 85868 92306 85874 92308
rect 86125 92306 86191 92309
rect 85868 92304 86191 92306
rect 85868 92248 86130 92304
rect 86186 92248 86191 92304
rect 85868 92246 86191 92248
rect 85868 92244 85874 92246
rect 86125 92243 86191 92246
rect 122046 92244 122052 92308
rect 122116 92306 122122 92308
rect 189717 92306 189783 92309
rect 122116 92304 189783 92306
rect 122116 92248 189722 92304
rect 189778 92248 189783 92304
rect 122116 92246 189783 92248
rect 122116 92244 122122 92246
rect 189717 92243 189783 92246
rect 115422 92108 115428 92172
rect 115492 92170 115498 92172
rect 177573 92170 177639 92173
rect 115492 92168 177639 92170
rect 115492 92112 177578 92168
rect 177634 92112 177639 92168
rect 115492 92110 177639 92112
rect 115492 92108 115498 92110
rect 177573 92107 177639 92110
rect 244917 91898 244983 91901
rect 255814 91898 255820 91900
rect 244917 91896 255820 91898
rect 244917 91840 244922 91896
rect 244978 91840 255820 91896
rect 244917 91838 255820 91840
rect 244917 91835 244983 91838
rect 255814 91836 255820 91838
rect 255884 91836 255890 91900
rect 99046 91700 99052 91764
rect 99116 91762 99122 91764
rect 106917 91762 106983 91765
rect 119705 91764 119771 91765
rect 121729 91764 121795 91765
rect 119654 91762 119660 91764
rect 99116 91760 106983 91762
rect 99116 91704 106922 91760
rect 106978 91704 106983 91760
rect 99116 91702 106983 91704
rect 119614 91702 119660 91762
rect 119724 91760 119771 91764
rect 121678 91762 121684 91764
rect 119766 91704 119771 91760
rect 99116 91700 99122 91702
rect 106917 91699 106983 91702
rect 119654 91700 119660 91702
rect 119724 91700 119771 91704
rect 121638 91702 121684 91762
rect 121748 91760 121795 91764
rect 121790 91704 121795 91760
rect 121678 91700 121684 91702
rect 121748 91700 121795 91704
rect 123150 91700 123156 91764
rect 123220 91762 123226 91764
rect 123753 91762 123819 91765
rect 123220 91760 123819 91762
rect 123220 91704 123758 91760
rect 123814 91704 123819 91760
rect 123220 91702 123819 91704
rect 123220 91700 123226 91702
rect 119705 91699 119771 91700
rect 121729 91699 121795 91700
rect 123753 91699 123819 91702
rect 178534 91700 178540 91764
rect 178604 91762 178610 91764
rect 273253 91762 273319 91765
rect 178604 91760 273319 91762
rect 178604 91704 273258 91760
rect 273314 91704 273319 91760
rect 178604 91702 273319 91704
rect 178604 91700 178610 91702
rect 273253 91699 273319 91702
rect 106406 91564 106412 91628
rect 106476 91626 106482 91628
rect 106641 91626 106707 91629
rect 106476 91624 106707 91626
rect 106476 91568 106646 91624
rect 106702 91568 106707 91624
rect 106476 91566 106707 91568
rect 106476 91564 106482 91566
rect 106641 91563 106707 91566
rect 106774 91564 106780 91628
rect 106844 91626 106850 91628
rect 209129 91626 209195 91629
rect 106844 91624 209195 91626
rect 106844 91568 209134 91624
rect 209190 91568 209195 91624
rect 106844 91566 209195 91568
rect 106844 91564 106850 91566
rect 209129 91563 209195 91566
rect 122782 91428 122788 91492
rect 122852 91490 122858 91492
rect 124029 91490 124095 91493
rect 122852 91488 124095 91490
rect 122852 91432 124034 91488
rect 124090 91432 124095 91488
rect 122852 91430 124095 91432
rect 122852 91428 122858 91430
rect 124029 91427 124095 91430
rect 125726 91428 125732 91492
rect 125796 91490 125802 91492
rect 126789 91490 126855 91493
rect 125796 91488 126855 91490
rect 125796 91432 126794 91488
rect 126850 91432 126855 91488
rect 125796 91430 126855 91432
rect 125796 91428 125802 91430
rect 126789 91427 126855 91430
rect 151537 91490 151603 91493
rect 151670 91490 151676 91492
rect 151537 91488 151676 91490
rect 151537 91432 151542 91488
rect 151598 91432 151676 91488
rect 151537 91430 151676 91432
rect 151537 91427 151603 91430
rect 151670 91428 151676 91430
rect 151740 91428 151746 91492
rect 96654 91292 96660 91356
rect 96724 91354 96730 91356
rect 97809 91354 97875 91357
rect 96724 91352 97875 91354
rect 96724 91296 97814 91352
rect 97870 91296 97875 91352
rect 96724 91294 97875 91296
rect 96724 91292 96730 91294
rect 97809 91291 97875 91294
rect 98126 91292 98132 91356
rect 98196 91354 98202 91356
rect 99281 91354 99347 91357
rect 98196 91352 99347 91354
rect 98196 91296 99286 91352
rect 99342 91296 99347 91352
rect 98196 91294 99347 91296
rect 98196 91292 98202 91294
rect 99281 91291 99347 91294
rect 100886 91292 100892 91356
rect 100956 91354 100962 91356
rect 101857 91354 101923 91357
rect 100956 91352 101923 91354
rect 100956 91296 101862 91352
rect 101918 91296 101923 91352
rect 100956 91294 101923 91296
rect 100956 91292 100962 91294
rect 101857 91291 101923 91294
rect 109166 91292 109172 91356
rect 109236 91354 109242 91356
rect 110229 91354 110295 91357
rect 111241 91356 111307 91357
rect 114369 91356 114435 91357
rect 111190 91354 111196 91356
rect 109236 91352 110295 91354
rect 109236 91296 110234 91352
rect 110290 91296 110295 91352
rect 109236 91294 110295 91296
rect 111150 91294 111196 91354
rect 111260 91352 111307 91356
rect 114318 91354 114324 91356
rect 111302 91296 111307 91352
rect 109236 91292 109242 91294
rect 110229 91291 110295 91294
rect 111190 91292 111196 91294
rect 111260 91292 111307 91296
rect 114278 91294 114324 91354
rect 114388 91352 114435 91356
rect 114430 91296 114435 91352
rect 114318 91292 114324 91294
rect 114388 91292 114435 91296
rect 124438 91292 124444 91356
rect 124508 91354 124514 91356
rect 125501 91354 125567 91357
rect 124508 91352 125567 91354
rect 124508 91296 125506 91352
rect 125562 91296 125567 91352
rect 124508 91294 125567 91296
rect 124508 91292 124514 91294
rect 111241 91291 111307 91292
rect 114369 91291 114435 91292
rect 125501 91291 125567 91294
rect 126646 91292 126652 91356
rect 126716 91354 126722 91356
rect 126881 91354 126947 91357
rect 126716 91352 126947 91354
rect 126716 91296 126886 91352
rect 126942 91296 126947 91352
rect 126716 91294 126947 91296
rect 126716 91292 126722 91294
rect 126881 91291 126947 91294
rect 151302 91292 151308 91356
rect 151372 91354 151378 91356
rect 151721 91354 151787 91357
rect 151372 91352 151787 91354
rect 151372 91296 151726 91352
rect 151782 91296 151787 91352
rect 151372 91294 151787 91296
rect 151372 91292 151378 91294
rect 151721 91291 151787 91294
rect 74758 91156 74764 91220
rect 74828 91218 74834 91220
rect 75729 91218 75795 91221
rect 74828 91216 75795 91218
rect 74828 91160 75734 91216
rect 75790 91160 75795 91216
rect 74828 91158 75795 91160
rect 74828 91156 74834 91158
rect 75729 91155 75795 91158
rect 84326 91156 84332 91220
rect 84396 91218 84402 91220
rect 85481 91218 85547 91221
rect 88057 91220 88123 91221
rect 88006 91218 88012 91220
rect 84396 91216 85547 91218
rect 84396 91160 85486 91216
rect 85542 91160 85547 91216
rect 84396 91158 85547 91160
rect 87966 91158 88012 91218
rect 88076 91216 88123 91220
rect 88118 91160 88123 91216
rect 84396 91156 84402 91158
rect 85481 91155 85547 91158
rect 88006 91156 88012 91158
rect 88076 91156 88123 91160
rect 90214 91156 90220 91220
rect 90284 91218 90290 91220
rect 91001 91218 91067 91221
rect 90284 91216 91067 91218
rect 90284 91160 91006 91216
rect 91062 91160 91067 91216
rect 90284 91158 91067 91160
rect 90284 91156 90290 91158
rect 88057 91155 88123 91156
rect 91001 91155 91067 91158
rect 92606 91156 92612 91220
rect 92676 91218 92682 91220
rect 93761 91218 93827 91221
rect 92676 91216 93827 91218
rect 92676 91160 93766 91216
rect 93822 91160 93827 91216
rect 92676 91158 93827 91160
rect 92676 91156 92682 91158
rect 93761 91155 93827 91158
rect 93894 91156 93900 91220
rect 93964 91218 93970 91220
rect 94681 91218 94747 91221
rect 93964 91216 94747 91218
rect 93964 91160 94686 91216
rect 94742 91160 94747 91216
rect 93964 91158 94747 91160
rect 93964 91156 93970 91158
rect 94681 91155 94747 91158
rect 96286 91156 96292 91220
rect 96356 91218 96362 91220
rect 96521 91218 96587 91221
rect 96356 91216 96587 91218
rect 96356 91160 96526 91216
rect 96582 91160 96587 91216
rect 96356 91158 96587 91160
rect 96356 91156 96362 91158
rect 96521 91155 96587 91158
rect 97206 91156 97212 91220
rect 97276 91218 97282 91220
rect 97901 91218 97967 91221
rect 97276 91216 97967 91218
rect 97276 91160 97906 91216
rect 97962 91160 97967 91216
rect 97276 91158 97967 91160
rect 97276 91156 97282 91158
rect 97901 91155 97967 91158
rect 98494 91156 98500 91220
rect 98564 91218 98570 91220
rect 99189 91218 99255 91221
rect 100569 91220 100635 91221
rect 100518 91218 100524 91220
rect 98564 91216 99255 91218
rect 98564 91160 99194 91216
rect 99250 91160 99255 91216
rect 98564 91158 99255 91160
rect 100478 91158 100524 91218
rect 100588 91216 100635 91220
rect 100630 91160 100635 91216
rect 98564 91156 98570 91158
rect 99189 91155 99255 91158
rect 100518 91156 100524 91158
rect 100588 91156 100635 91160
rect 101806 91156 101812 91220
rect 101876 91218 101882 91220
rect 101949 91218 102015 91221
rect 101876 91216 102015 91218
rect 101876 91160 101954 91216
rect 102010 91160 102015 91216
rect 101876 91158 102015 91160
rect 101876 91156 101882 91158
rect 100569 91155 100635 91156
rect 101949 91155 102015 91158
rect 102726 91156 102732 91220
rect 102796 91218 102802 91220
rect 103421 91218 103487 91221
rect 104249 91220 104315 91221
rect 104198 91218 104204 91220
rect 102796 91216 103487 91218
rect 102796 91160 103426 91216
rect 103482 91160 103487 91216
rect 102796 91158 103487 91160
rect 104158 91158 104204 91218
rect 104268 91216 104315 91220
rect 104310 91160 104315 91216
rect 102796 91156 102802 91158
rect 103421 91155 103487 91158
rect 104198 91156 104204 91158
rect 104268 91156 104315 91160
rect 104566 91156 104572 91220
rect 104636 91218 104642 91220
rect 104801 91218 104867 91221
rect 105537 91220 105603 91221
rect 105486 91218 105492 91220
rect 104636 91216 104867 91218
rect 104636 91160 104806 91216
rect 104862 91160 104867 91216
rect 104636 91158 104867 91160
rect 105446 91158 105492 91218
rect 105556 91216 105603 91220
rect 105598 91160 105603 91216
rect 104636 91156 104642 91158
rect 104249 91155 104315 91156
rect 104801 91155 104867 91158
rect 105486 91156 105492 91158
rect 105556 91156 105603 91160
rect 105670 91156 105676 91220
rect 105740 91218 105746 91220
rect 106089 91218 106155 91221
rect 105740 91216 106155 91218
rect 105740 91160 106094 91216
rect 106150 91160 106155 91216
rect 105740 91158 106155 91160
rect 105740 91156 105746 91158
rect 105537 91155 105603 91156
rect 106089 91155 106155 91158
rect 108062 91156 108068 91220
rect 108132 91218 108138 91220
rect 108941 91218 109007 91221
rect 108132 91216 109007 91218
rect 108132 91160 108946 91216
rect 109002 91160 109007 91216
rect 108132 91158 109007 91160
rect 108132 91156 108138 91158
rect 108941 91155 109007 91158
rect 109534 91156 109540 91220
rect 109604 91218 109610 91220
rect 110137 91218 110203 91221
rect 109604 91216 110203 91218
rect 109604 91160 110142 91216
rect 110198 91160 110203 91216
rect 109604 91158 110203 91160
rect 109604 91156 109610 91158
rect 110137 91155 110203 91158
rect 110638 91156 110644 91220
rect 110708 91218 110714 91220
rect 111701 91218 111767 91221
rect 110708 91216 111767 91218
rect 110708 91160 111706 91216
rect 111762 91160 111767 91216
rect 110708 91158 111767 91160
rect 110708 91156 110714 91158
rect 111701 91155 111767 91158
rect 111926 91156 111932 91220
rect 111996 91218 112002 91220
rect 112989 91218 113055 91221
rect 111996 91216 113055 91218
rect 111996 91160 112994 91216
rect 113050 91160 113055 91216
rect 111996 91158 113055 91160
rect 111996 91156 112002 91158
rect 112989 91155 113055 91158
rect 113214 91156 113220 91220
rect 113284 91218 113290 91220
rect 114461 91218 114527 91221
rect 113284 91216 114527 91218
rect 113284 91160 114466 91216
rect 114522 91160 114527 91216
rect 113284 91158 114527 91160
rect 113284 91156 113290 91158
rect 114461 91155 114527 91158
rect 114870 91156 114876 91220
rect 114940 91218 114946 91220
rect 115841 91218 115907 91221
rect 114940 91216 115907 91218
rect 114940 91160 115846 91216
rect 115902 91160 115907 91216
rect 114940 91158 115907 91160
rect 114940 91156 114946 91158
rect 115841 91155 115907 91158
rect 116710 91156 116716 91220
rect 116780 91218 116786 91220
rect 117221 91218 117287 91221
rect 118049 91220 118115 91221
rect 117998 91218 118004 91220
rect 116780 91216 117287 91218
rect 116780 91160 117226 91216
rect 117282 91160 117287 91216
rect 116780 91158 117287 91160
rect 117958 91158 118004 91218
rect 118068 91216 118115 91220
rect 118110 91160 118115 91216
rect 116780 91156 116786 91158
rect 117221 91155 117287 91158
rect 117998 91156 118004 91158
rect 118068 91156 118115 91160
rect 118182 91156 118188 91220
rect 118252 91218 118258 91220
rect 118601 91218 118667 91221
rect 118252 91216 118667 91218
rect 118252 91160 118606 91216
rect 118662 91160 118667 91216
rect 118252 91158 118667 91160
rect 118252 91156 118258 91158
rect 118049 91155 118115 91156
rect 118601 91155 118667 91158
rect 119286 91156 119292 91220
rect 119356 91218 119362 91220
rect 119889 91218 119955 91221
rect 119356 91216 119955 91218
rect 119356 91160 119894 91216
rect 119950 91160 119955 91216
rect 119356 91158 119955 91160
rect 119356 91156 119362 91158
rect 119889 91155 119955 91158
rect 120206 91156 120212 91220
rect 120276 91218 120282 91220
rect 120441 91218 120507 91221
rect 120276 91216 120507 91218
rect 120276 91160 120446 91216
rect 120502 91160 120507 91216
rect 120276 91158 120507 91160
rect 120276 91156 120282 91158
rect 120441 91155 120507 91158
rect 120574 91156 120580 91220
rect 120644 91218 120650 91220
rect 120809 91218 120875 91221
rect 120644 91216 120875 91218
rect 120644 91160 120814 91216
rect 120870 91160 120875 91216
rect 120644 91158 120875 91160
rect 120644 91156 120650 91158
rect 120809 91155 120875 91158
rect 123937 91218 124003 91221
rect 125409 91220 125475 91221
rect 124070 91218 124076 91220
rect 123937 91216 124076 91218
rect 123937 91160 123942 91216
rect 123998 91160 124076 91216
rect 123937 91158 124076 91160
rect 123937 91155 124003 91158
rect 124070 91156 124076 91158
rect 124140 91156 124146 91220
rect 125358 91218 125364 91220
rect 125318 91158 125364 91218
rect 125428 91216 125475 91220
rect 125470 91160 125475 91216
rect 125358 91156 125364 91158
rect 125428 91156 125475 91160
rect 126462 91156 126468 91220
rect 126532 91218 126538 91220
rect 126697 91218 126763 91221
rect 126532 91216 126763 91218
rect 126532 91160 126702 91216
rect 126758 91160 126763 91216
rect 126532 91158 126763 91160
rect 126532 91156 126538 91158
rect 125409 91155 125475 91156
rect 126697 91155 126763 91158
rect 127566 91156 127572 91220
rect 127636 91218 127642 91220
rect 128261 91218 128327 91221
rect 130745 91220 130811 91221
rect 130694 91218 130700 91220
rect 127636 91216 128327 91218
rect 127636 91160 128266 91216
rect 128322 91160 128327 91216
rect 127636 91158 128327 91160
rect 130654 91158 130700 91218
rect 130764 91216 130811 91220
rect 130806 91160 130811 91216
rect 127636 91156 127642 91158
rect 128261 91155 128327 91158
rect 130694 91156 130700 91158
rect 130764 91156 130811 91160
rect 133086 91156 133092 91220
rect 133156 91218 133162 91220
rect 133781 91218 133847 91221
rect 133156 91216 133847 91218
rect 133156 91160 133786 91216
rect 133842 91160 133847 91216
rect 133156 91158 133847 91160
rect 133156 91156 133162 91158
rect 130745 91155 130811 91156
rect 133781 91155 133847 91158
rect 151486 91156 151492 91220
rect 151556 91218 151562 91220
rect 151629 91218 151695 91221
rect 152089 91220 152155 91221
rect 152038 91218 152044 91220
rect 151556 91216 151695 91218
rect 151556 91160 151634 91216
rect 151690 91160 151695 91216
rect 151556 91158 151695 91160
rect 151998 91158 152044 91218
rect 152108 91216 152155 91220
rect 152150 91160 152155 91216
rect 151556 91156 151562 91158
rect 151629 91155 151695 91158
rect 152038 91156 152044 91158
rect 152108 91156 152155 91160
rect 152089 91155 152155 91156
rect 153101 91082 153167 91085
rect 184289 91082 184355 91085
rect 153101 91080 184355 91082
rect 153101 91024 153106 91080
rect 153162 91024 184294 91080
rect 184350 91024 184355 91080
rect 153101 91022 184355 91024
rect 153101 91019 153167 91022
rect 184289 91019 184355 91022
rect 191189 91082 191255 91085
rect 276013 91082 276079 91085
rect 276749 91082 276815 91085
rect 191189 91080 276815 91082
rect 191189 91024 191194 91080
rect 191250 91024 276018 91080
rect 276074 91024 276754 91080
rect 276810 91024 276815 91080
rect 191189 91022 276815 91024
rect 191189 91019 191255 91022
rect 276013 91019 276079 91022
rect 276749 91019 276815 91022
rect 230565 90946 230631 90949
rect 229050 90944 230631 90946
rect 229050 90888 230570 90944
rect 230626 90888 230631 90944
rect 229050 90886 230631 90888
rect 157977 90538 158043 90541
rect 165429 90538 165495 90541
rect 157977 90536 165495 90538
rect 157977 90480 157982 90536
rect 158038 90480 165434 90536
rect 165490 90480 165495 90536
rect 157977 90478 165495 90480
rect 157977 90475 158043 90478
rect 165429 90475 165495 90478
rect 86125 90402 86191 90405
rect 160093 90402 160159 90405
rect 86125 90400 160159 90402
rect 86125 90344 86130 90400
rect 86186 90344 160098 90400
rect 160154 90344 160159 90400
rect 86125 90342 160159 90344
rect 86125 90339 86191 90342
rect 160093 90339 160159 90342
rect 164969 90402 165035 90405
rect 211889 90402 211955 90405
rect 164969 90400 211955 90402
rect 164969 90344 164974 90400
rect 165030 90344 211894 90400
rect 211950 90344 211955 90400
rect 164969 90342 211955 90344
rect 164969 90339 165035 90342
rect 211889 90339 211955 90342
rect 215150 90340 215156 90404
rect 215220 90402 215226 90404
rect 227662 90402 227668 90404
rect 215220 90342 227668 90402
rect 215220 90340 215226 90342
rect 227662 90340 227668 90342
rect 227732 90402 227738 90404
rect 229050 90402 229110 90886
rect 230565 90883 230631 90886
rect 227732 90342 229110 90402
rect 227732 90340 227738 90342
rect 162117 89858 162183 89861
rect 166206 89858 166212 89860
rect 162117 89856 166212 89858
rect 162117 89800 162122 89856
rect 162178 89800 166212 89856
rect 162117 89798 166212 89800
rect 162117 89795 162183 89798
rect 166206 89796 166212 89798
rect 166276 89796 166282 89860
rect 123753 89722 123819 89725
rect 192569 89722 192635 89725
rect 123753 89720 192635 89722
rect 123753 89664 123758 89720
rect 123814 89664 192574 89720
rect 192630 89664 192635 89720
rect 123753 89662 192635 89664
rect 123753 89659 123819 89662
rect 192569 89659 192635 89662
rect 106641 89586 106707 89589
rect 171869 89586 171935 89589
rect 106641 89584 171935 89586
rect 106641 89528 106646 89584
rect 106702 89528 171874 89584
rect 171930 89528 171935 89584
rect 106641 89526 171935 89528
rect 106641 89523 106707 89526
rect 171869 89523 171935 89526
rect 67449 89042 67515 89045
rect 123477 89042 123543 89045
rect 67449 89040 123543 89042
rect 67449 88984 67454 89040
rect 67510 88984 123482 89040
rect 123538 88984 123543 89040
rect 67449 88982 123543 88984
rect 67449 88979 67515 88982
rect 123477 88979 123543 88982
rect 210417 89042 210483 89045
rect 247953 89042 248019 89045
rect 210417 89040 248019 89042
rect 210417 88984 210422 89040
rect 210478 88984 247958 89040
rect 248014 88984 248019 89040
rect 210417 88982 248019 88984
rect 210417 88979 210483 88982
rect 247953 88979 248019 88982
rect 160093 88226 160159 88229
rect 166533 88226 166599 88229
rect 160093 88224 166599 88226
rect 160093 88168 160098 88224
rect 160154 88168 166538 88224
rect 166594 88168 166599 88224
rect 160093 88166 166599 88168
rect 160093 88163 160159 88166
rect 166533 88163 166599 88166
rect 223430 88164 223436 88228
rect 223500 88226 223506 88228
rect 281533 88226 281599 88229
rect 223500 88224 281599 88226
rect 223500 88168 281538 88224
rect 281594 88168 281599 88224
rect 223500 88166 281599 88168
rect 223500 88164 223506 88166
rect 281533 88163 281599 88166
rect 130745 88090 130811 88093
rect 167637 88090 167703 88093
rect 130745 88088 167703 88090
rect 130745 88032 130750 88088
rect 130806 88032 167642 88088
rect 167698 88032 167703 88088
rect 130745 88030 167703 88032
rect 130745 88027 130811 88030
rect 167637 88027 167703 88030
rect 105537 87954 105603 87957
rect 187233 87954 187299 87957
rect 105537 87952 187299 87954
rect 105537 87896 105542 87952
rect 105598 87896 187238 87952
rect 187294 87896 187299 87952
rect 105537 87894 187299 87896
rect 105537 87891 105603 87894
rect 187233 87891 187299 87894
rect 100569 87546 100635 87549
rect 128997 87546 129063 87549
rect 100569 87544 129063 87546
rect 100569 87488 100574 87544
rect 100630 87488 129002 87544
rect 129058 87488 129063 87544
rect 100569 87486 129063 87488
rect 100569 87483 100635 87486
rect 128997 87483 129063 87486
rect 217225 87546 217291 87549
rect 277393 87546 277459 87549
rect 217225 87544 277459 87546
rect 217225 87488 217230 87544
rect 217286 87488 277398 87544
rect 277454 87488 277459 87544
rect 217225 87486 277459 87488
rect 217225 87483 217291 87486
rect 277393 87483 277459 87486
rect 88057 86866 88123 86869
rect 166441 86866 166507 86869
rect 88057 86864 166507 86866
rect 88057 86808 88062 86864
rect 88118 86808 166446 86864
rect 166502 86808 166507 86864
rect 88057 86806 166507 86808
rect 88057 86803 88123 86806
rect 166441 86803 166507 86806
rect 120073 86730 120139 86733
rect 180149 86730 180215 86733
rect 583753 86730 583819 86733
rect 120073 86728 180215 86730
rect 120073 86672 120078 86728
rect 120134 86672 180154 86728
rect 180210 86672 180215 86728
rect 120073 86670 180215 86672
rect 120073 86667 120139 86670
rect 180149 86667 180215 86670
rect 583710 86728 583819 86730
rect 583710 86672 583758 86728
rect 583814 86672 583819 86728
rect 583710 86667 583819 86672
rect 120441 86594 120507 86597
rect 176009 86594 176075 86597
rect 120441 86592 176075 86594
rect 120441 86536 120446 86592
rect 120502 86536 176014 86592
rect 176070 86536 176075 86592
rect 120441 86534 176075 86536
rect 120441 86531 120507 86534
rect 176009 86531 176075 86534
rect 583710 86322 583770 86667
rect 583342 86276 583770 86322
rect 583342 86262 584960 86276
rect 204989 86186 205055 86189
rect 280153 86186 280219 86189
rect 204989 86184 280219 86186
rect 204989 86128 204994 86184
rect 205050 86128 280158 86184
rect 280214 86128 280219 86184
rect 204989 86126 280219 86128
rect 583342 86186 583402 86262
rect 583520 86186 584960 86262
rect 583342 86126 584960 86186
rect 204989 86123 205055 86126
rect 280153 86123 280219 86126
rect 583520 86036 584960 86126
rect 94681 85506 94747 85509
rect 167913 85506 167979 85509
rect 94681 85504 167979 85506
rect 94681 85448 94686 85504
rect 94742 85448 167918 85504
rect 167974 85448 167979 85504
rect 94681 85446 167979 85448
rect 94681 85443 94747 85446
rect 167913 85443 167979 85446
rect 118049 85370 118115 85373
rect 169293 85370 169359 85373
rect 118049 85368 169359 85370
rect 118049 85312 118054 85368
rect 118110 85312 169298 85368
rect 169354 85312 169359 85368
rect 118049 85310 169359 85312
rect 118049 85307 118115 85310
rect 169293 85307 169359 85310
rect 126237 84826 126303 84829
rect 265617 84826 265683 84829
rect 126237 84824 265683 84826
rect -960 84690 480 84780
rect 126237 84768 126242 84824
rect 126298 84768 265622 84824
rect 265678 84768 265683 84824
rect 126237 84766 265683 84768
rect 126237 84763 126303 84766
rect 265617 84763 265683 84766
rect 3233 84690 3299 84693
rect -960 84688 3299 84690
rect -960 84632 3238 84688
rect 3294 84632 3299 84688
rect -960 84630 3299 84632
rect -960 84540 480 84630
rect 3233 84627 3299 84630
rect 96521 84146 96587 84149
rect 170673 84146 170739 84149
rect 96521 84144 170739 84146
rect 96521 84088 96526 84144
rect 96582 84088 170678 84144
rect 170734 84088 170739 84144
rect 96521 84086 170739 84088
rect 96521 84083 96587 84086
rect 170673 84083 170739 84086
rect 108941 84010 109007 84013
rect 181437 84010 181503 84013
rect 108941 84008 181503 84010
rect 108941 83952 108946 84008
rect 109002 83952 181442 84008
rect 181498 83952 181503 84008
rect 108941 83950 181503 83952
rect 108941 83947 109007 83950
rect 181437 83947 181503 83950
rect 30281 83466 30347 83469
rect 263041 83466 263107 83469
rect 30281 83464 263107 83466
rect 30281 83408 30286 83464
rect 30342 83408 263046 83464
rect 263102 83408 263107 83464
rect 30281 83406 263107 83408
rect 30281 83403 30347 83406
rect 263041 83403 263107 83406
rect 97809 82786 97875 82789
rect 203609 82786 203675 82789
rect 97809 82784 203675 82786
rect 97809 82728 97814 82784
rect 97870 82728 203614 82784
rect 203670 82728 203675 82784
rect 97809 82726 203675 82728
rect 97809 82723 97875 82726
rect 203609 82723 203675 82726
rect 67633 82650 67699 82653
rect 169109 82650 169175 82653
rect 67633 82648 169175 82650
rect 67633 82592 67638 82648
rect 67694 82592 169114 82648
rect 169170 82592 169175 82648
rect 67633 82590 169175 82592
rect 67633 82587 67699 82590
rect 169109 82587 169175 82590
rect 106181 82106 106247 82109
rect 267181 82106 267247 82109
rect 106181 82104 267247 82106
rect 106181 82048 106186 82104
rect 106242 82048 267186 82104
rect 267242 82048 267247 82104
rect 106181 82046 267247 82048
rect 106181 82043 106247 82046
rect 267181 82043 267247 82046
rect 66161 81426 66227 81429
rect 171777 81426 171843 81429
rect 66161 81424 171843 81426
rect 66161 81368 66166 81424
rect 66222 81368 171782 81424
rect 171838 81368 171843 81424
rect 66161 81366 171843 81368
rect 66161 81363 66227 81366
rect 171777 81363 171843 81366
rect 119981 80882 120047 80885
rect 261569 80882 261635 80885
rect 119981 80880 261635 80882
rect 119981 80824 119986 80880
rect 120042 80824 261574 80880
rect 261630 80824 261635 80880
rect 119981 80822 261635 80824
rect 119981 80819 120047 80822
rect 261569 80819 261635 80822
rect 15837 80746 15903 80749
rect 265709 80746 265775 80749
rect 15837 80744 265775 80746
rect 15837 80688 15842 80744
rect 15898 80688 265714 80744
rect 265770 80688 265775 80744
rect 15837 80686 265775 80688
rect 15837 80683 15903 80686
rect 265709 80683 265775 80686
rect 95141 79658 95207 79661
rect 256141 79658 256207 79661
rect 95141 79656 256207 79658
rect 95141 79600 95146 79656
rect 95202 79600 256146 79656
rect 256202 79600 256207 79656
rect 95141 79598 256207 79600
rect 95141 79595 95207 79598
rect 256141 79595 256207 79598
rect 61377 79522 61443 79525
rect 265985 79522 266051 79525
rect 61377 79520 266051 79522
rect 61377 79464 61382 79520
rect 61438 79464 265990 79520
rect 266046 79464 266051 79520
rect 61377 79462 266051 79464
rect 61377 79459 61443 79462
rect 265985 79459 266051 79462
rect 5441 79386 5507 79389
rect 225689 79386 225755 79389
rect 5441 79384 225755 79386
rect 5441 79328 5446 79384
rect 5502 79328 225694 79384
rect 225750 79328 225755 79384
rect 5441 79326 225755 79328
rect 5441 79323 5507 79326
rect 225689 79323 225755 79326
rect 104801 78570 104867 78573
rect 162117 78570 162183 78573
rect 104801 78568 162183 78570
rect 104801 78512 104806 78568
rect 104862 78512 162122 78568
rect 162178 78512 162183 78568
rect 104801 78510 162183 78512
rect 104801 78507 104867 78510
rect 162117 78507 162183 78510
rect 111057 78434 111123 78437
rect 168230 78434 168236 78436
rect 111057 78432 168236 78434
rect 111057 78376 111062 78432
rect 111118 78376 168236 78432
rect 111057 78374 168236 78376
rect 111057 78371 111123 78374
rect 168230 78372 168236 78374
rect 168300 78372 168306 78436
rect 41321 77890 41387 77893
rect 240869 77890 240935 77893
rect 41321 77888 240935 77890
rect 41321 77832 41326 77888
rect 41382 77832 240874 77888
rect 240930 77832 240935 77888
rect 41321 77830 240935 77832
rect 41321 77827 41387 77830
rect 240869 77827 240935 77830
rect 151077 76802 151143 76805
rect 250621 76802 250687 76805
rect 151077 76800 250687 76802
rect 151077 76744 151082 76800
rect 151138 76744 250626 76800
rect 250682 76744 250687 76800
rect 151077 76742 250687 76744
rect 151077 76739 151143 76742
rect 250621 76739 250687 76742
rect 93761 76666 93827 76669
rect 229737 76666 229803 76669
rect 93761 76664 229803 76666
rect 93761 76608 93766 76664
rect 93822 76608 229742 76664
rect 229798 76608 229803 76664
rect 93761 76606 229803 76608
rect 93761 76603 93827 76606
rect 229737 76603 229803 76606
rect 108941 76530 109007 76533
rect 249333 76530 249399 76533
rect 108941 76528 249399 76530
rect 108941 76472 108946 76528
rect 109002 76472 249338 76528
rect 249394 76472 249399 76528
rect 108941 76470 249399 76472
rect 108941 76467 109007 76470
rect 249333 76467 249399 76470
rect 19241 75306 19307 75309
rect 257613 75306 257679 75309
rect 19241 75304 257679 75306
rect 19241 75248 19246 75304
rect 19302 75248 257618 75304
rect 257674 75248 257679 75304
rect 19241 75246 257679 75248
rect 19241 75243 19307 75246
rect 257613 75243 257679 75246
rect 53598 75108 53604 75172
rect 53668 75170 53674 75172
rect 317505 75170 317571 75173
rect 53668 75168 317571 75170
rect 53668 75112 317510 75168
rect 317566 75112 317571 75168
rect 53668 75110 317571 75112
rect 53668 75108 53674 75110
rect 317505 75107 317571 75110
rect 122741 74082 122807 74085
rect 247861 74082 247927 74085
rect 122741 74080 247927 74082
rect 122741 74024 122746 74080
rect 122802 74024 247866 74080
rect 247922 74024 247927 74080
rect 122741 74022 247927 74024
rect 122741 74019 122807 74022
rect 247861 74019 247927 74022
rect 104801 73946 104867 73949
rect 235533 73946 235599 73949
rect 104801 73944 235599 73946
rect 104801 73888 104806 73944
rect 104862 73888 235538 73944
rect 235594 73888 235599 73944
rect 104801 73886 235599 73888
rect 104801 73883 104867 73886
rect 235533 73883 235599 73886
rect 50889 73810 50955 73813
rect 254669 73810 254735 73813
rect 50889 73808 254735 73810
rect 50889 73752 50894 73808
rect 50950 73752 254674 73808
rect 254730 73752 254735 73808
rect 50889 73750 254735 73752
rect 50889 73747 50955 73750
rect 254669 73747 254735 73750
rect 582557 72994 582623 72997
rect 583520 72994 584960 73084
rect 582557 72992 584960 72994
rect 582557 72936 582562 72992
rect 582618 72936 584960 72992
rect 582557 72934 584960 72936
rect 582557 72931 582623 72934
rect 583520 72844 584960 72934
rect 57881 72586 57947 72589
rect 253289 72586 253355 72589
rect 57881 72584 253355 72586
rect 57881 72528 57886 72584
rect 57942 72528 253294 72584
rect 253350 72528 253355 72584
rect 57881 72526 253355 72528
rect 57881 72523 57947 72526
rect 253289 72523 253355 72526
rect 59261 72450 59327 72453
rect 342253 72450 342319 72453
rect 59261 72448 342319 72450
rect 59261 72392 59266 72448
rect 59322 72392 342258 72448
rect 342314 72392 342319 72448
rect 59261 72390 342319 72392
rect 59261 72387 59327 72390
rect 342253 72387 342319 72390
rect -960 71634 480 71724
rect 3509 71634 3575 71637
rect -960 71632 3575 71634
rect -960 71576 3514 71632
rect 3570 71576 3575 71632
rect -960 71574 3575 71576
rect -960 71484 480 71574
rect 3509 71571 3575 71574
rect 55857 71226 55923 71229
rect 248413 71226 248479 71229
rect 55857 71224 248479 71226
rect 55857 71168 55862 71224
rect 55918 71168 248418 71224
rect 248474 71168 248479 71224
rect 55857 71166 248479 71168
rect 55857 71163 55923 71166
rect 248413 71163 248479 71166
rect 53741 71090 53807 71093
rect 262806 71090 262812 71092
rect 53741 71088 262812 71090
rect 53741 71032 53746 71088
rect 53802 71032 262812 71088
rect 53741 71030 262812 71032
rect 53741 71027 53807 71030
rect 262806 71028 262812 71030
rect 262876 71028 262882 71092
rect 130377 69730 130443 69733
rect 168414 69730 168420 69732
rect 130377 69728 168420 69730
rect 130377 69672 130382 69728
rect 130438 69672 168420 69728
rect 130377 69670 168420 69672
rect 130377 69667 130443 69670
rect 168414 69668 168420 69670
rect 168484 69668 168490 69732
rect 177389 69730 177455 69733
rect 242341 69730 242407 69733
rect 177389 69728 242407 69730
rect 177389 69672 177394 69728
rect 177450 69672 242346 69728
rect 242402 69672 242407 69728
rect 177389 69670 242407 69672
rect 177389 69667 177455 69670
rect 242341 69667 242407 69670
rect 60641 69594 60707 69597
rect 252001 69594 252067 69597
rect 60641 69592 252067 69594
rect 60641 69536 60646 69592
rect 60702 69536 252006 69592
rect 252062 69536 252067 69592
rect 60641 69534 252067 69536
rect 60641 69531 60707 69534
rect 252001 69531 252067 69534
rect 64781 68370 64847 68373
rect 257337 68370 257403 68373
rect 64781 68368 257403 68370
rect 64781 68312 64786 68368
rect 64842 68312 257342 68368
rect 257398 68312 257403 68368
rect 64781 68310 257403 68312
rect 64781 68307 64847 68310
rect 257337 68307 257403 68310
rect 67541 68234 67607 68237
rect 276105 68234 276171 68237
rect 67541 68232 276171 68234
rect 67541 68176 67546 68232
rect 67602 68176 276110 68232
rect 276166 68176 276171 68232
rect 67541 68174 276171 68176
rect 67541 68171 67607 68174
rect 276105 68171 276171 68174
rect 276105 67554 276171 67557
rect 277301 67554 277367 67557
rect 362902 67554 362908 67556
rect 276105 67552 362908 67554
rect 276105 67496 276110 67552
rect 276166 67496 277306 67552
rect 277362 67496 362908 67552
rect 276105 67494 362908 67496
rect 276105 67491 276171 67494
rect 277301 67491 277367 67494
rect 362902 67492 362908 67494
rect 362972 67492 362978 67556
rect 75821 67010 75887 67013
rect 239489 67010 239555 67013
rect 75821 67008 239555 67010
rect 75821 66952 75826 67008
rect 75882 66952 239494 67008
rect 239550 66952 239555 67008
rect 75821 66950 239555 66952
rect 75821 66947 75887 66950
rect 239489 66947 239555 66950
rect 61878 66812 61884 66876
rect 61948 66874 61954 66876
rect 307753 66874 307819 66877
rect 61948 66872 307819 66874
rect 61948 66816 307758 66872
rect 307814 66816 307819 66872
rect 61948 66814 307819 66816
rect 61948 66812 61954 66814
rect 307753 66811 307819 66814
rect 78581 65650 78647 65653
rect 267089 65650 267155 65653
rect 78581 65648 267155 65650
rect 78581 65592 78586 65648
rect 78642 65592 267094 65648
rect 267150 65592 267155 65648
rect 78581 65590 267155 65592
rect 78581 65587 78647 65590
rect 267089 65587 267155 65590
rect 48129 65514 48195 65517
rect 258901 65514 258967 65517
rect 48129 65512 258967 65514
rect 48129 65456 48134 65512
rect 48190 65456 258906 65512
rect 258962 65456 258967 65512
rect 48129 65454 258967 65456
rect 48129 65451 48195 65454
rect 258901 65451 258967 65454
rect 58617 64154 58683 64157
rect 222929 64154 222995 64157
rect 58617 64152 222995 64154
rect 58617 64096 58622 64152
rect 58678 64096 222934 64152
rect 222990 64096 222995 64152
rect 58617 64094 222995 64096
rect 58617 64091 58683 64094
rect 222929 64091 222995 64094
rect 89621 62930 89687 62933
rect 243629 62930 243695 62933
rect 89621 62928 243695 62930
rect 89621 62872 89626 62928
rect 89682 62872 243634 62928
rect 243690 62872 243695 62928
rect 89621 62870 243695 62872
rect 89621 62867 89687 62870
rect 243629 62867 243695 62870
rect 70301 62794 70367 62797
rect 260281 62794 260347 62797
rect 70301 62792 260347 62794
rect 70301 62736 70306 62792
rect 70362 62736 260286 62792
rect 260342 62736 260347 62792
rect 70301 62734 260347 62736
rect 70301 62731 70367 62734
rect 260281 62731 260347 62734
rect 79961 61570 80027 61573
rect 249241 61570 249307 61573
rect 79961 61568 249307 61570
rect 79961 61512 79966 61568
rect 80022 61512 249246 61568
rect 249302 61512 249307 61568
rect 79961 61510 249307 61512
rect 79961 61507 80027 61510
rect 249241 61507 249307 61510
rect 15101 61434 15167 61437
rect 242014 61434 242020 61436
rect 15101 61432 242020 61434
rect 15101 61376 15106 61432
rect 15162 61376 242020 61432
rect 15101 61374 242020 61376
rect 15101 61371 15167 61374
rect 242014 61372 242020 61374
rect 242084 61372 242090 61436
rect 45461 59938 45527 59941
rect 236729 59938 236795 59941
rect 45461 59936 236795 59938
rect 45461 59880 45466 59936
rect 45522 59880 236734 59936
rect 236790 59880 236795 59936
rect 45461 59878 236795 59880
rect 45461 59875 45527 59878
rect 236729 59875 236795 59878
rect 582925 59666 582991 59669
rect 583520 59666 584960 59756
rect 582925 59664 584960 59666
rect 582925 59608 582930 59664
rect 582986 59608 584960 59664
rect 582925 59606 584960 59608
rect 582925 59603 582991 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 3325 58578 3391 58581
rect -960 58576 3391 58578
rect -960 58520 3330 58576
rect 3386 58520 3391 58576
rect -960 58518 3391 58520
rect -960 58428 480 58518
rect 3325 58515 3391 58518
rect 38561 58578 38627 58581
rect 235257 58578 235323 58581
rect 38561 58576 235323 58578
rect 38561 58520 38566 58576
rect 38622 58520 235262 58576
rect 235318 58520 235323 58576
rect 38561 58518 235323 58520
rect 38561 58515 38627 58518
rect 235257 58515 235323 58518
rect 35801 57218 35867 57221
rect 229686 57218 229692 57220
rect 35801 57216 229692 57218
rect 35801 57160 35806 57216
rect 35862 57160 229692 57216
rect 35801 57158 229692 57160
rect 35801 57155 35867 57158
rect 229686 57156 229692 57158
rect 229756 57156 229762 57220
rect 31661 55858 31727 55861
rect 257429 55858 257495 55861
rect 31661 55856 257495 55858
rect 31661 55800 31666 55856
rect 31722 55800 257434 55856
rect 257490 55800 257495 55856
rect 31661 55798 257495 55800
rect 31661 55795 31727 55798
rect 257429 55795 257495 55798
rect 23381 54498 23447 54501
rect 232681 54498 232747 54501
rect 23381 54496 232747 54498
rect 23381 54440 23386 54496
rect 23442 54440 232686 54496
rect 232742 54440 232747 54496
rect 23381 54438 232747 54440
rect 23381 54435 23447 54438
rect 232681 54435 232747 54438
rect 111609 53138 111675 53141
rect 266997 53138 267063 53141
rect 111609 53136 267063 53138
rect 111609 53080 111614 53136
rect 111670 53080 267002 53136
rect 267058 53080 267063 53136
rect 111609 53078 267063 53080
rect 111609 53075 111675 53078
rect 266997 53075 267063 53078
rect 22001 51778 22067 51781
rect 269205 51778 269271 51781
rect 22001 51776 269271 51778
rect 22001 51720 22006 51776
rect 22062 51720 269210 51776
rect 269266 51720 269271 51776
rect 22001 51718 269271 51720
rect 22001 51715 22067 51718
rect 269205 51715 269271 51718
rect 44081 50282 44147 50285
rect 250294 50282 250300 50284
rect 44081 50280 250300 50282
rect 44081 50224 44086 50280
rect 44142 50224 250300 50280
rect 44081 50222 250300 50224
rect 44081 50219 44147 50222
rect 250294 50220 250300 50222
rect 250364 50220 250370 50284
rect 39941 48922 40007 48925
rect 261477 48922 261543 48925
rect 39941 48920 261543 48922
rect 39941 48864 39946 48920
rect 40002 48864 261482 48920
rect 261538 48864 261543 48920
rect 39941 48862 261543 48864
rect 39941 48859 40007 48862
rect 261477 48859 261543 48862
rect 582741 46338 582807 46341
rect 583520 46338 584960 46428
rect 582741 46336 584960 46338
rect 582741 46280 582746 46336
rect 582802 46280 584960 46336
rect 582741 46278 584960 46280
rect 582741 46275 582807 46278
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect 3509 45522 3575 45525
rect -960 45520 3575 45522
rect -960 45464 3514 45520
rect 3570 45464 3575 45520
rect -960 45462 3575 45464
rect -960 45372 480 45462
rect 3509 45459 3575 45462
rect 68921 44842 68987 44845
rect 264094 44842 264100 44844
rect 68921 44840 264100 44842
rect 68921 44784 68926 44840
rect 68982 44784 264100 44840
rect 68921 44782 264100 44784
rect 68921 44779 68987 44782
rect 264094 44780 264100 44782
rect 264164 44780 264170 44844
rect 200757 43482 200823 43485
rect 268377 43482 268443 43485
rect 200757 43480 268443 43482
rect 200757 43424 200762 43480
rect 200818 43424 268382 43480
rect 268438 43424 268443 43480
rect 200757 43422 268443 43424
rect 200757 43419 200823 43422
rect 268377 43419 268443 43422
rect 10961 42122 11027 42125
rect 230974 42122 230980 42124
rect 10961 42120 230980 42122
rect 10961 42064 10966 42120
rect 11022 42064 230980 42120
rect 10961 42062 230980 42064
rect 10961 42059 11027 42062
rect 230974 42060 230980 42062
rect 231044 42060 231050 42124
rect 65374 37844 65380 37908
rect 65444 37906 65450 37908
rect 278773 37906 278839 37909
rect 65444 37904 278839 37906
rect 65444 37848 278778 37904
rect 278834 37848 278839 37904
rect 65444 37846 278839 37848
rect 65444 37844 65450 37846
rect 278773 37843 278839 37846
rect 258574 37164 258580 37228
rect 258644 37226 258650 37228
rect 266353 37226 266419 37229
rect 258644 37224 266419 37226
rect 258644 37168 266358 37224
rect 266414 37168 266419 37224
rect 258644 37166 266419 37168
rect 258644 37164 258650 37166
rect 266353 37163 266419 37166
rect 33041 36546 33107 36549
rect 236637 36546 236703 36549
rect 33041 36544 236703 36546
rect 33041 36488 33046 36544
rect 33102 36488 236642 36544
rect 236698 36488 236703 36544
rect 33041 36486 236703 36488
rect 33041 36483 33107 36486
rect 236637 36483 236703 36486
rect 4061 35186 4127 35189
rect 266854 35186 266860 35188
rect 4061 35184 266860 35186
rect 4061 35128 4066 35184
rect 4122 35128 266860 35184
rect 4061 35126 266860 35128
rect 4061 35123 4127 35126
rect 266854 35124 266860 35126
rect 266924 35124 266930 35188
rect 67766 33900 67772 33964
rect 67836 33962 67842 33964
rect 256049 33962 256115 33965
rect 67836 33960 256115 33962
rect 67836 33904 256054 33960
rect 256110 33904 256115 33960
rect 67836 33902 256115 33904
rect 67836 33900 67842 33902
rect 256049 33899 256115 33902
rect 16481 33826 16547 33829
rect 219198 33826 219204 33828
rect 16481 33824 219204 33826
rect 16481 33768 16486 33824
rect 16542 33768 219204 33824
rect 16481 33766 219204 33768
rect 16481 33763 16547 33766
rect 219198 33764 219204 33766
rect 219268 33764 219274 33828
rect 583385 33146 583451 33149
rect 583520 33146 584960 33236
rect 583385 33144 584960 33146
rect 583385 33088 583390 33144
rect 583446 33088 584960 33144
rect 583385 33086 584960 33088
rect 583385 33083 583451 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 2865 32466 2931 32469
rect -960 32464 2931 32466
rect -960 32408 2870 32464
rect 2926 32408 2931 32464
rect -960 32406 2931 32408
rect -960 32316 480 32406
rect 2865 32403 2931 32406
rect 182817 30970 182883 30973
rect 269113 30970 269179 30973
rect 182817 30968 269179 30970
rect 182817 30912 182822 30968
rect 182878 30912 269118 30968
rect 269174 30912 269179 30968
rect 182817 30910 269179 30912
rect 182817 30907 182883 30910
rect 269113 30907 269179 30910
rect 188429 28250 188495 28253
rect 259453 28250 259519 28253
rect 188429 28248 259519 28250
rect 188429 28192 188434 28248
rect 188490 28192 259458 28248
rect 259514 28192 259519 28248
rect 188429 28190 259519 28192
rect 188429 28187 188495 28190
rect 259453 28187 259519 28190
rect 82721 26890 82787 26893
rect 233734 26890 233740 26892
rect 82721 26888 233740 26890
rect 82721 26832 82726 26888
rect 82782 26832 233740 26888
rect 82721 26830 233740 26832
rect 82721 26827 82787 26830
rect 233734 26828 233740 26830
rect 233804 26828 233810 26892
rect 213177 22674 213243 22677
rect 253197 22674 253263 22677
rect 213177 22672 253263 22674
rect 213177 22616 213182 22672
rect 213238 22616 253202 22672
rect 253258 22616 253263 22672
rect 213177 22614 253263 22616
rect 213177 22611 213243 22614
rect 253197 22611 253263 22614
rect 264973 22674 265039 22677
rect 295374 22674 295380 22676
rect 264973 22672 295380 22674
rect 264973 22616 264978 22672
rect 265034 22616 295380 22672
rect 264973 22614 295380 22616
rect 264973 22611 265039 22614
rect 295374 22612 295380 22614
rect 295444 22612 295450 22676
rect 253054 22068 253060 22132
rect 253124 22130 253130 22132
rect 253933 22130 253999 22133
rect 253124 22128 253999 22130
rect 253124 22072 253938 22128
rect 253994 22072 253999 22128
rect 253124 22070 253999 22072
rect 253124 22068 253130 22070
rect 253933 22067 253999 22070
rect 132493 21314 132559 21317
rect 165654 21314 165660 21316
rect 132493 21312 165660 21314
rect 132493 21256 132498 21312
rect 132554 21256 165660 21312
rect 132493 21254 165660 21256
rect 132493 21251 132559 21254
rect 165654 21252 165660 21254
rect 165724 21252 165730 21316
rect 175917 21314 175983 21317
rect 260833 21314 260899 21317
rect 175917 21312 260899 21314
rect 175917 21256 175922 21312
rect 175978 21256 260838 21312
rect 260894 21256 260899 21312
rect 175917 21254 260899 21256
rect 175917 21251 175983 21254
rect 260833 21251 260899 21254
rect 142797 20090 142863 20093
rect 188337 20090 188403 20093
rect 142797 20088 188403 20090
rect 142797 20032 142802 20088
rect 142858 20032 188342 20088
rect 188398 20032 188403 20088
rect 142797 20030 188403 20032
rect 142797 20027 142863 20030
rect 188337 20027 188403 20030
rect 174537 19954 174603 19957
rect 280797 19954 280863 19957
rect 174537 19952 280863 19954
rect 174537 19896 174542 19952
rect 174598 19896 280802 19952
rect 280858 19896 280863 19952
rect 174537 19894 280863 19896
rect 174537 19891 174603 19894
rect 280797 19891 280863 19894
rect 289813 19954 289879 19957
rect 303654 19954 303660 19956
rect 289813 19952 303660 19954
rect 289813 19896 289818 19952
rect 289874 19896 303660 19952
rect 289813 19894 303660 19896
rect 289813 19891 289879 19894
rect 303654 19892 303660 19894
rect 303724 19892 303730 19956
rect 582465 19818 582531 19821
rect 583520 19818 584960 19908
rect 582465 19816 584960 19818
rect 582465 19760 582470 19816
rect 582526 19760 584960 19816
rect 582465 19758 584960 19760
rect 582465 19755 582531 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 3417 19410 3483 19413
rect -960 19408 3483 19410
rect -960 19352 3422 19408
rect 3478 19352 3483 19408
rect -960 19350 3483 19352
rect -960 19260 480 19350
rect 3417 19347 3483 19350
rect 173750 18532 173756 18596
rect 173820 18594 173826 18596
rect 338757 18594 338823 18597
rect 173820 18592 338823 18594
rect 173820 18536 338762 18592
rect 338818 18536 338823 18592
rect 173820 18534 338823 18536
rect 173820 18532 173826 18534
rect 338757 18531 338823 18534
rect 189942 17308 189948 17372
rect 190012 17370 190018 17372
rect 263593 17370 263659 17373
rect 190012 17368 263659 17370
rect 190012 17312 263598 17368
rect 263654 17312 263659 17368
rect 190012 17310 263659 17312
rect 190012 17308 190018 17310
rect 263593 17307 263659 17310
rect 3969 17234 4035 17237
rect 223614 17234 223620 17236
rect 3969 17232 223620 17234
rect 3969 17176 3974 17232
rect 4030 17176 223620 17232
rect 3969 17174 223620 17176
rect 3969 17171 4035 17174
rect 223614 17172 223620 17174
rect 223684 17172 223690 17236
rect 186957 14514 187023 14517
rect 302877 14514 302943 14517
rect 186957 14512 302943 14514
rect 186957 14456 186962 14512
rect 187018 14456 302882 14512
rect 302938 14456 302943 14512
rect 186957 14454 302943 14456
rect 186957 14451 187023 14454
rect 302877 14451 302943 14454
rect 185342 12956 185348 13020
rect 185412 13018 185418 13020
rect 268285 13018 268351 13021
rect 185412 13016 268351 13018
rect 185412 12960 268290 13016
rect 268346 12960 268351 13016
rect 185412 12958 268351 12960
rect 185412 12956 185418 12958
rect 268285 12955 268351 12958
rect 112437 11658 112503 11661
rect 136449 11658 136515 11661
rect 112437 11656 136515 11658
rect 112437 11600 112442 11656
rect 112498 11600 136454 11656
rect 136510 11600 136515 11656
rect 112437 11598 136515 11600
rect 112437 11595 112503 11598
rect 136449 11595 136515 11598
rect 195329 11658 195395 11661
rect 270769 11658 270835 11661
rect 195329 11656 270835 11658
rect 195329 11600 195334 11656
rect 195390 11600 270774 11656
rect 270830 11600 270835 11656
rect 195329 11598 270835 11600
rect 195329 11595 195395 11598
rect 270769 11595 270835 11598
rect 268469 10298 268535 10301
rect 363086 10298 363092 10300
rect 268469 10296 363092 10298
rect 268469 10240 268474 10296
rect 268530 10240 363092 10296
rect 268469 10238 363092 10240
rect 268469 10235 268535 10238
rect 363086 10236 363092 10238
rect 363156 10236 363162 10300
rect 180558 9012 180564 9076
rect 180628 9074 180634 9076
rect 242893 9074 242959 9077
rect 180628 9072 242959 9074
rect 180628 9016 242898 9072
rect 242954 9016 242959 9072
rect 180628 9014 242959 9016
rect 180628 9012 180634 9014
rect 242893 9011 242959 9014
rect 565 8938 631 8941
rect 227662 8938 227668 8940
rect 565 8936 227668 8938
rect 565 8880 570 8936
rect 626 8880 227668 8936
rect 565 8878 227668 8880
rect 565 8875 631 8878
rect 227662 8876 227668 8878
rect 227732 8876 227738 8940
rect 170438 7516 170444 7580
rect 170508 7578 170514 7580
rect 244089 7578 244155 7581
rect 170508 7576 244155 7578
rect 170508 7520 244094 7576
rect 244150 7520 244155 7576
rect 170508 7518 244155 7520
rect 170508 7516 170514 7518
rect 244089 7515 244155 7518
rect 13 6898 79 6901
rect 326337 6898 326403 6901
rect 326797 6898 326863 6901
rect 385033 6898 385099 6901
rect 13 6896 122 6898
rect 13 6840 18 6896
rect 74 6840 122 6896
rect 13 6835 122 6840
rect 326337 6896 385099 6898
rect 326337 6840 326342 6896
rect 326398 6840 326802 6896
rect 326858 6840 385038 6896
rect 385094 6840 385099 6896
rect 326337 6838 385099 6840
rect 326337 6835 326403 6838
rect 326797 6835 326863 6838
rect 385033 6835 385099 6838
rect 62 6626 122 6835
rect 580165 6626 580231 6629
rect 583520 6626 584960 6716
rect 62 6580 674 6626
rect -960 6566 674 6580
rect -960 6490 480 6566
rect 614 6490 674 6566
rect 580165 6624 584960 6626
rect 580165 6568 580170 6624
rect 580226 6568 584960 6624
rect 580165 6566 584960 6568
rect 580165 6563 580231 6566
rect -960 6430 674 6490
rect 583520 6476 584960 6566
rect -960 6340 480 6430
rect 239305 5674 239371 5677
rect 244917 5674 244983 5677
rect 239305 5672 244983 5674
rect 239305 5616 239310 5672
rect 239366 5616 244922 5672
rect 244978 5616 244983 5672
rect 239305 5614 244983 5616
rect 239305 5611 239371 5614
rect 244917 5611 244983 5614
rect 191097 4858 191163 4861
rect 281901 4858 281967 4861
rect 191097 4856 281967 4858
rect 191097 4800 191102 4856
rect 191158 4800 281906 4856
rect 281962 4800 281967 4856
rect 191097 4798 281967 4800
rect 191097 4795 191163 4798
rect 281901 4795 281967 4798
rect 298461 4858 298527 4861
rect 356094 4858 356100 4860
rect 298461 4856 356100 4858
rect 298461 4800 298466 4856
rect 298522 4800 356100 4856
rect 298461 4798 356100 4800
rect 298461 4795 298527 4798
rect 356094 4796 356100 4798
rect 356164 4796 356170 4860
rect 197997 4042 198063 4045
rect 267733 4042 267799 4045
rect 268469 4042 268535 4045
rect 197997 4040 268535 4042
rect 197997 3984 198002 4040
rect 198058 3984 267738 4040
rect 267794 3984 268474 4040
rect 268530 3984 268535 4040
rect 197997 3982 268535 3984
rect 197997 3979 198063 3982
rect 267733 3979 267799 3982
rect 268469 3979 268535 3982
rect 342989 4042 343055 4045
rect 346945 4042 347011 4045
rect 342989 4040 347011 4042
rect 342989 3984 342994 4040
rect 343050 3984 346950 4040
rect 347006 3984 347011 4040
rect 342989 3982 347011 3984
rect 342989 3979 343055 3982
rect 346945 3979 347011 3982
rect 125869 3498 125935 3501
rect 196617 3498 196683 3501
rect 125869 3496 196683 3498
rect 125869 3440 125874 3496
rect 125930 3440 196622 3496
rect 196678 3440 196683 3496
rect 125869 3438 196683 3440
rect 125869 3435 125935 3438
rect 196617 3435 196683 3438
rect 246246 3436 246252 3500
rect 246316 3498 246322 3500
rect 247585 3498 247651 3501
rect 246316 3496 247651 3498
rect 246316 3440 247590 3496
rect 247646 3440 247651 3496
rect 246316 3438 247651 3440
rect 246316 3436 246322 3438
rect 247585 3435 247651 3438
rect 251766 3436 251772 3500
rect 251836 3498 251842 3500
rect 253473 3498 253539 3501
rect 251836 3496 253539 3498
rect 251836 3440 253478 3496
rect 253534 3440 253539 3496
rect 251836 3438 253539 3440
rect 251836 3436 251842 3438
rect 253473 3435 253539 3438
rect 277117 3498 277183 3501
rect 285622 3498 285628 3500
rect 277117 3496 285628 3498
rect 277117 3440 277122 3496
rect 277178 3440 285628 3496
rect 277117 3438 285628 3440
rect 277117 3435 277183 3438
rect 285622 3436 285628 3438
rect 285692 3436 285698 3500
rect 287646 3436 287652 3500
rect 287716 3498 287722 3500
rect 287789 3498 287855 3501
rect 287716 3496 287855 3498
rect 287716 3440 287794 3496
rect 287850 3440 287855 3496
rect 287716 3438 287855 3440
rect 287716 3436 287722 3438
rect 287789 3435 287855 3438
rect 291142 3436 291148 3500
rect 291212 3498 291218 3500
rect 291377 3498 291443 3501
rect 291212 3496 291443 3498
rect 291212 3440 291382 3496
rect 291438 3440 291443 3496
rect 291212 3438 291443 3440
rect 291212 3436 291218 3438
rect 291377 3435 291443 3438
rect 293166 3436 293172 3500
rect 293236 3498 293242 3500
rect 293677 3498 293743 3501
rect 293236 3496 293743 3498
rect 293236 3440 293682 3496
rect 293738 3440 293743 3496
rect 293236 3438 293743 3440
rect 293236 3436 293242 3438
rect 293677 3435 293743 3438
rect 299606 3436 299612 3500
rect 299676 3498 299682 3500
rect 300761 3498 300827 3501
rect 299676 3496 300827 3498
rect 299676 3440 300766 3496
rect 300822 3440 300827 3496
rect 299676 3438 300827 3440
rect 299676 3436 299682 3438
rect 300761 3435 300827 3438
rect 7649 3362 7715 3365
rect 177389 3362 177455 3365
rect 7649 3360 177455 3362
rect 7649 3304 7654 3360
rect 7710 3304 177394 3360
rect 177450 3304 177455 3360
rect 7649 3302 177455 3304
rect 7649 3299 7715 3302
rect 177389 3299 177455 3302
rect 241278 3300 241284 3364
rect 241348 3362 241354 3364
rect 252369 3362 252435 3365
rect 241348 3360 252435 3362
rect 241348 3304 252374 3360
rect 252430 3304 252435 3360
rect 241348 3302 252435 3304
rect 241348 3300 241354 3302
rect 252369 3299 252435 3302
rect 277301 3362 277367 3365
rect 284293 3362 284359 3365
rect 277301 3360 284359 3362
rect 277301 3304 277306 3360
rect 277362 3304 284298 3360
rect 284354 3304 284359 3360
rect 277301 3302 284359 3304
rect 277301 3299 277367 3302
rect 284293 3299 284359 3302
rect 285397 3362 285463 3365
rect 298134 3362 298140 3364
rect 285397 3360 298140 3362
rect 285397 3304 285402 3360
rect 285458 3304 298140 3360
rect 285397 3302 298140 3304
rect 285397 3299 285463 3302
rect 298134 3300 298140 3302
rect 298204 3300 298210 3364
rect 302734 3300 302740 3364
rect 302804 3362 302810 3364
rect 317321 3362 317387 3365
rect 302804 3360 317387 3362
rect 302804 3304 317326 3360
rect 317382 3304 317387 3360
rect 302804 3302 317387 3304
rect 302804 3300 302810 3302
rect 317321 3299 317387 3302
rect 330385 3362 330451 3365
rect 353293 3362 353359 3365
rect 330385 3360 353359 3362
rect 330385 3304 330390 3360
rect 330446 3304 353298 3360
rect 353354 3304 353359 3360
rect 330385 3302 353359 3304
rect 330385 3299 330451 3302
rect 353293 3299 353359 3302
rect 140037 2682 140103 2685
rect 142797 2682 142863 2685
rect 140037 2680 142863 2682
rect 140037 2624 140042 2680
rect 140098 2624 142802 2680
rect 142858 2624 142863 2680
rect 140037 2622 142863 2624
rect 140037 2619 140103 2622
rect 142797 2619 142863 2622
<< via3 >>
rect 69612 702476 69676 702540
rect 88012 590684 88076 590748
rect 93900 588644 93964 588708
rect 88196 588508 88260 588572
rect 88196 585652 88260 585716
rect 88196 582796 88260 582860
rect 69428 582252 69492 582316
rect 91508 578036 91572 578100
rect 124260 577492 124324 577556
rect 121684 572732 121748 572796
rect 67404 556820 67468 556884
rect 170260 552060 170324 552124
rect 66668 551380 66732 551444
rect 173020 550700 173084 550764
rect 197860 546620 197924 546684
rect 199516 546484 199580 546548
rect 67772 545940 67836 546004
rect 200620 545260 200684 545324
rect 67772 545124 67836 545188
rect 353340 545124 353404 545188
rect 161980 543900 162044 543964
rect 69428 542268 69492 542332
rect 188844 541180 188908 541244
rect 160692 539820 160756 539884
rect 362908 539684 362972 539748
rect 352052 538188 352116 538252
rect 67404 537372 67468 537436
rect 357572 537100 357636 537164
rect 68140 535468 68204 535532
rect 69612 535528 69676 535532
rect 69612 535472 69626 535528
rect 69626 535472 69676 535528
rect 69612 535468 69676 535472
rect 67772 535332 67836 535396
rect 191604 535332 191668 535396
rect 106412 534652 106476 534716
rect 183324 534108 183388 534172
rect 200068 533428 200132 533492
rect 179276 530572 179340 530636
rect 197860 526356 197924 526420
rect 66484 523772 66548 523836
rect 66668 523636 66732 523700
rect 195100 514932 195164 514996
rect 198596 512484 198660 512548
rect 356284 507044 356348 507108
rect 155724 504324 155788 504388
rect 184796 502420 184860 502484
rect 177804 496844 177868 496908
rect 198780 485556 198844 485620
rect 360148 480388 360212 480452
rect 122604 479436 122668 479500
rect 115980 473996 116044 474060
rect 104940 470596 105004 470660
rect 118188 469780 118252 469844
rect 70164 467876 70228 467940
rect 113220 467740 113284 467804
rect 107700 467060 107764 467124
rect 102180 464340 102244 464404
rect 71820 462844 71884 462908
rect 92980 462844 93044 462908
rect 89668 460124 89732 460188
rect 111748 460124 111812 460188
rect 94084 459580 94148 459644
rect 118740 458764 118804 458828
rect 358860 458356 358924 458420
rect 96660 457404 96724 457468
rect 108988 457404 109052 457468
rect 172468 456860 172532 456924
rect 90220 456180 90284 456244
rect 100708 456044 100772 456108
rect 98132 454684 98196 454748
rect 122972 453188 123036 453252
rect 91508 450468 91572 450532
rect 120028 450468 120092 450532
rect 172100 449924 172164 449988
rect 91508 447204 91572 447268
rect 115796 447204 115860 447268
rect 70164 447128 70228 447132
rect 70164 447072 70214 447128
rect 70214 447072 70228 447128
rect 70164 447068 70228 447072
rect 72372 446388 72436 446452
rect 68324 445844 68388 445908
rect 71820 445904 71884 445908
rect 71820 445848 71834 445904
rect 71834 445848 71884 445904
rect 71820 445844 71884 445848
rect 72740 445844 72804 445908
rect 93900 445708 93964 445772
rect 96292 445708 96356 445772
rect 100524 445708 100588 445772
rect 114324 445768 114388 445772
rect 114324 445712 114374 445768
rect 114374 445712 114388 445768
rect 114324 445708 114388 445712
rect 118004 445708 118068 445772
rect 108804 444620 108868 444684
rect 111564 444620 111628 444684
rect 124260 443804 124324 443868
rect 154068 442172 154132 442236
rect 197124 438908 197188 438972
rect 160876 436052 160940 436116
rect 122972 435372 123036 435436
rect 186820 430612 186884 430676
rect 120028 425988 120092 426052
rect 197860 421636 197924 421700
rect 121500 420820 121564 420884
rect 66668 419596 66732 419660
rect 121500 419596 121564 419660
rect 69244 407764 69308 407828
rect 165660 407764 165724 407828
rect 69244 407084 69308 407148
rect 192708 404500 192772 404564
rect 122604 403684 122668 403748
rect 356468 394436 356532 394500
rect 198596 393348 198660 393412
rect 72372 391852 72436 391916
rect 73108 391852 73172 391916
rect 92980 391096 93044 391100
rect 92980 391040 92994 391096
rect 92994 391040 93044 391096
rect 92980 391036 93044 391040
rect 121500 390628 121564 390692
rect 69612 390356 69676 390420
rect 89668 390356 89732 390420
rect 94084 390356 94148 390420
rect 96660 390356 96724 390420
rect 98132 390356 98196 390420
rect 102180 390416 102244 390420
rect 102180 390360 102194 390416
rect 102194 390360 102244 390416
rect 102180 390356 102244 390360
rect 104940 390416 105004 390420
rect 104940 390360 104990 390416
rect 104990 390360 105004 390416
rect 104940 390356 105004 390360
rect 106412 390356 106476 390420
rect 107700 390356 107764 390420
rect 108988 390356 109052 390420
rect 115980 390416 116044 390420
rect 115980 390360 115994 390416
rect 115994 390360 116044 390416
rect 115980 390356 116044 390360
rect 118188 390356 118252 390420
rect 118740 390416 118804 390420
rect 118740 390360 118790 390416
rect 118790 390360 118804 390416
rect 118740 390356 118804 390360
rect 100708 390280 100772 390284
rect 100708 390224 100758 390280
rect 100758 390224 100772 390280
rect 100708 390220 100772 390224
rect 70900 389268 70964 389332
rect 169708 389268 169772 389332
rect 356100 389268 356164 389332
rect 68140 388996 68204 389060
rect 73108 389056 73172 389060
rect 73108 389000 73122 389056
rect 73122 389000 73172 389056
rect 73108 388996 73172 389000
rect 90220 388996 90284 389060
rect 91508 388860 91572 388924
rect 111748 388996 111812 389060
rect 113220 389056 113284 389060
rect 113220 389000 113234 389056
rect 113234 389000 113284 389056
rect 113220 388996 113284 389000
rect 356100 386548 356164 386612
rect 195836 384780 195900 384844
rect 363092 384644 363156 384708
rect 356284 383964 356348 384028
rect 356284 383692 356348 383756
rect 356100 381516 356164 381580
rect 356468 381516 356532 381580
rect 200068 381108 200132 381172
rect 111564 380972 111628 381036
rect 115796 379204 115860 379268
rect 111748 378660 111812 378724
rect 114324 378116 114388 378180
rect 196572 378116 196636 378180
rect 357572 377980 357636 378044
rect 198780 377572 198844 377636
rect 67772 377436 67836 377500
rect 68324 377300 68388 377364
rect 195836 376484 195900 376548
rect 354812 376348 354876 376412
rect 353340 375940 353404 376004
rect 241652 375260 241716 375324
rect 288388 375260 288452 375324
rect 354444 375260 354508 375324
rect 244780 374580 244844 374644
rect 303660 374036 303724 374100
rect 96292 373356 96356 373420
rect 356100 371316 356164 371380
rect 69796 370500 69860 370564
rect 100524 369956 100588 370020
rect 195284 368596 195348 368660
rect 69612 368460 69676 368524
rect 224908 367780 224972 367844
rect 157932 367644 157996 367708
rect 285628 365740 285692 365804
rect 64644 364652 64708 364716
rect 196572 362340 196636 362404
rect 357572 362204 357636 362268
rect 71084 361796 71148 361860
rect 157748 360028 157812 360092
rect 356284 359348 356348 359412
rect 159956 356628 160020 356692
rect 358860 356628 358924 356692
rect 352052 355404 352116 355468
rect 180564 354044 180628 354108
rect 180564 353500 180628 353564
rect 199516 353500 199580 353564
rect 234476 352548 234540 352612
rect 211660 351324 211724 351388
rect 240732 351188 240796 351252
rect 108804 349148 108868 349212
rect 72740 349012 72804 349076
rect 68876 348468 68940 348532
rect 187004 347712 187068 347716
rect 187004 347656 187018 347712
rect 187018 347656 187068 347712
rect 187004 347652 187068 347656
rect 248460 347108 248524 347172
rect 66668 346972 66732 347036
rect 187004 346428 187068 346492
rect 245700 345748 245764 345812
rect 155724 345068 155788 345132
rect 295380 343708 295444 343772
rect 360148 344252 360212 344316
rect 168972 342892 169036 342956
rect 159404 341532 159468 341596
rect 78444 341396 78508 341460
rect 251772 341396 251836 341460
rect 73476 340036 73540 340100
rect 212580 339628 212644 339692
rect 230428 339492 230492 339556
rect 67956 339356 68020 339420
rect 68876 339356 68940 339420
rect 118004 339356 118068 339420
rect 156644 339356 156708 339420
rect 210740 338676 210804 338740
rect 67956 338268 68020 338332
rect 202644 337588 202708 337652
rect 83964 337452 84028 337516
rect 81020 335956 81084 336020
rect 69796 335412 69860 335476
rect 154620 334596 154684 334660
rect 214420 334596 214484 334660
rect 222332 334188 222396 334252
rect 155724 331876 155788 331940
rect 189948 331876 190012 331940
rect 232084 331740 232148 331804
rect 156828 331332 156892 331396
rect 158484 331332 158548 331396
rect 75684 331196 75748 331260
rect 93900 330108 93964 330172
rect 168236 329700 168300 329764
rect 69428 329156 69492 329220
rect 71084 329156 71148 329220
rect 77156 329156 77220 329220
rect 82676 329156 82740 329220
rect 255268 328476 255332 328540
rect 69428 328340 69492 328404
rect 169524 327116 169588 327180
rect 156828 326300 156892 326364
rect 61884 325756 61948 325820
rect 69428 325484 69492 325548
rect 69428 323988 69492 324052
rect 291148 323580 291212 323644
rect 195100 322220 195164 322284
rect 253060 322084 253124 322148
rect 176516 318004 176580 318068
rect 185348 315284 185412 315348
rect 249748 315284 249812 315348
rect 198596 314740 198660 314804
rect 277900 314740 277964 314804
rect 174676 314196 174740 314260
rect 215340 314060 215404 314124
rect 200620 312428 200684 312492
rect 213868 312428 213932 312492
rect 160692 311884 160756 311948
rect 159220 309708 159284 309772
rect 159956 309028 160020 309092
rect 159956 308348 160020 308412
rect 281580 307668 281644 307732
rect 263548 306444 263612 306508
rect 207980 305764 208044 305828
rect 159404 303724 159468 303788
rect 168972 303724 169036 303788
rect 247724 303588 247788 303652
rect 227668 302772 227732 302836
rect 195836 300928 195900 300932
rect 195836 300872 195850 300928
rect 195850 300872 195900 300928
rect 195836 300868 195900 300872
rect 157932 300052 157996 300116
rect 158484 300052 158548 300116
rect 66668 298752 66732 298756
rect 66668 298696 66682 298752
rect 66682 298696 66732 298752
rect 66668 298692 66732 298696
rect 242940 298692 243004 298756
rect 240364 298420 240428 298484
rect 244412 298148 244476 298212
rect 184060 297468 184124 297532
rect 172468 296652 172532 296716
rect 357572 296652 357636 296716
rect 157012 296244 157076 296308
rect 172468 296244 172532 296308
rect 206876 296244 206940 296308
rect 219204 296108 219268 296172
rect 357572 295972 357636 296036
rect 173756 295292 173820 295356
rect 203196 295292 203260 295356
rect 200620 294476 200684 294540
rect 163452 293116 163516 293180
rect 249932 292708 249996 292772
rect 217548 291756 217612 291820
rect 196940 290396 197004 290460
rect 156828 289172 156892 289236
rect 160876 288628 160940 288692
rect 240732 288356 240796 288420
rect 199332 287404 199396 287468
rect 221044 287268 221108 287332
rect 231900 287268 231964 287332
rect 228220 287132 228284 287196
rect 238708 287132 238772 287196
rect 53604 285696 53668 285700
rect 234660 285908 234724 285972
rect 244044 285908 244108 285972
rect 226932 285772 226996 285836
rect 53604 285640 53618 285696
rect 53618 285640 53668 285696
rect 53604 285636 53668 285640
rect 200620 285636 200684 285700
rect 209636 285636 209700 285700
rect 215340 285636 215404 285700
rect 226196 285636 226260 285700
rect 249012 285772 249076 285836
rect 198780 284412 198844 284476
rect 208164 284140 208228 284204
rect 216444 284004 216508 284068
rect 201356 283868 201420 283932
rect 215524 283868 215588 283932
rect 220860 283868 220924 283932
rect 224724 283928 224788 283932
rect 224724 283872 224738 283928
rect 224738 283872 224788 283928
rect 224724 283868 224788 283872
rect 227668 283868 227732 283932
rect 228772 283868 228836 283932
rect 229692 283868 229756 283932
rect 230980 283928 231044 283932
rect 230980 283872 231030 283928
rect 231030 283872 231044 283928
rect 230980 283868 231044 283872
rect 236500 283868 236564 283932
rect 237972 283868 238036 283932
rect 67772 280196 67836 280260
rect 244780 280060 244844 280124
rect 255268 280060 255332 280124
rect 198780 279380 198844 279444
rect 198780 279244 198844 279308
rect 249932 278760 249996 278764
rect 249932 278704 249982 278760
rect 249982 278704 249996 278760
rect 249932 278700 249996 278704
rect 198596 278020 198660 278084
rect 157748 277748 157812 277812
rect 160692 276660 160756 276724
rect 66852 276116 66916 276180
rect 245700 275300 245764 275364
rect 178540 272444 178604 272508
rect 199332 271084 199396 271148
rect 67956 269588 68020 269652
rect 244228 269860 244292 269924
rect 160140 269316 160204 269380
rect 169524 269180 169588 269244
rect 243492 269044 243556 269108
rect 66852 268364 66916 268428
rect 281764 268364 281828 268428
rect 170444 267608 170508 267612
rect 170444 267552 170494 267608
rect 170494 267552 170508 267608
rect 170444 267548 170508 267552
rect 67404 267412 67468 267476
rect 195836 267276 195900 267340
rect 170444 266460 170508 266524
rect 169708 266324 169772 266388
rect 168972 265508 169036 265572
rect 198780 265508 198844 265572
rect 199332 263060 199396 263124
rect 249012 261428 249076 261492
rect 162164 260068 162228 260132
rect 161980 259524 162044 259588
rect 244412 259524 244476 259588
rect 195284 259388 195348 259452
rect 65380 257892 65444 257956
rect 69428 257076 69492 257140
rect 247724 255988 247788 256052
rect 67956 254356 68020 254420
rect 195100 254356 195164 254420
rect 197860 252588 197924 252652
rect 66668 252180 66732 252244
rect 248460 252180 248524 252244
rect 168420 251228 168484 251292
rect 160140 251092 160204 251156
rect 248460 249868 248524 249932
rect 67772 248916 67836 248980
rect 159404 247556 159468 247620
rect 160876 247556 160940 247620
rect 158116 245788 158180 245852
rect 186820 245788 186884 245852
rect 156828 244972 156892 245036
rect 168972 244972 169036 245036
rect 64644 242932 64708 242996
rect 245700 242932 245764 242996
rect 67404 242796 67468 242860
rect 195284 242856 195348 242860
rect 195284 242800 195334 242856
rect 195334 242800 195348 242856
rect 195284 242796 195348 242800
rect 157932 242116 157996 242180
rect 81020 242040 81084 242044
rect 81020 241984 81034 242040
rect 81034 241984 81084 242040
rect 81020 241980 81084 241984
rect 154620 242040 154684 242044
rect 154620 241984 154670 242040
rect 154670 241984 154684 242040
rect 154620 241980 154684 241984
rect 195284 241844 195348 241908
rect 170260 241572 170324 241636
rect 156460 241436 156524 241500
rect 243492 241300 243556 241364
rect 168236 240076 168300 240140
rect 202644 240136 202708 240140
rect 202644 240080 202658 240136
rect 202658 240080 202708 240136
rect 202644 240076 202708 240080
rect 203196 240076 203260 240140
rect 208164 240136 208228 240140
rect 208164 240080 208214 240136
rect 208214 240080 208228 240136
rect 208164 240076 208228 240080
rect 210740 240136 210804 240140
rect 210740 240080 210754 240136
rect 210754 240080 210804 240136
rect 210740 240076 210804 240080
rect 213868 240136 213932 240140
rect 213868 240080 213918 240136
rect 213918 240080 213932 240136
rect 213868 240076 213932 240080
rect 214420 240076 214484 240140
rect 217548 240136 217612 240140
rect 217548 240080 217562 240136
rect 217562 240080 217612 240136
rect 217548 240076 217612 240080
rect 219204 240076 219268 240140
rect 221044 240076 221108 240140
rect 230428 240076 230492 240140
rect 230980 240076 231044 240140
rect 232084 240076 232148 240140
rect 234476 240076 234540 240140
rect 238708 240076 238772 240140
rect 207980 239940 208044 240004
rect 248460 239532 248524 239596
rect 206876 238580 206940 238644
rect 212580 238580 212644 238644
rect 222332 238580 222396 238644
rect 243860 238580 243924 238644
rect 196940 238444 197004 238508
rect 224908 238444 224972 238508
rect 226196 238444 226260 238508
rect 78444 237280 78508 237284
rect 78444 237224 78494 237280
rect 78494 237224 78508 237280
rect 78444 237220 78508 237224
rect 83964 237220 84028 237284
rect 73476 236676 73540 236740
rect 154068 235860 154132 235924
rect 184060 235588 184124 235652
rect 239260 235648 239324 235652
rect 239260 235592 239274 235648
rect 239274 235592 239324 235648
rect 239260 235588 239324 235592
rect 158116 235180 158180 235244
rect 159220 233820 159284 233884
rect 156644 231780 156708 231844
rect 245700 231372 245764 231436
rect 195284 229740 195348 229804
rect 70900 228788 70964 228852
rect 173020 228652 173084 228716
rect 82676 227564 82740 227628
rect 184796 226264 184860 226268
rect 184796 226208 184810 226264
rect 184810 226208 184860 226264
rect 184796 226204 184860 226208
rect 242940 226068 243004 226132
rect 69612 225660 69676 225724
rect 160876 224572 160940 224636
rect 233188 223544 233252 223548
rect 233188 223488 233238 223544
rect 233238 223488 233252 223544
rect 233188 223484 233252 223488
rect 215156 222320 215220 222324
rect 215156 222264 215170 222320
rect 215170 222264 215220 222320
rect 215156 222260 215220 222264
rect 195100 220764 195164 220828
rect 75684 220084 75748 220148
rect 228220 219540 228284 219604
rect 172100 218996 172164 219060
rect 177988 217636 178052 217700
rect 177988 217228 178052 217292
rect 298140 217228 298204 217292
rect 176516 216004 176580 216068
rect 241652 215868 241716 215932
rect 188844 215188 188908 215252
rect 249932 215112 249996 215116
rect 249932 215056 249946 215112
rect 249946 215056 249996 215112
rect 249932 215052 249996 215056
rect 302740 214644 302804 214708
rect 215524 214508 215588 214572
rect 183324 213888 183388 213892
rect 183324 213832 183338 213888
rect 183338 213832 183388 213888
rect 183324 213828 183388 213832
rect 66668 213148 66732 213212
rect 237972 212468 238036 212532
rect 174676 211788 174740 211852
rect 209636 211304 209700 211308
rect 209636 211248 209686 211304
rect 209686 211248 209700 211304
rect 209636 211244 209700 211248
rect 162164 210836 162228 210900
rect 163452 210700 163516 210764
rect 179276 209476 179340 209540
rect 179276 208932 179340 208996
rect 192708 208252 192772 208316
rect 293172 207572 293236 207636
rect 192708 207164 192772 207228
rect 191604 206348 191668 206412
rect 197124 205532 197188 205596
rect 199332 202268 199396 202332
rect 67956 201316 68020 201380
rect 224908 199548 224972 199612
rect 246252 199276 246316 199340
rect 248460 197916 248524 197980
rect 211660 197236 211724 197300
rect 212396 197236 212460 197300
rect 173020 196692 173084 196756
rect 212396 196556 212460 196620
rect 258580 196556 258644 196620
rect 220860 192476 220924 192540
rect 287652 189620 287716 189684
rect 288388 189620 288452 189684
rect 242940 189076 243004 189140
rect 237420 188532 237484 188596
rect 216444 188396 216508 188460
rect 284524 188396 284588 188460
rect 77156 188260 77220 188324
rect 233372 185812 233436 185876
rect 232084 185676 232148 185740
rect 299612 184996 299676 185060
rect 280476 183092 280540 183156
rect 187004 182956 187068 183020
rect 288572 182956 288636 183020
rect 280292 181460 280356 181524
rect 224908 181188 224972 181252
rect 226932 180236 226996 180300
rect 287100 180236 287164 180300
rect 224724 180100 224788 180164
rect 237972 180100 238036 180164
rect 290596 180100 290660 180164
rect 241652 178740 241716 178804
rect 284340 178740 284404 178804
rect 228772 178604 228836 178668
rect 279004 178604 279068 178668
rect 116900 178196 116964 178260
rect 110644 177924 110708 177988
rect 109540 177788 109604 177852
rect 98316 177516 98380 177580
rect 100708 177576 100772 177580
rect 100708 177520 100758 177576
rect 100758 177520 100772 177576
rect 100708 177516 100772 177520
rect 105676 177516 105740 177580
rect 106964 177516 107028 177580
rect 113220 177516 113284 177580
rect 115796 177576 115860 177580
rect 115796 177520 115846 177576
rect 115846 177520 115860 177576
rect 115796 177516 115860 177520
rect 118372 177516 118436 177580
rect 121868 177576 121932 177580
rect 121868 177520 121918 177576
rect 121918 177520 121932 177576
rect 121868 177516 121932 177520
rect 124444 177516 124508 177580
rect 127020 177516 127084 177580
rect 132356 177576 132420 177580
rect 132356 177520 132406 177576
rect 132406 177520 132420 177576
rect 132356 177516 132420 177520
rect 133092 177516 133156 177580
rect 283788 177380 283852 177444
rect 240548 177244 240612 177308
rect 255820 177244 255884 177308
rect 279372 177244 279436 177308
rect 112116 177108 112180 177172
rect 114324 177168 114388 177172
rect 114324 177112 114374 177168
rect 114374 177112 114388 177168
rect 114324 177108 114388 177112
rect 119476 177108 119540 177172
rect 134380 177108 134444 177172
rect 104572 176972 104636 177036
rect 229140 176972 229204 177036
rect 97028 176836 97092 176900
rect 101996 176836 102060 176900
rect 230612 176836 230676 176900
rect 285812 176836 285876 176900
rect 123156 176700 123220 176764
rect 125732 176700 125796 176764
rect 129412 176760 129476 176764
rect 129412 176704 129462 176760
rect 129462 176704 129476 176760
rect 129412 176700 129476 176704
rect 148180 176760 148244 176764
rect 148180 176704 148230 176760
rect 148230 176704 148244 176760
rect 148180 176700 148244 176704
rect 158852 176700 158916 176764
rect 99420 176428 99484 176492
rect 103284 176428 103348 176492
rect 128124 176488 128188 176492
rect 128124 176432 128174 176488
rect 128174 176432 128188 176488
rect 128124 176428 128188 176432
rect 244412 175884 244476 175948
rect 130700 175672 130764 175676
rect 130700 175616 130750 175672
rect 130750 175616 130764 175672
rect 130700 175612 130764 175616
rect 135668 175672 135732 175676
rect 135668 175616 135718 175672
rect 135718 175616 135732 175672
rect 135668 175612 135732 175616
rect 120764 175476 120828 175540
rect 108068 175340 108132 175404
rect 236684 175204 236748 175268
rect 241284 175204 241348 175268
rect 279372 175204 279436 175268
rect 236500 175068 236564 175132
rect 240364 174252 240428 174316
rect 247724 173844 247788 173908
rect 279372 173708 279436 173772
rect 244228 172756 244292 172820
rect 280108 172348 280172 172412
rect 280476 172348 280540 172412
rect 233372 171124 233436 171188
rect 279556 170580 279620 170644
rect 230612 169492 230676 169556
rect 231900 167588 231964 167652
rect 230980 167180 231044 167244
rect 287100 167044 287164 167108
rect 237420 161468 237484 161532
rect 230980 159564 231044 159628
rect 281764 157252 281828 157316
rect 239260 156572 239324 156636
rect 281580 156436 281644 156500
rect 234660 154804 234724 154868
rect 233188 153036 233252 153100
rect 240548 152492 240612 152556
rect 172100 152356 172164 152420
rect 244412 150996 244476 151060
rect 249748 150452 249812 150516
rect 247724 150044 247788 150108
rect 229140 149636 229204 149700
rect 242940 149092 243004 149156
rect 229140 148004 229204 148068
rect 230428 147868 230492 147932
rect 232084 147188 232148 147252
rect 249932 147052 249996 147116
rect 231716 146916 231780 146980
rect 283788 146508 283852 146572
rect 231716 145828 231780 145892
rect 236684 145284 236748 145348
rect 230428 144060 230492 144124
rect 248460 144060 248524 144124
rect 288572 143516 288636 143580
rect 170260 142700 170324 142764
rect 237972 142428 238036 142492
rect 230428 141612 230492 141676
rect 232452 141612 232516 141676
rect 230980 141476 231044 141540
rect 231716 141340 231780 141404
rect 229140 141068 229204 141132
rect 266860 140388 266924 140452
rect 284524 140388 284588 140452
rect 244780 139980 244844 140044
rect 241652 138756 241716 138820
rect 237972 138620 238036 138684
rect 267780 138620 267844 138684
rect 229692 137260 229756 137324
rect 279372 135220 279436 135284
rect 231716 134948 231780 135012
rect 233740 134132 233804 134196
rect 264100 133044 264164 133108
rect 230980 132092 231044 132156
rect 262812 131412 262876 131476
rect 250300 129916 250364 129980
rect 231164 128964 231228 129028
rect 267596 128420 267660 128484
rect 242020 127060 242084 127124
rect 280292 126788 280356 126852
rect 244964 126244 245028 126308
rect 230980 125972 231044 126036
rect 231164 119716 231228 119780
rect 166212 119308 166276 119372
rect 290596 117328 290660 117332
rect 290596 117272 290646 117328
rect 290646 117272 290660 117328
rect 290596 117268 290660 117272
rect 229692 114820 229756 114884
rect 263548 109108 263612 109172
rect 244964 105436 245028 105500
rect 260052 103804 260116 103868
rect 168236 103532 168300 103596
rect 263548 102988 263612 103052
rect 285812 102308 285876 102372
rect 244780 100676 244844 100740
rect 232452 98500 232516 98564
rect 237972 97956 238036 98020
rect 229140 97880 229204 97884
rect 229140 97824 229154 97880
rect 229154 97824 229204 97880
rect 229140 97820 229204 97824
rect 229140 97200 229204 97204
rect 229140 97144 229190 97200
rect 229190 97144 229204 97200
rect 229140 97140 229204 97144
rect 284340 97004 284404 97068
rect 268516 96732 268580 96796
rect 263548 95780 263612 95844
rect 223620 95508 223684 95572
rect 228956 95508 229020 95572
rect 223436 95372 223500 95436
rect 228772 95372 228836 95436
rect 201356 95100 201420 95164
rect 268516 94964 268580 95028
rect 107702 94752 107766 94756
rect 107702 94696 107750 94752
rect 107750 94696 107766 94752
rect 107702 94692 107766 94696
rect 117086 94752 117150 94756
rect 117086 94696 117134 94752
rect 117134 94696 117150 94752
rect 117086 94692 117150 94696
rect 151492 94692 151556 94756
rect 151766 94692 151830 94756
rect 99604 94012 99668 94076
rect 219388 94012 219452 94076
rect 91324 93876 91388 93940
rect 114324 93740 114388 93804
rect 129412 93604 129476 93668
rect 95004 93528 95068 93532
rect 95004 93472 95054 93528
rect 95054 93472 95068 93528
rect 95004 93468 95068 93472
rect 115796 93528 115860 93532
rect 115796 93472 115846 93528
rect 115846 93472 115860 93528
rect 115796 93468 115860 93472
rect 103284 93256 103348 93260
rect 103284 93200 103334 93256
rect 103334 93200 103348 93256
rect 103284 93196 103348 93200
rect 110276 93256 110340 93260
rect 110276 93200 110326 93256
rect 110326 93200 110340 93256
rect 110276 93196 110340 93200
rect 260052 93196 260116 93260
rect 267596 93196 267660 93260
rect 267780 92516 267844 92580
rect 86724 92440 86788 92444
rect 86724 92384 86774 92440
rect 86774 92384 86788 92440
rect 86724 92380 86788 92384
rect 88932 92380 88996 92444
rect 101996 92440 102060 92444
rect 101996 92384 102046 92440
rect 102046 92384 102060 92440
rect 101996 92380 102060 92384
rect 112300 92440 112364 92444
rect 112300 92384 112350 92440
rect 112350 92384 112364 92440
rect 112300 92380 112364 92384
rect 132356 92440 132420 92444
rect 132356 92384 132406 92440
rect 132406 92384 132420 92440
rect 132356 92380 132420 92384
rect 134380 92380 134444 92444
rect 136036 92440 136100 92444
rect 136036 92384 136086 92440
rect 136086 92384 136100 92440
rect 136036 92380 136100 92384
rect 85804 92244 85868 92308
rect 122052 92244 122116 92308
rect 115428 92108 115492 92172
rect 255820 91836 255884 91900
rect 99052 91700 99116 91764
rect 119660 91760 119724 91764
rect 119660 91704 119710 91760
rect 119710 91704 119724 91760
rect 119660 91700 119724 91704
rect 121684 91760 121748 91764
rect 121684 91704 121734 91760
rect 121734 91704 121748 91760
rect 121684 91700 121748 91704
rect 123156 91700 123220 91764
rect 178540 91700 178604 91764
rect 106412 91564 106476 91628
rect 106780 91564 106844 91628
rect 122788 91428 122852 91492
rect 125732 91428 125796 91492
rect 151676 91428 151740 91492
rect 96660 91292 96724 91356
rect 98132 91292 98196 91356
rect 100892 91292 100956 91356
rect 109172 91292 109236 91356
rect 111196 91352 111260 91356
rect 111196 91296 111246 91352
rect 111246 91296 111260 91352
rect 111196 91292 111260 91296
rect 114324 91352 114388 91356
rect 114324 91296 114374 91352
rect 114374 91296 114388 91352
rect 114324 91292 114388 91296
rect 124444 91292 124508 91356
rect 126652 91292 126716 91356
rect 151308 91292 151372 91356
rect 74764 91156 74828 91220
rect 84332 91156 84396 91220
rect 88012 91216 88076 91220
rect 88012 91160 88062 91216
rect 88062 91160 88076 91216
rect 88012 91156 88076 91160
rect 90220 91156 90284 91220
rect 92612 91156 92676 91220
rect 93900 91156 93964 91220
rect 96292 91156 96356 91220
rect 97212 91156 97276 91220
rect 98500 91156 98564 91220
rect 100524 91216 100588 91220
rect 100524 91160 100574 91216
rect 100574 91160 100588 91216
rect 100524 91156 100588 91160
rect 101812 91156 101876 91220
rect 102732 91156 102796 91220
rect 104204 91216 104268 91220
rect 104204 91160 104254 91216
rect 104254 91160 104268 91216
rect 104204 91156 104268 91160
rect 104572 91156 104636 91220
rect 105492 91216 105556 91220
rect 105492 91160 105542 91216
rect 105542 91160 105556 91216
rect 105492 91156 105556 91160
rect 105676 91156 105740 91220
rect 108068 91156 108132 91220
rect 109540 91156 109604 91220
rect 110644 91156 110708 91220
rect 111932 91156 111996 91220
rect 113220 91156 113284 91220
rect 114876 91156 114940 91220
rect 116716 91156 116780 91220
rect 118004 91216 118068 91220
rect 118004 91160 118054 91216
rect 118054 91160 118068 91216
rect 118004 91156 118068 91160
rect 118188 91156 118252 91220
rect 119292 91156 119356 91220
rect 120212 91156 120276 91220
rect 120580 91156 120644 91220
rect 124076 91156 124140 91220
rect 125364 91216 125428 91220
rect 125364 91160 125414 91216
rect 125414 91160 125428 91216
rect 125364 91156 125428 91160
rect 126468 91156 126532 91220
rect 127572 91156 127636 91220
rect 130700 91216 130764 91220
rect 130700 91160 130750 91216
rect 130750 91160 130764 91216
rect 130700 91156 130764 91160
rect 133092 91156 133156 91220
rect 151492 91156 151556 91220
rect 152044 91216 152108 91220
rect 152044 91160 152094 91216
rect 152094 91160 152108 91216
rect 152044 91156 152108 91160
rect 215156 90340 215220 90404
rect 227668 90340 227732 90404
rect 166212 89796 166276 89860
rect 223436 88164 223500 88228
rect 168236 78372 168300 78436
rect 53604 75108 53668 75172
rect 262812 71028 262876 71092
rect 168420 69668 168484 69732
rect 362908 67492 362972 67556
rect 61884 66812 61948 66876
rect 242020 61372 242084 61436
rect 229692 57156 229756 57220
rect 250300 50220 250364 50284
rect 264100 44780 264164 44844
rect 230980 42060 231044 42124
rect 65380 37844 65444 37908
rect 258580 37164 258644 37228
rect 266860 35124 266924 35188
rect 67772 33900 67836 33964
rect 219204 33764 219268 33828
rect 233740 26828 233804 26892
rect 295380 22612 295444 22676
rect 253060 22068 253124 22132
rect 165660 21252 165724 21316
rect 303660 19892 303724 19956
rect 173756 18532 173820 18596
rect 189948 17308 190012 17372
rect 223620 17172 223684 17236
rect 185348 12956 185412 13020
rect 363092 10236 363156 10300
rect 180564 9012 180628 9076
rect 227668 8876 227732 8940
rect 170444 7516 170508 7580
rect 356100 4796 356164 4860
rect 246252 3436 246316 3500
rect 251772 3436 251836 3500
rect 285628 3436 285692 3500
rect 287652 3436 287716 3500
rect 291148 3436 291212 3500
rect 293172 3436 293236 3500
rect 299612 3436 299676 3500
rect 241284 3300 241348 3364
rect 298140 3300 298204 3364
rect 302740 3300 302804 3364
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 680614 -8106 711002
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 -8106 680614
rect -8726 680294 -8106 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 -8106 680294
rect -8726 644614 -8106 680058
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 -8106 644614
rect -8726 644294 -8106 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 -8106 644294
rect -8726 608614 -8106 644058
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 -8106 608614
rect -8726 608294 -8106 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 -8106 608294
rect -8726 572614 -8106 608058
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 -8106 572614
rect -8726 572294 -8106 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 -8106 572294
rect -8726 536614 -8106 572058
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 -8106 536614
rect -8726 536294 -8106 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 -8106 536294
rect -8726 500614 -8106 536058
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 -8106 500614
rect -8726 500294 -8106 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 -8106 500294
rect -8726 464614 -8106 500058
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 -8106 464614
rect -8726 464294 -8106 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 -8106 464294
rect -8726 428614 -8106 464058
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 -8106 428614
rect -8726 428294 -8106 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 -8106 428294
rect -8726 392614 -8106 428058
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 -8106 392614
rect -8726 392294 -8106 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 -8106 392294
rect -8726 356614 -8106 392058
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 -8106 356614
rect -8726 356294 -8106 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 -8106 356294
rect -8726 320614 -8106 356058
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 -8106 320614
rect -8726 320294 -8106 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 -8106 320294
rect -8726 284614 -8106 320058
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 -8106 284614
rect -8726 284294 -8106 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 -8106 284294
rect -8726 248614 -8106 284058
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 -8106 248614
rect -8726 248294 -8106 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 -8106 248294
rect -8726 212614 -8106 248058
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 -8106 212614
rect -8726 212294 -8106 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 -8106 212294
rect -8726 176614 -8106 212058
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 -8106 176614
rect -8726 176294 -8106 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 -8106 176294
rect -8726 140614 -8106 176058
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 -8106 140614
rect -8726 140294 -8106 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 -8106 140294
rect -8726 104614 -8106 140058
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 -8106 104614
rect -8726 104294 -8106 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 -8106 104294
rect -8726 68614 -8106 104058
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 -8106 68614
rect -8726 68294 -8106 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 -8106 68294
rect -8726 32614 -8106 68058
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 -8106 32614
rect -8726 32294 -8106 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 -8106 32294
rect -8726 -7066 -8106 32058
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 698614 -7146 710042
rect 12954 710598 13574 711590
rect 12954 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 13574 710598
rect 12954 710278 13574 710362
rect 12954 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 13574 710278
rect -7766 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 -7146 698614
rect -7766 698294 -7146 698378
rect -7766 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 -7146 698294
rect -7766 662614 -7146 698058
rect -7766 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 -7146 662614
rect -7766 662294 -7146 662378
rect -7766 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 -7146 662294
rect -7766 626614 -7146 662058
rect -7766 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 -7146 626614
rect -7766 626294 -7146 626378
rect -7766 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 -7146 626294
rect -7766 590614 -7146 626058
rect -7766 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 -7146 590614
rect -7766 590294 -7146 590378
rect -7766 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 -7146 590294
rect -7766 554614 -7146 590058
rect -7766 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 -7146 554614
rect -7766 554294 -7146 554378
rect -7766 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 -7146 554294
rect -7766 518614 -7146 554058
rect -7766 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 -7146 518614
rect -7766 518294 -7146 518378
rect -7766 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 -7146 518294
rect -7766 482614 -7146 518058
rect -7766 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 -7146 482614
rect -7766 482294 -7146 482378
rect -7766 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 -7146 482294
rect -7766 446614 -7146 482058
rect -7766 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 -7146 446614
rect -7766 446294 -7146 446378
rect -7766 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 -7146 446294
rect -7766 410614 -7146 446058
rect -7766 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 -7146 410614
rect -7766 410294 -7146 410378
rect -7766 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 -7146 410294
rect -7766 374614 -7146 410058
rect -7766 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 -7146 374614
rect -7766 374294 -7146 374378
rect -7766 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 -7146 374294
rect -7766 338614 -7146 374058
rect -7766 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 -7146 338614
rect -7766 338294 -7146 338378
rect -7766 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 -7146 338294
rect -7766 302614 -7146 338058
rect -7766 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 -7146 302614
rect -7766 302294 -7146 302378
rect -7766 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 -7146 302294
rect -7766 266614 -7146 302058
rect -7766 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 -7146 266614
rect -7766 266294 -7146 266378
rect -7766 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 -7146 266294
rect -7766 230614 -7146 266058
rect -7766 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 -7146 230614
rect -7766 230294 -7146 230378
rect -7766 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 -7146 230294
rect -7766 194614 -7146 230058
rect -7766 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 -7146 194614
rect -7766 194294 -7146 194378
rect -7766 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 -7146 194294
rect -7766 158614 -7146 194058
rect -7766 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 -7146 158614
rect -7766 158294 -7146 158378
rect -7766 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 -7146 158294
rect -7766 122614 -7146 158058
rect -7766 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 -7146 122614
rect -7766 122294 -7146 122378
rect -7766 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 -7146 122294
rect -7766 86614 -7146 122058
rect -7766 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 -7146 86614
rect -7766 86294 -7146 86378
rect -7766 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 -7146 86294
rect -7766 50614 -7146 86058
rect -7766 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 -7146 50614
rect -7766 50294 -7146 50378
rect -7766 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 -7146 50294
rect -7766 14614 -7146 50058
rect -7766 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 -7146 14614
rect -7766 14294 -7146 14378
rect -7766 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 -7146 14294
rect -7766 -6106 -7146 14058
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 676894 -6186 709082
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 -6186 676894
rect -6806 676574 -6186 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 -6186 676574
rect -6806 640894 -6186 676338
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 -6186 640894
rect -6806 640574 -6186 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 -6186 640574
rect -6806 604894 -6186 640338
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 -6186 604894
rect -6806 604574 -6186 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 -6186 604574
rect -6806 568894 -6186 604338
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 -6186 568894
rect -6806 568574 -6186 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 -6186 568574
rect -6806 532894 -6186 568338
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 -6186 532894
rect -6806 532574 -6186 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 -6186 532574
rect -6806 496894 -6186 532338
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 -6186 496894
rect -6806 496574 -6186 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 -6186 496574
rect -6806 460894 -6186 496338
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 -6186 460894
rect -6806 460574 -6186 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 -6186 460574
rect -6806 424894 -6186 460338
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 -6186 424894
rect -6806 424574 -6186 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 -6186 424574
rect -6806 388894 -6186 424338
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 -6186 388894
rect -6806 388574 -6186 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 -6186 388574
rect -6806 352894 -6186 388338
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 -6186 352894
rect -6806 352574 -6186 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 -6186 352574
rect -6806 316894 -6186 352338
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 -6186 316894
rect -6806 316574 -6186 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 -6186 316574
rect -6806 280894 -6186 316338
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 -6186 280894
rect -6806 280574 -6186 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 -6186 280574
rect -6806 244894 -6186 280338
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 -6186 244894
rect -6806 244574 -6186 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 -6186 244574
rect -6806 208894 -6186 244338
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 -6186 208894
rect -6806 208574 -6186 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 -6186 208574
rect -6806 172894 -6186 208338
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 -6186 172894
rect -6806 172574 -6186 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 -6186 172574
rect -6806 136894 -6186 172338
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 -6186 136894
rect -6806 136574 -6186 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 -6186 136574
rect -6806 100894 -6186 136338
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 -6186 100894
rect -6806 100574 -6186 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 -6186 100574
rect -6806 64894 -6186 100338
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 -6186 64894
rect -6806 64574 -6186 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 -6186 64574
rect -6806 28894 -6186 64338
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 -6186 28894
rect -6806 28574 -6186 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 -6186 28574
rect -6806 -5146 -6186 28338
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 694894 -5226 708122
rect 9234 708678 9854 709670
rect 9234 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 9854 708678
rect 9234 708358 9854 708442
rect 9234 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 9854 708358
rect -5846 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 -5226 694894
rect -5846 694574 -5226 694658
rect -5846 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 -5226 694574
rect -5846 658894 -5226 694338
rect -5846 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 -5226 658894
rect -5846 658574 -5226 658658
rect -5846 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 -5226 658574
rect -5846 622894 -5226 658338
rect -5846 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 -5226 622894
rect -5846 622574 -5226 622658
rect -5846 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 -5226 622574
rect -5846 586894 -5226 622338
rect -5846 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 -5226 586894
rect -5846 586574 -5226 586658
rect -5846 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 -5226 586574
rect -5846 550894 -5226 586338
rect -5846 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 -5226 550894
rect -5846 550574 -5226 550658
rect -5846 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 -5226 550574
rect -5846 514894 -5226 550338
rect -5846 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 -5226 514894
rect -5846 514574 -5226 514658
rect -5846 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 -5226 514574
rect -5846 478894 -5226 514338
rect -5846 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 -5226 478894
rect -5846 478574 -5226 478658
rect -5846 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 -5226 478574
rect -5846 442894 -5226 478338
rect -5846 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 -5226 442894
rect -5846 442574 -5226 442658
rect -5846 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 -5226 442574
rect -5846 406894 -5226 442338
rect -5846 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 -5226 406894
rect -5846 406574 -5226 406658
rect -5846 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 -5226 406574
rect -5846 370894 -5226 406338
rect -5846 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 -5226 370894
rect -5846 370574 -5226 370658
rect -5846 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 -5226 370574
rect -5846 334894 -5226 370338
rect -5846 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 -5226 334894
rect -5846 334574 -5226 334658
rect -5846 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 -5226 334574
rect -5846 298894 -5226 334338
rect -5846 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 -5226 298894
rect -5846 298574 -5226 298658
rect -5846 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 -5226 298574
rect -5846 262894 -5226 298338
rect -5846 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 -5226 262894
rect -5846 262574 -5226 262658
rect -5846 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 -5226 262574
rect -5846 226894 -5226 262338
rect -5846 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 -5226 226894
rect -5846 226574 -5226 226658
rect -5846 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 -5226 226574
rect -5846 190894 -5226 226338
rect -5846 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 -5226 190894
rect -5846 190574 -5226 190658
rect -5846 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 -5226 190574
rect -5846 154894 -5226 190338
rect -5846 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 -5226 154894
rect -5846 154574 -5226 154658
rect -5846 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 -5226 154574
rect -5846 118894 -5226 154338
rect -5846 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 -5226 118894
rect -5846 118574 -5226 118658
rect -5846 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 -5226 118574
rect -5846 82894 -5226 118338
rect -5846 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 -5226 82894
rect -5846 82574 -5226 82658
rect -5846 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 -5226 82574
rect -5846 46894 -5226 82338
rect -5846 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 -5226 46894
rect -5846 46574 -5226 46658
rect -5846 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 -5226 46574
rect -5846 10894 -5226 46338
rect -5846 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 -5226 10894
rect -5846 10574 -5226 10658
rect -5846 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 -5226 10574
rect -5846 -4186 -5226 10338
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 673174 -4266 707162
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 -4266 673174
rect -4886 672854 -4266 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 -4266 672854
rect -4886 637174 -4266 672618
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 -4266 637174
rect -4886 636854 -4266 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 -4266 636854
rect -4886 601174 -4266 636618
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 -4266 601174
rect -4886 600854 -4266 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 -4266 600854
rect -4886 565174 -4266 600618
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 -4266 565174
rect -4886 564854 -4266 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 -4266 564854
rect -4886 529174 -4266 564618
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 -4266 529174
rect -4886 528854 -4266 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 -4266 528854
rect -4886 493174 -4266 528618
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 -4266 493174
rect -4886 492854 -4266 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 -4266 492854
rect -4886 457174 -4266 492618
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 -4266 457174
rect -4886 456854 -4266 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 -4266 456854
rect -4886 421174 -4266 456618
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 -4266 421174
rect -4886 420854 -4266 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 -4266 420854
rect -4886 385174 -4266 420618
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 -4266 385174
rect -4886 384854 -4266 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 -4266 384854
rect -4886 349174 -4266 384618
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 -4266 349174
rect -4886 348854 -4266 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 -4266 348854
rect -4886 313174 -4266 348618
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 -4266 313174
rect -4886 312854 -4266 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 -4266 312854
rect -4886 277174 -4266 312618
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 -4266 277174
rect -4886 276854 -4266 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 -4266 276854
rect -4886 241174 -4266 276618
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 -4266 241174
rect -4886 240854 -4266 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 -4266 240854
rect -4886 205174 -4266 240618
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 -4266 205174
rect -4886 204854 -4266 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 -4266 204854
rect -4886 169174 -4266 204618
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 -4266 169174
rect -4886 168854 -4266 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 -4266 168854
rect -4886 133174 -4266 168618
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 -4266 133174
rect -4886 132854 -4266 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 -4266 132854
rect -4886 97174 -4266 132618
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 -4266 97174
rect -4886 96854 -4266 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 -4266 96854
rect -4886 61174 -4266 96618
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 -4266 61174
rect -4886 60854 -4266 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 -4266 60854
rect -4886 25174 -4266 60618
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 -4266 25174
rect -4886 24854 -4266 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 -4266 24854
rect -4886 -3226 -4266 24618
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 691174 -3306 706202
rect 5514 706758 6134 707750
rect 5514 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 6134 706758
rect 5514 706438 6134 706522
rect 5514 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 6134 706438
rect -3926 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 -3306 691174
rect -3926 690854 -3306 690938
rect -3926 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 -3306 690854
rect -3926 655174 -3306 690618
rect -3926 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 -3306 655174
rect -3926 654854 -3306 654938
rect -3926 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 -3306 654854
rect -3926 619174 -3306 654618
rect -3926 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 -3306 619174
rect -3926 618854 -3306 618938
rect -3926 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 -3306 618854
rect -3926 583174 -3306 618618
rect -3926 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 -3306 583174
rect -3926 582854 -3306 582938
rect -3926 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 -3306 582854
rect -3926 547174 -3306 582618
rect -3926 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 -3306 547174
rect -3926 546854 -3306 546938
rect -3926 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 -3306 546854
rect -3926 511174 -3306 546618
rect -3926 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 -3306 511174
rect -3926 510854 -3306 510938
rect -3926 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 -3306 510854
rect -3926 475174 -3306 510618
rect -3926 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 -3306 475174
rect -3926 474854 -3306 474938
rect -3926 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 -3306 474854
rect -3926 439174 -3306 474618
rect -3926 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 -3306 439174
rect -3926 438854 -3306 438938
rect -3926 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 -3306 438854
rect -3926 403174 -3306 438618
rect -3926 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 -3306 403174
rect -3926 402854 -3306 402938
rect -3926 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 -3306 402854
rect -3926 367174 -3306 402618
rect -3926 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 -3306 367174
rect -3926 366854 -3306 366938
rect -3926 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 -3306 366854
rect -3926 331174 -3306 366618
rect -3926 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 -3306 331174
rect -3926 330854 -3306 330938
rect -3926 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 -3306 330854
rect -3926 295174 -3306 330618
rect -3926 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 -3306 295174
rect -3926 294854 -3306 294938
rect -3926 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 -3306 294854
rect -3926 259174 -3306 294618
rect -3926 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 -3306 259174
rect -3926 258854 -3306 258938
rect -3926 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 -3306 258854
rect -3926 223174 -3306 258618
rect -3926 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 -3306 223174
rect -3926 222854 -3306 222938
rect -3926 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 -3306 222854
rect -3926 187174 -3306 222618
rect -3926 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 -3306 187174
rect -3926 186854 -3306 186938
rect -3926 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 -3306 186854
rect -3926 151174 -3306 186618
rect -3926 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 -3306 151174
rect -3926 150854 -3306 150938
rect -3926 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 -3306 150854
rect -3926 115174 -3306 150618
rect -3926 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 -3306 115174
rect -3926 114854 -3306 114938
rect -3926 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 -3306 114854
rect -3926 79174 -3306 114618
rect -3926 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 -3306 79174
rect -3926 78854 -3306 78938
rect -3926 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 -3306 78854
rect -3926 43174 -3306 78618
rect -3926 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 -3306 43174
rect -3926 42854 -3306 42938
rect -3926 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 -3306 42854
rect -3926 7174 -3306 42618
rect -3926 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 -3306 7174
rect -3926 6854 -3306 6938
rect -3926 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 -3306 6854
rect -3926 -2266 -3306 6618
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 669454 -2346 705242
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 -2346 669454
rect -2966 669134 -2346 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 -2346 669134
rect -2966 633454 -2346 668898
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 -2346 633454
rect -2966 633134 -2346 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 -2346 633134
rect -2966 597454 -2346 632898
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 -2346 597454
rect -2966 597134 -2346 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 -2346 597134
rect -2966 561454 -2346 596898
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 -2346 561454
rect -2966 561134 -2346 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 -2346 561134
rect -2966 525454 -2346 560898
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 -2346 525454
rect -2966 525134 -2346 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 -2346 525134
rect -2966 489454 -2346 524898
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 -2346 489454
rect -2966 489134 -2346 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 -2346 489134
rect -2966 453454 -2346 488898
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 -2346 453454
rect -2966 453134 -2346 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 -2346 453134
rect -2966 417454 -2346 452898
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 -2346 417454
rect -2966 417134 -2346 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 -2346 417134
rect -2966 381454 -2346 416898
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 -2346 381454
rect -2966 381134 -2346 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 -2346 381134
rect -2966 345454 -2346 380898
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 -2346 345454
rect -2966 345134 -2346 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 -2346 345134
rect -2966 309454 -2346 344898
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 -2346 309454
rect -2966 309134 -2346 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 -2346 309134
rect -2966 273454 -2346 308898
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 -2346 273454
rect -2966 273134 -2346 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 -2346 273134
rect -2966 237454 -2346 272898
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 -2346 237454
rect -2966 237134 -2346 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 -2346 237134
rect -2966 201454 -2346 236898
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 -2346 201454
rect -2966 201134 -2346 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 -2346 201134
rect -2966 165454 -2346 200898
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 -2346 165454
rect -2966 165134 -2346 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 -2346 165134
rect -2966 129454 -2346 164898
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 -2346 129454
rect -2966 129134 -2346 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 -2346 129134
rect -2966 93454 -2346 128898
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 -2346 93454
rect -2966 93134 -2346 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 -2346 93134
rect -2966 57454 -2346 92898
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 -2346 57454
rect -2966 57134 -2346 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 -2346 57134
rect -2966 21454 -2346 56898
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 -2346 21454
rect -2966 21134 -2346 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 -2346 21134
rect -2966 -1306 -2346 20898
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 705830
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect 1794 -1894 2414 -902
rect 5514 691174 6134 706202
rect 5514 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 6134 691174
rect 5514 690854 6134 690938
rect 5514 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 6134 690854
rect 5514 655174 6134 690618
rect 5514 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 6134 655174
rect 5514 654854 6134 654938
rect 5514 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 6134 654854
rect 5514 619174 6134 654618
rect 5514 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 6134 619174
rect 5514 618854 6134 618938
rect 5514 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 6134 618854
rect 5514 583174 6134 618618
rect 5514 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 6134 583174
rect 5514 582854 6134 582938
rect 5514 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 6134 582854
rect 5514 547174 6134 582618
rect 5514 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 6134 547174
rect 5514 546854 6134 546938
rect 5514 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 6134 546854
rect 5514 511174 6134 546618
rect 5514 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 6134 511174
rect 5514 510854 6134 510938
rect 5514 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 6134 510854
rect 5514 475174 6134 510618
rect 5514 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 6134 475174
rect 5514 474854 6134 474938
rect 5514 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 6134 474854
rect 5514 439174 6134 474618
rect 5514 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 6134 439174
rect 5514 438854 6134 438938
rect 5514 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 6134 438854
rect 5514 403174 6134 438618
rect 5514 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 6134 403174
rect 5514 402854 6134 402938
rect 5514 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 6134 402854
rect 5514 367174 6134 402618
rect 5514 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 6134 367174
rect 5514 366854 6134 366938
rect 5514 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 6134 366854
rect 5514 331174 6134 366618
rect 5514 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 6134 331174
rect 5514 330854 6134 330938
rect 5514 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 6134 330854
rect 5514 295174 6134 330618
rect 5514 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 6134 295174
rect 5514 294854 6134 294938
rect 5514 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 6134 294854
rect 5514 259174 6134 294618
rect 5514 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 6134 259174
rect 5514 258854 6134 258938
rect 5514 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 6134 258854
rect 5514 223174 6134 258618
rect 5514 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 6134 223174
rect 5514 222854 6134 222938
rect 5514 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 6134 222854
rect 5514 187174 6134 222618
rect 5514 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 6134 187174
rect 5514 186854 6134 186938
rect 5514 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 6134 186854
rect 5514 151174 6134 186618
rect 5514 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 6134 151174
rect 5514 150854 6134 150938
rect 5514 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 6134 150854
rect 5514 115174 6134 150618
rect 5514 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 6134 115174
rect 5514 114854 6134 114938
rect 5514 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 6134 114854
rect 5514 79174 6134 114618
rect 5514 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 6134 79174
rect 5514 78854 6134 78938
rect 5514 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 6134 78854
rect 5514 43174 6134 78618
rect 5514 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 6134 43174
rect 5514 42854 6134 42938
rect 5514 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 6134 42854
rect 5514 7174 6134 42618
rect 5514 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 6134 7174
rect 5514 6854 6134 6938
rect 5514 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 6134 6854
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect 5514 -2266 6134 6618
rect 5514 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 6134 -2266
rect 5514 -2586 6134 -2502
rect 5514 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 6134 -2586
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect 5514 -3814 6134 -2822
rect 9234 694894 9854 708122
rect 9234 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 9854 694894
rect 9234 694574 9854 694658
rect 9234 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 9854 694574
rect 9234 658894 9854 694338
rect 9234 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 9854 658894
rect 9234 658574 9854 658658
rect 9234 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 9854 658574
rect 9234 622894 9854 658338
rect 9234 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 9854 622894
rect 9234 622574 9854 622658
rect 9234 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 9854 622574
rect 9234 586894 9854 622338
rect 9234 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 9854 586894
rect 9234 586574 9854 586658
rect 9234 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 9854 586574
rect 9234 550894 9854 586338
rect 9234 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 9854 550894
rect 9234 550574 9854 550658
rect 9234 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 9854 550574
rect 9234 514894 9854 550338
rect 9234 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 9854 514894
rect 9234 514574 9854 514658
rect 9234 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 9854 514574
rect 9234 478894 9854 514338
rect 9234 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 9854 478894
rect 9234 478574 9854 478658
rect 9234 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 9854 478574
rect 9234 442894 9854 478338
rect 9234 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 9854 442894
rect 9234 442574 9854 442658
rect 9234 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 9854 442574
rect 9234 406894 9854 442338
rect 9234 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 9854 406894
rect 9234 406574 9854 406658
rect 9234 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 9854 406574
rect 9234 370894 9854 406338
rect 9234 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 9854 370894
rect 9234 370574 9854 370658
rect 9234 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 9854 370574
rect 9234 334894 9854 370338
rect 9234 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 9854 334894
rect 9234 334574 9854 334658
rect 9234 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 9854 334574
rect 9234 298894 9854 334338
rect 9234 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 9854 298894
rect 9234 298574 9854 298658
rect 9234 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 9854 298574
rect 9234 262894 9854 298338
rect 9234 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 9854 262894
rect 9234 262574 9854 262658
rect 9234 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 9854 262574
rect 9234 226894 9854 262338
rect 9234 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 9854 226894
rect 9234 226574 9854 226658
rect 9234 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 9854 226574
rect 9234 190894 9854 226338
rect 9234 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 9854 190894
rect 9234 190574 9854 190658
rect 9234 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 9854 190574
rect 9234 154894 9854 190338
rect 9234 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 9854 154894
rect 9234 154574 9854 154658
rect 9234 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 9854 154574
rect 9234 118894 9854 154338
rect 9234 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 9854 118894
rect 9234 118574 9854 118658
rect 9234 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 9854 118574
rect 9234 82894 9854 118338
rect 9234 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 9854 82894
rect 9234 82574 9854 82658
rect 9234 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 9854 82574
rect 9234 46894 9854 82338
rect 9234 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 9854 46894
rect 9234 46574 9854 46658
rect 9234 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 9854 46574
rect 9234 10894 9854 46338
rect 9234 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 9854 10894
rect 9234 10574 9854 10658
rect 9234 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 9854 10574
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect 9234 -4186 9854 10338
rect 9234 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 9854 -4186
rect 9234 -4506 9854 -4422
rect 9234 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 9854 -4506
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect 9234 -5734 9854 -4742
rect 12954 698614 13574 710042
rect 30954 711558 31574 711590
rect 30954 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 31574 711558
rect 30954 711238 31574 711322
rect 30954 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 31574 711238
rect 27234 709638 27854 709670
rect 27234 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 27854 709638
rect 27234 709318 27854 709402
rect 27234 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 27854 709318
rect 23514 707718 24134 707750
rect 23514 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 24134 707718
rect 23514 707398 24134 707482
rect 23514 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 24134 707398
rect 12954 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 13574 698614
rect 12954 698294 13574 698378
rect 12954 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 13574 698294
rect 12954 662614 13574 698058
rect 12954 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 13574 662614
rect 12954 662294 13574 662378
rect 12954 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 13574 662294
rect 12954 626614 13574 662058
rect 12954 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 13574 626614
rect 12954 626294 13574 626378
rect 12954 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 13574 626294
rect 12954 590614 13574 626058
rect 12954 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 13574 590614
rect 12954 590294 13574 590378
rect 12954 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 13574 590294
rect 12954 554614 13574 590058
rect 12954 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 13574 554614
rect 12954 554294 13574 554378
rect 12954 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 13574 554294
rect 12954 518614 13574 554058
rect 12954 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 13574 518614
rect 12954 518294 13574 518378
rect 12954 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 13574 518294
rect 12954 482614 13574 518058
rect 12954 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 13574 482614
rect 12954 482294 13574 482378
rect 12954 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 13574 482294
rect 12954 446614 13574 482058
rect 12954 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 13574 446614
rect 12954 446294 13574 446378
rect 12954 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 13574 446294
rect 12954 410614 13574 446058
rect 12954 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 13574 410614
rect 12954 410294 13574 410378
rect 12954 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 13574 410294
rect 12954 374614 13574 410058
rect 12954 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 13574 374614
rect 12954 374294 13574 374378
rect 12954 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 13574 374294
rect 12954 338614 13574 374058
rect 12954 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 13574 338614
rect 12954 338294 13574 338378
rect 12954 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 13574 338294
rect 12954 302614 13574 338058
rect 12954 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 13574 302614
rect 12954 302294 13574 302378
rect 12954 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 13574 302294
rect 12954 266614 13574 302058
rect 12954 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 13574 266614
rect 12954 266294 13574 266378
rect 12954 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 13574 266294
rect 12954 230614 13574 266058
rect 12954 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 13574 230614
rect 12954 230294 13574 230378
rect 12954 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 13574 230294
rect 12954 194614 13574 230058
rect 12954 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 13574 194614
rect 12954 194294 13574 194378
rect 12954 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 13574 194294
rect 12954 158614 13574 194058
rect 12954 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 13574 158614
rect 12954 158294 13574 158378
rect 12954 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 13574 158294
rect 12954 122614 13574 158058
rect 12954 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 13574 122614
rect 12954 122294 13574 122378
rect 12954 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 13574 122294
rect 12954 86614 13574 122058
rect 12954 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 13574 86614
rect 12954 86294 13574 86378
rect 12954 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 13574 86294
rect 12954 50614 13574 86058
rect 12954 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 13574 50614
rect 12954 50294 13574 50378
rect 12954 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 13574 50294
rect 12954 14614 13574 50058
rect 12954 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 13574 14614
rect 12954 14294 13574 14378
rect 12954 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 13574 14294
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect 12954 -6106 13574 14058
rect 19794 705798 20414 705830
rect 19794 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 20414 705798
rect 19794 705478 20414 705562
rect 19794 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 20414 705478
rect 19794 669454 20414 705242
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -1306 20414 20898
rect 19794 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 20414 -1306
rect 19794 -1626 20414 -1542
rect 19794 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 20414 -1626
rect 19794 -1894 20414 -1862
rect 23514 673174 24134 707162
rect 23514 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 24134 673174
rect 23514 672854 24134 672938
rect 23514 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 24134 672854
rect 23514 637174 24134 672618
rect 23514 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 24134 637174
rect 23514 636854 24134 636938
rect 23514 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 24134 636854
rect 23514 601174 24134 636618
rect 23514 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 24134 601174
rect 23514 600854 24134 600938
rect 23514 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 24134 600854
rect 23514 565174 24134 600618
rect 23514 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 24134 565174
rect 23514 564854 24134 564938
rect 23514 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 24134 564854
rect 23514 529174 24134 564618
rect 23514 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 24134 529174
rect 23514 528854 24134 528938
rect 23514 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 24134 528854
rect 23514 493174 24134 528618
rect 23514 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 24134 493174
rect 23514 492854 24134 492938
rect 23514 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 24134 492854
rect 23514 457174 24134 492618
rect 23514 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 24134 457174
rect 23514 456854 24134 456938
rect 23514 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 24134 456854
rect 23514 421174 24134 456618
rect 23514 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 24134 421174
rect 23514 420854 24134 420938
rect 23514 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 24134 420854
rect 23514 385174 24134 420618
rect 23514 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 24134 385174
rect 23514 384854 24134 384938
rect 23514 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 24134 384854
rect 23514 349174 24134 384618
rect 23514 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 24134 349174
rect 23514 348854 24134 348938
rect 23514 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 24134 348854
rect 23514 313174 24134 348618
rect 23514 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 24134 313174
rect 23514 312854 24134 312938
rect 23514 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 24134 312854
rect 23514 277174 24134 312618
rect 23514 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 24134 277174
rect 23514 276854 24134 276938
rect 23514 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 24134 276854
rect 23514 241174 24134 276618
rect 23514 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 24134 241174
rect 23514 240854 24134 240938
rect 23514 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 24134 240854
rect 23514 205174 24134 240618
rect 23514 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 24134 205174
rect 23514 204854 24134 204938
rect 23514 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 24134 204854
rect 23514 169174 24134 204618
rect 23514 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 24134 169174
rect 23514 168854 24134 168938
rect 23514 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 24134 168854
rect 23514 133174 24134 168618
rect 23514 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 24134 133174
rect 23514 132854 24134 132938
rect 23514 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 24134 132854
rect 23514 97174 24134 132618
rect 23514 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 24134 97174
rect 23514 96854 24134 96938
rect 23514 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 24134 96854
rect 23514 61174 24134 96618
rect 23514 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 24134 61174
rect 23514 60854 24134 60938
rect 23514 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 24134 60854
rect 23514 25174 24134 60618
rect 23514 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 24134 25174
rect 23514 24854 24134 24938
rect 23514 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 24134 24854
rect 23514 -3226 24134 24618
rect 23514 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 24134 -3226
rect 23514 -3546 24134 -3462
rect 23514 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 24134 -3546
rect 23514 -3814 24134 -3782
rect 27234 676894 27854 709082
rect 27234 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 27854 676894
rect 27234 676574 27854 676658
rect 27234 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 27854 676574
rect 27234 640894 27854 676338
rect 27234 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 27854 640894
rect 27234 640574 27854 640658
rect 27234 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 27854 640574
rect 27234 604894 27854 640338
rect 27234 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 27854 604894
rect 27234 604574 27854 604658
rect 27234 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 27854 604574
rect 27234 568894 27854 604338
rect 27234 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 27854 568894
rect 27234 568574 27854 568658
rect 27234 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 27854 568574
rect 27234 532894 27854 568338
rect 27234 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 27854 532894
rect 27234 532574 27854 532658
rect 27234 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 27854 532574
rect 27234 496894 27854 532338
rect 27234 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 27854 496894
rect 27234 496574 27854 496658
rect 27234 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 27854 496574
rect 27234 460894 27854 496338
rect 27234 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 27854 460894
rect 27234 460574 27854 460658
rect 27234 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 27854 460574
rect 27234 424894 27854 460338
rect 27234 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 27854 424894
rect 27234 424574 27854 424658
rect 27234 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 27854 424574
rect 27234 388894 27854 424338
rect 27234 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 27854 388894
rect 27234 388574 27854 388658
rect 27234 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 27854 388574
rect 27234 352894 27854 388338
rect 27234 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 27854 352894
rect 27234 352574 27854 352658
rect 27234 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 27854 352574
rect 27234 316894 27854 352338
rect 27234 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 27854 316894
rect 27234 316574 27854 316658
rect 27234 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 27854 316574
rect 27234 280894 27854 316338
rect 27234 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 27854 280894
rect 27234 280574 27854 280658
rect 27234 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 27854 280574
rect 27234 244894 27854 280338
rect 27234 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 27854 244894
rect 27234 244574 27854 244658
rect 27234 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 27854 244574
rect 27234 208894 27854 244338
rect 27234 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 27854 208894
rect 27234 208574 27854 208658
rect 27234 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 27854 208574
rect 27234 172894 27854 208338
rect 27234 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 27854 172894
rect 27234 172574 27854 172658
rect 27234 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 27854 172574
rect 27234 136894 27854 172338
rect 27234 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 27854 136894
rect 27234 136574 27854 136658
rect 27234 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 27854 136574
rect 27234 100894 27854 136338
rect 27234 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 27854 100894
rect 27234 100574 27854 100658
rect 27234 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 27854 100574
rect 27234 64894 27854 100338
rect 27234 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 27854 64894
rect 27234 64574 27854 64658
rect 27234 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 27854 64574
rect 27234 28894 27854 64338
rect 27234 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 27854 28894
rect 27234 28574 27854 28658
rect 27234 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 27854 28574
rect 27234 -5146 27854 28338
rect 27234 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 27854 -5146
rect 27234 -5466 27854 -5382
rect 27234 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 27854 -5466
rect 27234 -5734 27854 -5702
rect 30954 680614 31574 711002
rect 48954 710598 49574 711590
rect 48954 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 49574 710598
rect 48954 710278 49574 710362
rect 48954 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 49574 710278
rect 45234 708678 45854 709670
rect 45234 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 45854 708678
rect 45234 708358 45854 708442
rect 45234 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 45854 708358
rect 41514 706758 42134 707750
rect 41514 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 42134 706758
rect 41514 706438 42134 706522
rect 41514 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 42134 706438
rect 30954 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 31574 680614
rect 30954 680294 31574 680378
rect 30954 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 31574 680294
rect 30954 644614 31574 680058
rect 30954 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 31574 644614
rect 30954 644294 31574 644378
rect 30954 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 31574 644294
rect 30954 608614 31574 644058
rect 30954 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 31574 608614
rect 30954 608294 31574 608378
rect 30954 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 31574 608294
rect 30954 572614 31574 608058
rect 30954 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 31574 572614
rect 30954 572294 31574 572378
rect 30954 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 31574 572294
rect 30954 536614 31574 572058
rect 30954 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 31574 536614
rect 30954 536294 31574 536378
rect 30954 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 31574 536294
rect 30954 500614 31574 536058
rect 30954 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 31574 500614
rect 30954 500294 31574 500378
rect 30954 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 31574 500294
rect 30954 464614 31574 500058
rect 30954 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 31574 464614
rect 30954 464294 31574 464378
rect 30954 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 31574 464294
rect 30954 428614 31574 464058
rect 30954 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 31574 428614
rect 30954 428294 31574 428378
rect 30954 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 31574 428294
rect 30954 392614 31574 428058
rect 30954 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 31574 392614
rect 30954 392294 31574 392378
rect 30954 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 31574 392294
rect 30954 356614 31574 392058
rect 30954 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 31574 356614
rect 30954 356294 31574 356378
rect 30954 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 31574 356294
rect 30954 320614 31574 356058
rect 30954 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 31574 320614
rect 30954 320294 31574 320378
rect 30954 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 31574 320294
rect 30954 284614 31574 320058
rect 30954 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 31574 284614
rect 30954 284294 31574 284378
rect 30954 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 31574 284294
rect 30954 248614 31574 284058
rect 30954 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 31574 248614
rect 30954 248294 31574 248378
rect 30954 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 31574 248294
rect 30954 212614 31574 248058
rect 30954 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 31574 212614
rect 30954 212294 31574 212378
rect 30954 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 31574 212294
rect 30954 176614 31574 212058
rect 30954 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 31574 176614
rect 30954 176294 31574 176378
rect 30954 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 31574 176294
rect 30954 140614 31574 176058
rect 30954 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 31574 140614
rect 30954 140294 31574 140378
rect 30954 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 31574 140294
rect 30954 104614 31574 140058
rect 30954 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 31574 104614
rect 30954 104294 31574 104378
rect 30954 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 31574 104294
rect 30954 68614 31574 104058
rect 30954 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 31574 68614
rect 30954 68294 31574 68378
rect 30954 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 31574 68294
rect 30954 32614 31574 68058
rect 30954 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 31574 32614
rect 30954 32294 31574 32378
rect 30954 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 31574 32294
rect 12954 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 13574 -6106
rect 12954 -6426 13574 -6342
rect 12954 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 13574 -6426
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 12954 -7654 13574 -6662
rect 30954 -7066 31574 32058
rect 37794 704838 38414 705830
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -1894 38414 -902
rect 41514 691174 42134 706202
rect 41514 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 42134 691174
rect 41514 690854 42134 690938
rect 41514 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 42134 690854
rect 41514 655174 42134 690618
rect 41514 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 42134 655174
rect 41514 654854 42134 654938
rect 41514 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 42134 654854
rect 41514 619174 42134 654618
rect 41514 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 42134 619174
rect 41514 618854 42134 618938
rect 41514 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 42134 618854
rect 41514 583174 42134 618618
rect 41514 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 42134 583174
rect 41514 582854 42134 582938
rect 41514 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 42134 582854
rect 41514 547174 42134 582618
rect 41514 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 42134 547174
rect 41514 546854 42134 546938
rect 41514 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 42134 546854
rect 41514 511174 42134 546618
rect 41514 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 42134 511174
rect 41514 510854 42134 510938
rect 41514 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 42134 510854
rect 41514 475174 42134 510618
rect 41514 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 42134 475174
rect 41514 474854 42134 474938
rect 41514 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 42134 474854
rect 41514 439174 42134 474618
rect 41514 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 42134 439174
rect 41514 438854 42134 438938
rect 41514 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 42134 438854
rect 41514 403174 42134 438618
rect 41514 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 42134 403174
rect 41514 402854 42134 402938
rect 41514 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 42134 402854
rect 41514 367174 42134 402618
rect 41514 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 42134 367174
rect 41514 366854 42134 366938
rect 41514 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 42134 366854
rect 41514 331174 42134 366618
rect 41514 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 42134 331174
rect 41514 330854 42134 330938
rect 41514 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 42134 330854
rect 41514 295174 42134 330618
rect 41514 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 42134 295174
rect 41514 294854 42134 294938
rect 41514 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 42134 294854
rect 41514 259174 42134 294618
rect 41514 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 42134 259174
rect 41514 258854 42134 258938
rect 41514 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 42134 258854
rect 41514 223174 42134 258618
rect 41514 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 42134 223174
rect 41514 222854 42134 222938
rect 41514 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 42134 222854
rect 41514 187174 42134 222618
rect 41514 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 42134 187174
rect 41514 186854 42134 186938
rect 41514 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 42134 186854
rect 41514 151174 42134 186618
rect 41514 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 42134 151174
rect 41514 150854 42134 150938
rect 41514 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 42134 150854
rect 41514 115174 42134 150618
rect 41514 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 42134 115174
rect 41514 114854 42134 114938
rect 41514 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 42134 114854
rect 41514 79174 42134 114618
rect 41514 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 42134 79174
rect 41514 78854 42134 78938
rect 41514 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 42134 78854
rect 41514 43174 42134 78618
rect 41514 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 42134 43174
rect 41514 42854 42134 42938
rect 41514 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 42134 42854
rect 41514 7174 42134 42618
rect 41514 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 42134 7174
rect 41514 6854 42134 6938
rect 41514 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 42134 6854
rect 41514 -2266 42134 6618
rect 41514 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 42134 -2266
rect 41514 -2586 42134 -2502
rect 41514 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 42134 -2586
rect 41514 -3814 42134 -2822
rect 45234 694894 45854 708122
rect 45234 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 45854 694894
rect 45234 694574 45854 694658
rect 45234 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 45854 694574
rect 45234 658894 45854 694338
rect 45234 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 45854 658894
rect 45234 658574 45854 658658
rect 45234 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 45854 658574
rect 45234 622894 45854 658338
rect 45234 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 45854 622894
rect 45234 622574 45854 622658
rect 45234 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 45854 622574
rect 45234 586894 45854 622338
rect 45234 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 45854 586894
rect 45234 586574 45854 586658
rect 45234 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 45854 586574
rect 45234 550894 45854 586338
rect 45234 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 45854 550894
rect 45234 550574 45854 550658
rect 45234 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 45854 550574
rect 45234 514894 45854 550338
rect 45234 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 45854 514894
rect 45234 514574 45854 514658
rect 45234 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 45854 514574
rect 45234 478894 45854 514338
rect 45234 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 45854 478894
rect 45234 478574 45854 478658
rect 45234 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 45854 478574
rect 45234 442894 45854 478338
rect 45234 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 45854 442894
rect 45234 442574 45854 442658
rect 45234 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 45854 442574
rect 45234 406894 45854 442338
rect 45234 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 45854 406894
rect 45234 406574 45854 406658
rect 45234 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 45854 406574
rect 45234 370894 45854 406338
rect 45234 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 45854 370894
rect 45234 370574 45854 370658
rect 45234 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 45854 370574
rect 45234 334894 45854 370338
rect 45234 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 45854 334894
rect 45234 334574 45854 334658
rect 45234 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 45854 334574
rect 45234 298894 45854 334338
rect 45234 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 45854 298894
rect 45234 298574 45854 298658
rect 45234 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 45854 298574
rect 45234 262894 45854 298338
rect 45234 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 45854 262894
rect 45234 262574 45854 262658
rect 45234 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 45854 262574
rect 45234 226894 45854 262338
rect 45234 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 45854 226894
rect 45234 226574 45854 226658
rect 45234 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 45854 226574
rect 45234 190894 45854 226338
rect 45234 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 45854 190894
rect 45234 190574 45854 190658
rect 45234 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 45854 190574
rect 45234 154894 45854 190338
rect 45234 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 45854 154894
rect 45234 154574 45854 154658
rect 45234 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 45854 154574
rect 45234 118894 45854 154338
rect 45234 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 45854 118894
rect 45234 118574 45854 118658
rect 45234 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 45854 118574
rect 45234 82894 45854 118338
rect 45234 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 45854 82894
rect 45234 82574 45854 82658
rect 45234 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 45854 82574
rect 45234 46894 45854 82338
rect 45234 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 45854 46894
rect 45234 46574 45854 46658
rect 45234 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 45854 46574
rect 45234 10894 45854 46338
rect 45234 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 45854 10894
rect 45234 10574 45854 10658
rect 45234 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 45854 10574
rect 45234 -4186 45854 10338
rect 45234 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 45854 -4186
rect 45234 -4506 45854 -4422
rect 45234 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 45854 -4506
rect 45234 -5734 45854 -4742
rect 48954 698614 49574 710042
rect 66954 711558 67574 711590
rect 66954 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 67574 711558
rect 66954 711238 67574 711322
rect 66954 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 67574 711238
rect 63234 709638 63854 709670
rect 63234 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 63854 709638
rect 63234 709318 63854 709402
rect 63234 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 63854 709318
rect 59514 707718 60134 707750
rect 59514 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 60134 707718
rect 59514 707398 60134 707482
rect 59514 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 60134 707398
rect 48954 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 49574 698614
rect 48954 698294 49574 698378
rect 48954 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 49574 698294
rect 48954 662614 49574 698058
rect 48954 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 49574 662614
rect 48954 662294 49574 662378
rect 48954 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 49574 662294
rect 48954 626614 49574 662058
rect 48954 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 49574 626614
rect 48954 626294 49574 626378
rect 48954 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 49574 626294
rect 48954 590614 49574 626058
rect 48954 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 49574 590614
rect 48954 590294 49574 590378
rect 48954 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 49574 590294
rect 48954 554614 49574 590058
rect 48954 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 49574 554614
rect 48954 554294 49574 554378
rect 48954 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 49574 554294
rect 48954 518614 49574 554058
rect 48954 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 49574 518614
rect 48954 518294 49574 518378
rect 48954 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 49574 518294
rect 48954 482614 49574 518058
rect 48954 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 49574 482614
rect 48954 482294 49574 482378
rect 48954 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 49574 482294
rect 48954 446614 49574 482058
rect 48954 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 49574 446614
rect 48954 446294 49574 446378
rect 48954 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 49574 446294
rect 48954 410614 49574 446058
rect 48954 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 49574 410614
rect 48954 410294 49574 410378
rect 48954 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 49574 410294
rect 48954 374614 49574 410058
rect 48954 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 49574 374614
rect 48954 374294 49574 374378
rect 48954 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 49574 374294
rect 48954 338614 49574 374058
rect 48954 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 49574 338614
rect 48954 338294 49574 338378
rect 48954 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 49574 338294
rect 48954 302614 49574 338058
rect 48954 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 49574 302614
rect 48954 302294 49574 302378
rect 48954 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 49574 302294
rect 48954 266614 49574 302058
rect 55794 705798 56414 705830
rect 55794 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 56414 705798
rect 55794 705478 56414 705562
rect 55794 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 56414 705478
rect 55794 669454 56414 705242
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55794 525454 56414 560898
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55794 453454 56414 488898
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55794 417454 56414 452898
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55794 381454 56414 416898
rect 55794 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 56414 381454
rect 55794 381134 56414 381218
rect 55794 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 56414 381134
rect 55794 345454 56414 380898
rect 55794 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 56414 345454
rect 55794 345134 56414 345218
rect 55794 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 56414 345134
rect 55794 309454 56414 344898
rect 55794 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 56414 309454
rect 55794 309134 56414 309218
rect 55794 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 56414 309134
rect 53603 285700 53669 285701
rect 53603 285636 53604 285700
rect 53668 285636 53669 285700
rect 53603 285635 53669 285636
rect 48954 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 49574 266614
rect 48954 266294 49574 266378
rect 48954 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 49574 266294
rect 48954 230614 49574 266058
rect 48954 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 49574 230614
rect 48954 230294 49574 230378
rect 48954 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 49574 230294
rect 48954 194614 49574 230058
rect 48954 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 49574 194614
rect 48954 194294 49574 194378
rect 48954 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 49574 194294
rect 48954 158614 49574 194058
rect 48954 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 49574 158614
rect 48954 158294 49574 158378
rect 48954 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 49574 158294
rect 48954 122614 49574 158058
rect 48954 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 49574 122614
rect 48954 122294 49574 122378
rect 48954 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 49574 122294
rect 48954 86614 49574 122058
rect 48954 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 49574 86614
rect 48954 86294 49574 86378
rect 48954 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 49574 86294
rect 48954 50614 49574 86058
rect 53606 75173 53666 285635
rect 55794 273454 56414 308898
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 55794 237454 56414 272898
rect 55794 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 56414 237454
rect 55794 237134 56414 237218
rect 55794 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 56414 237134
rect 55794 201454 56414 236898
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 55794 165454 56414 200898
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 129454 56414 164898
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 53603 75172 53669 75173
rect 53603 75108 53604 75172
rect 53668 75108 53669 75172
rect 53603 75107 53669 75108
rect 48954 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 49574 50614
rect 48954 50294 49574 50378
rect 48954 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 49574 50294
rect 48954 14614 49574 50058
rect 48954 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 49574 14614
rect 48954 14294 49574 14378
rect 48954 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 49574 14294
rect 30954 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 31574 -7066
rect 30954 -7386 31574 -7302
rect 30954 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 31574 -7386
rect 30954 -7654 31574 -7622
rect 48954 -6106 49574 14058
rect 55794 57454 56414 92898
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55794 21454 56414 56898
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -1306 56414 20898
rect 55794 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 56414 -1306
rect 55794 -1626 56414 -1542
rect 55794 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 56414 -1626
rect 55794 -1894 56414 -1862
rect 59514 673174 60134 707162
rect 59514 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 60134 673174
rect 59514 672854 60134 672938
rect 59514 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 60134 672854
rect 59514 637174 60134 672618
rect 59514 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 60134 637174
rect 59514 636854 60134 636938
rect 59514 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 60134 636854
rect 59514 601174 60134 636618
rect 59514 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 60134 601174
rect 59514 600854 60134 600938
rect 59514 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 60134 600854
rect 59514 565174 60134 600618
rect 59514 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 60134 565174
rect 59514 564854 60134 564938
rect 59514 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 60134 564854
rect 59514 529174 60134 564618
rect 59514 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 60134 529174
rect 59514 528854 60134 528938
rect 59514 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 60134 528854
rect 59514 493174 60134 528618
rect 59514 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 60134 493174
rect 59514 492854 60134 492938
rect 59514 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 60134 492854
rect 59514 457174 60134 492618
rect 59514 456938 59546 457174
rect 59782 456938 59866 457174
rect 60102 456938 60134 457174
rect 59514 456854 60134 456938
rect 59514 456618 59546 456854
rect 59782 456618 59866 456854
rect 60102 456618 60134 456854
rect 59514 421174 60134 456618
rect 59514 420938 59546 421174
rect 59782 420938 59866 421174
rect 60102 420938 60134 421174
rect 59514 420854 60134 420938
rect 59514 420618 59546 420854
rect 59782 420618 59866 420854
rect 60102 420618 60134 420854
rect 59514 385174 60134 420618
rect 59514 384938 59546 385174
rect 59782 384938 59866 385174
rect 60102 384938 60134 385174
rect 59514 384854 60134 384938
rect 59514 384618 59546 384854
rect 59782 384618 59866 384854
rect 60102 384618 60134 384854
rect 59514 349174 60134 384618
rect 59514 348938 59546 349174
rect 59782 348938 59866 349174
rect 60102 348938 60134 349174
rect 59514 348854 60134 348938
rect 59514 348618 59546 348854
rect 59782 348618 59866 348854
rect 60102 348618 60134 348854
rect 59514 313174 60134 348618
rect 63234 676894 63854 709082
rect 63234 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 63854 676894
rect 63234 676574 63854 676658
rect 63234 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 63854 676574
rect 63234 640894 63854 676338
rect 63234 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 63854 640894
rect 63234 640574 63854 640658
rect 63234 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 63854 640574
rect 63234 604894 63854 640338
rect 63234 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 63854 604894
rect 63234 604574 63854 604658
rect 63234 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 63854 604574
rect 63234 568894 63854 604338
rect 66954 680614 67574 711002
rect 84954 710598 85574 711590
rect 84954 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 85574 710598
rect 84954 710278 85574 710362
rect 84954 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 85574 710278
rect 81234 708678 81854 709670
rect 81234 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 81854 708678
rect 81234 708358 81854 708442
rect 81234 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 81854 708358
rect 77514 706758 78134 707750
rect 77514 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 78134 706758
rect 77514 706438 78134 706522
rect 77514 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 78134 706438
rect 73794 704838 74414 705830
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 69611 702540 69677 702541
rect 69611 702476 69612 702540
rect 69676 702476 69677 702540
rect 69611 702475 69677 702476
rect 66954 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 67574 680614
rect 66954 680294 67574 680378
rect 66954 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 67574 680294
rect 66954 644614 67574 680058
rect 66954 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 67574 644614
rect 66954 644294 67574 644378
rect 66954 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 67574 644294
rect 66954 608614 67574 644058
rect 66954 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 67574 608614
rect 66954 608294 67574 608378
rect 66954 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 67574 608294
rect 66954 591166 67574 608058
rect 69614 586530 69674 702475
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73794 591166 74414 614898
rect 77514 691174 78134 706202
rect 77514 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 78134 691174
rect 77514 690854 78134 690938
rect 77514 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 78134 690854
rect 77514 655174 78134 690618
rect 77514 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 78134 655174
rect 77514 654854 78134 654938
rect 77514 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 78134 654854
rect 77514 619174 78134 654618
rect 77514 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 78134 619174
rect 77514 618854 78134 618938
rect 77514 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 78134 618854
rect 77514 591166 78134 618618
rect 81234 694894 81854 708122
rect 81234 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 81854 694894
rect 81234 694574 81854 694658
rect 81234 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 81854 694574
rect 81234 658894 81854 694338
rect 81234 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 81854 658894
rect 81234 658574 81854 658658
rect 81234 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 81854 658574
rect 81234 622894 81854 658338
rect 81234 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 81854 622894
rect 81234 622574 81854 622658
rect 81234 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 81854 622574
rect 81234 591166 81854 622338
rect 84954 698614 85574 710042
rect 102954 711558 103574 711590
rect 102954 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 103574 711558
rect 102954 711238 103574 711322
rect 102954 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 103574 711238
rect 99234 709638 99854 709670
rect 99234 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 99854 709638
rect 99234 709318 99854 709402
rect 99234 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 99854 709318
rect 95514 707718 96134 707750
rect 95514 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 96134 707718
rect 95514 707398 96134 707482
rect 95514 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 96134 707398
rect 84954 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 85574 698614
rect 84954 698294 85574 698378
rect 84954 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 85574 698294
rect 84954 662614 85574 698058
rect 84954 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 85574 662614
rect 84954 662294 85574 662378
rect 84954 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 85574 662294
rect 84954 626614 85574 662058
rect 84954 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 85574 626614
rect 84954 626294 85574 626378
rect 84954 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 85574 626294
rect 84954 591166 85574 626058
rect 91794 705798 92414 705830
rect 91794 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 92414 705798
rect 91794 705478 92414 705562
rect 91794 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 92414 705478
rect 91794 669454 92414 705242
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 633454 92414 668898
rect 91794 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 92414 633454
rect 91794 633134 92414 633218
rect 91794 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 92414 633134
rect 91794 597454 92414 632898
rect 91794 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 92414 597454
rect 91794 597134 92414 597218
rect 91794 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 92414 597134
rect 88011 590748 88077 590749
rect 88011 590684 88012 590748
rect 88076 590684 88077 590748
rect 88011 590683 88077 590684
rect 69430 586470 69674 586530
rect 69430 582317 69490 586470
rect 88014 583130 88074 590683
rect 88195 588572 88261 588573
rect 88195 588508 88196 588572
rect 88260 588508 88261 588572
rect 88195 588507 88261 588508
rect 88198 585717 88258 588507
rect 88195 585716 88261 585717
rect 88195 585652 88196 585716
rect 88260 585652 88261 585716
rect 88195 585651 88261 585652
rect 88014 583070 88258 583130
rect 88198 582861 88258 583070
rect 88195 582860 88261 582861
rect 88195 582796 88196 582860
rect 88260 582796 88261 582860
rect 88195 582795 88261 582796
rect 69427 582316 69493 582317
rect 69427 582252 69428 582316
rect 69492 582252 69493 582316
rect 69427 582251 69493 582252
rect 72679 579454 72999 579486
rect 72679 579218 72721 579454
rect 72957 579218 72999 579454
rect 72679 579134 72999 579218
rect 72679 578898 72721 579134
rect 72957 578898 72999 579134
rect 72679 578866 72999 578898
rect 78609 579454 78929 579486
rect 78609 579218 78651 579454
rect 78887 579218 78929 579454
rect 78609 579134 78929 579218
rect 78609 578898 78651 579134
rect 78887 578898 78929 579134
rect 78609 578866 78929 578898
rect 84540 579454 84860 579486
rect 84540 579218 84582 579454
rect 84818 579218 84860 579454
rect 84540 579134 84860 579218
rect 84540 578898 84582 579134
rect 84818 578898 84860 579134
rect 84540 578866 84860 578898
rect 91507 578100 91573 578101
rect 91507 578036 91508 578100
rect 91572 578036 91573 578100
rect 91507 578035 91573 578036
rect 63234 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 63854 568894
rect 63234 568574 63854 568658
rect 63234 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 63854 568574
rect 63234 532894 63854 568338
rect 75644 561454 75964 561486
rect 75644 561218 75686 561454
rect 75922 561218 75964 561454
rect 75644 561134 75964 561218
rect 75644 560898 75686 561134
rect 75922 560898 75964 561134
rect 75644 560866 75964 560898
rect 81575 561454 81895 561486
rect 81575 561218 81617 561454
rect 81853 561218 81895 561454
rect 81575 561134 81895 561218
rect 81575 560898 81617 561134
rect 81853 560898 81895 561134
rect 81575 560866 81895 560898
rect 67403 556884 67469 556885
rect 67403 556820 67404 556884
rect 67468 556820 67469 556884
rect 67403 556819 67469 556820
rect 66667 551444 66733 551445
rect 66667 551380 66668 551444
rect 66732 551380 66733 551444
rect 66667 551379 66733 551380
rect 63234 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 63854 532894
rect 63234 532574 63854 532658
rect 63234 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 63854 532574
rect 63234 496894 63854 532338
rect 66670 528570 66730 551379
rect 67406 537437 67466 556819
rect 67771 546004 67837 546005
rect 67771 545940 67772 546004
rect 67836 545940 67837 546004
rect 67771 545939 67837 545940
rect 67774 545189 67834 545939
rect 67771 545188 67837 545189
rect 67771 545124 67772 545188
rect 67836 545124 67837 545188
rect 67771 545123 67837 545124
rect 67403 537436 67469 537437
rect 67403 537372 67404 537436
rect 67468 537372 67469 537436
rect 67403 537371 67469 537372
rect 66486 528510 66730 528570
rect 66954 536614 67574 537166
rect 66954 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 67574 536614
rect 66954 536294 67574 536378
rect 66954 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 67574 536294
rect 66486 523837 66546 528510
rect 66483 523836 66549 523837
rect 66483 523772 66484 523836
rect 66548 523772 66549 523836
rect 66483 523771 66549 523772
rect 66667 523700 66733 523701
rect 66667 523636 66668 523700
rect 66732 523636 66733 523700
rect 66667 523635 66733 523636
rect 63234 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 63854 496894
rect 63234 496574 63854 496658
rect 63234 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 63854 496574
rect 63234 460894 63854 496338
rect 63234 460658 63266 460894
rect 63502 460658 63586 460894
rect 63822 460658 63854 460894
rect 63234 460574 63854 460658
rect 63234 460338 63266 460574
rect 63502 460338 63586 460574
rect 63822 460338 63854 460574
rect 63234 424894 63854 460338
rect 63234 424658 63266 424894
rect 63502 424658 63586 424894
rect 63822 424658 63854 424894
rect 63234 424574 63854 424658
rect 63234 424338 63266 424574
rect 63502 424338 63586 424574
rect 63822 424338 63854 424574
rect 63234 388894 63854 424338
rect 66670 419661 66730 523635
rect 66954 500614 67574 536058
rect 67774 535397 67834 545123
rect 72679 543454 72999 543486
rect 72679 543218 72721 543454
rect 72957 543218 72999 543454
rect 72679 543134 72999 543218
rect 72679 542898 72721 543134
rect 72957 542898 72999 543134
rect 72679 542866 72999 542898
rect 78609 543454 78929 543486
rect 78609 543218 78651 543454
rect 78887 543218 78929 543454
rect 78609 543134 78929 543218
rect 78609 542898 78651 543134
rect 78887 542898 78929 543134
rect 78609 542866 78929 542898
rect 84540 543454 84860 543486
rect 84540 543218 84582 543454
rect 84818 543218 84860 543454
rect 84540 543134 84860 543218
rect 84540 542898 84582 543134
rect 84818 542898 84860 543134
rect 84540 542866 84860 542898
rect 69427 542332 69493 542333
rect 69427 542268 69428 542332
rect 69492 542268 69493 542332
rect 69427 542267 69493 542268
rect 69430 538230 69490 542267
rect 69430 538170 69858 538230
rect 68139 535532 68205 535533
rect 68139 535468 68140 535532
rect 68204 535468 68205 535532
rect 68139 535467 68205 535468
rect 69611 535532 69677 535533
rect 69611 535468 69612 535532
rect 69676 535468 69677 535532
rect 69611 535467 69677 535468
rect 67771 535396 67837 535397
rect 67771 535332 67772 535396
rect 67836 535332 67837 535396
rect 67771 535331 67837 535332
rect 66954 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 67574 500614
rect 66954 500294 67574 500378
rect 66954 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 67574 500294
rect 66954 464614 67574 500058
rect 66954 464378 66986 464614
rect 67222 464378 67306 464614
rect 67542 464378 67574 464614
rect 66954 464294 67574 464378
rect 66954 464058 66986 464294
rect 67222 464058 67306 464294
rect 67542 464058 67574 464294
rect 66954 446407 67574 464058
rect 66667 419660 66733 419661
rect 66667 419596 66668 419660
rect 66732 419596 66733 419660
rect 66667 419595 66733 419596
rect 68142 389061 68202 535467
rect 68323 445908 68389 445909
rect 68323 445844 68324 445908
rect 68388 445844 68389 445908
rect 68323 445843 68389 445844
rect 68139 389060 68205 389061
rect 68139 388996 68140 389060
rect 68204 388996 68205 389060
rect 68139 388995 68205 388996
rect 63234 388658 63266 388894
rect 63502 388658 63586 388894
rect 63822 388658 63854 388894
rect 63234 388574 63854 388658
rect 63234 388338 63266 388574
rect 63502 388338 63586 388574
rect 63822 388338 63854 388574
rect 63234 352894 63854 388338
rect 64643 364716 64709 364717
rect 64643 364652 64644 364716
rect 64708 364652 64709 364716
rect 64643 364651 64709 364652
rect 63234 352658 63266 352894
rect 63502 352658 63586 352894
rect 63822 352658 63854 352894
rect 63234 352574 63854 352658
rect 63234 352338 63266 352574
rect 63502 352338 63586 352574
rect 63822 352338 63854 352574
rect 61883 325820 61949 325821
rect 61883 325756 61884 325820
rect 61948 325756 61949 325820
rect 61883 325755 61949 325756
rect 59514 312938 59546 313174
rect 59782 312938 59866 313174
rect 60102 312938 60134 313174
rect 59514 312854 60134 312938
rect 59514 312618 59546 312854
rect 59782 312618 59866 312854
rect 60102 312618 60134 312854
rect 59514 277174 60134 312618
rect 59514 276938 59546 277174
rect 59782 276938 59866 277174
rect 60102 276938 60134 277174
rect 59514 276854 60134 276938
rect 59514 276618 59546 276854
rect 59782 276618 59866 276854
rect 60102 276618 60134 276854
rect 59514 241174 60134 276618
rect 59514 240938 59546 241174
rect 59782 240938 59866 241174
rect 60102 240938 60134 241174
rect 59514 240854 60134 240938
rect 59514 240618 59546 240854
rect 59782 240618 59866 240854
rect 60102 240618 60134 240854
rect 59514 205174 60134 240618
rect 59514 204938 59546 205174
rect 59782 204938 59866 205174
rect 60102 204938 60134 205174
rect 59514 204854 60134 204938
rect 59514 204618 59546 204854
rect 59782 204618 59866 204854
rect 60102 204618 60134 204854
rect 59514 169174 60134 204618
rect 59514 168938 59546 169174
rect 59782 168938 59866 169174
rect 60102 168938 60134 169174
rect 59514 168854 60134 168938
rect 59514 168618 59546 168854
rect 59782 168618 59866 168854
rect 60102 168618 60134 168854
rect 59514 133174 60134 168618
rect 59514 132938 59546 133174
rect 59782 132938 59866 133174
rect 60102 132938 60134 133174
rect 59514 132854 60134 132938
rect 59514 132618 59546 132854
rect 59782 132618 59866 132854
rect 60102 132618 60134 132854
rect 59514 97174 60134 132618
rect 59514 96938 59546 97174
rect 59782 96938 59866 97174
rect 60102 96938 60134 97174
rect 59514 96854 60134 96938
rect 59514 96618 59546 96854
rect 59782 96618 59866 96854
rect 60102 96618 60134 96854
rect 59514 61174 60134 96618
rect 61886 66877 61946 325755
rect 63234 316894 63854 352338
rect 63234 316658 63266 316894
rect 63502 316658 63586 316894
rect 63822 316658 63854 316894
rect 63234 316574 63854 316658
rect 63234 316338 63266 316574
rect 63502 316338 63586 316574
rect 63822 316338 63854 316574
rect 63234 280894 63854 316338
rect 63234 280658 63266 280894
rect 63502 280658 63586 280894
rect 63822 280658 63854 280894
rect 63234 280574 63854 280658
rect 63234 280338 63266 280574
rect 63502 280338 63586 280574
rect 63822 280338 63854 280574
rect 63234 244894 63854 280338
rect 63234 244658 63266 244894
rect 63502 244658 63586 244894
rect 63822 244658 63854 244894
rect 63234 244574 63854 244658
rect 63234 244338 63266 244574
rect 63502 244338 63586 244574
rect 63822 244338 63854 244574
rect 63234 208894 63854 244338
rect 64646 242997 64706 364651
rect 66954 356614 67574 388356
rect 67771 377500 67837 377501
rect 67771 377436 67772 377500
rect 67836 377436 67837 377500
rect 67771 377435 67837 377436
rect 66954 356378 66986 356614
rect 67222 356378 67306 356614
rect 67542 356378 67574 356614
rect 66954 356294 67574 356378
rect 66954 356058 66986 356294
rect 67222 356058 67306 356294
rect 67542 356058 67574 356294
rect 66667 347036 66733 347037
rect 66667 346972 66668 347036
rect 66732 346972 66733 347036
rect 66667 346971 66733 346972
rect 66670 298757 66730 346971
rect 66954 331592 67574 356058
rect 66667 298756 66733 298757
rect 66667 298692 66668 298756
rect 66732 298692 66733 298756
rect 66667 298691 66733 298692
rect 67774 280261 67834 377435
rect 68326 377365 68386 445843
rect 69614 414030 69674 535467
rect 69798 480270 69858 538170
rect 73794 507454 74414 537166
rect 73794 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 74414 507454
rect 73794 507134 74414 507218
rect 73794 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 74414 507134
rect 69798 480210 70226 480270
rect 70166 467941 70226 480210
rect 73794 471454 74414 506898
rect 73794 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 74414 471454
rect 73794 471134 74414 471218
rect 73794 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 74414 471134
rect 70163 467940 70229 467941
rect 70163 467876 70164 467940
rect 70228 467876 70229 467940
rect 70163 467875 70229 467876
rect 70166 447133 70226 467875
rect 71819 462908 71885 462909
rect 71819 462844 71820 462908
rect 71884 462844 71885 462908
rect 71819 462843 71885 462844
rect 70163 447132 70229 447133
rect 70163 447068 70164 447132
rect 70228 447068 70229 447132
rect 70163 447067 70229 447068
rect 71822 445909 71882 462843
rect 72371 446452 72437 446453
rect 72371 446388 72372 446452
rect 72436 446388 72437 446452
rect 73794 446407 74414 470898
rect 77514 511174 78134 537166
rect 77514 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 78134 511174
rect 77514 510854 78134 510938
rect 77514 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 78134 510854
rect 77514 475174 78134 510618
rect 77514 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 78134 475174
rect 77514 474854 78134 474938
rect 77514 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 78134 474854
rect 77514 446407 78134 474618
rect 81234 514894 81854 537166
rect 81234 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 81854 514894
rect 81234 514574 81854 514658
rect 81234 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 81854 514574
rect 81234 478894 81854 514338
rect 81234 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 81854 478894
rect 81234 478574 81854 478658
rect 81234 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 81854 478574
rect 81234 446407 81854 478338
rect 84954 518614 85574 537166
rect 84954 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 85574 518614
rect 84954 518294 85574 518378
rect 84954 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 85574 518294
rect 84954 482614 85574 518058
rect 84954 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 85574 482614
rect 84954 482294 85574 482378
rect 84954 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 85574 482294
rect 84954 446407 85574 482058
rect 89667 460188 89733 460189
rect 89667 460124 89668 460188
rect 89732 460124 89733 460188
rect 89667 460123 89733 460124
rect 72371 446387 72437 446388
rect 71819 445908 71885 445909
rect 71819 445844 71820 445908
rect 71884 445844 71885 445908
rect 71819 445843 71885 445844
rect 69062 413970 69674 414030
rect 69062 404370 69122 413970
rect 69243 407828 69309 407829
rect 69243 407764 69244 407828
rect 69308 407826 69309 407828
rect 69308 407766 69490 407826
rect 69308 407764 69309 407766
rect 69243 407763 69309 407764
rect 69246 407149 69306 407763
rect 69243 407148 69309 407149
rect 69243 407084 69244 407148
rect 69308 407084 69309 407148
rect 69243 407083 69309 407084
rect 69430 404370 69490 407766
rect 69062 404310 69306 404370
rect 69430 404310 69858 404370
rect 69246 396130 69306 404310
rect 69798 404290 69858 404310
rect 69798 404230 70042 404290
rect 69982 396130 70042 404230
rect 69246 396070 69674 396130
rect 69614 390421 69674 396070
rect 69798 396070 70042 396130
rect 69611 390420 69677 390421
rect 69611 390356 69612 390420
rect 69676 390356 69677 390420
rect 69611 390355 69677 390356
rect 68323 377364 68389 377365
rect 68323 377300 68324 377364
rect 68388 377300 68389 377364
rect 68323 377299 68389 377300
rect 69798 370565 69858 396070
rect 72374 391917 72434 446387
rect 72739 445908 72805 445909
rect 72739 445844 72740 445908
rect 72804 445844 72805 445908
rect 72739 445843 72805 445844
rect 72371 391916 72437 391917
rect 72371 391852 72372 391916
rect 72436 391852 72437 391916
rect 72371 391851 72437 391852
rect 70899 389332 70965 389333
rect 70899 389268 70900 389332
rect 70964 389268 70965 389332
rect 70899 389267 70965 389268
rect 69795 370564 69861 370565
rect 69795 370500 69796 370564
rect 69860 370500 69861 370564
rect 69795 370499 69861 370500
rect 69611 368524 69677 368525
rect 69611 368460 69612 368524
rect 69676 368460 69677 368524
rect 69611 368459 69677 368460
rect 68875 348532 68941 348533
rect 68875 348468 68876 348532
rect 68940 348468 68941 348532
rect 68875 348467 68941 348468
rect 68878 339421 68938 348467
rect 67955 339420 68021 339421
rect 67955 339356 67956 339420
rect 68020 339356 68021 339420
rect 67955 339355 68021 339356
rect 68875 339420 68941 339421
rect 68875 339356 68876 339420
rect 68940 339356 68941 339420
rect 68875 339355 68941 339356
rect 67958 338333 68018 339355
rect 67955 338332 68021 338333
rect 67955 338268 67956 338332
rect 68020 338268 68021 338332
rect 67955 338267 68021 338268
rect 67771 280260 67837 280261
rect 67771 280196 67772 280260
rect 67836 280196 67837 280260
rect 67771 280195 67837 280196
rect 66851 276180 66917 276181
rect 66851 276116 66852 276180
rect 66916 276116 66917 276180
rect 66851 276115 66917 276116
rect 66854 268429 66914 276115
rect 67958 269653 68018 338267
rect 69427 329220 69493 329221
rect 69427 329156 69428 329220
rect 69492 329156 69493 329220
rect 69427 329155 69493 329156
rect 69430 328405 69490 329155
rect 69427 328404 69493 328405
rect 69427 328340 69428 328404
rect 69492 328340 69493 328404
rect 69427 328339 69493 328340
rect 69614 325710 69674 368459
rect 69795 335476 69861 335477
rect 69795 335412 69796 335476
rect 69860 335412 69861 335476
rect 69795 335411 69861 335412
rect 69430 325650 69674 325710
rect 69430 325549 69490 325650
rect 69427 325548 69493 325549
rect 69427 325484 69428 325548
rect 69492 325484 69493 325548
rect 69427 325483 69493 325484
rect 69427 324052 69493 324053
rect 69427 323988 69428 324052
rect 69492 324050 69493 324052
rect 69798 324050 69858 335411
rect 69492 323990 69858 324050
rect 69492 323988 69493 323990
rect 69427 323987 69493 323988
rect 67955 269652 68021 269653
rect 67955 269588 67956 269652
rect 68020 269588 68021 269652
rect 67955 269587 68021 269588
rect 66851 268428 66917 268429
rect 66851 268364 66852 268428
rect 66916 268364 66917 268428
rect 66851 268363 66917 268364
rect 67403 267476 67469 267477
rect 67403 267412 67404 267476
rect 67468 267412 67469 267476
rect 67403 267411 67469 267412
rect 65379 257956 65445 257957
rect 65379 257892 65380 257956
rect 65444 257892 65445 257956
rect 65379 257891 65445 257892
rect 64643 242996 64709 242997
rect 64643 242932 64644 242996
rect 64708 242932 64709 242996
rect 64643 242931 64709 242932
rect 63234 208658 63266 208894
rect 63502 208658 63586 208894
rect 63822 208658 63854 208894
rect 63234 208574 63854 208658
rect 63234 208338 63266 208574
rect 63502 208338 63586 208574
rect 63822 208338 63854 208574
rect 63234 172894 63854 208338
rect 63234 172658 63266 172894
rect 63502 172658 63586 172894
rect 63822 172658 63854 172894
rect 63234 172574 63854 172658
rect 63234 172338 63266 172574
rect 63502 172338 63586 172574
rect 63822 172338 63854 172574
rect 63234 136894 63854 172338
rect 63234 136658 63266 136894
rect 63502 136658 63586 136894
rect 63822 136658 63854 136894
rect 63234 136574 63854 136658
rect 63234 136338 63266 136574
rect 63502 136338 63586 136574
rect 63822 136338 63854 136574
rect 63234 100894 63854 136338
rect 63234 100658 63266 100894
rect 63502 100658 63586 100894
rect 63822 100658 63854 100894
rect 63234 100574 63854 100658
rect 63234 100338 63266 100574
rect 63502 100338 63586 100574
rect 63822 100338 63854 100574
rect 61883 66876 61949 66877
rect 61883 66812 61884 66876
rect 61948 66812 61949 66876
rect 61883 66811 61949 66812
rect 59514 60938 59546 61174
rect 59782 60938 59866 61174
rect 60102 60938 60134 61174
rect 59514 60854 60134 60938
rect 59514 60618 59546 60854
rect 59782 60618 59866 60854
rect 60102 60618 60134 60854
rect 59514 25174 60134 60618
rect 59514 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 60134 25174
rect 59514 24854 60134 24938
rect 59514 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 60134 24854
rect 59514 -3226 60134 24618
rect 59514 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 60134 -3226
rect 59514 -3546 60134 -3462
rect 59514 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 60134 -3546
rect 59514 -3814 60134 -3782
rect 63234 64894 63854 100338
rect 63234 64658 63266 64894
rect 63502 64658 63586 64894
rect 63822 64658 63854 64894
rect 63234 64574 63854 64658
rect 63234 64338 63266 64574
rect 63502 64338 63586 64574
rect 63822 64338 63854 64574
rect 63234 28894 63854 64338
rect 65382 37909 65442 257891
rect 66667 252244 66733 252245
rect 66667 252180 66668 252244
rect 66732 252180 66733 252244
rect 66667 252179 66733 252180
rect 66670 213213 66730 252179
rect 67406 242861 67466 267411
rect 69427 257140 69493 257141
rect 69427 257076 69428 257140
rect 69492 257076 69493 257140
rect 69427 257075 69493 257076
rect 67955 254420 68021 254421
rect 67955 254356 67956 254420
rect 68020 254356 68021 254420
rect 67955 254355 68021 254356
rect 67771 248980 67837 248981
rect 67771 248916 67772 248980
rect 67836 248916 67837 248980
rect 67771 248915 67837 248916
rect 67403 242860 67469 242861
rect 67403 242796 67404 242860
rect 67468 242796 67469 242860
rect 67403 242795 67469 242796
rect 66667 213212 66733 213213
rect 66667 213148 66668 213212
rect 66732 213148 66733 213212
rect 66667 213147 66733 213148
rect 66954 212614 67574 239592
rect 66954 212378 66986 212614
rect 67222 212378 67306 212614
rect 67542 212378 67574 212614
rect 66954 212294 67574 212378
rect 66954 212058 66986 212294
rect 67222 212058 67306 212294
rect 67542 212058 67574 212294
rect 66954 176600 67574 212058
rect 66954 68614 67574 93100
rect 66954 68378 66986 68614
rect 67222 68378 67306 68614
rect 67542 68378 67574 68614
rect 66954 68294 67574 68378
rect 66954 68058 66986 68294
rect 67222 68058 67306 68294
rect 67542 68058 67574 68294
rect 65379 37908 65445 37909
rect 65379 37844 65380 37908
rect 65444 37844 65445 37908
rect 65379 37843 65445 37844
rect 63234 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 63854 28894
rect 63234 28574 63854 28658
rect 63234 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 63854 28574
rect 63234 -5146 63854 28338
rect 63234 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 63854 -5146
rect 63234 -5466 63854 -5382
rect 63234 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 63854 -5466
rect 63234 -5734 63854 -5702
rect 66954 32614 67574 68058
rect 67774 33965 67834 248915
rect 67958 201381 68018 254355
rect 69430 248430 69490 257075
rect 69430 248370 69674 248430
rect 69614 225725 69674 248370
rect 70902 228853 70962 389267
rect 71083 361860 71149 361861
rect 71083 361796 71084 361860
rect 71148 361796 71149 361860
rect 71083 361795 71149 361796
rect 71086 329221 71146 361795
rect 72742 349077 72802 445843
rect 72978 435454 73298 435486
rect 72978 435218 73020 435454
rect 73256 435218 73298 435454
rect 72978 435134 73298 435218
rect 72978 434898 73020 435134
rect 73256 434898 73298 435134
rect 72978 434866 73298 434898
rect 88338 417454 88658 417486
rect 88338 417218 88380 417454
rect 88616 417218 88658 417454
rect 88338 417134 88658 417218
rect 88338 416898 88380 417134
rect 88616 416898 88658 417134
rect 88338 416866 88658 416898
rect 72978 399454 73298 399486
rect 72978 399218 73020 399454
rect 73256 399218 73298 399454
rect 72978 399134 73298 399218
rect 72978 398898 73020 399134
rect 73256 398898 73298 399134
rect 72978 398866 73298 398898
rect 73107 391916 73173 391917
rect 73107 391852 73108 391916
rect 73172 391852 73173 391916
rect 73107 391851 73173 391852
rect 73110 389061 73170 391851
rect 89670 390421 89730 460123
rect 90219 456244 90285 456245
rect 90219 456180 90220 456244
rect 90284 456180 90285 456244
rect 90219 456179 90285 456180
rect 89667 390420 89733 390421
rect 89667 390356 89668 390420
rect 89732 390356 89733 390420
rect 89667 390355 89733 390356
rect 90222 389061 90282 456179
rect 91510 450533 91570 578035
rect 91794 561454 92414 596898
rect 95514 673174 96134 707162
rect 95514 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 96134 673174
rect 95514 672854 96134 672938
rect 95514 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 96134 672854
rect 95514 637174 96134 672618
rect 95514 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 96134 637174
rect 95514 636854 96134 636938
rect 95514 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 96134 636854
rect 95514 601174 96134 636618
rect 95514 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 96134 601174
rect 95514 600854 96134 600938
rect 95514 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 96134 600854
rect 93899 588708 93965 588709
rect 93899 588644 93900 588708
rect 93964 588644 93965 588708
rect 93899 588643 93965 588644
rect 91794 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 92414 561454
rect 91794 561134 92414 561218
rect 91794 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 92414 561134
rect 91794 525454 92414 560898
rect 91794 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 92414 525454
rect 91794 525134 92414 525218
rect 91794 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 92414 525134
rect 91794 489454 92414 524898
rect 91794 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 92414 489454
rect 91794 489134 92414 489218
rect 91794 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 92414 489134
rect 91794 453454 92414 488898
rect 92979 462908 93045 462909
rect 92979 462844 92980 462908
rect 93044 462844 93045 462908
rect 92979 462843 93045 462844
rect 91794 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 92414 453454
rect 91794 453134 92414 453218
rect 91794 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 92414 453134
rect 91507 450532 91573 450533
rect 91507 450468 91508 450532
rect 91572 450468 91573 450532
rect 91507 450467 91573 450468
rect 91507 447268 91573 447269
rect 91507 447204 91508 447268
rect 91572 447204 91573 447268
rect 91507 447203 91573 447204
rect 73107 389060 73173 389061
rect 73107 388996 73108 389060
rect 73172 388996 73173 389060
rect 73107 388995 73173 388996
rect 90219 389060 90285 389061
rect 90219 388996 90220 389060
rect 90284 388996 90285 389060
rect 90219 388995 90285 388996
rect 91510 388925 91570 447203
rect 91794 446407 92414 452898
rect 92982 391101 93042 462843
rect 93902 445773 93962 588643
rect 95514 565174 96134 600618
rect 95514 564938 95546 565174
rect 95782 564938 95866 565174
rect 96102 564938 96134 565174
rect 95514 564854 96134 564938
rect 95514 564618 95546 564854
rect 95782 564618 95866 564854
rect 96102 564618 96134 564854
rect 95514 529174 96134 564618
rect 95514 528938 95546 529174
rect 95782 528938 95866 529174
rect 96102 528938 96134 529174
rect 95514 528854 96134 528938
rect 95514 528618 95546 528854
rect 95782 528618 95866 528854
rect 96102 528618 96134 528854
rect 95514 493174 96134 528618
rect 95514 492938 95546 493174
rect 95782 492938 95866 493174
rect 96102 492938 96134 493174
rect 95514 492854 96134 492938
rect 95514 492618 95546 492854
rect 95782 492618 95866 492854
rect 96102 492618 96134 492854
rect 94083 459644 94149 459645
rect 94083 459580 94084 459644
rect 94148 459580 94149 459644
rect 94083 459579 94149 459580
rect 93899 445772 93965 445773
rect 93899 445708 93900 445772
rect 93964 445708 93965 445772
rect 93899 445707 93965 445708
rect 92979 391100 93045 391101
rect 92979 391036 92980 391100
rect 93044 391036 93045 391100
rect 92979 391035 93045 391036
rect 91507 388924 91573 388925
rect 91507 388860 91508 388924
rect 91572 388860 91573 388924
rect 91507 388859 91573 388860
rect 73794 363454 74414 388356
rect 73794 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 74414 363454
rect 73794 363134 74414 363218
rect 73794 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 74414 363134
rect 72739 349076 72805 349077
rect 72739 349012 72740 349076
rect 72804 349012 72805 349076
rect 72739 349011 72805 349012
rect 73475 340100 73541 340101
rect 73475 340036 73476 340100
rect 73540 340036 73541 340100
rect 73475 340035 73541 340036
rect 71083 329220 71149 329221
rect 71083 329156 71084 329220
rect 71148 329156 71149 329220
rect 71083 329155 71149 329156
rect 72978 291454 73298 291486
rect 72978 291218 73020 291454
rect 73256 291218 73298 291454
rect 72978 291134 73298 291218
rect 72978 290898 73020 291134
rect 73256 290898 73298 291134
rect 72978 290866 73298 290898
rect 72978 255454 73298 255486
rect 72978 255218 73020 255454
rect 73256 255218 73298 255454
rect 72978 255134 73298 255218
rect 72978 254898 73020 255134
rect 73256 254898 73298 255134
rect 72978 254866 73298 254898
rect 73478 236741 73538 340035
rect 73794 331592 74414 362898
rect 77514 367174 78134 388356
rect 77514 366938 77546 367174
rect 77782 366938 77866 367174
rect 78102 366938 78134 367174
rect 77514 366854 78134 366938
rect 77514 366618 77546 366854
rect 77782 366618 77866 366854
rect 78102 366618 78134 366854
rect 77514 331592 78134 366618
rect 81234 370894 81854 388356
rect 81234 370658 81266 370894
rect 81502 370658 81586 370894
rect 81822 370658 81854 370894
rect 81234 370574 81854 370658
rect 81234 370338 81266 370574
rect 81502 370338 81586 370574
rect 81822 370338 81854 370574
rect 78443 341460 78509 341461
rect 78443 341396 78444 341460
rect 78508 341396 78509 341460
rect 78443 341395 78509 341396
rect 75683 331260 75749 331261
rect 75683 331196 75684 331260
rect 75748 331196 75749 331260
rect 75683 331195 75749 331196
rect 73475 236740 73541 236741
rect 73475 236676 73476 236740
rect 73540 236676 73541 236740
rect 73475 236675 73541 236676
rect 70899 228852 70965 228853
rect 70899 228788 70900 228852
rect 70964 228788 70965 228852
rect 70899 228787 70965 228788
rect 69611 225724 69677 225725
rect 69611 225660 69612 225724
rect 69676 225660 69677 225724
rect 69611 225659 69677 225660
rect 73794 219454 74414 239592
rect 75686 220149 75746 331195
rect 77155 329220 77221 329221
rect 77155 329156 77156 329220
rect 77220 329156 77221 329220
rect 77155 329155 77221 329156
rect 75683 220148 75749 220149
rect 75683 220084 75684 220148
rect 75748 220084 75749 220148
rect 75683 220083 75749 220084
rect 73794 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 74414 219454
rect 73794 219134 74414 219218
rect 73794 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 74414 219134
rect 67955 201380 68021 201381
rect 67955 201316 67956 201380
rect 68020 201316 68021 201380
rect 67955 201315 68021 201316
rect 73794 183454 74414 218898
rect 77158 188325 77218 329155
rect 77514 223174 78134 239592
rect 78446 237285 78506 341395
rect 81019 336020 81085 336021
rect 81019 335956 81020 336020
rect 81084 335956 81085 336020
rect 81019 335955 81085 335956
rect 81022 242045 81082 335955
rect 81234 334894 81854 370338
rect 84954 374614 85574 388356
rect 84954 374378 84986 374614
rect 85222 374378 85306 374614
rect 85542 374378 85574 374614
rect 84954 374294 85574 374378
rect 84954 374058 84986 374294
rect 85222 374058 85306 374294
rect 85542 374058 85574 374294
rect 84954 338614 85574 374058
rect 84954 338378 84986 338614
rect 85222 338378 85306 338614
rect 85542 338378 85574 338614
rect 84954 338294 85574 338378
rect 84954 338058 84986 338294
rect 85222 338058 85306 338294
rect 85542 338058 85574 338294
rect 83963 337516 84029 337517
rect 83963 337452 83964 337516
rect 84028 337452 84029 337516
rect 83963 337451 84029 337452
rect 81234 334658 81266 334894
rect 81502 334658 81586 334894
rect 81822 334658 81854 334894
rect 81234 334574 81854 334658
rect 81234 334338 81266 334574
rect 81502 334338 81586 334574
rect 81822 334338 81854 334574
rect 81234 331592 81854 334338
rect 82675 329220 82741 329221
rect 82675 329156 82676 329220
rect 82740 329156 82741 329220
rect 82675 329155 82741 329156
rect 81019 242044 81085 242045
rect 81019 241980 81020 242044
rect 81084 241980 81085 242044
rect 81019 241979 81085 241980
rect 78443 237284 78509 237285
rect 78443 237220 78444 237284
rect 78508 237220 78509 237284
rect 78443 237219 78509 237220
rect 77514 222938 77546 223174
rect 77782 222938 77866 223174
rect 78102 222938 78134 223174
rect 77514 222854 78134 222938
rect 77514 222618 77546 222854
rect 77782 222618 77866 222854
rect 78102 222618 78134 222854
rect 77155 188324 77221 188325
rect 77155 188260 77156 188324
rect 77220 188260 77221 188324
rect 77155 188259 77221 188260
rect 73794 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 74414 183454
rect 73794 183134 74414 183218
rect 73794 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 74414 183134
rect 73794 176600 74414 182898
rect 77514 187174 78134 222618
rect 77514 186938 77546 187174
rect 77782 186938 77866 187174
rect 78102 186938 78134 187174
rect 77514 186854 78134 186938
rect 77514 186618 77546 186854
rect 77782 186618 77866 186854
rect 78102 186618 78134 186854
rect 77514 176600 78134 186618
rect 81234 226894 81854 239592
rect 82678 227629 82738 329155
rect 83966 237285 84026 337451
rect 84954 331592 85574 338058
rect 91794 381454 92414 388356
rect 91794 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 92414 381454
rect 91794 381134 92414 381218
rect 91794 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 92414 381134
rect 91794 345454 92414 380898
rect 91794 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 92414 345454
rect 91794 345134 92414 345218
rect 91794 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 92414 345134
rect 91794 331592 92414 344898
rect 93902 330173 93962 445707
rect 94086 390421 94146 459579
rect 95514 457174 96134 492618
rect 99234 676894 99854 709082
rect 99234 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 99854 676894
rect 99234 676574 99854 676658
rect 99234 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 99854 676574
rect 99234 640894 99854 676338
rect 99234 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 99854 640894
rect 99234 640574 99854 640658
rect 99234 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 99854 640574
rect 99234 604894 99854 640338
rect 99234 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 99854 604894
rect 99234 604574 99854 604658
rect 99234 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 99854 604574
rect 99234 568894 99854 604338
rect 99234 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 99854 568894
rect 99234 568574 99854 568658
rect 99234 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 99854 568574
rect 99234 532894 99854 568338
rect 99234 532658 99266 532894
rect 99502 532658 99586 532894
rect 99822 532658 99854 532894
rect 99234 532574 99854 532658
rect 99234 532338 99266 532574
rect 99502 532338 99586 532574
rect 99822 532338 99854 532574
rect 99234 496894 99854 532338
rect 99234 496658 99266 496894
rect 99502 496658 99586 496894
rect 99822 496658 99854 496894
rect 99234 496574 99854 496658
rect 99234 496338 99266 496574
rect 99502 496338 99586 496574
rect 99822 496338 99854 496574
rect 99234 460894 99854 496338
rect 102954 680614 103574 711002
rect 120954 710598 121574 711590
rect 120954 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 121574 710598
rect 120954 710278 121574 710362
rect 120954 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 121574 710278
rect 117234 708678 117854 709670
rect 117234 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 117854 708678
rect 117234 708358 117854 708442
rect 117234 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 117854 708358
rect 113514 706758 114134 707750
rect 113514 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 114134 706758
rect 113514 706438 114134 706522
rect 113514 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 114134 706438
rect 102954 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 103574 680614
rect 102954 680294 103574 680378
rect 102954 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 103574 680294
rect 102954 644614 103574 680058
rect 102954 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 103574 644614
rect 102954 644294 103574 644378
rect 102954 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 103574 644294
rect 102954 608614 103574 644058
rect 102954 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 103574 608614
rect 102954 608294 103574 608378
rect 102954 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 103574 608294
rect 102954 572614 103574 608058
rect 102954 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 103574 572614
rect 102954 572294 103574 572378
rect 102954 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 103574 572294
rect 102954 536614 103574 572058
rect 102954 536378 102986 536614
rect 103222 536378 103306 536614
rect 103542 536378 103574 536614
rect 102954 536294 103574 536378
rect 102954 536058 102986 536294
rect 103222 536058 103306 536294
rect 103542 536058 103574 536294
rect 102954 500614 103574 536058
rect 109794 704838 110414 705830
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 615454 110414 650898
rect 109794 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 110414 615454
rect 109794 615134 110414 615218
rect 109794 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 110414 615134
rect 109794 579454 110414 614898
rect 109794 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 110414 579454
rect 109794 579134 110414 579218
rect 109794 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 110414 579134
rect 109794 543454 110414 578898
rect 109794 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 110414 543454
rect 109794 543134 110414 543218
rect 109794 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 110414 543134
rect 106411 534716 106477 534717
rect 106411 534652 106412 534716
rect 106476 534652 106477 534716
rect 106411 534651 106477 534652
rect 102954 500378 102986 500614
rect 103222 500378 103306 500614
rect 103542 500378 103574 500614
rect 102954 500294 103574 500378
rect 102954 500058 102986 500294
rect 103222 500058 103306 500294
rect 103542 500058 103574 500294
rect 102954 464614 103574 500058
rect 104939 470660 105005 470661
rect 104939 470596 104940 470660
rect 105004 470596 105005 470660
rect 104939 470595 105005 470596
rect 102179 464404 102245 464405
rect 102179 464340 102180 464404
rect 102244 464340 102245 464404
rect 102179 464339 102245 464340
rect 102954 464378 102986 464614
rect 103222 464378 103306 464614
rect 103542 464378 103574 464614
rect 99234 460658 99266 460894
rect 99502 460658 99586 460894
rect 99822 460658 99854 460894
rect 99234 460574 99854 460658
rect 99234 460338 99266 460574
rect 99502 460338 99586 460574
rect 99822 460338 99854 460574
rect 96659 457468 96725 457469
rect 96659 457404 96660 457468
rect 96724 457404 96725 457468
rect 96659 457403 96725 457404
rect 95514 456938 95546 457174
rect 95782 456938 95866 457174
rect 96102 456938 96134 457174
rect 95514 456854 96134 456938
rect 95514 456618 95546 456854
rect 95782 456618 95866 456854
rect 96102 456618 96134 456854
rect 95514 446407 96134 456618
rect 96291 445772 96357 445773
rect 96291 445708 96292 445772
rect 96356 445708 96357 445772
rect 96291 445707 96357 445708
rect 94083 390420 94149 390421
rect 94083 390356 94084 390420
rect 94148 390356 94149 390420
rect 94083 390355 94149 390356
rect 95514 385174 96134 388356
rect 95514 384938 95546 385174
rect 95782 384938 95866 385174
rect 96102 384938 96134 385174
rect 95514 384854 96134 384938
rect 95514 384618 95546 384854
rect 95782 384618 95866 384854
rect 96102 384618 96134 384854
rect 95514 349174 96134 384618
rect 96294 373421 96354 445707
rect 96662 390421 96722 457403
rect 98131 454748 98197 454749
rect 98131 454684 98132 454748
rect 98196 454684 98197 454748
rect 98131 454683 98197 454684
rect 98134 390421 98194 454683
rect 99234 446407 99854 460338
rect 100707 456108 100773 456109
rect 100707 456044 100708 456108
rect 100772 456044 100773 456108
rect 100707 456043 100773 456044
rect 100523 445772 100589 445773
rect 100523 445708 100524 445772
rect 100588 445708 100589 445772
rect 100523 445707 100589 445708
rect 96659 390420 96725 390421
rect 96659 390356 96660 390420
rect 96724 390356 96725 390420
rect 96659 390355 96725 390356
rect 98131 390420 98197 390421
rect 98131 390356 98132 390420
rect 98196 390356 98197 390420
rect 98131 390355 98197 390356
rect 96291 373420 96357 373421
rect 96291 373356 96292 373420
rect 96356 373356 96357 373420
rect 96291 373355 96357 373356
rect 95514 348938 95546 349174
rect 95782 348938 95866 349174
rect 96102 348938 96134 349174
rect 95514 348854 96134 348938
rect 95514 348618 95546 348854
rect 95782 348618 95866 348854
rect 96102 348618 96134 348854
rect 95514 331592 96134 348618
rect 99234 352894 99854 388356
rect 100526 370021 100586 445707
rect 100710 390285 100770 456043
rect 102182 390421 102242 464339
rect 102954 464294 103574 464378
rect 102954 464058 102986 464294
rect 103222 464058 103306 464294
rect 103542 464058 103574 464294
rect 102954 446407 103574 464058
rect 103698 435454 104018 435486
rect 103698 435218 103740 435454
rect 103976 435218 104018 435454
rect 103698 435134 104018 435218
rect 103698 434898 103740 435134
rect 103976 434898 104018 435134
rect 103698 434866 104018 434898
rect 103698 399454 104018 399486
rect 103698 399218 103740 399454
rect 103976 399218 104018 399454
rect 103698 399134 104018 399218
rect 103698 398898 103740 399134
rect 103976 398898 104018 399134
rect 103698 398866 104018 398898
rect 104942 390421 105002 470595
rect 106414 390421 106474 534651
rect 109794 507454 110414 542898
rect 109794 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 110414 507454
rect 109794 507134 110414 507218
rect 109794 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 110414 507134
rect 109794 471454 110414 506898
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 107699 467124 107765 467125
rect 107699 467060 107700 467124
rect 107764 467060 107765 467124
rect 107699 467059 107765 467060
rect 107702 390421 107762 467059
rect 108987 457468 109053 457469
rect 108987 457404 108988 457468
rect 109052 457404 109053 457468
rect 108987 457403 109053 457404
rect 108803 444684 108869 444685
rect 108803 444620 108804 444684
rect 108868 444620 108869 444684
rect 108803 444619 108869 444620
rect 102179 390420 102245 390421
rect 102179 390356 102180 390420
rect 102244 390356 102245 390420
rect 102179 390355 102245 390356
rect 104939 390420 105005 390421
rect 104939 390356 104940 390420
rect 105004 390356 105005 390420
rect 104939 390355 105005 390356
rect 106411 390420 106477 390421
rect 106411 390356 106412 390420
rect 106476 390356 106477 390420
rect 106411 390355 106477 390356
rect 107699 390420 107765 390421
rect 107699 390356 107700 390420
rect 107764 390356 107765 390420
rect 107699 390355 107765 390356
rect 100707 390284 100773 390285
rect 100707 390220 100708 390284
rect 100772 390220 100773 390284
rect 100707 390219 100773 390220
rect 100523 370020 100589 370021
rect 100523 369956 100524 370020
rect 100588 369956 100589 370020
rect 100523 369955 100589 369956
rect 99234 352658 99266 352894
rect 99502 352658 99586 352894
rect 99822 352658 99854 352894
rect 99234 352574 99854 352658
rect 99234 352338 99266 352574
rect 99502 352338 99586 352574
rect 99822 352338 99854 352574
rect 99234 331592 99854 352338
rect 102954 356614 103574 388356
rect 102954 356378 102986 356614
rect 103222 356378 103306 356614
rect 103542 356378 103574 356614
rect 102954 356294 103574 356378
rect 102954 356058 102986 356294
rect 103222 356058 103306 356294
rect 103542 356058 103574 356294
rect 102954 331592 103574 356058
rect 108806 349213 108866 444619
rect 108990 390421 109050 457403
rect 109794 446407 110414 470898
rect 113514 691174 114134 706202
rect 113514 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 114134 691174
rect 113514 690854 114134 690938
rect 113514 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 114134 690854
rect 113514 655174 114134 690618
rect 113514 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 114134 655174
rect 113514 654854 114134 654938
rect 113514 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 114134 654854
rect 113514 619174 114134 654618
rect 113514 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 114134 619174
rect 113514 618854 114134 618938
rect 113514 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 114134 618854
rect 113514 583174 114134 618618
rect 113514 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 114134 583174
rect 113514 582854 114134 582938
rect 113514 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 114134 582854
rect 113514 547174 114134 582618
rect 113514 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 114134 547174
rect 113514 546854 114134 546938
rect 113514 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 114134 546854
rect 113514 511174 114134 546618
rect 113514 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 114134 511174
rect 113514 510854 114134 510938
rect 113514 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 114134 510854
rect 113514 475174 114134 510618
rect 113514 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 114134 475174
rect 113514 474854 114134 474938
rect 113514 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 114134 474854
rect 113219 467804 113285 467805
rect 113219 467740 113220 467804
rect 113284 467740 113285 467804
rect 113219 467739 113285 467740
rect 111747 460188 111813 460189
rect 111747 460124 111748 460188
rect 111812 460124 111813 460188
rect 111747 460123 111813 460124
rect 111563 444684 111629 444685
rect 111563 444620 111564 444684
rect 111628 444620 111629 444684
rect 111563 444619 111629 444620
rect 108987 390420 109053 390421
rect 108987 390356 108988 390420
rect 109052 390356 109053 390420
rect 108987 390355 109053 390356
rect 109794 363454 110414 388356
rect 111566 381037 111626 444619
rect 111750 389061 111810 460123
rect 113222 389061 113282 467739
rect 113514 446407 114134 474618
rect 117234 694894 117854 708122
rect 117234 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 117854 694894
rect 117234 694574 117854 694658
rect 117234 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 117854 694574
rect 117234 658894 117854 694338
rect 117234 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 117854 658894
rect 117234 658574 117854 658658
rect 117234 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 117854 658574
rect 117234 622894 117854 658338
rect 117234 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 117854 622894
rect 117234 622574 117854 622658
rect 117234 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 117854 622574
rect 117234 586894 117854 622338
rect 117234 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 117854 586894
rect 117234 586574 117854 586658
rect 117234 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 117854 586574
rect 117234 550894 117854 586338
rect 117234 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 117854 550894
rect 117234 550574 117854 550658
rect 117234 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 117854 550574
rect 117234 514894 117854 550338
rect 117234 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 117854 514894
rect 117234 514574 117854 514658
rect 117234 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 117854 514574
rect 117234 478894 117854 514338
rect 117234 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 117854 478894
rect 117234 478574 117854 478658
rect 117234 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 117854 478574
rect 115979 474060 116045 474061
rect 115979 473996 115980 474060
rect 116044 473996 116045 474060
rect 115979 473995 116045 473996
rect 115795 447268 115861 447269
rect 115795 447204 115796 447268
rect 115860 447204 115861 447268
rect 115795 447203 115861 447204
rect 114323 445772 114389 445773
rect 114323 445708 114324 445772
rect 114388 445708 114389 445772
rect 114323 445707 114389 445708
rect 111747 389060 111813 389061
rect 111747 388996 111748 389060
rect 111812 388996 111813 389060
rect 111747 388995 111813 388996
rect 113219 389060 113285 389061
rect 113219 388996 113220 389060
rect 113284 388996 113285 389060
rect 113219 388995 113285 388996
rect 111563 381036 111629 381037
rect 111563 380972 111564 381036
rect 111628 380972 111629 381036
rect 111563 380971 111629 380972
rect 111750 378725 111810 388995
rect 111747 378724 111813 378725
rect 111747 378660 111748 378724
rect 111812 378660 111813 378724
rect 111747 378659 111813 378660
rect 109794 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 110414 363454
rect 109794 363134 110414 363218
rect 109794 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 110414 363134
rect 108803 349212 108869 349213
rect 108803 349148 108804 349212
rect 108868 349148 108869 349212
rect 108803 349147 108869 349148
rect 109794 331592 110414 362898
rect 113514 367174 114134 388356
rect 114326 378181 114386 445707
rect 115798 379269 115858 447203
rect 115982 390421 116042 473995
rect 117234 446407 117854 478338
rect 120954 698614 121574 710042
rect 138954 711558 139574 711590
rect 138954 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 139574 711558
rect 138954 711238 139574 711322
rect 138954 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 139574 711238
rect 135234 709638 135854 709670
rect 135234 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 135854 709638
rect 135234 709318 135854 709402
rect 135234 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 135854 709318
rect 131514 707718 132134 707750
rect 131514 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 132134 707718
rect 131514 707398 132134 707482
rect 131514 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 132134 707398
rect 120954 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 121574 698614
rect 120954 698294 121574 698378
rect 120954 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 121574 698294
rect 120954 662614 121574 698058
rect 120954 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 121574 662614
rect 120954 662294 121574 662378
rect 120954 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 121574 662294
rect 120954 626614 121574 662058
rect 120954 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 121574 626614
rect 120954 626294 121574 626378
rect 120954 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 121574 626294
rect 120954 590614 121574 626058
rect 120954 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 121574 590614
rect 120954 590294 121574 590378
rect 120954 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 121574 590294
rect 120954 554614 121574 590058
rect 127794 705798 128414 705830
rect 127794 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 128414 705798
rect 127794 705478 128414 705562
rect 127794 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 128414 705478
rect 127794 669454 128414 705242
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 633454 128414 668898
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 127794 597454 128414 632898
rect 127794 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 128414 597454
rect 127794 597134 128414 597218
rect 127794 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 128414 597134
rect 124259 577556 124325 577557
rect 124259 577492 124260 577556
rect 124324 577492 124325 577556
rect 124259 577491 124325 577492
rect 121683 572796 121749 572797
rect 121683 572732 121684 572796
rect 121748 572732 121749 572796
rect 121683 572731 121749 572732
rect 120954 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 121574 554614
rect 120954 554294 121574 554378
rect 120954 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 121574 554294
rect 120954 518614 121574 554058
rect 120954 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 121574 518614
rect 120954 518294 121574 518378
rect 120954 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 121574 518294
rect 120954 482614 121574 518058
rect 120954 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 121574 482614
rect 120954 482294 121574 482378
rect 120954 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 121574 482294
rect 118187 469844 118253 469845
rect 118187 469780 118188 469844
rect 118252 469780 118253 469844
rect 118187 469779 118253 469780
rect 118003 445772 118069 445773
rect 118003 445708 118004 445772
rect 118068 445708 118069 445772
rect 118003 445707 118069 445708
rect 115979 390420 116045 390421
rect 115979 390356 115980 390420
rect 116044 390356 116045 390420
rect 115979 390355 116045 390356
rect 115795 379268 115861 379269
rect 115795 379204 115796 379268
rect 115860 379204 115861 379268
rect 115795 379203 115861 379204
rect 114323 378180 114389 378181
rect 114323 378116 114324 378180
rect 114388 378116 114389 378180
rect 114323 378115 114389 378116
rect 113514 366938 113546 367174
rect 113782 366938 113866 367174
rect 114102 366938 114134 367174
rect 113514 366854 114134 366938
rect 113514 366618 113546 366854
rect 113782 366618 113866 366854
rect 114102 366618 114134 366854
rect 113514 331592 114134 366618
rect 117234 370894 117854 388356
rect 117234 370658 117266 370894
rect 117502 370658 117586 370894
rect 117822 370658 117854 370894
rect 117234 370574 117854 370658
rect 117234 370338 117266 370574
rect 117502 370338 117586 370574
rect 117822 370338 117854 370574
rect 117234 334894 117854 370338
rect 118006 339421 118066 445707
rect 118190 390421 118250 469779
rect 118739 458828 118805 458829
rect 118739 458764 118740 458828
rect 118804 458764 118805 458828
rect 118739 458763 118805 458764
rect 118742 390421 118802 458763
rect 120027 450532 120093 450533
rect 120027 450468 120028 450532
rect 120092 450468 120093 450532
rect 120027 450467 120093 450468
rect 120030 426053 120090 450467
rect 120954 446407 121574 482058
rect 120027 426052 120093 426053
rect 120027 425988 120028 426052
rect 120092 425988 120093 426052
rect 120027 425987 120093 425988
rect 121686 422310 121746 572731
rect 122603 479500 122669 479501
rect 122603 479436 122604 479500
rect 122668 479436 122669 479500
rect 122603 479435 122669 479436
rect 121502 422250 121746 422310
rect 121502 420885 121562 422250
rect 121499 420884 121565 420885
rect 121499 420820 121500 420884
rect 121564 420820 121565 420884
rect 121499 420819 121565 420820
rect 121502 419661 121562 420819
rect 121499 419660 121565 419661
rect 121499 419596 121500 419660
rect 121564 419596 121565 419660
rect 121499 419595 121565 419596
rect 119058 417454 119378 417486
rect 119058 417218 119100 417454
rect 119336 417218 119378 417454
rect 119058 417134 119378 417218
rect 119058 416898 119100 417134
rect 119336 416898 119378 417134
rect 119058 416866 119378 416898
rect 121502 390693 121562 419595
rect 122606 403749 122666 479435
rect 122971 453252 123037 453253
rect 122971 453188 122972 453252
rect 123036 453188 123037 453252
rect 122971 453187 123037 453188
rect 122974 435437 123034 453187
rect 124262 443869 124322 577491
rect 127794 561454 128414 596898
rect 127794 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 128414 561454
rect 127794 561134 128414 561218
rect 127794 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 128414 561134
rect 127794 525454 128414 560898
rect 127794 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 128414 525454
rect 127794 525134 128414 525218
rect 127794 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 128414 525134
rect 127794 489454 128414 524898
rect 127794 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 128414 489454
rect 127794 489134 128414 489218
rect 127794 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 128414 489134
rect 127794 453454 128414 488898
rect 127794 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 128414 453454
rect 127794 453134 128414 453218
rect 127794 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 128414 453134
rect 124259 443868 124325 443869
rect 124259 443804 124260 443868
rect 124324 443804 124325 443868
rect 124259 443803 124325 443804
rect 122971 435436 123037 435437
rect 122971 435372 122972 435436
rect 123036 435372 123037 435436
rect 122971 435371 123037 435372
rect 127794 417454 128414 452898
rect 127794 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 128414 417454
rect 127794 417134 128414 417218
rect 127794 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 128414 417134
rect 122603 403748 122669 403749
rect 122603 403684 122604 403748
rect 122668 403684 122669 403748
rect 122603 403683 122669 403684
rect 121499 390692 121565 390693
rect 121499 390628 121500 390692
rect 121564 390628 121565 390692
rect 121499 390627 121565 390628
rect 118187 390420 118253 390421
rect 118187 390356 118188 390420
rect 118252 390356 118253 390420
rect 118187 390355 118253 390356
rect 118739 390420 118805 390421
rect 118739 390356 118740 390420
rect 118804 390356 118805 390420
rect 118739 390355 118805 390356
rect 120954 374614 121574 388356
rect 120954 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 121574 374614
rect 120954 374294 121574 374378
rect 120954 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 121574 374294
rect 118003 339420 118069 339421
rect 118003 339356 118004 339420
rect 118068 339356 118069 339420
rect 118003 339355 118069 339356
rect 117234 334658 117266 334894
rect 117502 334658 117586 334894
rect 117822 334658 117854 334894
rect 117234 334574 117854 334658
rect 117234 334338 117266 334574
rect 117502 334338 117586 334574
rect 117822 334338 117854 334574
rect 117234 331592 117854 334338
rect 120954 338614 121574 374058
rect 120954 338378 120986 338614
rect 121222 338378 121306 338614
rect 121542 338378 121574 338614
rect 120954 338294 121574 338378
rect 120954 338058 120986 338294
rect 121222 338058 121306 338294
rect 121542 338058 121574 338294
rect 120954 331592 121574 338058
rect 127794 381454 128414 416898
rect 127794 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 128414 381454
rect 127794 381134 128414 381218
rect 127794 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 128414 381134
rect 127794 345454 128414 380898
rect 127794 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 128414 345454
rect 127794 345134 128414 345218
rect 127794 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 128414 345134
rect 127794 331592 128414 344898
rect 131514 673174 132134 707162
rect 131514 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 132134 673174
rect 131514 672854 132134 672938
rect 131514 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 132134 672854
rect 131514 637174 132134 672618
rect 131514 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 132134 637174
rect 131514 636854 132134 636938
rect 131514 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 132134 636854
rect 131514 601174 132134 636618
rect 131514 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 132134 601174
rect 131514 600854 132134 600938
rect 131514 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 132134 600854
rect 131514 565174 132134 600618
rect 131514 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 132134 565174
rect 131514 564854 132134 564938
rect 131514 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 132134 564854
rect 131514 529174 132134 564618
rect 131514 528938 131546 529174
rect 131782 528938 131866 529174
rect 132102 528938 132134 529174
rect 131514 528854 132134 528938
rect 131514 528618 131546 528854
rect 131782 528618 131866 528854
rect 132102 528618 132134 528854
rect 131514 493174 132134 528618
rect 131514 492938 131546 493174
rect 131782 492938 131866 493174
rect 132102 492938 132134 493174
rect 131514 492854 132134 492938
rect 131514 492618 131546 492854
rect 131782 492618 131866 492854
rect 132102 492618 132134 492854
rect 131514 457174 132134 492618
rect 131514 456938 131546 457174
rect 131782 456938 131866 457174
rect 132102 456938 132134 457174
rect 131514 456854 132134 456938
rect 131514 456618 131546 456854
rect 131782 456618 131866 456854
rect 132102 456618 132134 456854
rect 131514 421174 132134 456618
rect 131514 420938 131546 421174
rect 131782 420938 131866 421174
rect 132102 420938 132134 421174
rect 131514 420854 132134 420938
rect 131514 420618 131546 420854
rect 131782 420618 131866 420854
rect 132102 420618 132134 420854
rect 131514 385174 132134 420618
rect 131514 384938 131546 385174
rect 131782 384938 131866 385174
rect 132102 384938 132134 385174
rect 131514 384854 132134 384938
rect 131514 384618 131546 384854
rect 131782 384618 131866 384854
rect 132102 384618 132134 384854
rect 131514 349174 132134 384618
rect 131514 348938 131546 349174
rect 131782 348938 131866 349174
rect 132102 348938 132134 349174
rect 131514 348854 132134 348938
rect 131514 348618 131546 348854
rect 131782 348618 131866 348854
rect 132102 348618 132134 348854
rect 131514 331592 132134 348618
rect 135234 676894 135854 709082
rect 135234 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 135854 676894
rect 135234 676574 135854 676658
rect 135234 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 135854 676574
rect 135234 640894 135854 676338
rect 135234 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 135854 640894
rect 135234 640574 135854 640658
rect 135234 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 135854 640574
rect 135234 604894 135854 640338
rect 135234 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 135854 604894
rect 135234 604574 135854 604658
rect 135234 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 135854 604574
rect 135234 568894 135854 604338
rect 135234 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 135854 568894
rect 135234 568574 135854 568658
rect 135234 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 135854 568574
rect 135234 532894 135854 568338
rect 135234 532658 135266 532894
rect 135502 532658 135586 532894
rect 135822 532658 135854 532894
rect 135234 532574 135854 532658
rect 135234 532338 135266 532574
rect 135502 532338 135586 532574
rect 135822 532338 135854 532574
rect 135234 496894 135854 532338
rect 135234 496658 135266 496894
rect 135502 496658 135586 496894
rect 135822 496658 135854 496894
rect 135234 496574 135854 496658
rect 135234 496338 135266 496574
rect 135502 496338 135586 496574
rect 135822 496338 135854 496574
rect 135234 460894 135854 496338
rect 135234 460658 135266 460894
rect 135502 460658 135586 460894
rect 135822 460658 135854 460894
rect 135234 460574 135854 460658
rect 135234 460338 135266 460574
rect 135502 460338 135586 460574
rect 135822 460338 135854 460574
rect 135234 424894 135854 460338
rect 135234 424658 135266 424894
rect 135502 424658 135586 424894
rect 135822 424658 135854 424894
rect 135234 424574 135854 424658
rect 135234 424338 135266 424574
rect 135502 424338 135586 424574
rect 135822 424338 135854 424574
rect 135234 388894 135854 424338
rect 135234 388658 135266 388894
rect 135502 388658 135586 388894
rect 135822 388658 135854 388894
rect 135234 388574 135854 388658
rect 135234 388338 135266 388574
rect 135502 388338 135586 388574
rect 135822 388338 135854 388574
rect 135234 352894 135854 388338
rect 135234 352658 135266 352894
rect 135502 352658 135586 352894
rect 135822 352658 135854 352894
rect 135234 352574 135854 352658
rect 135234 352338 135266 352574
rect 135502 352338 135586 352574
rect 135822 352338 135854 352574
rect 135234 331592 135854 352338
rect 138954 680614 139574 711002
rect 156954 710598 157574 711590
rect 156954 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 157574 710598
rect 156954 710278 157574 710362
rect 156954 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 157574 710278
rect 153234 708678 153854 709670
rect 153234 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 153854 708678
rect 153234 708358 153854 708442
rect 153234 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 153854 708358
rect 149514 706758 150134 707750
rect 149514 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 150134 706758
rect 149514 706438 150134 706522
rect 149514 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 150134 706438
rect 138954 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 139574 680614
rect 138954 680294 139574 680378
rect 138954 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 139574 680294
rect 138954 644614 139574 680058
rect 138954 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 139574 644614
rect 138954 644294 139574 644378
rect 138954 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 139574 644294
rect 138954 608614 139574 644058
rect 138954 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 139574 608614
rect 138954 608294 139574 608378
rect 138954 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 139574 608294
rect 138954 572614 139574 608058
rect 138954 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 139574 572614
rect 138954 572294 139574 572378
rect 138954 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 139574 572294
rect 138954 536614 139574 572058
rect 138954 536378 138986 536614
rect 139222 536378 139306 536614
rect 139542 536378 139574 536614
rect 138954 536294 139574 536378
rect 138954 536058 138986 536294
rect 139222 536058 139306 536294
rect 139542 536058 139574 536294
rect 138954 500614 139574 536058
rect 138954 500378 138986 500614
rect 139222 500378 139306 500614
rect 139542 500378 139574 500614
rect 138954 500294 139574 500378
rect 138954 500058 138986 500294
rect 139222 500058 139306 500294
rect 139542 500058 139574 500294
rect 138954 464614 139574 500058
rect 138954 464378 138986 464614
rect 139222 464378 139306 464614
rect 139542 464378 139574 464614
rect 138954 464294 139574 464378
rect 138954 464058 138986 464294
rect 139222 464058 139306 464294
rect 139542 464058 139574 464294
rect 138954 428614 139574 464058
rect 138954 428378 138986 428614
rect 139222 428378 139306 428614
rect 139542 428378 139574 428614
rect 138954 428294 139574 428378
rect 138954 428058 138986 428294
rect 139222 428058 139306 428294
rect 139542 428058 139574 428294
rect 138954 392614 139574 428058
rect 138954 392378 138986 392614
rect 139222 392378 139306 392614
rect 139542 392378 139574 392614
rect 138954 392294 139574 392378
rect 138954 392058 138986 392294
rect 139222 392058 139306 392294
rect 139542 392058 139574 392294
rect 138954 356614 139574 392058
rect 138954 356378 138986 356614
rect 139222 356378 139306 356614
rect 139542 356378 139574 356614
rect 138954 356294 139574 356378
rect 138954 356058 138986 356294
rect 139222 356058 139306 356294
rect 139542 356058 139574 356294
rect 138954 331592 139574 356058
rect 145794 704838 146414 705830
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 579454 146414 614898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 543454 146414 578898
rect 145794 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 146414 543454
rect 145794 543134 146414 543218
rect 145794 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 146414 543134
rect 145794 507454 146414 542898
rect 145794 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 146414 507454
rect 145794 507134 146414 507218
rect 145794 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 146414 507134
rect 145794 471454 146414 506898
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 145794 435454 146414 470898
rect 145794 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 146414 435454
rect 145794 435134 146414 435218
rect 145794 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 146414 435134
rect 145794 399454 146414 434898
rect 145794 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 146414 399454
rect 145794 399134 146414 399218
rect 145794 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 146414 399134
rect 145794 363454 146414 398898
rect 145794 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 146414 363454
rect 145794 363134 146414 363218
rect 145794 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 146414 363134
rect 145794 331592 146414 362898
rect 149514 691174 150134 706202
rect 149514 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 150134 691174
rect 149514 690854 150134 690938
rect 149514 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 150134 690854
rect 149514 655174 150134 690618
rect 149514 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 150134 655174
rect 149514 654854 150134 654938
rect 149514 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 150134 654854
rect 149514 619174 150134 654618
rect 149514 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 150134 619174
rect 149514 618854 150134 618938
rect 149514 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 150134 618854
rect 149514 583174 150134 618618
rect 149514 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 150134 583174
rect 149514 582854 150134 582938
rect 149514 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 150134 582854
rect 149514 547174 150134 582618
rect 149514 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 150134 547174
rect 149514 546854 150134 546938
rect 149514 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 150134 546854
rect 149514 511174 150134 546618
rect 149514 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 150134 511174
rect 149514 510854 150134 510938
rect 149514 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 150134 510854
rect 149514 475174 150134 510618
rect 149514 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 150134 475174
rect 149514 474854 150134 474938
rect 149514 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 150134 474854
rect 149514 439174 150134 474618
rect 149514 438938 149546 439174
rect 149782 438938 149866 439174
rect 150102 438938 150134 439174
rect 149514 438854 150134 438938
rect 149514 438618 149546 438854
rect 149782 438618 149866 438854
rect 150102 438618 150134 438854
rect 149514 403174 150134 438618
rect 149514 402938 149546 403174
rect 149782 402938 149866 403174
rect 150102 402938 150134 403174
rect 149514 402854 150134 402938
rect 149514 402618 149546 402854
rect 149782 402618 149866 402854
rect 150102 402618 150134 402854
rect 149514 367174 150134 402618
rect 149514 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 150134 367174
rect 149514 366854 150134 366938
rect 149514 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 150134 366854
rect 149514 331592 150134 366618
rect 153234 694894 153854 708122
rect 153234 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 153854 694894
rect 153234 694574 153854 694658
rect 153234 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 153854 694574
rect 153234 658894 153854 694338
rect 153234 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 153854 658894
rect 153234 658574 153854 658658
rect 153234 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 153854 658574
rect 153234 622894 153854 658338
rect 153234 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 153854 622894
rect 153234 622574 153854 622658
rect 153234 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 153854 622574
rect 153234 586894 153854 622338
rect 153234 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 153854 586894
rect 153234 586574 153854 586658
rect 153234 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 153854 586574
rect 153234 550894 153854 586338
rect 153234 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 153854 550894
rect 153234 550574 153854 550658
rect 153234 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 153854 550574
rect 153234 514894 153854 550338
rect 153234 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 153854 514894
rect 153234 514574 153854 514658
rect 153234 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 153854 514574
rect 153234 478894 153854 514338
rect 156954 698614 157574 710042
rect 174954 711558 175574 711590
rect 174954 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 175574 711558
rect 174954 711238 175574 711322
rect 174954 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 175574 711238
rect 171234 709638 171854 709670
rect 171234 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 171854 709638
rect 171234 709318 171854 709402
rect 171234 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 171854 709318
rect 167514 707718 168134 707750
rect 167514 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 168134 707718
rect 167514 707398 168134 707482
rect 167514 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 168134 707398
rect 156954 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 157574 698614
rect 156954 698294 157574 698378
rect 156954 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 157574 698294
rect 156954 662614 157574 698058
rect 156954 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 157574 662614
rect 156954 662294 157574 662378
rect 156954 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 157574 662294
rect 156954 626614 157574 662058
rect 156954 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 157574 626614
rect 156954 626294 157574 626378
rect 156954 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 157574 626294
rect 156954 590614 157574 626058
rect 156954 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 157574 590614
rect 156954 590294 157574 590378
rect 156954 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 157574 590294
rect 156954 554614 157574 590058
rect 156954 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 157574 554614
rect 156954 554294 157574 554378
rect 156954 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 157574 554294
rect 156954 518614 157574 554058
rect 163794 705798 164414 705830
rect 163794 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 164414 705798
rect 163794 705478 164414 705562
rect 163794 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 164414 705478
rect 163794 669454 164414 705242
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 633454 164414 668898
rect 163794 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 164414 633454
rect 163794 633134 164414 633218
rect 163794 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 164414 633134
rect 163794 597454 164414 632898
rect 163794 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 164414 597454
rect 163794 597134 164414 597218
rect 163794 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 164414 597134
rect 163794 561454 164414 596898
rect 163794 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 164414 561454
rect 163794 561134 164414 561218
rect 163794 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 164414 561134
rect 161979 543964 162045 543965
rect 161979 543900 161980 543964
rect 162044 543900 162045 543964
rect 161979 543899 162045 543900
rect 160691 539884 160757 539885
rect 160691 539820 160692 539884
rect 160756 539820 160757 539884
rect 160691 539819 160757 539820
rect 156954 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 157574 518614
rect 156954 518294 157574 518378
rect 156954 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 157574 518294
rect 155723 504388 155789 504389
rect 155723 504324 155724 504388
rect 155788 504324 155789 504388
rect 155723 504323 155789 504324
rect 153234 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 153854 478894
rect 153234 478574 153854 478658
rect 153234 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 153854 478574
rect 153234 442894 153854 478338
rect 153234 442658 153266 442894
rect 153502 442658 153586 442894
rect 153822 442658 153854 442894
rect 153234 442574 153854 442658
rect 153234 442338 153266 442574
rect 153502 442338 153586 442574
rect 153822 442338 153854 442574
rect 153234 406894 153854 442338
rect 154067 442236 154133 442237
rect 154067 442172 154068 442236
rect 154132 442172 154133 442236
rect 154067 442171 154133 442172
rect 153234 406658 153266 406894
rect 153502 406658 153586 406894
rect 153822 406658 153854 406894
rect 153234 406574 153854 406658
rect 153234 406338 153266 406574
rect 153502 406338 153586 406574
rect 153822 406338 153854 406574
rect 153234 370894 153854 406338
rect 153234 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 153854 370894
rect 153234 370574 153854 370658
rect 153234 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 153854 370574
rect 153234 334894 153854 370338
rect 153234 334658 153266 334894
rect 153502 334658 153586 334894
rect 153822 334658 153854 334894
rect 153234 334574 153854 334658
rect 153234 334338 153266 334574
rect 153502 334338 153586 334574
rect 153822 334338 153854 334574
rect 153234 331592 153854 334338
rect 93899 330172 93965 330173
rect 93899 330108 93900 330172
rect 93964 330108 93965 330172
rect 93899 330107 93965 330108
rect 88338 309454 88658 309486
rect 88338 309218 88380 309454
rect 88616 309218 88658 309454
rect 88338 309134 88658 309218
rect 88338 308898 88380 309134
rect 88616 308898 88658 309134
rect 88338 308866 88658 308898
rect 119058 309454 119378 309486
rect 119058 309218 119100 309454
rect 119336 309218 119378 309454
rect 119058 309134 119378 309218
rect 119058 308898 119100 309134
rect 119336 308898 119378 309134
rect 119058 308866 119378 308898
rect 149778 309454 150098 309486
rect 149778 309218 149820 309454
rect 150056 309218 150098 309454
rect 149778 309134 150098 309218
rect 149778 308898 149820 309134
rect 150056 308898 150098 309134
rect 149778 308866 150098 308898
rect 103698 291454 104018 291486
rect 103698 291218 103740 291454
rect 103976 291218 104018 291454
rect 103698 291134 104018 291218
rect 103698 290898 103740 291134
rect 103976 290898 104018 291134
rect 103698 290866 104018 290898
rect 134418 291454 134738 291486
rect 134418 291218 134460 291454
rect 134696 291218 134738 291454
rect 134418 291134 134738 291218
rect 134418 290898 134460 291134
rect 134696 290898 134738 291134
rect 134418 290866 134738 290898
rect 88338 273454 88658 273486
rect 88338 273218 88380 273454
rect 88616 273218 88658 273454
rect 88338 273134 88658 273218
rect 88338 272898 88380 273134
rect 88616 272898 88658 273134
rect 88338 272866 88658 272898
rect 119058 273454 119378 273486
rect 119058 273218 119100 273454
rect 119336 273218 119378 273454
rect 119058 273134 119378 273218
rect 119058 272898 119100 273134
rect 119336 272898 119378 273134
rect 119058 272866 119378 272898
rect 149778 273454 150098 273486
rect 149778 273218 149820 273454
rect 150056 273218 150098 273454
rect 149778 273134 150098 273218
rect 149778 272898 149820 273134
rect 150056 272898 150098 273134
rect 149778 272866 150098 272898
rect 103698 255454 104018 255486
rect 103698 255218 103740 255454
rect 103976 255218 104018 255454
rect 103698 255134 104018 255218
rect 103698 254898 103740 255134
rect 103976 254898 104018 255134
rect 103698 254866 104018 254898
rect 134418 255454 134738 255486
rect 134418 255218 134460 255454
rect 134696 255218 134738 255454
rect 134418 255134 134738 255218
rect 134418 254898 134460 255134
rect 134696 254898 134738 255134
rect 134418 254866 134738 254898
rect 83963 237284 84029 237285
rect 83963 237220 83964 237284
rect 84028 237220 84029 237284
rect 83963 237219 84029 237220
rect 84954 230614 85574 239592
rect 84954 230378 84986 230614
rect 85222 230378 85306 230614
rect 85542 230378 85574 230614
rect 84954 230294 85574 230378
rect 84954 230058 84986 230294
rect 85222 230058 85306 230294
rect 85542 230058 85574 230294
rect 82675 227628 82741 227629
rect 82675 227564 82676 227628
rect 82740 227564 82741 227628
rect 82675 227563 82741 227564
rect 81234 226658 81266 226894
rect 81502 226658 81586 226894
rect 81822 226658 81854 226894
rect 81234 226574 81854 226658
rect 81234 226338 81266 226574
rect 81502 226338 81586 226574
rect 81822 226338 81854 226574
rect 81234 190894 81854 226338
rect 81234 190658 81266 190894
rect 81502 190658 81586 190894
rect 81822 190658 81854 190894
rect 81234 190574 81854 190658
rect 81234 190338 81266 190574
rect 81502 190338 81586 190574
rect 81822 190338 81854 190574
rect 81234 176600 81854 190338
rect 84954 194614 85574 230058
rect 84954 194378 84986 194614
rect 85222 194378 85306 194614
rect 85542 194378 85574 194614
rect 84954 194294 85574 194378
rect 84954 194058 84986 194294
rect 85222 194058 85306 194294
rect 85542 194058 85574 194294
rect 84954 176600 85574 194058
rect 91794 237454 92414 239592
rect 91794 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 92414 237454
rect 91794 237134 92414 237218
rect 91794 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 92414 237134
rect 91794 201454 92414 236898
rect 91794 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 92414 201454
rect 91794 201134 92414 201218
rect 91794 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 92414 201134
rect 91794 176600 92414 200898
rect 95514 205174 96134 239592
rect 95514 204938 95546 205174
rect 95782 204938 95866 205174
rect 96102 204938 96134 205174
rect 95514 204854 96134 204938
rect 95514 204618 95546 204854
rect 95782 204618 95866 204854
rect 96102 204618 96134 204854
rect 95514 176600 96134 204618
rect 99234 208894 99854 239592
rect 99234 208658 99266 208894
rect 99502 208658 99586 208894
rect 99822 208658 99854 208894
rect 99234 208574 99854 208658
rect 99234 208338 99266 208574
rect 99502 208338 99586 208574
rect 99822 208338 99854 208574
rect 98315 177580 98381 177581
rect 98315 177516 98316 177580
rect 98380 177516 98381 177580
rect 98315 177515 98381 177516
rect 97027 176900 97093 176901
rect 97027 176836 97028 176900
rect 97092 176836 97093 176900
rect 97027 176835 97093 176836
rect 97030 175130 97090 176835
rect 96960 175070 97090 175130
rect 98318 175130 98378 177515
rect 99234 176600 99854 208338
rect 102954 212614 103574 239592
rect 102954 212378 102986 212614
rect 103222 212378 103306 212614
rect 103542 212378 103574 212614
rect 102954 212294 103574 212378
rect 102954 212058 102986 212294
rect 103222 212058 103306 212294
rect 103542 212058 103574 212294
rect 100707 177580 100773 177581
rect 100707 177516 100708 177580
rect 100772 177516 100773 177580
rect 100707 177515 100773 177516
rect 99419 176492 99485 176493
rect 99419 176428 99420 176492
rect 99484 176428 99485 176492
rect 99419 176427 99485 176428
rect 99422 175130 99482 176427
rect 98318 175070 98380 175130
rect 96960 174494 97020 175070
rect 98320 174494 98380 175070
rect 99408 175070 99482 175130
rect 100710 175130 100770 177515
rect 101995 176900 102061 176901
rect 101995 176836 101996 176900
rect 102060 176836 102061 176900
rect 101995 176835 102061 176836
rect 101998 175130 102058 176835
rect 102954 176600 103574 212058
rect 109794 219454 110414 239592
rect 109794 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 110414 219454
rect 109794 219134 110414 219218
rect 109794 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 110414 219134
rect 109794 183454 110414 218898
rect 109794 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 110414 183454
rect 109794 183134 110414 183218
rect 109794 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 110414 183134
rect 109539 177852 109605 177853
rect 109539 177788 109540 177852
rect 109604 177788 109605 177852
rect 109539 177787 109605 177788
rect 105675 177580 105741 177581
rect 105675 177516 105676 177580
rect 105740 177516 105741 177580
rect 105675 177515 105741 177516
rect 106963 177580 107029 177581
rect 106963 177516 106964 177580
rect 107028 177516 107029 177580
rect 106963 177515 107029 177516
rect 104571 177036 104637 177037
rect 104571 176972 104572 177036
rect 104636 176972 104637 177036
rect 104571 176971 104637 176972
rect 103283 176492 103349 176493
rect 103283 176428 103284 176492
rect 103348 176428 103349 176492
rect 103283 176427 103349 176428
rect 100710 175070 100828 175130
rect 99408 174494 99468 175070
rect 100768 174494 100828 175070
rect 101992 175070 102058 175130
rect 103286 175130 103346 176427
rect 104574 175130 104634 176971
rect 105678 175130 105738 177515
rect 103286 175070 103412 175130
rect 104574 175070 104636 175130
rect 101992 174494 102052 175070
rect 103352 174494 103412 175070
rect 104576 174494 104636 175070
rect 105664 175070 105738 175130
rect 106966 175130 107026 177515
rect 108067 175404 108133 175405
rect 108067 175340 108068 175404
rect 108132 175340 108133 175404
rect 108067 175339 108133 175340
rect 108070 175130 108130 175339
rect 109542 175130 109602 177787
rect 109794 176600 110414 182898
rect 113514 223174 114134 239592
rect 113514 222938 113546 223174
rect 113782 222938 113866 223174
rect 114102 222938 114134 223174
rect 113514 222854 114134 222938
rect 113514 222618 113546 222854
rect 113782 222618 113866 222854
rect 114102 222618 114134 222854
rect 113514 187174 114134 222618
rect 113514 186938 113546 187174
rect 113782 186938 113866 187174
rect 114102 186938 114134 187174
rect 113514 186854 114134 186938
rect 113514 186618 113546 186854
rect 113782 186618 113866 186854
rect 114102 186618 114134 186854
rect 110643 177988 110709 177989
rect 110643 177924 110644 177988
rect 110708 177924 110709 177988
rect 110643 177923 110709 177924
rect 106966 175070 107084 175130
rect 108070 175070 108172 175130
rect 105664 174494 105724 175070
rect 107024 174494 107084 175070
rect 108112 174494 108172 175070
rect 109472 175070 109602 175130
rect 110646 175130 110706 177923
rect 113219 177580 113285 177581
rect 113219 177516 113220 177580
rect 113284 177516 113285 177580
rect 113219 177515 113285 177516
rect 112115 177172 112181 177173
rect 112115 177108 112116 177172
rect 112180 177108 112181 177172
rect 112115 177107 112181 177108
rect 112118 175130 112178 177107
rect 113222 175130 113282 177515
rect 113514 176600 114134 186618
rect 117234 226894 117854 239592
rect 117234 226658 117266 226894
rect 117502 226658 117586 226894
rect 117822 226658 117854 226894
rect 117234 226574 117854 226658
rect 117234 226338 117266 226574
rect 117502 226338 117586 226574
rect 117822 226338 117854 226574
rect 117234 190894 117854 226338
rect 117234 190658 117266 190894
rect 117502 190658 117586 190894
rect 117822 190658 117854 190894
rect 117234 190574 117854 190658
rect 117234 190338 117266 190574
rect 117502 190338 117586 190574
rect 117822 190338 117854 190574
rect 116899 178260 116965 178261
rect 116899 178196 116900 178260
rect 116964 178196 116965 178260
rect 116899 178195 116965 178196
rect 115795 177580 115861 177581
rect 115795 177516 115796 177580
rect 115860 177516 115861 177580
rect 115795 177515 115861 177516
rect 114323 177172 114389 177173
rect 114323 177108 114324 177172
rect 114388 177108 114389 177172
rect 114323 177107 114389 177108
rect 110646 175070 110756 175130
rect 109472 174494 109532 175070
rect 110696 174494 110756 175070
rect 112056 175070 112178 175130
rect 113144 175070 113282 175130
rect 114326 175130 114386 177107
rect 115798 175130 115858 177515
rect 114326 175070 114428 175130
rect 112056 174494 112116 175070
rect 113144 174494 113204 175070
rect 114368 174494 114428 175070
rect 115728 175070 115858 175130
rect 116902 175130 116962 178195
rect 117234 176600 117854 190338
rect 120954 230614 121574 239592
rect 120954 230378 120986 230614
rect 121222 230378 121306 230614
rect 121542 230378 121574 230614
rect 120954 230294 121574 230378
rect 120954 230058 120986 230294
rect 121222 230058 121306 230294
rect 121542 230058 121574 230294
rect 120954 194614 121574 230058
rect 120954 194378 120986 194614
rect 121222 194378 121306 194614
rect 121542 194378 121574 194614
rect 120954 194294 121574 194378
rect 120954 194058 120986 194294
rect 121222 194058 121306 194294
rect 121542 194058 121574 194294
rect 118371 177580 118437 177581
rect 118371 177516 118372 177580
rect 118436 177516 118437 177580
rect 118371 177515 118437 177516
rect 118374 175130 118434 177515
rect 119475 177172 119541 177173
rect 119475 177108 119476 177172
rect 119540 177108 119541 177172
rect 119475 177107 119541 177108
rect 119478 175130 119538 177107
rect 120954 176600 121574 194058
rect 127794 237454 128414 239592
rect 127794 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 128414 237454
rect 127794 237134 128414 237218
rect 127794 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 128414 237134
rect 127794 201454 128414 236898
rect 127794 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 128414 201454
rect 127794 201134 128414 201218
rect 127794 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 128414 201134
rect 121867 177580 121933 177581
rect 121867 177516 121868 177580
rect 121932 177516 121933 177580
rect 121867 177515 121933 177516
rect 124443 177580 124509 177581
rect 124443 177516 124444 177580
rect 124508 177516 124509 177580
rect 124443 177515 124509 177516
rect 127019 177580 127085 177581
rect 127019 177516 127020 177580
rect 127084 177516 127085 177580
rect 127019 177515 127085 177516
rect 120763 175540 120829 175541
rect 120763 175476 120764 175540
rect 120828 175476 120829 175540
rect 120763 175475 120829 175476
rect 120766 175130 120826 175475
rect 121870 175130 121930 177515
rect 123155 176764 123221 176765
rect 123155 176700 123156 176764
rect 123220 176700 123221 176764
rect 123155 176699 123221 176700
rect 123158 175130 123218 176699
rect 124446 175130 124506 177515
rect 125731 176764 125797 176765
rect 125731 176700 125732 176764
rect 125796 176700 125797 176764
rect 125731 176699 125797 176700
rect 125734 175130 125794 176699
rect 127022 175130 127082 177515
rect 127794 176600 128414 200898
rect 131514 205174 132134 239592
rect 131514 204938 131546 205174
rect 131782 204938 131866 205174
rect 132102 204938 132134 205174
rect 131514 204854 132134 204938
rect 131514 204618 131546 204854
rect 131782 204618 131866 204854
rect 132102 204618 132134 204854
rect 129411 176764 129477 176765
rect 129411 176700 129412 176764
rect 129476 176700 129477 176764
rect 129411 176699 129477 176700
rect 128123 176492 128189 176493
rect 128123 176428 128124 176492
rect 128188 176428 128189 176492
rect 128123 176427 128189 176428
rect 128126 175130 128186 176427
rect 116902 175070 117012 175130
rect 115728 174494 115788 175070
rect 116952 174494 117012 175070
rect 118312 175070 118434 175130
rect 119400 175070 119538 175130
rect 120760 175070 120826 175130
rect 121848 175070 121930 175130
rect 123072 175070 123218 175130
rect 124432 175070 124506 175130
rect 125656 175070 125794 175130
rect 127016 175070 127082 175130
rect 128104 175070 128186 175130
rect 129414 175130 129474 176699
rect 131514 176600 132134 204618
rect 135234 208894 135854 239592
rect 135234 208658 135266 208894
rect 135502 208658 135586 208894
rect 135822 208658 135854 208894
rect 135234 208574 135854 208658
rect 135234 208338 135266 208574
rect 135502 208338 135586 208574
rect 135822 208338 135854 208574
rect 132355 177580 132421 177581
rect 132355 177516 132356 177580
rect 132420 177516 132421 177580
rect 132355 177515 132421 177516
rect 133091 177580 133157 177581
rect 133091 177516 133092 177580
rect 133156 177516 133157 177580
rect 133091 177515 133157 177516
rect 130699 175676 130765 175677
rect 130699 175612 130700 175676
rect 130764 175612 130765 175676
rect 130699 175611 130765 175612
rect 130702 175130 130762 175611
rect 132358 175130 132418 177515
rect 129414 175070 129524 175130
rect 118312 174494 118372 175070
rect 119400 174494 119460 175070
rect 120760 174494 120820 175070
rect 121848 174494 121908 175070
rect 123072 174494 123132 175070
rect 124432 174494 124492 175070
rect 125656 174494 125716 175070
rect 127016 174494 127076 175070
rect 128104 174494 128164 175070
rect 129464 174494 129524 175070
rect 130688 175070 130762 175130
rect 132048 175070 132418 175130
rect 133094 175130 133154 177515
rect 134379 177172 134445 177173
rect 134379 177108 134380 177172
rect 134444 177108 134445 177172
rect 134379 177107 134445 177108
rect 134382 175130 134442 177107
rect 135234 176600 135854 208338
rect 138954 212614 139574 239592
rect 138954 212378 138986 212614
rect 139222 212378 139306 212614
rect 139542 212378 139574 212614
rect 138954 212294 139574 212378
rect 138954 212058 138986 212294
rect 139222 212058 139306 212294
rect 139542 212058 139574 212294
rect 138954 176600 139574 212058
rect 145794 219454 146414 239592
rect 145794 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 146414 219454
rect 145794 219134 146414 219218
rect 145794 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 146414 219134
rect 145794 183454 146414 218898
rect 145794 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 146414 183454
rect 145794 183134 146414 183218
rect 145794 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 146414 183134
rect 145794 176600 146414 182898
rect 149514 223174 150134 239592
rect 149514 222938 149546 223174
rect 149782 222938 149866 223174
rect 150102 222938 150134 223174
rect 149514 222854 150134 222938
rect 149514 222618 149546 222854
rect 149782 222618 149866 222854
rect 150102 222618 150134 222854
rect 149514 187174 150134 222618
rect 149514 186938 149546 187174
rect 149782 186938 149866 187174
rect 150102 186938 150134 187174
rect 149514 186854 150134 186938
rect 149514 186618 149546 186854
rect 149782 186618 149866 186854
rect 150102 186618 150134 186854
rect 148179 176764 148245 176765
rect 148179 176700 148180 176764
rect 148244 176700 148245 176764
rect 148179 176699 148245 176700
rect 135667 175676 135733 175677
rect 135667 175612 135668 175676
rect 135732 175612 135733 175676
rect 135667 175611 135733 175612
rect 133094 175070 133196 175130
rect 130688 174494 130748 175070
rect 132048 174494 132108 175070
rect 133136 174494 133196 175070
rect 134360 175070 134442 175130
rect 135670 175130 135730 175611
rect 148182 175130 148242 176699
rect 149514 176600 150134 186618
rect 153234 226894 153854 239592
rect 154070 235925 154130 442171
rect 155726 345133 155786 504323
rect 156954 482614 157574 518058
rect 156954 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 157574 482614
rect 156954 482294 157574 482378
rect 156954 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 157574 482294
rect 156954 446614 157574 482058
rect 156954 446378 156986 446614
rect 157222 446378 157306 446614
rect 157542 446378 157574 446614
rect 156954 446294 157574 446378
rect 156954 446058 156986 446294
rect 157222 446058 157306 446294
rect 157542 446058 157574 446294
rect 156954 410614 157574 446058
rect 156954 410378 156986 410614
rect 157222 410378 157306 410614
rect 157542 410378 157574 410614
rect 156954 410294 157574 410378
rect 156954 410058 156986 410294
rect 157222 410058 157306 410294
rect 157542 410058 157574 410294
rect 156954 374614 157574 410058
rect 156954 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 157574 374614
rect 156954 374294 157574 374378
rect 156954 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 157574 374294
rect 155723 345132 155789 345133
rect 155723 345068 155724 345132
rect 155788 345068 155789 345132
rect 155723 345067 155789 345068
rect 154619 334660 154685 334661
rect 154619 334596 154620 334660
rect 154684 334596 154685 334660
rect 154619 334595 154685 334596
rect 154622 242045 154682 334595
rect 155726 331941 155786 345067
rect 156643 339420 156709 339421
rect 156643 339356 156644 339420
rect 156708 339356 156709 339420
rect 156643 339355 156709 339356
rect 155723 331940 155789 331941
rect 155723 331876 155724 331940
rect 155788 331876 155789 331940
rect 155723 331875 155789 331876
rect 156646 306390 156706 339355
rect 156954 338614 157574 374058
rect 157931 367708 157997 367709
rect 157931 367644 157932 367708
rect 157996 367644 157997 367708
rect 157931 367643 157997 367644
rect 157934 364350 157994 367643
rect 157750 364290 157994 364350
rect 157750 360093 157810 364290
rect 157747 360092 157813 360093
rect 157747 360028 157748 360092
rect 157812 360028 157813 360092
rect 157747 360027 157813 360028
rect 156954 338378 156986 338614
rect 157222 338378 157306 338614
rect 157542 338378 157574 338614
rect 156954 338294 157574 338378
rect 156954 338058 156986 338294
rect 157222 338058 157306 338294
rect 157542 338058 157574 338294
rect 156954 331592 157574 338058
rect 156827 331396 156893 331397
rect 156827 331332 156828 331396
rect 156892 331332 156893 331396
rect 156827 331331 156893 331332
rect 156830 326365 156890 331331
rect 156827 326364 156893 326365
rect 156827 326300 156828 326364
rect 156892 326300 156893 326364
rect 156827 326299 156893 326300
rect 156646 306330 156890 306390
rect 156830 289237 156890 306330
rect 157011 296308 157077 296309
rect 157011 296244 157012 296308
rect 157076 296244 157077 296308
rect 157011 296243 157077 296244
rect 156827 289236 156893 289237
rect 156827 289172 156828 289236
rect 156892 289172 156893 289236
rect 156827 289171 156893 289172
rect 157014 277410 157074 296243
rect 157750 277813 157810 360027
rect 159955 356692 160021 356693
rect 159955 356628 159956 356692
rect 160020 356628 160021 356692
rect 159955 356627 160021 356628
rect 159403 341596 159469 341597
rect 159403 341532 159404 341596
rect 159468 341532 159469 341596
rect 159403 341531 159469 341532
rect 158483 331396 158549 331397
rect 158483 331332 158484 331396
rect 158548 331332 158549 331396
rect 158483 331331 158549 331332
rect 158486 300117 158546 331331
rect 159219 309772 159285 309773
rect 159219 309708 159220 309772
rect 159284 309708 159285 309772
rect 159219 309707 159285 309708
rect 157931 300116 157997 300117
rect 157931 300052 157932 300116
rect 157996 300052 157997 300116
rect 157931 300051 157997 300052
rect 158483 300116 158549 300117
rect 158483 300052 158484 300116
rect 158548 300052 158549 300116
rect 158483 300051 158549 300052
rect 157747 277812 157813 277813
rect 157747 277748 157748 277812
rect 157812 277748 157813 277812
rect 157747 277747 157813 277748
rect 156462 277350 157074 277410
rect 154619 242044 154685 242045
rect 154619 241980 154620 242044
rect 154684 241980 154685 242044
rect 154619 241979 154685 241980
rect 156462 241501 156522 277350
rect 156827 245036 156893 245037
rect 156827 244972 156828 245036
rect 156892 244972 156893 245036
rect 156827 244971 156893 244972
rect 156830 241770 156890 244971
rect 157934 242181 157994 300051
rect 158115 245852 158181 245853
rect 158115 245788 158116 245852
rect 158180 245788 158181 245852
rect 158115 245787 158181 245788
rect 157931 242180 157997 242181
rect 157931 242116 157932 242180
rect 157996 242116 157997 242180
rect 157931 242115 157997 242116
rect 156646 241710 156890 241770
rect 156459 241500 156525 241501
rect 156459 241436 156460 241500
rect 156524 241436 156525 241500
rect 156459 241435 156525 241436
rect 154067 235924 154133 235925
rect 154067 235860 154068 235924
rect 154132 235860 154133 235924
rect 154067 235859 154133 235860
rect 156646 231845 156706 241710
rect 156643 231844 156709 231845
rect 156643 231780 156644 231844
rect 156708 231780 156709 231844
rect 156643 231779 156709 231780
rect 153234 226658 153266 226894
rect 153502 226658 153586 226894
rect 153822 226658 153854 226894
rect 153234 226574 153854 226658
rect 153234 226338 153266 226574
rect 153502 226338 153586 226574
rect 153822 226338 153854 226574
rect 153234 190894 153854 226338
rect 153234 190658 153266 190894
rect 153502 190658 153586 190894
rect 153822 190658 153854 190894
rect 153234 190574 153854 190658
rect 153234 190338 153266 190574
rect 153502 190338 153586 190574
rect 153822 190338 153854 190574
rect 153234 176600 153854 190338
rect 156954 230614 157574 239592
rect 158118 235245 158178 245787
rect 158115 235244 158181 235245
rect 158115 235180 158116 235244
rect 158180 235180 158181 235244
rect 158115 235179 158181 235180
rect 159222 233885 159282 309707
rect 159406 303789 159466 341531
rect 159958 309093 160018 356627
rect 160694 311949 160754 539819
rect 160875 436116 160941 436117
rect 160875 436052 160876 436116
rect 160940 436052 160941 436116
rect 160875 436051 160941 436052
rect 160691 311948 160757 311949
rect 160691 311884 160692 311948
rect 160756 311884 160757 311948
rect 160691 311883 160757 311884
rect 159955 309092 160021 309093
rect 159955 309028 159956 309092
rect 160020 309028 160021 309092
rect 159955 309027 160021 309028
rect 159958 308413 160018 309027
rect 159955 308412 160021 308413
rect 159955 308348 159956 308412
rect 160020 308348 160021 308412
rect 159955 308347 160021 308348
rect 159403 303788 159469 303789
rect 159403 303724 159404 303788
rect 159468 303724 159469 303788
rect 159403 303723 159469 303724
rect 159406 247621 159466 303723
rect 160878 288693 160938 436051
rect 160875 288692 160941 288693
rect 160875 288628 160876 288692
rect 160940 288628 160941 288692
rect 160875 288627 160941 288628
rect 160878 277410 160938 288627
rect 160694 277350 160938 277410
rect 160694 276725 160754 277350
rect 160691 276724 160757 276725
rect 160691 276660 160692 276724
rect 160756 276660 160757 276724
rect 160691 276659 160757 276660
rect 160139 269380 160205 269381
rect 160139 269316 160140 269380
rect 160204 269316 160205 269380
rect 160139 269315 160205 269316
rect 160142 251157 160202 269315
rect 161982 259589 162042 543899
rect 163794 525454 164414 560898
rect 163794 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 164414 525454
rect 163794 525134 164414 525218
rect 163794 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 164414 525134
rect 163794 489454 164414 524898
rect 163794 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 164414 489454
rect 163794 489134 164414 489218
rect 163794 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 164414 489134
rect 163794 453454 164414 488898
rect 163794 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 164414 453454
rect 163794 453134 164414 453218
rect 163794 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 164414 453134
rect 163794 417454 164414 452898
rect 163794 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 164414 417454
rect 163794 417134 164414 417218
rect 163794 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 164414 417134
rect 163794 381454 164414 416898
rect 167514 673174 168134 707162
rect 167514 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 168134 673174
rect 167514 672854 168134 672938
rect 167514 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 168134 672854
rect 167514 637174 168134 672618
rect 167514 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 168134 637174
rect 167514 636854 168134 636938
rect 167514 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 168134 636854
rect 167514 601174 168134 636618
rect 167514 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 168134 601174
rect 167514 600854 168134 600938
rect 167514 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 168134 600854
rect 167514 565174 168134 600618
rect 167514 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 168134 565174
rect 167514 564854 168134 564938
rect 167514 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 168134 564854
rect 167514 529174 168134 564618
rect 171234 676894 171854 709082
rect 171234 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 171854 676894
rect 171234 676574 171854 676658
rect 171234 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 171854 676574
rect 171234 640894 171854 676338
rect 171234 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 171854 640894
rect 171234 640574 171854 640658
rect 171234 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 171854 640574
rect 171234 604894 171854 640338
rect 171234 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 171854 604894
rect 171234 604574 171854 604658
rect 171234 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 171854 604574
rect 171234 568894 171854 604338
rect 171234 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 171854 568894
rect 171234 568574 171854 568658
rect 171234 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 171854 568574
rect 170259 552124 170325 552125
rect 170259 552060 170260 552124
rect 170324 552060 170325 552124
rect 170259 552059 170325 552060
rect 167514 528938 167546 529174
rect 167782 528938 167866 529174
rect 168102 528938 168134 529174
rect 167514 528854 168134 528938
rect 167514 528618 167546 528854
rect 167782 528618 167866 528854
rect 168102 528618 168134 528854
rect 167514 493174 168134 528618
rect 167514 492938 167546 493174
rect 167782 492938 167866 493174
rect 168102 492938 168134 493174
rect 167514 492854 168134 492938
rect 167514 492618 167546 492854
rect 167782 492618 167866 492854
rect 168102 492618 168134 492854
rect 167514 457174 168134 492618
rect 167514 456938 167546 457174
rect 167782 456938 167866 457174
rect 168102 456938 168134 457174
rect 167514 456854 168134 456938
rect 167514 456618 167546 456854
rect 167782 456618 167866 456854
rect 168102 456618 168134 456854
rect 167514 421174 168134 456618
rect 167514 420938 167546 421174
rect 167782 420938 167866 421174
rect 168102 420938 168134 421174
rect 167514 420854 168134 420938
rect 167514 420618 167546 420854
rect 167782 420618 167866 420854
rect 168102 420618 168134 420854
rect 165659 407828 165725 407829
rect 165659 407764 165660 407828
rect 165724 407764 165725 407828
rect 165659 407763 165725 407764
rect 163794 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 164414 381454
rect 163794 381134 164414 381218
rect 163794 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 164414 381134
rect 163794 345454 164414 380898
rect 163794 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 164414 345454
rect 163794 345134 164414 345218
rect 163794 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 164414 345134
rect 163794 309454 164414 344898
rect 163794 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 164414 309454
rect 163794 309134 164414 309218
rect 163794 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 164414 309134
rect 163451 293180 163517 293181
rect 163451 293116 163452 293180
rect 163516 293116 163517 293180
rect 163451 293115 163517 293116
rect 162163 260132 162229 260133
rect 162163 260068 162164 260132
rect 162228 260068 162229 260132
rect 162163 260067 162229 260068
rect 161979 259588 162045 259589
rect 161979 259524 161980 259588
rect 162044 259524 162045 259588
rect 161979 259523 162045 259524
rect 160139 251156 160205 251157
rect 160139 251092 160140 251156
rect 160204 251092 160205 251156
rect 160139 251091 160205 251092
rect 159403 247620 159469 247621
rect 159403 247556 159404 247620
rect 159468 247556 159469 247620
rect 159403 247555 159469 247556
rect 160875 247620 160941 247621
rect 160875 247556 160876 247620
rect 160940 247556 160941 247620
rect 160875 247555 160941 247556
rect 159219 233884 159285 233885
rect 159219 233820 159220 233884
rect 159284 233820 159285 233884
rect 159219 233819 159285 233820
rect 156954 230378 156986 230614
rect 157222 230378 157306 230614
rect 157542 230378 157574 230614
rect 156954 230294 157574 230378
rect 156954 230058 156986 230294
rect 157222 230058 157306 230294
rect 157542 230058 157574 230294
rect 156954 194614 157574 230058
rect 160878 224637 160938 247555
rect 160875 224636 160941 224637
rect 160875 224572 160876 224636
rect 160940 224572 160941 224636
rect 160875 224571 160941 224572
rect 162166 210901 162226 260067
rect 162163 210900 162229 210901
rect 162163 210836 162164 210900
rect 162228 210836 162229 210900
rect 162163 210835 162229 210836
rect 163454 210765 163514 293115
rect 163794 273454 164414 308898
rect 163794 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 164414 273454
rect 163794 273134 164414 273218
rect 163794 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 164414 273134
rect 163794 237454 164414 272898
rect 163794 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 164414 237454
rect 163794 237134 164414 237218
rect 163794 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 164414 237134
rect 163451 210764 163517 210765
rect 163451 210700 163452 210764
rect 163516 210700 163517 210764
rect 163451 210699 163517 210700
rect 156954 194378 156986 194614
rect 157222 194378 157306 194614
rect 157542 194378 157574 194614
rect 156954 194294 157574 194378
rect 156954 194058 156986 194294
rect 157222 194058 157306 194294
rect 157542 194058 157574 194294
rect 156954 176600 157574 194058
rect 163794 201454 164414 236898
rect 163794 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 164414 201454
rect 163794 201134 164414 201218
rect 163794 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 164414 201134
rect 158851 176764 158917 176765
rect 158851 176700 158852 176764
rect 158916 176700 158917 176764
rect 158851 176699 158917 176700
rect 158854 175130 158914 176699
rect 163794 176600 164414 200898
rect 135670 175070 135780 175130
rect 148182 175070 148292 175130
rect 134360 174494 134420 175070
rect 135720 174494 135780 175070
rect 148232 174494 148292 175070
rect 158840 175070 158914 175130
rect 158840 174494 158900 175070
rect 69072 165454 69420 165486
rect 69072 165218 69128 165454
rect 69364 165218 69420 165454
rect 69072 165134 69420 165218
rect 69072 164898 69128 165134
rect 69364 164898 69420 165134
rect 69072 164866 69420 164898
rect 164136 165454 164484 165486
rect 164136 165218 164192 165454
rect 164428 165218 164484 165454
rect 164136 165134 164484 165218
rect 164136 164898 164192 165134
rect 164428 164898 164484 165134
rect 164136 164866 164484 164898
rect 69752 147454 70100 147486
rect 69752 147218 69808 147454
rect 70044 147218 70100 147454
rect 69752 147134 70100 147218
rect 69752 146898 69808 147134
rect 70044 146898 70100 147134
rect 69752 146866 70100 146898
rect 163456 147454 163804 147486
rect 163456 147218 163512 147454
rect 163748 147218 163804 147454
rect 163456 147134 163804 147218
rect 163456 146898 163512 147134
rect 163748 146898 163804 147134
rect 163456 146866 163804 146898
rect 69072 129454 69420 129486
rect 69072 129218 69128 129454
rect 69364 129218 69420 129454
rect 69072 129134 69420 129218
rect 69072 128898 69128 129134
rect 69364 128898 69420 129134
rect 69072 128866 69420 128898
rect 164136 129454 164484 129486
rect 164136 129218 164192 129454
rect 164428 129218 164484 129454
rect 164136 129134 164484 129218
rect 164136 128898 164192 129134
rect 164428 128898 164484 129134
rect 164136 128866 164484 128898
rect 69752 111454 70100 111486
rect 69752 111218 69808 111454
rect 70044 111218 70100 111454
rect 69752 111134 70100 111218
rect 69752 110898 69808 111134
rect 70044 110898 70100 111134
rect 69752 110866 70100 110898
rect 163456 111454 163804 111486
rect 163456 111218 163512 111454
rect 163748 111218 163804 111454
rect 163456 111134 163804 111218
rect 163456 110898 163512 111134
rect 163748 110898 163804 111134
rect 163456 110866 163804 110898
rect 74656 94890 74716 95200
rect 84312 94890 84372 95200
rect 85536 94890 85596 95200
rect 86624 94890 86684 95200
rect 87984 94890 88044 95200
rect 88936 94890 88996 95200
rect 74656 94830 74826 94890
rect 84312 94830 84394 94890
rect 85536 94830 85866 94890
rect 86624 94830 86786 94890
rect 87984 94830 88074 94890
rect 73794 75454 74414 93100
rect 74766 91221 74826 94830
rect 74763 91220 74829 91221
rect 74763 91156 74764 91220
rect 74828 91156 74829 91220
rect 74763 91155 74829 91156
rect 73794 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 74414 75454
rect 73794 75134 74414 75218
rect 73794 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 74414 75134
rect 73794 39454 74414 74898
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 67771 33964 67837 33965
rect 67771 33900 67772 33964
rect 67836 33900 67837 33964
rect 67771 33899 67837 33900
rect 66954 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 67574 32614
rect 66954 32294 67574 32378
rect 66954 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 67574 32294
rect 48954 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 49574 -6106
rect 48954 -6426 49574 -6342
rect 48954 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 49574 -6426
rect 48954 -7654 49574 -6662
rect 66954 -7066 67574 32058
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -1894 74414 -902
rect 77514 79174 78134 93100
rect 77514 78938 77546 79174
rect 77782 78938 77866 79174
rect 78102 78938 78134 79174
rect 77514 78854 78134 78938
rect 77514 78618 77546 78854
rect 77782 78618 77866 78854
rect 78102 78618 78134 78854
rect 77514 43174 78134 78618
rect 77514 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 78134 43174
rect 77514 42854 78134 42938
rect 77514 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 78134 42854
rect 77514 7174 78134 42618
rect 77514 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 78134 7174
rect 77514 6854 78134 6938
rect 77514 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 78134 6854
rect 77514 -2266 78134 6618
rect 77514 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 78134 -2266
rect 77514 -2586 78134 -2502
rect 77514 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 78134 -2586
rect 77514 -3814 78134 -2822
rect 81234 82894 81854 93100
rect 84334 91221 84394 94830
rect 84331 91220 84397 91221
rect 84331 91156 84332 91220
rect 84396 91156 84397 91220
rect 84331 91155 84397 91156
rect 81234 82658 81266 82894
rect 81502 82658 81586 82894
rect 81822 82658 81854 82894
rect 81234 82574 81854 82658
rect 81234 82338 81266 82574
rect 81502 82338 81586 82574
rect 81822 82338 81854 82574
rect 81234 46894 81854 82338
rect 81234 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 81854 46894
rect 81234 46574 81854 46658
rect 81234 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 81854 46574
rect 81234 10894 81854 46338
rect 81234 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 81854 10894
rect 81234 10574 81854 10658
rect 81234 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 81854 10574
rect 81234 -4186 81854 10338
rect 81234 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 81854 -4186
rect 81234 -4506 81854 -4422
rect 81234 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 81854 -4506
rect 81234 -5734 81854 -4742
rect 84954 86614 85574 93100
rect 85806 92309 85866 94830
rect 86726 92445 86786 94830
rect 86723 92444 86789 92445
rect 86723 92380 86724 92444
rect 86788 92380 86789 92444
rect 86723 92379 86789 92380
rect 85803 92308 85869 92309
rect 85803 92244 85804 92308
rect 85868 92244 85869 92308
rect 85803 92243 85869 92244
rect 88014 91221 88074 94830
rect 88934 94830 88996 94890
rect 90160 94890 90220 95200
rect 91384 94890 91444 95200
rect 90160 94830 90282 94890
rect 88934 92445 88994 94830
rect 88931 92444 88997 92445
rect 88931 92380 88932 92444
rect 88996 92380 88997 92444
rect 88931 92379 88997 92380
rect 90222 91221 90282 94830
rect 91326 94830 91444 94890
rect 92472 94890 92532 95200
rect 93832 94890 93892 95200
rect 94920 94890 94980 95200
rect 96008 94890 96068 95200
rect 96688 94890 96748 95200
rect 92472 94830 92674 94890
rect 93832 94830 93962 94890
rect 94920 94830 95066 94890
rect 96008 94830 96354 94890
rect 91326 93941 91386 94830
rect 91323 93940 91389 93941
rect 91323 93876 91324 93940
rect 91388 93876 91389 93940
rect 91323 93875 91389 93876
rect 88011 91220 88077 91221
rect 88011 91156 88012 91220
rect 88076 91156 88077 91220
rect 88011 91155 88077 91156
rect 90219 91220 90285 91221
rect 90219 91156 90220 91220
rect 90284 91156 90285 91220
rect 90219 91155 90285 91156
rect 84954 86378 84986 86614
rect 85222 86378 85306 86614
rect 85542 86378 85574 86614
rect 84954 86294 85574 86378
rect 84954 86058 84986 86294
rect 85222 86058 85306 86294
rect 85542 86058 85574 86294
rect 84954 50614 85574 86058
rect 84954 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 85574 50614
rect 84954 50294 85574 50378
rect 84954 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 85574 50294
rect 84954 14614 85574 50058
rect 84954 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 85574 14614
rect 84954 14294 85574 14378
rect 84954 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 85574 14294
rect 66954 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 67574 -7066
rect 66954 -7386 67574 -7302
rect 66954 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 67574 -7386
rect 66954 -7654 67574 -7622
rect 84954 -6106 85574 14058
rect 91794 57454 92414 93100
rect 92614 91221 92674 94830
rect 93902 91221 93962 94830
rect 95006 93533 95066 94830
rect 95003 93532 95069 93533
rect 95003 93468 95004 93532
rect 95068 93468 95069 93532
rect 95003 93467 95069 93468
rect 92611 91220 92677 91221
rect 92611 91156 92612 91220
rect 92676 91156 92677 91220
rect 92611 91155 92677 91156
rect 93899 91220 93965 91221
rect 93899 91156 93900 91220
rect 93964 91156 93965 91220
rect 93899 91155 93965 91156
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -1306 92414 20898
rect 91794 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 92414 -1306
rect 91794 -1626 92414 -1542
rect 91794 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 92414 -1626
rect 91794 -1894 92414 -1862
rect 95514 61174 96134 93100
rect 96294 91221 96354 94830
rect 96662 94830 96748 94890
rect 97096 94890 97156 95200
rect 98048 94890 98108 95200
rect 98456 94890 98516 95200
rect 99136 94890 99196 95200
rect 97096 94830 97274 94890
rect 98048 94830 98194 94890
rect 98456 94830 98562 94890
rect 96662 91357 96722 94830
rect 96659 91356 96725 91357
rect 96659 91292 96660 91356
rect 96724 91292 96725 91356
rect 96659 91291 96725 91292
rect 97214 91221 97274 94830
rect 98134 91357 98194 94830
rect 98131 91356 98197 91357
rect 98131 91292 98132 91356
rect 98196 91292 98197 91356
rect 98131 91291 98197 91292
rect 98502 91221 98562 94830
rect 99054 94830 99196 94890
rect 99544 94890 99604 95200
rect 100632 94890 100692 95200
rect 99544 94830 99666 94890
rect 99054 91765 99114 94830
rect 99606 94077 99666 94830
rect 100526 94830 100692 94890
rect 100768 94890 100828 95200
rect 101856 94890 101916 95200
rect 100768 94830 100954 94890
rect 99603 94076 99669 94077
rect 99603 94012 99604 94076
rect 99668 94012 99669 94076
rect 99603 94011 99669 94012
rect 99051 91764 99117 91765
rect 99051 91700 99052 91764
rect 99116 91700 99117 91764
rect 99051 91699 99117 91700
rect 96291 91220 96357 91221
rect 96291 91156 96292 91220
rect 96356 91156 96357 91220
rect 96291 91155 96357 91156
rect 97211 91220 97277 91221
rect 97211 91156 97212 91220
rect 97276 91156 97277 91220
rect 97211 91155 97277 91156
rect 98499 91220 98565 91221
rect 98499 91156 98500 91220
rect 98564 91156 98565 91220
rect 98499 91155 98565 91156
rect 95514 60938 95546 61174
rect 95782 60938 95866 61174
rect 96102 60938 96134 61174
rect 95514 60854 96134 60938
rect 95514 60618 95546 60854
rect 95782 60618 95866 60854
rect 96102 60618 96134 60854
rect 95514 25174 96134 60618
rect 95514 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 96134 25174
rect 95514 24854 96134 24938
rect 95514 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 96134 24854
rect 95514 -3226 96134 24618
rect 95514 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 96134 -3226
rect 95514 -3546 96134 -3462
rect 95514 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 96134 -3546
rect 95514 -3814 96134 -3782
rect 99234 64894 99854 93100
rect 100526 91221 100586 94830
rect 100894 91357 100954 94830
rect 101814 94830 101916 94890
rect 101992 94890 102052 95200
rect 102944 94890 103004 95200
rect 101992 94830 102058 94890
rect 100891 91356 100957 91357
rect 100891 91292 100892 91356
rect 100956 91292 100957 91356
rect 100891 91291 100957 91292
rect 101814 91221 101874 94830
rect 101998 92445 102058 94830
rect 102734 94830 103004 94890
rect 103216 94890 103276 95200
rect 104304 94890 104364 95200
rect 103216 94830 103346 94890
rect 101995 92444 102061 92445
rect 101995 92380 101996 92444
rect 102060 92380 102061 92444
rect 101995 92379 102061 92380
rect 102734 91221 102794 94830
rect 103286 93261 103346 94830
rect 104206 94830 104364 94890
rect 104440 94890 104500 95200
rect 105392 94890 105452 95200
rect 105664 94890 105724 95200
rect 106480 94890 106540 95200
rect 104440 94830 104634 94890
rect 105392 94830 105554 94890
rect 105664 94830 105738 94890
rect 103283 93260 103349 93261
rect 103283 93196 103284 93260
rect 103348 93196 103349 93260
rect 103283 93195 103349 93196
rect 100523 91220 100589 91221
rect 100523 91156 100524 91220
rect 100588 91156 100589 91220
rect 100523 91155 100589 91156
rect 101811 91220 101877 91221
rect 101811 91156 101812 91220
rect 101876 91156 101877 91220
rect 101811 91155 101877 91156
rect 102731 91220 102797 91221
rect 102731 91156 102732 91220
rect 102796 91156 102797 91220
rect 102731 91155 102797 91156
rect 99234 64658 99266 64894
rect 99502 64658 99586 64894
rect 99822 64658 99854 64894
rect 99234 64574 99854 64658
rect 99234 64338 99266 64574
rect 99502 64338 99586 64574
rect 99822 64338 99854 64574
rect 99234 28894 99854 64338
rect 99234 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 99854 28894
rect 99234 28574 99854 28658
rect 99234 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 99854 28574
rect 99234 -5146 99854 28338
rect 99234 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 99854 -5146
rect 99234 -5466 99854 -5382
rect 99234 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 99854 -5466
rect 99234 -5734 99854 -5702
rect 102954 68614 103574 93100
rect 104206 91221 104266 94830
rect 104574 91221 104634 94830
rect 105494 91221 105554 94830
rect 105678 91221 105738 94830
rect 106414 94830 106540 94890
rect 106616 94890 106676 95200
rect 106616 94830 106842 94890
rect 106414 91629 106474 94830
rect 106782 91629 106842 94830
rect 107704 94757 107764 95200
rect 108112 94890 108172 95200
rect 108070 94830 108172 94890
rect 109064 94890 109124 95200
rect 109472 94890 109532 95200
rect 110152 94890 110212 95200
rect 110696 94890 110756 95200
rect 111240 94890 111300 95200
rect 109064 94830 109234 94890
rect 109472 94830 109602 94890
rect 110152 94830 110338 94890
rect 107701 94756 107767 94757
rect 107701 94692 107702 94756
rect 107766 94692 107767 94756
rect 107701 94691 107767 94692
rect 106411 91628 106477 91629
rect 106411 91564 106412 91628
rect 106476 91564 106477 91628
rect 106411 91563 106477 91564
rect 106779 91628 106845 91629
rect 106779 91564 106780 91628
rect 106844 91564 106845 91628
rect 106779 91563 106845 91564
rect 108070 91221 108130 94830
rect 109174 91357 109234 94830
rect 109171 91356 109237 91357
rect 109171 91292 109172 91356
rect 109236 91292 109237 91356
rect 109171 91291 109237 91292
rect 109542 91221 109602 94830
rect 110278 93261 110338 94830
rect 110646 94830 110756 94890
rect 111198 94830 111300 94890
rect 111920 94890 111980 95200
rect 112328 94890 112388 95200
rect 111920 94830 111994 94890
rect 110275 93260 110341 93261
rect 110275 93196 110276 93260
rect 110340 93196 110341 93260
rect 110275 93195 110341 93196
rect 104203 91220 104269 91221
rect 104203 91156 104204 91220
rect 104268 91156 104269 91220
rect 104203 91155 104269 91156
rect 104571 91220 104637 91221
rect 104571 91156 104572 91220
rect 104636 91156 104637 91220
rect 104571 91155 104637 91156
rect 105491 91220 105557 91221
rect 105491 91156 105492 91220
rect 105556 91156 105557 91220
rect 105491 91155 105557 91156
rect 105675 91220 105741 91221
rect 105675 91156 105676 91220
rect 105740 91156 105741 91220
rect 105675 91155 105741 91156
rect 108067 91220 108133 91221
rect 108067 91156 108068 91220
rect 108132 91156 108133 91220
rect 108067 91155 108133 91156
rect 109539 91220 109605 91221
rect 109539 91156 109540 91220
rect 109604 91156 109605 91220
rect 109539 91155 109605 91156
rect 102954 68378 102986 68614
rect 103222 68378 103306 68614
rect 103542 68378 103574 68614
rect 102954 68294 103574 68378
rect 102954 68058 102986 68294
rect 103222 68058 103306 68294
rect 103542 68058 103574 68294
rect 102954 32614 103574 68058
rect 102954 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 103574 32614
rect 102954 32294 103574 32378
rect 102954 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 103574 32294
rect 84954 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 85574 -6106
rect 84954 -6426 85574 -6342
rect 84954 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 85574 -6426
rect 84954 -7654 85574 -6662
rect 102954 -7066 103574 32058
rect 109794 75454 110414 93100
rect 110646 91221 110706 94830
rect 111198 91357 111258 94830
rect 111195 91356 111261 91357
rect 111195 91292 111196 91356
rect 111260 91292 111261 91356
rect 111195 91291 111261 91292
rect 111934 91221 111994 94830
rect 112302 94830 112388 94890
rect 113144 94890 113204 95200
rect 113688 94890 113748 95200
rect 114368 94890 114428 95200
rect 113144 94830 113282 94890
rect 113688 94830 114202 94890
rect 112302 92445 112362 94830
rect 112299 92444 112365 92445
rect 112299 92380 112300 92444
rect 112364 92380 112365 92444
rect 112299 92379 112365 92380
rect 113222 91221 113282 94830
rect 114142 93530 114202 94830
rect 114326 94830 114428 94890
rect 114776 94890 114836 95200
rect 115456 94890 115516 95200
rect 115864 94890 115924 95200
rect 114776 94830 114938 94890
rect 114326 93805 114386 94830
rect 114323 93804 114389 93805
rect 114323 93740 114324 93804
rect 114388 93740 114389 93804
rect 114323 93739 114389 93740
rect 114142 93470 114386 93530
rect 110643 91220 110709 91221
rect 110643 91156 110644 91220
rect 110708 91156 110709 91220
rect 110643 91155 110709 91156
rect 111931 91220 111997 91221
rect 111931 91156 111932 91220
rect 111996 91156 111997 91220
rect 111931 91155 111997 91156
rect 113219 91220 113285 91221
rect 113219 91156 113220 91220
rect 113284 91156 113285 91220
rect 113219 91155 113285 91156
rect 109794 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 110414 75454
rect 109794 75134 110414 75218
rect 109794 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 110414 75134
rect 109794 39454 110414 74898
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -1894 110414 -902
rect 113514 79174 114134 93100
rect 114326 91357 114386 93470
rect 114323 91356 114389 91357
rect 114323 91292 114324 91356
rect 114388 91292 114389 91356
rect 114323 91291 114389 91292
rect 114878 91221 114938 94830
rect 115430 94830 115516 94890
rect 115798 94830 115924 94890
rect 116680 94890 116740 95200
rect 116680 94830 116778 94890
rect 115430 92173 115490 94830
rect 115798 93533 115858 94830
rect 115795 93532 115861 93533
rect 115795 93468 115796 93532
rect 115860 93468 115861 93532
rect 115795 93467 115861 93468
rect 115427 92172 115493 92173
rect 115427 92108 115428 92172
rect 115492 92108 115493 92172
rect 115427 92107 115493 92108
rect 116718 91221 116778 94830
rect 117088 94757 117148 95200
rect 117904 94890 117964 95200
rect 118176 94890 118236 95200
rect 119400 94890 119460 95200
rect 117904 94830 118066 94890
rect 118176 94830 118250 94890
rect 117085 94756 117151 94757
rect 117085 94692 117086 94756
rect 117150 94692 117151 94756
rect 117085 94691 117151 94692
rect 114875 91220 114941 91221
rect 114875 91156 114876 91220
rect 114940 91156 114941 91220
rect 114875 91155 114941 91156
rect 116715 91220 116781 91221
rect 116715 91156 116716 91220
rect 116780 91156 116781 91220
rect 116715 91155 116781 91156
rect 113514 78938 113546 79174
rect 113782 78938 113866 79174
rect 114102 78938 114134 79174
rect 113514 78854 114134 78938
rect 113514 78618 113546 78854
rect 113782 78618 113866 78854
rect 114102 78618 114134 78854
rect 113514 43174 114134 78618
rect 113514 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 114134 43174
rect 113514 42854 114134 42938
rect 113514 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 114134 42854
rect 113514 7174 114134 42618
rect 113514 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 114134 7174
rect 113514 6854 114134 6938
rect 113514 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 114134 6854
rect 113514 -2266 114134 6618
rect 113514 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 114134 -2266
rect 113514 -2586 114134 -2502
rect 113514 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 114134 -2586
rect 113514 -3814 114134 -2822
rect 117234 82894 117854 93100
rect 118006 91221 118066 94830
rect 118190 91221 118250 94830
rect 119294 94830 119460 94890
rect 119536 94890 119596 95200
rect 120216 94890 120276 95200
rect 120624 94890 120684 95200
rect 121712 94890 121772 95200
rect 119536 94830 119722 94890
rect 119294 91221 119354 94830
rect 119662 91765 119722 94830
rect 120214 94830 120276 94890
rect 120582 94830 120684 94890
rect 121686 94830 121772 94890
rect 121984 94890 122044 95200
rect 122800 94890 122860 95200
rect 123208 94890 123268 95200
rect 121984 94830 122114 94890
rect 122800 94830 123034 94890
rect 119659 91764 119725 91765
rect 119659 91700 119660 91764
rect 119724 91700 119725 91764
rect 119659 91699 119725 91700
rect 120214 91221 120274 94830
rect 120582 91221 120642 94830
rect 118003 91220 118069 91221
rect 118003 91156 118004 91220
rect 118068 91156 118069 91220
rect 118003 91155 118069 91156
rect 118187 91220 118253 91221
rect 118187 91156 118188 91220
rect 118252 91156 118253 91220
rect 118187 91155 118253 91156
rect 119291 91220 119357 91221
rect 119291 91156 119292 91220
rect 119356 91156 119357 91220
rect 119291 91155 119357 91156
rect 120211 91220 120277 91221
rect 120211 91156 120212 91220
rect 120276 91156 120277 91220
rect 120211 91155 120277 91156
rect 120579 91220 120645 91221
rect 120579 91156 120580 91220
rect 120644 91156 120645 91220
rect 120579 91155 120645 91156
rect 117234 82658 117266 82894
rect 117502 82658 117586 82894
rect 117822 82658 117854 82894
rect 117234 82574 117854 82658
rect 117234 82338 117266 82574
rect 117502 82338 117586 82574
rect 117822 82338 117854 82574
rect 117234 46894 117854 82338
rect 117234 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 117854 46894
rect 117234 46574 117854 46658
rect 117234 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 117854 46574
rect 117234 10894 117854 46338
rect 117234 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 117854 10894
rect 117234 10574 117854 10658
rect 117234 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 117854 10574
rect 117234 -4186 117854 10338
rect 117234 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 117854 -4186
rect 117234 -4506 117854 -4422
rect 117234 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 117854 -4506
rect 117234 -5734 117854 -4742
rect 120954 86614 121574 93100
rect 121686 91765 121746 94830
rect 122054 92309 122114 94830
rect 122974 93870 123034 94830
rect 122606 93810 123034 93870
rect 123158 94830 123268 94890
rect 124024 94890 124084 95200
rect 124432 94890 124492 95200
rect 125384 94890 125444 95200
rect 124024 94830 124138 94890
rect 124432 94830 124506 94890
rect 122051 92308 122117 92309
rect 122051 92244 122052 92308
rect 122116 92244 122117 92308
rect 122051 92243 122117 92244
rect 121683 91764 121749 91765
rect 121683 91700 121684 91764
rect 121748 91700 121749 91764
rect 121683 91699 121749 91700
rect 122606 91490 122666 93810
rect 123158 91765 123218 94830
rect 123155 91764 123221 91765
rect 123155 91700 123156 91764
rect 123220 91700 123221 91764
rect 123155 91699 123221 91700
rect 122787 91492 122853 91493
rect 122787 91490 122788 91492
rect 122606 91430 122788 91490
rect 122787 91428 122788 91430
rect 122852 91428 122853 91492
rect 122787 91427 122853 91428
rect 124078 91221 124138 94830
rect 124446 91357 124506 94830
rect 125366 94830 125444 94890
rect 125656 94890 125716 95200
rect 126472 94890 126532 95200
rect 125656 94830 125794 94890
rect 124443 91356 124509 91357
rect 124443 91292 124444 91356
rect 124508 91292 124509 91356
rect 124443 91291 124509 91292
rect 125366 91221 125426 94830
rect 125734 91493 125794 94830
rect 126470 94830 126532 94890
rect 126608 94890 126668 95200
rect 128104 94890 128164 95200
rect 126608 94830 126714 94890
rect 125731 91492 125797 91493
rect 125731 91428 125732 91492
rect 125796 91428 125797 91492
rect 125731 91427 125797 91428
rect 126470 91221 126530 94830
rect 126654 91357 126714 94830
rect 127574 94830 128164 94890
rect 129328 94890 129388 95200
rect 130688 94890 130748 95200
rect 131912 94890 131972 95200
rect 133136 94890 133196 95200
rect 129328 94830 129474 94890
rect 130688 94830 130762 94890
rect 131912 94830 132418 94890
rect 126651 91356 126717 91357
rect 126651 91292 126652 91356
rect 126716 91292 126717 91356
rect 126651 91291 126717 91292
rect 127574 91221 127634 94830
rect 129414 93669 129474 94830
rect 129411 93668 129477 93669
rect 129411 93604 129412 93668
rect 129476 93604 129477 93668
rect 129411 93603 129477 93604
rect 124075 91220 124141 91221
rect 124075 91156 124076 91220
rect 124140 91156 124141 91220
rect 124075 91155 124141 91156
rect 125363 91220 125429 91221
rect 125363 91156 125364 91220
rect 125428 91156 125429 91220
rect 125363 91155 125429 91156
rect 126467 91220 126533 91221
rect 126467 91156 126468 91220
rect 126532 91156 126533 91220
rect 126467 91155 126533 91156
rect 127571 91220 127637 91221
rect 127571 91156 127572 91220
rect 127636 91156 127637 91220
rect 127571 91155 127637 91156
rect 120954 86378 120986 86614
rect 121222 86378 121306 86614
rect 121542 86378 121574 86614
rect 120954 86294 121574 86378
rect 120954 86058 120986 86294
rect 121222 86058 121306 86294
rect 121542 86058 121574 86294
rect 120954 50614 121574 86058
rect 120954 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 121574 50614
rect 120954 50294 121574 50378
rect 120954 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 121574 50294
rect 120954 14614 121574 50058
rect 120954 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 121574 14614
rect 120954 14294 121574 14378
rect 120954 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 121574 14294
rect 102954 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 103574 -7066
rect 102954 -7386 103574 -7302
rect 102954 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 103574 -7386
rect 102954 -7654 103574 -7622
rect 120954 -6106 121574 14058
rect 127794 57454 128414 93100
rect 130702 91221 130762 94830
rect 130699 91220 130765 91221
rect 130699 91156 130700 91220
rect 130764 91156 130765 91220
rect 130699 91155 130765 91156
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -1306 128414 20898
rect 127794 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 128414 -1306
rect 127794 -1626 128414 -1542
rect 127794 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 128414 -1626
rect 127794 -1894 128414 -1862
rect 131514 61174 132134 93100
rect 132358 92445 132418 94830
rect 133094 94830 133196 94890
rect 134360 94890 134420 95200
rect 135584 94890 135644 95200
rect 151496 94890 151556 95200
rect 134360 94830 134442 94890
rect 135584 94830 136098 94890
rect 132355 92444 132421 92445
rect 132355 92380 132356 92444
rect 132420 92380 132421 92444
rect 132355 92379 132421 92380
rect 133094 91221 133154 94830
rect 134382 92445 134442 94830
rect 134379 92444 134445 92445
rect 134379 92380 134380 92444
rect 134444 92380 134445 92444
rect 134379 92379 134445 92380
rect 133091 91220 133157 91221
rect 133091 91156 133092 91220
rect 133156 91156 133157 91220
rect 133091 91155 133157 91156
rect 131514 60938 131546 61174
rect 131782 60938 131866 61174
rect 132102 60938 132134 61174
rect 131514 60854 132134 60938
rect 131514 60618 131546 60854
rect 131782 60618 131866 60854
rect 132102 60618 132134 60854
rect 131514 25174 132134 60618
rect 131514 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 132134 25174
rect 131514 24854 132134 24938
rect 131514 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 132134 24854
rect 131514 -3226 132134 24618
rect 131514 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 132134 -3226
rect 131514 -3546 132134 -3462
rect 131514 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 132134 -3546
rect 131514 -3814 132134 -3782
rect 135234 64894 135854 93100
rect 136038 92445 136098 94830
rect 151310 94830 151556 94890
rect 136035 92444 136101 92445
rect 136035 92380 136036 92444
rect 136100 92380 136101 92444
rect 136035 92379 136101 92380
rect 135234 64658 135266 64894
rect 135502 64658 135586 64894
rect 135822 64658 135854 64894
rect 135234 64574 135854 64658
rect 135234 64338 135266 64574
rect 135502 64338 135586 64574
rect 135822 64338 135854 64574
rect 135234 28894 135854 64338
rect 135234 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 135854 28894
rect 135234 28574 135854 28658
rect 135234 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 135854 28574
rect 135234 -5146 135854 28338
rect 135234 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 135854 -5146
rect 135234 -5466 135854 -5382
rect 135234 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 135854 -5466
rect 135234 -5734 135854 -5702
rect 138954 68614 139574 93100
rect 138954 68378 138986 68614
rect 139222 68378 139306 68614
rect 139542 68378 139574 68614
rect 138954 68294 139574 68378
rect 138954 68058 138986 68294
rect 139222 68058 139306 68294
rect 139542 68058 139574 68294
rect 138954 32614 139574 68058
rect 138954 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 139574 32614
rect 138954 32294 139574 32378
rect 138954 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 139574 32294
rect 120954 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 121574 -6106
rect 120954 -6426 121574 -6342
rect 120954 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 121574 -6426
rect 120954 -7654 121574 -6662
rect 138954 -7066 139574 32058
rect 145794 75454 146414 93100
rect 145794 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 146414 75454
rect 145794 75134 146414 75218
rect 145794 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 146414 75134
rect 145794 39454 146414 74898
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -1894 146414 -902
rect 149514 79174 150134 93100
rect 151310 91357 151370 94830
rect 151491 94756 151557 94757
rect 151491 94692 151492 94756
rect 151556 94692 151557 94756
rect 151491 94691 151557 94692
rect 151307 91356 151373 91357
rect 151307 91292 151308 91356
rect 151372 91292 151373 91356
rect 151307 91291 151373 91292
rect 151494 91221 151554 94691
rect 151632 94210 151692 95200
rect 151768 94757 151828 95200
rect 151904 94890 151964 95200
rect 151904 94830 152106 94890
rect 151765 94756 151831 94757
rect 151765 94692 151766 94756
rect 151830 94692 151831 94756
rect 151765 94691 151831 94692
rect 151632 94150 151738 94210
rect 151678 91493 151738 94150
rect 151675 91492 151741 91493
rect 151675 91428 151676 91492
rect 151740 91428 151741 91492
rect 151675 91427 151741 91428
rect 152046 91221 152106 94830
rect 151491 91220 151557 91221
rect 151491 91156 151492 91220
rect 151556 91156 151557 91220
rect 151491 91155 151557 91156
rect 152043 91220 152109 91221
rect 152043 91156 152044 91220
rect 152108 91156 152109 91220
rect 152043 91155 152109 91156
rect 149514 78938 149546 79174
rect 149782 78938 149866 79174
rect 150102 78938 150134 79174
rect 149514 78854 150134 78938
rect 149514 78618 149546 78854
rect 149782 78618 149866 78854
rect 150102 78618 150134 78854
rect 149514 43174 150134 78618
rect 149514 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 150134 43174
rect 149514 42854 150134 42938
rect 149514 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 150134 42854
rect 149514 7174 150134 42618
rect 149514 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 150134 7174
rect 149514 6854 150134 6938
rect 149514 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 150134 6854
rect 149514 -2266 150134 6618
rect 149514 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 150134 -2266
rect 149514 -2586 150134 -2502
rect 149514 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 150134 -2586
rect 149514 -3814 150134 -2822
rect 153234 82894 153854 93100
rect 153234 82658 153266 82894
rect 153502 82658 153586 82894
rect 153822 82658 153854 82894
rect 153234 82574 153854 82658
rect 153234 82338 153266 82574
rect 153502 82338 153586 82574
rect 153822 82338 153854 82574
rect 153234 46894 153854 82338
rect 153234 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 153854 46894
rect 153234 46574 153854 46658
rect 153234 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 153854 46574
rect 153234 10894 153854 46338
rect 153234 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 153854 10894
rect 153234 10574 153854 10658
rect 153234 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 153854 10574
rect 153234 -4186 153854 10338
rect 153234 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 153854 -4186
rect 153234 -4506 153854 -4422
rect 153234 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 153854 -4506
rect 153234 -5734 153854 -4742
rect 156954 86614 157574 93100
rect 156954 86378 156986 86614
rect 157222 86378 157306 86614
rect 157542 86378 157574 86614
rect 156954 86294 157574 86378
rect 156954 86058 156986 86294
rect 157222 86058 157306 86294
rect 157542 86058 157574 86294
rect 156954 50614 157574 86058
rect 156954 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 157574 50614
rect 156954 50294 157574 50378
rect 156954 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 157574 50294
rect 156954 14614 157574 50058
rect 156954 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 157574 14614
rect 156954 14294 157574 14378
rect 156954 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 157574 14294
rect 138954 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 139574 -7066
rect 138954 -7386 139574 -7302
rect 138954 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 139574 -7386
rect 138954 -7654 139574 -7622
rect 156954 -6106 157574 14058
rect 163794 57454 164414 93100
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163794 21454 164414 56898
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 165662 21317 165722 407763
rect 167514 385174 168134 420618
rect 169707 389332 169773 389333
rect 169707 389268 169708 389332
rect 169772 389268 169773 389332
rect 169707 389267 169773 389268
rect 167514 384938 167546 385174
rect 167782 384938 167866 385174
rect 168102 384938 168134 385174
rect 167514 384854 168134 384938
rect 167514 384618 167546 384854
rect 167782 384618 167866 384854
rect 168102 384618 168134 384854
rect 167514 349174 168134 384618
rect 167514 348938 167546 349174
rect 167782 348938 167866 349174
rect 168102 348938 168134 349174
rect 167514 348854 168134 348938
rect 167514 348618 167546 348854
rect 167782 348618 167866 348854
rect 168102 348618 168134 348854
rect 167514 313174 168134 348618
rect 168971 342956 169037 342957
rect 168971 342892 168972 342956
rect 169036 342892 169037 342956
rect 168971 342891 169037 342892
rect 168235 329764 168301 329765
rect 168235 329700 168236 329764
rect 168300 329700 168301 329764
rect 168235 329699 168301 329700
rect 167514 312938 167546 313174
rect 167782 312938 167866 313174
rect 168102 312938 168134 313174
rect 167514 312854 168134 312938
rect 167514 312618 167546 312854
rect 167782 312618 167866 312854
rect 168102 312618 168134 312854
rect 167514 277174 168134 312618
rect 167514 276938 167546 277174
rect 167782 276938 167866 277174
rect 168102 276938 168134 277174
rect 167514 276854 168134 276938
rect 167514 276618 167546 276854
rect 167782 276618 167866 276854
rect 168102 276618 168134 276854
rect 167514 241174 168134 276618
rect 167514 240938 167546 241174
rect 167782 240938 167866 241174
rect 168102 240938 168134 241174
rect 167514 240854 168134 240938
rect 167514 240618 167546 240854
rect 167782 240618 167866 240854
rect 168102 240618 168134 240854
rect 167514 205174 168134 240618
rect 168238 240141 168298 329699
rect 168974 303789 169034 342891
rect 169523 327180 169589 327181
rect 169523 327116 169524 327180
rect 169588 327116 169589 327180
rect 169523 327115 169589 327116
rect 168971 303788 169037 303789
rect 168971 303724 168972 303788
rect 169036 303724 169037 303788
rect 168971 303723 169037 303724
rect 169526 269245 169586 327115
rect 169523 269244 169589 269245
rect 169523 269180 169524 269244
rect 169588 269180 169589 269244
rect 169523 269179 169589 269180
rect 169710 266389 169770 389267
rect 169707 266388 169773 266389
rect 169707 266324 169708 266388
rect 169772 266324 169773 266388
rect 169707 266323 169773 266324
rect 168971 265572 169037 265573
rect 168971 265508 168972 265572
rect 169036 265508 169037 265572
rect 168971 265507 169037 265508
rect 168419 251292 168485 251293
rect 168419 251228 168420 251292
rect 168484 251228 168485 251292
rect 168419 251227 168485 251228
rect 168235 240140 168301 240141
rect 168235 240076 168236 240140
rect 168300 240076 168301 240140
rect 168235 240075 168301 240076
rect 167514 204938 167546 205174
rect 167782 204938 167866 205174
rect 168102 204938 168134 205174
rect 167514 204854 168134 204938
rect 167514 204618 167546 204854
rect 167782 204618 167866 204854
rect 168102 204618 168134 204854
rect 167514 169174 168134 204618
rect 167514 168938 167546 169174
rect 167782 168938 167866 169174
rect 168102 168938 168134 169174
rect 167514 168854 168134 168938
rect 167514 168618 167546 168854
rect 167782 168618 167866 168854
rect 168102 168618 168134 168854
rect 167514 133174 168134 168618
rect 167514 132938 167546 133174
rect 167782 132938 167866 133174
rect 168102 132938 168134 133174
rect 167514 132854 168134 132938
rect 167514 132618 167546 132854
rect 167782 132618 167866 132854
rect 168102 132618 168134 132854
rect 166211 119372 166277 119373
rect 166211 119308 166212 119372
rect 166276 119308 166277 119372
rect 166211 119307 166277 119308
rect 166214 89861 166274 119307
rect 167514 97174 168134 132618
rect 168235 103596 168301 103597
rect 168235 103532 168236 103596
rect 168300 103532 168301 103596
rect 168235 103531 168301 103532
rect 167514 96938 167546 97174
rect 167782 96938 167866 97174
rect 168102 96938 168134 97174
rect 167514 96854 168134 96938
rect 167514 96618 167546 96854
rect 167782 96618 167866 96854
rect 168102 96618 168134 96854
rect 166211 89860 166277 89861
rect 166211 89796 166212 89860
rect 166276 89796 166277 89860
rect 166211 89795 166277 89796
rect 167514 61174 168134 96618
rect 168238 78437 168298 103531
rect 168235 78436 168301 78437
rect 168235 78372 168236 78436
rect 168300 78372 168301 78436
rect 168235 78371 168301 78372
rect 168422 69733 168482 251227
rect 168974 245037 169034 265507
rect 168971 245036 169037 245037
rect 168971 244972 168972 245036
rect 169036 244972 169037 245036
rect 168971 244971 169037 244972
rect 170262 241637 170322 552059
rect 171234 532894 171854 568338
rect 174954 680614 175574 711002
rect 192954 710598 193574 711590
rect 192954 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 193574 710598
rect 192954 710278 193574 710362
rect 192954 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 193574 710278
rect 189234 708678 189854 709670
rect 189234 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 189854 708678
rect 189234 708358 189854 708442
rect 189234 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 189854 708358
rect 185514 706758 186134 707750
rect 185514 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 186134 706758
rect 185514 706438 186134 706522
rect 185514 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 186134 706438
rect 174954 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 175574 680614
rect 174954 680294 175574 680378
rect 174954 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 175574 680294
rect 174954 644614 175574 680058
rect 174954 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 175574 644614
rect 174954 644294 175574 644378
rect 174954 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 175574 644294
rect 174954 608614 175574 644058
rect 174954 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 175574 608614
rect 174954 608294 175574 608378
rect 174954 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 175574 608294
rect 174954 572614 175574 608058
rect 174954 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 175574 572614
rect 174954 572294 175574 572378
rect 174954 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 175574 572294
rect 173019 550764 173085 550765
rect 173019 550700 173020 550764
rect 173084 550700 173085 550764
rect 173019 550699 173085 550700
rect 171234 532658 171266 532894
rect 171502 532658 171586 532894
rect 171822 532658 171854 532894
rect 171234 532574 171854 532658
rect 171234 532338 171266 532574
rect 171502 532338 171586 532574
rect 171822 532338 171854 532574
rect 171234 496894 171854 532338
rect 171234 496658 171266 496894
rect 171502 496658 171586 496894
rect 171822 496658 171854 496894
rect 171234 496574 171854 496658
rect 171234 496338 171266 496574
rect 171502 496338 171586 496574
rect 171822 496338 171854 496574
rect 171234 460894 171854 496338
rect 171234 460658 171266 460894
rect 171502 460658 171586 460894
rect 171822 460658 171854 460894
rect 171234 460574 171854 460658
rect 171234 460338 171266 460574
rect 171502 460338 171586 460574
rect 171822 460338 171854 460574
rect 171234 424894 171854 460338
rect 172467 456924 172533 456925
rect 172467 456860 172468 456924
rect 172532 456860 172533 456924
rect 172467 456859 172533 456860
rect 172099 449988 172165 449989
rect 172099 449924 172100 449988
rect 172164 449924 172165 449988
rect 172099 449923 172165 449924
rect 171234 424658 171266 424894
rect 171502 424658 171586 424894
rect 171822 424658 171854 424894
rect 171234 424574 171854 424658
rect 171234 424338 171266 424574
rect 171502 424338 171586 424574
rect 171822 424338 171854 424574
rect 171234 388894 171854 424338
rect 171234 388658 171266 388894
rect 171502 388658 171586 388894
rect 171822 388658 171854 388894
rect 171234 388574 171854 388658
rect 171234 388338 171266 388574
rect 171502 388338 171586 388574
rect 171822 388338 171854 388574
rect 171234 352894 171854 388338
rect 171234 352658 171266 352894
rect 171502 352658 171586 352894
rect 171822 352658 171854 352894
rect 171234 352574 171854 352658
rect 171234 352338 171266 352574
rect 171502 352338 171586 352574
rect 171822 352338 171854 352574
rect 171234 316894 171854 352338
rect 171234 316658 171266 316894
rect 171502 316658 171586 316894
rect 171822 316658 171854 316894
rect 171234 316574 171854 316658
rect 171234 316338 171266 316574
rect 171502 316338 171586 316574
rect 171822 316338 171854 316574
rect 171234 280894 171854 316338
rect 171234 280658 171266 280894
rect 171502 280658 171586 280894
rect 171822 280658 171854 280894
rect 171234 280574 171854 280658
rect 171234 280338 171266 280574
rect 171502 280338 171586 280574
rect 171822 280338 171854 280574
rect 170443 267612 170509 267613
rect 170443 267548 170444 267612
rect 170508 267548 170509 267612
rect 170443 267547 170509 267548
rect 170446 266525 170506 267547
rect 170443 266524 170509 266525
rect 170443 266460 170444 266524
rect 170508 266460 170509 266524
rect 170443 266459 170509 266460
rect 170259 241636 170325 241637
rect 170259 241572 170260 241636
rect 170324 241572 170325 241636
rect 170259 241571 170325 241572
rect 170262 142765 170322 241571
rect 170259 142764 170325 142765
rect 170259 142700 170260 142764
rect 170324 142700 170325 142764
rect 170259 142699 170325 142700
rect 168419 69732 168485 69733
rect 168419 69668 168420 69732
rect 168484 69668 168485 69732
rect 168419 69667 168485 69668
rect 167514 60938 167546 61174
rect 167782 60938 167866 61174
rect 168102 60938 168134 61174
rect 167514 60854 168134 60938
rect 167514 60618 167546 60854
rect 167782 60618 167866 60854
rect 168102 60618 168134 60854
rect 167514 25174 168134 60618
rect 167514 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 168134 25174
rect 167514 24854 168134 24938
rect 167514 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 168134 24854
rect 165659 21316 165725 21317
rect 165659 21252 165660 21316
rect 165724 21252 165725 21316
rect 165659 21251 165725 21252
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -1306 164414 20898
rect 163794 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 164414 -1306
rect 163794 -1626 164414 -1542
rect 163794 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 164414 -1626
rect 163794 -1894 164414 -1862
rect 167514 -3226 168134 24618
rect 170446 7581 170506 266459
rect 171234 244894 171854 280338
rect 171234 244658 171266 244894
rect 171502 244658 171586 244894
rect 171822 244658 171854 244894
rect 171234 244574 171854 244658
rect 171234 244338 171266 244574
rect 171502 244338 171586 244574
rect 171822 244338 171854 244574
rect 171234 208894 171854 244338
rect 172102 219061 172162 449923
rect 172470 296717 172530 456859
rect 172467 296716 172533 296717
rect 172467 296652 172468 296716
rect 172532 296652 172533 296716
rect 172467 296651 172533 296652
rect 172470 296309 172530 296651
rect 172467 296308 172533 296309
rect 172467 296244 172468 296308
rect 172532 296244 172533 296308
rect 172467 296243 172533 296244
rect 173022 228717 173082 550699
rect 174954 536614 175574 572058
rect 174954 536378 174986 536614
rect 175222 536378 175306 536614
rect 175542 536378 175574 536614
rect 174954 536294 175574 536378
rect 174954 536058 174986 536294
rect 175222 536058 175306 536294
rect 175542 536058 175574 536294
rect 174954 500614 175574 536058
rect 181794 704838 182414 705830
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 181794 543454 182414 578898
rect 181794 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 182414 543454
rect 181794 543134 182414 543218
rect 181794 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 182414 543134
rect 179275 530636 179341 530637
rect 179275 530572 179276 530636
rect 179340 530572 179341 530636
rect 179275 530571 179341 530572
rect 174954 500378 174986 500614
rect 175222 500378 175306 500614
rect 175542 500378 175574 500614
rect 174954 500294 175574 500378
rect 174954 500058 174986 500294
rect 175222 500058 175306 500294
rect 175542 500058 175574 500294
rect 174954 464614 175574 500058
rect 177803 496908 177869 496909
rect 177803 496844 177804 496908
rect 177868 496844 177869 496908
rect 177803 496843 177869 496844
rect 174954 464378 174986 464614
rect 175222 464378 175306 464614
rect 175542 464378 175574 464614
rect 174954 464294 175574 464378
rect 174954 464058 174986 464294
rect 175222 464058 175306 464294
rect 175542 464058 175574 464294
rect 174954 428614 175574 464058
rect 174954 428378 174986 428614
rect 175222 428378 175306 428614
rect 175542 428378 175574 428614
rect 174954 428294 175574 428378
rect 174954 428058 174986 428294
rect 175222 428058 175306 428294
rect 175542 428058 175574 428294
rect 174954 392614 175574 428058
rect 174954 392378 174986 392614
rect 175222 392378 175306 392614
rect 175542 392378 175574 392614
rect 174954 392294 175574 392378
rect 174954 392058 174986 392294
rect 175222 392058 175306 392294
rect 175542 392058 175574 392294
rect 174954 356614 175574 392058
rect 174954 356378 174986 356614
rect 175222 356378 175306 356614
rect 175542 356378 175574 356614
rect 174954 356294 175574 356378
rect 174954 356058 174986 356294
rect 175222 356058 175306 356294
rect 175542 356058 175574 356294
rect 174954 320614 175574 356058
rect 174954 320378 174986 320614
rect 175222 320378 175306 320614
rect 175542 320378 175574 320614
rect 174954 320294 175574 320378
rect 174954 320058 174986 320294
rect 175222 320058 175306 320294
rect 175542 320058 175574 320294
rect 174675 314260 174741 314261
rect 174675 314196 174676 314260
rect 174740 314196 174741 314260
rect 174675 314195 174741 314196
rect 173755 295356 173821 295357
rect 173755 295292 173756 295356
rect 173820 295292 173821 295356
rect 173755 295291 173821 295292
rect 173019 228716 173085 228717
rect 173019 228652 173020 228716
rect 173084 228652 173085 228716
rect 173019 228651 173085 228652
rect 172099 219060 172165 219061
rect 172099 218996 172100 219060
rect 172164 218996 172165 219060
rect 172099 218995 172165 218996
rect 171234 208658 171266 208894
rect 171502 208658 171586 208894
rect 171822 208658 171854 208894
rect 171234 208574 171854 208658
rect 171234 208338 171266 208574
rect 171502 208338 171586 208574
rect 171822 208338 171854 208574
rect 171234 172894 171854 208338
rect 171234 172658 171266 172894
rect 171502 172658 171586 172894
rect 171822 172658 171854 172894
rect 171234 172574 171854 172658
rect 171234 172338 171266 172574
rect 171502 172338 171586 172574
rect 171822 172338 171854 172574
rect 171234 136894 171854 172338
rect 172102 152421 172162 218995
rect 173022 196757 173082 228651
rect 173019 196756 173085 196757
rect 173019 196692 173020 196756
rect 173084 196692 173085 196756
rect 173019 196691 173085 196692
rect 172099 152420 172165 152421
rect 172099 152356 172100 152420
rect 172164 152356 172165 152420
rect 172099 152355 172165 152356
rect 171234 136658 171266 136894
rect 171502 136658 171586 136894
rect 171822 136658 171854 136894
rect 171234 136574 171854 136658
rect 171234 136338 171266 136574
rect 171502 136338 171586 136574
rect 171822 136338 171854 136574
rect 171234 100894 171854 136338
rect 171234 100658 171266 100894
rect 171502 100658 171586 100894
rect 171822 100658 171854 100894
rect 171234 100574 171854 100658
rect 171234 100338 171266 100574
rect 171502 100338 171586 100574
rect 171822 100338 171854 100574
rect 171234 64894 171854 100338
rect 171234 64658 171266 64894
rect 171502 64658 171586 64894
rect 171822 64658 171854 64894
rect 171234 64574 171854 64658
rect 171234 64338 171266 64574
rect 171502 64338 171586 64574
rect 171822 64338 171854 64574
rect 171234 28894 171854 64338
rect 171234 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 171854 28894
rect 171234 28574 171854 28658
rect 171234 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 171854 28574
rect 170443 7580 170509 7581
rect 170443 7516 170444 7580
rect 170508 7516 170509 7580
rect 170443 7515 170509 7516
rect 167514 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 168134 -3226
rect 167514 -3546 168134 -3462
rect 167514 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 168134 -3546
rect 167514 -3814 168134 -3782
rect 171234 -5146 171854 28338
rect 173758 18597 173818 295291
rect 174678 211853 174738 314195
rect 174954 284614 175574 320058
rect 176515 318068 176581 318069
rect 176515 318004 176516 318068
rect 176580 318004 176581 318068
rect 176515 318003 176581 318004
rect 174954 284378 174986 284614
rect 175222 284378 175306 284614
rect 175542 284378 175574 284614
rect 174954 284294 175574 284378
rect 174954 284058 174986 284294
rect 175222 284058 175306 284294
rect 175542 284058 175574 284294
rect 174954 248614 175574 284058
rect 174954 248378 174986 248614
rect 175222 248378 175306 248614
rect 175542 248378 175574 248614
rect 174954 248294 175574 248378
rect 174954 248058 174986 248294
rect 175222 248058 175306 248294
rect 175542 248058 175574 248294
rect 174954 212614 175574 248058
rect 176518 216069 176578 318003
rect 177806 229110 177866 496843
rect 178539 272508 178605 272509
rect 178539 272444 178540 272508
rect 178604 272444 178605 272508
rect 178539 272443 178605 272444
rect 177806 229050 178050 229110
rect 177990 217701 178050 229050
rect 177987 217700 178053 217701
rect 177987 217636 177988 217700
rect 178052 217636 178053 217700
rect 177987 217635 178053 217636
rect 177990 217293 178050 217635
rect 177987 217292 178053 217293
rect 177987 217228 177988 217292
rect 178052 217228 178053 217292
rect 177987 217227 178053 217228
rect 176515 216068 176581 216069
rect 176515 216004 176516 216068
rect 176580 216004 176581 216068
rect 176515 216003 176581 216004
rect 174954 212378 174986 212614
rect 175222 212378 175306 212614
rect 175542 212378 175574 212614
rect 174954 212294 175574 212378
rect 174954 212058 174986 212294
rect 175222 212058 175306 212294
rect 175542 212058 175574 212294
rect 174675 211852 174741 211853
rect 174675 211788 174676 211852
rect 174740 211788 174741 211852
rect 174675 211787 174741 211788
rect 174954 176614 175574 212058
rect 174954 176378 174986 176614
rect 175222 176378 175306 176614
rect 175542 176378 175574 176614
rect 174954 176294 175574 176378
rect 174954 176058 174986 176294
rect 175222 176058 175306 176294
rect 175542 176058 175574 176294
rect 174954 140614 175574 176058
rect 174954 140378 174986 140614
rect 175222 140378 175306 140614
rect 175542 140378 175574 140614
rect 174954 140294 175574 140378
rect 174954 140058 174986 140294
rect 175222 140058 175306 140294
rect 175542 140058 175574 140294
rect 174954 104614 175574 140058
rect 174954 104378 174986 104614
rect 175222 104378 175306 104614
rect 175542 104378 175574 104614
rect 174954 104294 175574 104378
rect 174954 104058 174986 104294
rect 175222 104058 175306 104294
rect 175542 104058 175574 104294
rect 174954 68614 175574 104058
rect 178542 91765 178602 272443
rect 179278 209541 179338 530571
rect 181794 507454 182414 542898
rect 185514 691174 186134 706202
rect 185514 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 186134 691174
rect 185514 690854 186134 690938
rect 185514 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 186134 690854
rect 185514 655174 186134 690618
rect 185514 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 186134 655174
rect 185514 654854 186134 654938
rect 185514 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 186134 654854
rect 185514 619174 186134 654618
rect 185514 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 186134 619174
rect 185514 618854 186134 618938
rect 185514 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 186134 618854
rect 185514 583174 186134 618618
rect 185514 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 186134 583174
rect 185514 582854 186134 582938
rect 185514 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 186134 582854
rect 185514 547174 186134 582618
rect 185514 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 186134 547174
rect 185514 546854 186134 546938
rect 185514 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 186134 546854
rect 183323 534172 183389 534173
rect 183323 534108 183324 534172
rect 183388 534108 183389 534172
rect 183323 534107 183389 534108
rect 181794 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 182414 507454
rect 181794 507134 182414 507218
rect 181794 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 182414 507134
rect 181794 471454 182414 506898
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 181794 435454 182414 470898
rect 181794 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 182414 435454
rect 181794 435134 182414 435218
rect 181794 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 182414 435134
rect 181794 399454 182414 434898
rect 181794 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 182414 399454
rect 181794 399134 182414 399218
rect 181794 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 182414 399134
rect 181794 363454 182414 398898
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 180563 354108 180629 354109
rect 180563 354044 180564 354108
rect 180628 354044 180629 354108
rect 180563 354043 180629 354044
rect 180566 353565 180626 354043
rect 180563 353564 180629 353565
rect 180563 353500 180564 353564
rect 180628 353500 180629 353564
rect 180563 353499 180629 353500
rect 179275 209540 179341 209541
rect 179275 209476 179276 209540
rect 179340 209476 179341 209540
rect 179275 209475 179341 209476
rect 179278 208997 179338 209475
rect 179275 208996 179341 208997
rect 179275 208932 179276 208996
rect 179340 208932 179341 208996
rect 179275 208931 179341 208932
rect 178539 91764 178605 91765
rect 178539 91700 178540 91764
rect 178604 91700 178605 91764
rect 178539 91699 178605 91700
rect 174954 68378 174986 68614
rect 175222 68378 175306 68614
rect 175542 68378 175574 68614
rect 174954 68294 175574 68378
rect 174954 68058 174986 68294
rect 175222 68058 175306 68294
rect 175542 68058 175574 68294
rect 174954 32614 175574 68058
rect 174954 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 175574 32614
rect 174954 32294 175574 32378
rect 174954 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 175574 32294
rect 173755 18596 173821 18597
rect 173755 18532 173756 18596
rect 173820 18532 173821 18596
rect 173755 18531 173821 18532
rect 171234 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 171854 -5146
rect 171234 -5466 171854 -5382
rect 171234 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 171854 -5466
rect 171234 -5734 171854 -5702
rect 156954 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 157574 -6106
rect 156954 -6426 157574 -6342
rect 156954 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 157574 -6426
rect 156954 -7654 157574 -6662
rect 174954 -7066 175574 32058
rect 180566 9077 180626 353499
rect 181794 327454 182414 362898
rect 181794 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 182414 327454
rect 181794 327134 182414 327218
rect 181794 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 182414 327134
rect 181794 291454 182414 326898
rect 181794 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 182414 291454
rect 181794 291134 182414 291218
rect 181794 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 182414 291134
rect 181794 255454 182414 290898
rect 181794 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 182414 255454
rect 181794 255134 182414 255218
rect 181794 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 182414 255134
rect 181794 219454 182414 254898
rect 181794 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 182414 219454
rect 181794 219134 182414 219218
rect 181794 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 182414 219134
rect 181794 183454 182414 218898
rect 183326 213893 183386 534107
rect 185514 511174 186134 546618
rect 189234 694894 189854 708122
rect 189234 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 189854 694894
rect 189234 694574 189854 694658
rect 189234 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 189854 694574
rect 189234 658894 189854 694338
rect 189234 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 189854 658894
rect 189234 658574 189854 658658
rect 189234 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 189854 658574
rect 189234 622894 189854 658338
rect 189234 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 189854 622894
rect 189234 622574 189854 622658
rect 189234 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 189854 622574
rect 189234 586894 189854 622338
rect 189234 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 189854 586894
rect 189234 586574 189854 586658
rect 189234 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 189854 586574
rect 189234 550894 189854 586338
rect 189234 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 189854 550894
rect 189234 550574 189854 550658
rect 189234 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 189854 550574
rect 188843 541244 188909 541245
rect 188843 541180 188844 541244
rect 188908 541180 188909 541244
rect 188843 541179 188909 541180
rect 185514 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 186134 511174
rect 185514 510854 186134 510938
rect 185514 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 186134 510854
rect 184795 502484 184861 502485
rect 184795 502420 184796 502484
rect 184860 502420 184861 502484
rect 184795 502419 184861 502420
rect 184059 297532 184125 297533
rect 184059 297468 184060 297532
rect 184124 297468 184125 297532
rect 184059 297467 184125 297468
rect 184062 235653 184122 297467
rect 184059 235652 184125 235653
rect 184059 235588 184060 235652
rect 184124 235588 184125 235652
rect 184059 235587 184125 235588
rect 184798 226269 184858 502419
rect 185514 475174 186134 510618
rect 185514 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 186134 475174
rect 185514 474854 186134 474938
rect 185514 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 186134 474854
rect 185514 439174 186134 474618
rect 185514 438938 185546 439174
rect 185782 438938 185866 439174
rect 186102 438938 186134 439174
rect 185514 438854 186134 438938
rect 185514 438618 185546 438854
rect 185782 438618 185866 438854
rect 186102 438618 186134 438854
rect 185514 403174 186134 438618
rect 186819 430676 186885 430677
rect 186819 430612 186820 430676
rect 186884 430612 186885 430676
rect 186819 430611 186885 430612
rect 185514 402938 185546 403174
rect 185782 402938 185866 403174
rect 186102 402938 186134 403174
rect 185514 402854 186134 402938
rect 185514 402618 185546 402854
rect 185782 402618 185866 402854
rect 186102 402618 186134 402854
rect 185514 367174 186134 402618
rect 185514 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 186134 367174
rect 185514 366854 186134 366938
rect 185514 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 186134 366854
rect 185514 331174 186134 366618
rect 185514 330938 185546 331174
rect 185782 330938 185866 331174
rect 186102 330938 186134 331174
rect 185514 330854 186134 330938
rect 185514 330618 185546 330854
rect 185782 330618 185866 330854
rect 186102 330618 186134 330854
rect 185347 315348 185413 315349
rect 185347 315284 185348 315348
rect 185412 315284 185413 315348
rect 185347 315283 185413 315284
rect 184795 226268 184861 226269
rect 184795 226204 184796 226268
rect 184860 226204 184861 226268
rect 184795 226203 184861 226204
rect 183323 213892 183389 213893
rect 183323 213828 183324 213892
rect 183388 213828 183389 213892
rect 183323 213827 183389 213828
rect 181794 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 182414 183454
rect 181794 183134 182414 183218
rect 181794 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 182414 183134
rect 181794 147454 182414 182898
rect 181794 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 182414 147454
rect 181794 147134 182414 147218
rect 181794 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 182414 147134
rect 181794 111454 182414 146898
rect 181794 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 182414 111454
rect 181794 111134 182414 111218
rect 181794 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 182414 111134
rect 181794 75454 182414 110898
rect 181794 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 182414 75454
rect 181794 75134 182414 75218
rect 181794 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 182414 75134
rect 181794 39454 182414 74898
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 180563 9076 180629 9077
rect 180563 9012 180564 9076
rect 180628 9012 180629 9076
rect 180563 9011 180629 9012
rect 181794 3454 182414 38898
rect 185350 13021 185410 315283
rect 185514 295174 186134 330618
rect 185514 294938 185546 295174
rect 185782 294938 185866 295174
rect 186102 294938 186134 295174
rect 185514 294854 186134 294938
rect 185514 294618 185546 294854
rect 185782 294618 185866 294854
rect 186102 294618 186134 294854
rect 185514 259174 186134 294618
rect 185514 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 186134 259174
rect 185514 258854 186134 258938
rect 185514 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 186134 258854
rect 185514 223174 186134 258618
rect 186822 245853 186882 430611
rect 187003 347716 187069 347717
rect 187003 347652 187004 347716
rect 187068 347652 187069 347716
rect 187003 347651 187069 347652
rect 187006 346493 187066 347651
rect 187003 346492 187069 346493
rect 187003 346428 187004 346492
rect 187068 346428 187069 346492
rect 187003 346427 187069 346428
rect 186819 245852 186885 245853
rect 186819 245788 186820 245852
rect 186884 245788 186885 245852
rect 186819 245787 186885 245788
rect 185514 222938 185546 223174
rect 185782 222938 185866 223174
rect 186102 222938 186134 223174
rect 185514 222854 186134 222938
rect 185514 222618 185546 222854
rect 185782 222618 185866 222854
rect 186102 222618 186134 222854
rect 185514 187174 186134 222618
rect 185514 186938 185546 187174
rect 185782 186938 185866 187174
rect 186102 186938 186134 187174
rect 185514 186854 186134 186938
rect 185514 186618 185546 186854
rect 185782 186618 185866 186854
rect 186102 186618 186134 186854
rect 185514 151174 186134 186618
rect 187006 183021 187066 346427
rect 188846 215253 188906 541179
rect 189234 514894 189854 550338
rect 192954 698614 193574 710042
rect 210954 711558 211574 711590
rect 210954 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 211574 711558
rect 210954 711238 211574 711322
rect 210954 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 211574 711238
rect 207234 709638 207854 709670
rect 207234 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 207854 709638
rect 207234 709318 207854 709402
rect 207234 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 207854 709318
rect 203514 707718 204134 707750
rect 203514 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 204134 707718
rect 203514 707398 204134 707482
rect 203514 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 204134 707398
rect 192954 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 193574 698614
rect 192954 698294 193574 698378
rect 192954 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 193574 698294
rect 192954 662614 193574 698058
rect 192954 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 193574 662614
rect 192954 662294 193574 662378
rect 192954 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 193574 662294
rect 192954 626614 193574 662058
rect 192954 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 193574 626614
rect 192954 626294 193574 626378
rect 192954 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 193574 626294
rect 192954 590614 193574 626058
rect 192954 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 193574 590614
rect 192954 590294 193574 590378
rect 192954 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 193574 590294
rect 192954 554614 193574 590058
rect 192954 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 193574 554614
rect 192954 554294 193574 554378
rect 192954 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 193574 554294
rect 191603 535396 191669 535397
rect 191603 535332 191604 535396
rect 191668 535332 191669 535396
rect 191603 535331 191669 535332
rect 189234 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 189854 514894
rect 189234 514574 189854 514658
rect 189234 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 189854 514574
rect 189234 478894 189854 514338
rect 189234 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 189854 478894
rect 189234 478574 189854 478658
rect 189234 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 189854 478574
rect 189234 442894 189854 478338
rect 189234 442658 189266 442894
rect 189502 442658 189586 442894
rect 189822 442658 189854 442894
rect 189234 442574 189854 442658
rect 189234 442338 189266 442574
rect 189502 442338 189586 442574
rect 189822 442338 189854 442574
rect 189234 406894 189854 442338
rect 189234 406658 189266 406894
rect 189502 406658 189586 406894
rect 189822 406658 189854 406894
rect 189234 406574 189854 406658
rect 189234 406338 189266 406574
rect 189502 406338 189586 406574
rect 189822 406338 189854 406574
rect 189234 370894 189854 406338
rect 189234 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 189854 370894
rect 189234 370574 189854 370658
rect 189234 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 189854 370574
rect 189234 334894 189854 370338
rect 189234 334658 189266 334894
rect 189502 334658 189586 334894
rect 189822 334658 189854 334894
rect 189234 334574 189854 334658
rect 189234 334338 189266 334574
rect 189502 334338 189586 334574
rect 189822 334338 189854 334574
rect 189234 298894 189854 334338
rect 189947 331940 190013 331941
rect 189947 331876 189948 331940
rect 190012 331876 190013 331940
rect 189947 331875 190013 331876
rect 189234 298658 189266 298894
rect 189502 298658 189586 298894
rect 189822 298658 189854 298894
rect 189234 298574 189854 298658
rect 189234 298338 189266 298574
rect 189502 298338 189586 298574
rect 189822 298338 189854 298574
rect 189234 262894 189854 298338
rect 189234 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 189854 262894
rect 189234 262574 189854 262658
rect 189234 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 189854 262574
rect 189234 226894 189854 262338
rect 189234 226658 189266 226894
rect 189502 226658 189586 226894
rect 189822 226658 189854 226894
rect 189234 226574 189854 226658
rect 189234 226338 189266 226574
rect 189502 226338 189586 226574
rect 189822 226338 189854 226574
rect 188843 215252 188909 215253
rect 188843 215188 188844 215252
rect 188908 215188 188909 215252
rect 188843 215187 188909 215188
rect 189234 190894 189854 226338
rect 189234 190658 189266 190894
rect 189502 190658 189586 190894
rect 189822 190658 189854 190894
rect 189234 190574 189854 190658
rect 189234 190338 189266 190574
rect 189502 190338 189586 190574
rect 189822 190338 189854 190574
rect 187003 183020 187069 183021
rect 187003 182956 187004 183020
rect 187068 182956 187069 183020
rect 187003 182955 187069 182956
rect 185514 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 186134 151174
rect 185514 150854 186134 150938
rect 185514 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 186134 150854
rect 185514 115174 186134 150618
rect 185514 114938 185546 115174
rect 185782 114938 185866 115174
rect 186102 114938 186134 115174
rect 185514 114854 186134 114938
rect 185514 114618 185546 114854
rect 185782 114618 185866 114854
rect 186102 114618 186134 114854
rect 185514 79174 186134 114618
rect 185514 78938 185546 79174
rect 185782 78938 185866 79174
rect 186102 78938 186134 79174
rect 185514 78854 186134 78938
rect 185514 78618 185546 78854
rect 185782 78618 185866 78854
rect 186102 78618 186134 78854
rect 185514 43174 186134 78618
rect 185514 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 186134 43174
rect 185514 42854 186134 42938
rect 185514 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 186134 42854
rect 185347 13020 185413 13021
rect 185347 12956 185348 13020
rect 185412 12956 185413 13020
rect 185347 12955 185413 12956
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -1894 182414 -902
rect 185514 7174 186134 42618
rect 185514 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 186134 7174
rect 185514 6854 186134 6938
rect 185514 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 186134 6854
rect 185514 -2266 186134 6618
rect 185514 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 186134 -2266
rect 185514 -2586 186134 -2502
rect 185514 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 186134 -2586
rect 185514 -3814 186134 -2822
rect 189234 154894 189854 190338
rect 189234 154658 189266 154894
rect 189502 154658 189586 154894
rect 189822 154658 189854 154894
rect 189234 154574 189854 154658
rect 189234 154338 189266 154574
rect 189502 154338 189586 154574
rect 189822 154338 189854 154574
rect 189234 118894 189854 154338
rect 189234 118658 189266 118894
rect 189502 118658 189586 118894
rect 189822 118658 189854 118894
rect 189234 118574 189854 118658
rect 189234 118338 189266 118574
rect 189502 118338 189586 118574
rect 189822 118338 189854 118574
rect 189234 82894 189854 118338
rect 189234 82658 189266 82894
rect 189502 82658 189586 82894
rect 189822 82658 189854 82894
rect 189234 82574 189854 82658
rect 189234 82338 189266 82574
rect 189502 82338 189586 82574
rect 189822 82338 189854 82574
rect 189234 46894 189854 82338
rect 189234 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 189854 46894
rect 189234 46574 189854 46658
rect 189234 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 189854 46574
rect 189234 10894 189854 46338
rect 189950 17373 190010 331875
rect 191606 206413 191666 535331
rect 192954 518614 193574 554058
rect 199794 705798 200414 705830
rect 199794 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 200414 705798
rect 199794 705478 200414 705562
rect 199794 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 200414 705478
rect 199794 669454 200414 705242
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 633454 200414 668898
rect 199794 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 200414 633454
rect 199794 633134 200414 633218
rect 199794 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 200414 633134
rect 199794 597454 200414 632898
rect 199794 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 200414 597454
rect 199794 597134 200414 597218
rect 199794 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 200414 597134
rect 199794 561454 200414 596898
rect 199794 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 200414 561454
rect 199794 561134 200414 561218
rect 199794 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 200414 561134
rect 197859 546684 197925 546685
rect 197859 546620 197860 546684
rect 197924 546620 197925 546684
rect 197859 546619 197925 546620
rect 197862 526421 197922 546619
rect 199515 546548 199581 546549
rect 199515 546484 199516 546548
rect 199580 546484 199581 546548
rect 199515 546483 199581 546484
rect 197859 526420 197925 526421
rect 197859 526356 197860 526420
rect 197924 526356 197925 526420
rect 197859 526355 197925 526356
rect 192954 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 193574 518614
rect 192954 518294 193574 518378
rect 192954 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 193574 518294
rect 192954 482614 193574 518058
rect 195099 514996 195165 514997
rect 195099 514932 195100 514996
rect 195164 514932 195165 514996
rect 195099 514931 195165 514932
rect 192954 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 193574 482614
rect 192954 482294 193574 482378
rect 192954 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 193574 482294
rect 192954 446614 193574 482058
rect 192954 446378 192986 446614
rect 193222 446378 193306 446614
rect 193542 446378 193574 446614
rect 192954 446294 193574 446378
rect 192954 446058 192986 446294
rect 193222 446058 193306 446294
rect 193542 446058 193574 446294
rect 192954 410614 193574 446058
rect 192954 410378 192986 410614
rect 193222 410378 193306 410614
rect 193542 410378 193574 410614
rect 192954 410294 193574 410378
rect 192954 410058 192986 410294
rect 193222 410058 193306 410294
rect 193542 410058 193574 410294
rect 192707 404564 192773 404565
rect 192707 404500 192708 404564
rect 192772 404500 192773 404564
rect 192707 404499 192773 404500
rect 192710 208317 192770 404499
rect 192954 374614 193574 410058
rect 192954 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 193574 374614
rect 192954 374294 193574 374378
rect 192954 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 193574 374294
rect 192954 338614 193574 374058
rect 192954 338378 192986 338614
rect 193222 338378 193306 338614
rect 193542 338378 193574 338614
rect 192954 338294 193574 338378
rect 192954 338058 192986 338294
rect 193222 338058 193306 338294
rect 193542 338058 193574 338294
rect 192954 302614 193574 338058
rect 195102 322285 195162 514931
rect 198595 512548 198661 512549
rect 198595 512484 198596 512548
rect 198660 512484 198661 512548
rect 198595 512483 198661 512484
rect 197123 438972 197189 438973
rect 197123 438908 197124 438972
rect 197188 438908 197189 438972
rect 197123 438907 197189 438908
rect 195835 384844 195901 384845
rect 195835 384780 195836 384844
rect 195900 384780 195901 384844
rect 195835 384779 195901 384780
rect 195838 376549 195898 384779
rect 196571 378180 196637 378181
rect 196571 378116 196572 378180
rect 196636 378116 196637 378180
rect 196571 378115 196637 378116
rect 195835 376548 195901 376549
rect 195835 376484 195836 376548
rect 195900 376484 195901 376548
rect 195835 376483 195901 376484
rect 195283 368660 195349 368661
rect 195283 368596 195284 368660
rect 195348 368596 195349 368660
rect 195283 368595 195349 368596
rect 195099 322284 195165 322285
rect 195099 322220 195100 322284
rect 195164 322220 195165 322284
rect 195099 322219 195165 322220
rect 192954 302378 192986 302614
rect 193222 302378 193306 302614
rect 193542 302378 193574 302614
rect 192954 302294 193574 302378
rect 192954 302058 192986 302294
rect 193222 302058 193306 302294
rect 193542 302058 193574 302294
rect 192954 266614 193574 302058
rect 192954 266378 192986 266614
rect 193222 266378 193306 266614
rect 193542 266378 193574 266614
rect 192954 266294 193574 266378
rect 192954 266058 192986 266294
rect 193222 266058 193306 266294
rect 193542 266058 193574 266294
rect 192954 230614 193574 266058
rect 195286 259453 195346 368595
rect 196574 362405 196634 378115
rect 196571 362404 196637 362405
rect 196571 362340 196572 362404
rect 196636 362340 196637 362404
rect 196571 362339 196637 362340
rect 195835 300932 195901 300933
rect 195835 300868 195836 300932
rect 195900 300868 195901 300932
rect 195835 300867 195901 300868
rect 195838 267341 195898 300867
rect 196939 290460 197005 290461
rect 196939 290396 196940 290460
rect 197004 290396 197005 290460
rect 196939 290395 197005 290396
rect 195835 267340 195901 267341
rect 195835 267276 195836 267340
rect 195900 267276 195901 267340
rect 195835 267275 195901 267276
rect 195283 259452 195349 259453
rect 195283 259388 195284 259452
rect 195348 259388 195349 259452
rect 195283 259387 195349 259388
rect 195099 254420 195165 254421
rect 195099 254356 195100 254420
rect 195164 254356 195165 254420
rect 195099 254355 195165 254356
rect 192954 230378 192986 230614
rect 193222 230378 193306 230614
rect 193542 230378 193574 230614
rect 192954 230294 193574 230378
rect 192954 230058 192986 230294
rect 193222 230058 193306 230294
rect 193542 230058 193574 230294
rect 192707 208316 192773 208317
rect 192707 208252 192708 208316
rect 192772 208252 192773 208316
rect 192707 208251 192773 208252
rect 192710 207229 192770 208251
rect 192707 207228 192773 207229
rect 192707 207164 192708 207228
rect 192772 207164 192773 207228
rect 192707 207163 192773 207164
rect 191603 206412 191669 206413
rect 191603 206348 191604 206412
rect 191668 206348 191669 206412
rect 191603 206347 191669 206348
rect 192954 194614 193574 230058
rect 195102 220829 195162 254355
rect 195283 242860 195349 242861
rect 195283 242796 195284 242860
rect 195348 242796 195349 242860
rect 195283 242795 195349 242796
rect 195286 241909 195346 242795
rect 195283 241908 195349 241909
rect 195283 241844 195284 241908
rect 195348 241844 195349 241908
rect 195283 241843 195349 241844
rect 195286 229805 195346 241843
rect 196942 238509 197002 290395
rect 196939 238508 197005 238509
rect 196939 238444 196940 238508
rect 197004 238444 197005 238508
rect 196939 238443 197005 238444
rect 195283 229804 195349 229805
rect 195283 229740 195284 229804
rect 195348 229740 195349 229804
rect 195283 229739 195349 229740
rect 195099 220828 195165 220829
rect 195099 220764 195100 220828
rect 195164 220764 195165 220828
rect 195099 220763 195165 220764
rect 197126 205597 197186 438907
rect 197859 421700 197925 421701
rect 197859 421636 197860 421700
rect 197924 421636 197925 421700
rect 197859 421635 197925 421636
rect 197862 252653 197922 421635
rect 198598 393413 198658 512483
rect 198779 485620 198845 485621
rect 198779 485556 198780 485620
rect 198844 485556 198845 485620
rect 198779 485555 198845 485556
rect 198595 393412 198661 393413
rect 198595 393348 198596 393412
rect 198660 393348 198661 393412
rect 198595 393347 198661 393348
rect 198598 314805 198658 393347
rect 198782 377637 198842 485555
rect 198779 377636 198845 377637
rect 198779 377572 198780 377636
rect 198844 377572 198845 377636
rect 198779 377571 198845 377572
rect 199518 353565 199578 546483
rect 199794 537993 200414 560898
rect 203514 673174 204134 707162
rect 203514 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 204134 673174
rect 203514 672854 204134 672938
rect 203514 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 204134 672854
rect 203514 637174 204134 672618
rect 203514 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 204134 637174
rect 203514 636854 204134 636938
rect 203514 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 204134 636854
rect 203514 601174 204134 636618
rect 203514 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 204134 601174
rect 203514 600854 204134 600938
rect 203514 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 204134 600854
rect 203514 565174 204134 600618
rect 203514 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 204134 565174
rect 203514 564854 204134 564938
rect 203514 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 204134 564854
rect 200619 545324 200685 545325
rect 200619 545260 200620 545324
rect 200684 545260 200685 545324
rect 200619 545259 200685 545260
rect 200067 533492 200133 533493
rect 200067 533428 200068 533492
rect 200132 533490 200133 533492
rect 200622 533490 200682 545259
rect 203514 537993 204134 564618
rect 207234 676894 207854 709082
rect 207234 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 207854 676894
rect 207234 676574 207854 676658
rect 207234 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 207854 676574
rect 207234 640894 207854 676338
rect 207234 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 207854 640894
rect 207234 640574 207854 640658
rect 207234 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 207854 640574
rect 207234 604894 207854 640338
rect 207234 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 207854 604894
rect 207234 604574 207854 604658
rect 207234 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 207854 604574
rect 207234 568894 207854 604338
rect 207234 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 207854 568894
rect 207234 568574 207854 568658
rect 207234 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 207854 568574
rect 207234 537993 207854 568338
rect 210954 680614 211574 711002
rect 228954 710598 229574 711590
rect 228954 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 229574 710598
rect 228954 710278 229574 710362
rect 228954 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 229574 710278
rect 225234 708678 225854 709670
rect 225234 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 225854 708678
rect 225234 708358 225854 708442
rect 225234 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 225854 708358
rect 221514 706758 222134 707750
rect 221514 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 222134 706758
rect 221514 706438 222134 706522
rect 221514 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 222134 706438
rect 210954 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 211574 680614
rect 210954 680294 211574 680378
rect 210954 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 211574 680294
rect 210954 644614 211574 680058
rect 210954 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 211574 644614
rect 210954 644294 211574 644378
rect 210954 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 211574 644294
rect 210954 608614 211574 644058
rect 210954 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 211574 608614
rect 210954 608294 211574 608378
rect 210954 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 211574 608294
rect 210954 572614 211574 608058
rect 210954 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 211574 572614
rect 210954 572294 211574 572378
rect 210954 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 211574 572294
rect 210954 537993 211574 572058
rect 217794 704838 218414 705830
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 579454 218414 614898
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 217794 543454 218414 578898
rect 217794 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 218414 543454
rect 217794 543134 218414 543218
rect 217794 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 218414 543134
rect 217794 537993 218414 542898
rect 221514 691174 222134 706202
rect 221514 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 222134 691174
rect 221514 690854 222134 690938
rect 221514 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 222134 690854
rect 221514 655174 222134 690618
rect 221514 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 222134 655174
rect 221514 654854 222134 654938
rect 221514 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 222134 654854
rect 221514 619174 222134 654618
rect 221514 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 222134 619174
rect 221514 618854 222134 618938
rect 221514 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 222134 618854
rect 221514 583174 222134 618618
rect 221514 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 222134 583174
rect 221514 582854 222134 582938
rect 221514 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 222134 582854
rect 221514 547174 222134 582618
rect 221514 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 222134 547174
rect 221514 546854 222134 546938
rect 221514 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 222134 546854
rect 221514 537993 222134 546618
rect 225234 694894 225854 708122
rect 225234 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 225854 694894
rect 225234 694574 225854 694658
rect 225234 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 225854 694574
rect 225234 658894 225854 694338
rect 225234 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 225854 658894
rect 225234 658574 225854 658658
rect 225234 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 225854 658574
rect 225234 622894 225854 658338
rect 225234 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 225854 622894
rect 225234 622574 225854 622658
rect 225234 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 225854 622574
rect 225234 586894 225854 622338
rect 225234 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 225854 586894
rect 225234 586574 225854 586658
rect 225234 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 225854 586574
rect 225234 550894 225854 586338
rect 225234 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 225854 550894
rect 225234 550574 225854 550658
rect 225234 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 225854 550574
rect 225234 537993 225854 550338
rect 228954 698614 229574 710042
rect 246954 711558 247574 711590
rect 246954 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 247574 711558
rect 246954 711238 247574 711322
rect 246954 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 247574 711238
rect 243234 709638 243854 709670
rect 243234 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 243854 709638
rect 243234 709318 243854 709402
rect 243234 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 243854 709318
rect 239514 707718 240134 707750
rect 239514 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 240134 707718
rect 239514 707398 240134 707482
rect 239514 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 240134 707398
rect 228954 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 229574 698614
rect 228954 698294 229574 698378
rect 228954 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 229574 698294
rect 228954 662614 229574 698058
rect 228954 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 229574 662614
rect 228954 662294 229574 662378
rect 228954 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 229574 662294
rect 228954 626614 229574 662058
rect 228954 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 229574 626614
rect 228954 626294 229574 626378
rect 228954 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 229574 626294
rect 228954 590614 229574 626058
rect 228954 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 229574 590614
rect 228954 590294 229574 590378
rect 228954 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 229574 590294
rect 228954 554614 229574 590058
rect 228954 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 229574 554614
rect 228954 554294 229574 554378
rect 228954 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 229574 554294
rect 228954 537993 229574 554058
rect 235794 705798 236414 705830
rect 235794 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 236414 705798
rect 235794 705478 236414 705562
rect 235794 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 236414 705478
rect 235794 669454 236414 705242
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 633454 236414 668898
rect 235794 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 236414 633454
rect 235794 633134 236414 633218
rect 235794 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 236414 633134
rect 235794 597454 236414 632898
rect 235794 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 236414 597454
rect 235794 597134 236414 597218
rect 235794 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 236414 597134
rect 235794 561454 236414 596898
rect 235794 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 236414 561454
rect 235794 561134 236414 561218
rect 235794 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 236414 561134
rect 235794 537993 236414 560898
rect 239514 673174 240134 707162
rect 239514 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 240134 673174
rect 239514 672854 240134 672938
rect 239514 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 240134 672854
rect 239514 637174 240134 672618
rect 239514 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 240134 637174
rect 239514 636854 240134 636938
rect 239514 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 240134 636854
rect 239514 601174 240134 636618
rect 239514 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 240134 601174
rect 239514 600854 240134 600938
rect 239514 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 240134 600854
rect 239514 565174 240134 600618
rect 239514 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 240134 565174
rect 239514 564854 240134 564938
rect 239514 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 240134 564854
rect 239514 537993 240134 564618
rect 243234 676894 243854 709082
rect 243234 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 243854 676894
rect 243234 676574 243854 676658
rect 243234 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 243854 676574
rect 243234 640894 243854 676338
rect 243234 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 243854 640894
rect 243234 640574 243854 640658
rect 243234 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 243854 640574
rect 243234 604894 243854 640338
rect 243234 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 243854 604894
rect 243234 604574 243854 604658
rect 243234 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 243854 604574
rect 243234 568894 243854 604338
rect 243234 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 243854 568894
rect 243234 568574 243854 568658
rect 243234 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 243854 568574
rect 243234 537993 243854 568338
rect 246954 680614 247574 711002
rect 264954 710598 265574 711590
rect 264954 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 265574 710598
rect 264954 710278 265574 710362
rect 264954 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 265574 710278
rect 261234 708678 261854 709670
rect 261234 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 261854 708678
rect 261234 708358 261854 708442
rect 261234 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 261854 708358
rect 257514 706758 258134 707750
rect 257514 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 258134 706758
rect 257514 706438 258134 706522
rect 257514 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 258134 706438
rect 246954 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 247574 680614
rect 246954 680294 247574 680378
rect 246954 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 247574 680294
rect 246954 644614 247574 680058
rect 246954 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 247574 644614
rect 246954 644294 247574 644378
rect 246954 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 247574 644294
rect 246954 608614 247574 644058
rect 246954 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 247574 608614
rect 246954 608294 247574 608378
rect 246954 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 247574 608294
rect 246954 572614 247574 608058
rect 246954 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 247574 572614
rect 246954 572294 247574 572378
rect 246954 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 247574 572294
rect 246954 537993 247574 572058
rect 253794 704838 254414 705830
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 615454 254414 650898
rect 253794 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 254414 615454
rect 253794 615134 254414 615218
rect 253794 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 254414 615134
rect 253794 579454 254414 614898
rect 253794 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 254414 579454
rect 253794 579134 254414 579218
rect 253794 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 254414 579134
rect 253794 543454 254414 578898
rect 253794 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 254414 543454
rect 253794 543134 254414 543218
rect 253794 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 254414 543134
rect 253794 537993 254414 542898
rect 257514 691174 258134 706202
rect 257514 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 258134 691174
rect 257514 690854 258134 690938
rect 257514 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 258134 690854
rect 257514 655174 258134 690618
rect 257514 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 258134 655174
rect 257514 654854 258134 654938
rect 257514 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 258134 654854
rect 257514 619174 258134 654618
rect 257514 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 258134 619174
rect 257514 618854 258134 618938
rect 257514 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 258134 618854
rect 257514 583174 258134 618618
rect 257514 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 258134 583174
rect 257514 582854 258134 582938
rect 257514 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 258134 582854
rect 257514 547174 258134 582618
rect 257514 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 258134 547174
rect 257514 546854 258134 546938
rect 257514 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 258134 546854
rect 257514 537993 258134 546618
rect 261234 694894 261854 708122
rect 261234 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 261854 694894
rect 261234 694574 261854 694658
rect 261234 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 261854 694574
rect 261234 658894 261854 694338
rect 261234 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 261854 658894
rect 261234 658574 261854 658658
rect 261234 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 261854 658574
rect 261234 622894 261854 658338
rect 261234 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 261854 622894
rect 261234 622574 261854 622658
rect 261234 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 261854 622574
rect 261234 586894 261854 622338
rect 261234 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 261854 586894
rect 261234 586574 261854 586658
rect 261234 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 261854 586574
rect 261234 550894 261854 586338
rect 261234 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 261854 550894
rect 261234 550574 261854 550658
rect 261234 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 261854 550574
rect 261234 537993 261854 550338
rect 264954 698614 265574 710042
rect 282954 711558 283574 711590
rect 282954 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 283574 711558
rect 282954 711238 283574 711322
rect 282954 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 283574 711238
rect 279234 709638 279854 709670
rect 279234 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 279854 709638
rect 279234 709318 279854 709402
rect 279234 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 279854 709318
rect 275514 707718 276134 707750
rect 275514 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 276134 707718
rect 275514 707398 276134 707482
rect 275514 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 276134 707398
rect 264954 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 265574 698614
rect 264954 698294 265574 698378
rect 264954 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 265574 698294
rect 264954 662614 265574 698058
rect 264954 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 265574 662614
rect 264954 662294 265574 662378
rect 264954 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 265574 662294
rect 264954 626614 265574 662058
rect 264954 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 265574 626614
rect 264954 626294 265574 626378
rect 264954 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 265574 626294
rect 264954 590614 265574 626058
rect 264954 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 265574 590614
rect 264954 590294 265574 590378
rect 264954 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 265574 590294
rect 264954 554614 265574 590058
rect 264954 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 265574 554614
rect 264954 554294 265574 554378
rect 264954 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 265574 554294
rect 264954 537993 265574 554058
rect 271794 705798 272414 705830
rect 271794 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 272414 705798
rect 271794 705478 272414 705562
rect 271794 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 272414 705478
rect 271794 669454 272414 705242
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 633454 272414 668898
rect 271794 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 272414 633454
rect 271794 633134 272414 633218
rect 271794 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 272414 633134
rect 271794 597454 272414 632898
rect 271794 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 272414 597454
rect 271794 597134 272414 597218
rect 271794 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 272414 597134
rect 271794 561454 272414 596898
rect 271794 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 272414 561454
rect 271794 561134 272414 561218
rect 271794 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 272414 561134
rect 271794 537993 272414 560898
rect 275514 673174 276134 707162
rect 275514 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 276134 673174
rect 275514 672854 276134 672938
rect 275514 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 276134 672854
rect 275514 637174 276134 672618
rect 275514 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 276134 637174
rect 275514 636854 276134 636938
rect 275514 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 276134 636854
rect 275514 601174 276134 636618
rect 275514 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 276134 601174
rect 275514 600854 276134 600938
rect 275514 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 276134 600854
rect 275514 565174 276134 600618
rect 275514 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 276134 565174
rect 275514 564854 276134 564938
rect 275514 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 276134 564854
rect 275514 537993 276134 564618
rect 279234 676894 279854 709082
rect 279234 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 279854 676894
rect 279234 676574 279854 676658
rect 279234 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 279854 676574
rect 279234 640894 279854 676338
rect 279234 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 279854 640894
rect 279234 640574 279854 640658
rect 279234 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 279854 640574
rect 279234 604894 279854 640338
rect 279234 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 279854 604894
rect 279234 604574 279854 604658
rect 279234 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 279854 604574
rect 279234 568894 279854 604338
rect 279234 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 279854 568894
rect 279234 568574 279854 568658
rect 279234 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 279854 568574
rect 279234 537993 279854 568338
rect 282954 680614 283574 711002
rect 300954 710598 301574 711590
rect 300954 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 301574 710598
rect 300954 710278 301574 710362
rect 300954 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 301574 710278
rect 297234 708678 297854 709670
rect 297234 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 297854 708678
rect 297234 708358 297854 708442
rect 297234 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 297854 708358
rect 293514 706758 294134 707750
rect 293514 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 294134 706758
rect 293514 706438 294134 706522
rect 293514 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 294134 706438
rect 282954 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 283574 680614
rect 282954 680294 283574 680378
rect 282954 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 283574 680294
rect 282954 644614 283574 680058
rect 282954 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 283574 644614
rect 282954 644294 283574 644378
rect 282954 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 283574 644294
rect 282954 608614 283574 644058
rect 282954 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 283574 608614
rect 282954 608294 283574 608378
rect 282954 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 283574 608294
rect 282954 572614 283574 608058
rect 282954 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 283574 572614
rect 282954 572294 283574 572378
rect 282954 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 283574 572294
rect 282954 537993 283574 572058
rect 289794 704838 290414 705830
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 543454 290414 578898
rect 289794 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 290414 543454
rect 289794 543134 290414 543218
rect 289794 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 290414 543134
rect 289794 537993 290414 542898
rect 293514 691174 294134 706202
rect 293514 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 294134 691174
rect 293514 690854 294134 690938
rect 293514 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 294134 690854
rect 293514 655174 294134 690618
rect 293514 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 294134 655174
rect 293514 654854 294134 654938
rect 293514 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 294134 654854
rect 293514 619174 294134 654618
rect 293514 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 294134 619174
rect 293514 618854 294134 618938
rect 293514 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 294134 618854
rect 293514 583174 294134 618618
rect 293514 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 294134 583174
rect 293514 582854 294134 582938
rect 293514 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 294134 582854
rect 293514 547174 294134 582618
rect 293514 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 294134 547174
rect 293514 546854 294134 546938
rect 293514 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 294134 546854
rect 293514 537993 294134 546618
rect 297234 694894 297854 708122
rect 297234 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 297854 694894
rect 297234 694574 297854 694658
rect 297234 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 297854 694574
rect 297234 658894 297854 694338
rect 297234 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 297854 658894
rect 297234 658574 297854 658658
rect 297234 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 297854 658574
rect 297234 622894 297854 658338
rect 297234 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 297854 622894
rect 297234 622574 297854 622658
rect 297234 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 297854 622574
rect 297234 586894 297854 622338
rect 297234 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 297854 586894
rect 297234 586574 297854 586658
rect 297234 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 297854 586574
rect 297234 550894 297854 586338
rect 297234 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 297854 550894
rect 297234 550574 297854 550658
rect 297234 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 297854 550574
rect 297234 537993 297854 550338
rect 300954 698614 301574 710042
rect 318954 711558 319574 711590
rect 318954 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 319574 711558
rect 318954 711238 319574 711322
rect 318954 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 319574 711238
rect 315234 709638 315854 709670
rect 315234 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 315854 709638
rect 315234 709318 315854 709402
rect 315234 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 315854 709318
rect 311514 707718 312134 707750
rect 311514 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 312134 707718
rect 311514 707398 312134 707482
rect 311514 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 312134 707398
rect 300954 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 301574 698614
rect 300954 698294 301574 698378
rect 300954 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 301574 698294
rect 300954 662614 301574 698058
rect 300954 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 301574 662614
rect 300954 662294 301574 662378
rect 300954 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 301574 662294
rect 300954 626614 301574 662058
rect 300954 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 301574 626614
rect 300954 626294 301574 626378
rect 300954 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 301574 626294
rect 300954 590614 301574 626058
rect 300954 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 301574 590614
rect 300954 590294 301574 590378
rect 300954 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 301574 590294
rect 300954 554614 301574 590058
rect 300954 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 301574 554614
rect 300954 554294 301574 554378
rect 300954 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 301574 554294
rect 300954 537993 301574 554058
rect 307794 705798 308414 705830
rect 307794 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 308414 705798
rect 307794 705478 308414 705562
rect 307794 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 308414 705478
rect 307794 669454 308414 705242
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 633454 308414 668898
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 307794 597454 308414 632898
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 307794 561454 308414 596898
rect 307794 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 308414 561454
rect 307794 561134 308414 561218
rect 307794 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 308414 561134
rect 307794 537993 308414 560898
rect 311514 673174 312134 707162
rect 311514 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 312134 673174
rect 311514 672854 312134 672938
rect 311514 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 312134 672854
rect 311514 637174 312134 672618
rect 311514 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 312134 637174
rect 311514 636854 312134 636938
rect 311514 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 312134 636854
rect 311514 601174 312134 636618
rect 311514 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 312134 601174
rect 311514 600854 312134 600938
rect 311514 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 312134 600854
rect 311514 565174 312134 600618
rect 311514 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 312134 565174
rect 311514 564854 312134 564938
rect 311514 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 312134 564854
rect 311514 537993 312134 564618
rect 315234 676894 315854 709082
rect 315234 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 315854 676894
rect 315234 676574 315854 676658
rect 315234 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 315854 676574
rect 315234 640894 315854 676338
rect 315234 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 315854 640894
rect 315234 640574 315854 640658
rect 315234 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 315854 640574
rect 315234 604894 315854 640338
rect 315234 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 315854 604894
rect 315234 604574 315854 604658
rect 315234 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 315854 604574
rect 315234 568894 315854 604338
rect 315234 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 315854 568894
rect 315234 568574 315854 568658
rect 315234 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 315854 568574
rect 315234 537993 315854 568338
rect 318954 680614 319574 711002
rect 336954 710598 337574 711590
rect 336954 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 337574 710598
rect 336954 710278 337574 710362
rect 336954 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 337574 710278
rect 333234 708678 333854 709670
rect 333234 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 333854 708678
rect 333234 708358 333854 708442
rect 333234 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 333854 708358
rect 329514 706758 330134 707750
rect 329514 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 330134 706758
rect 329514 706438 330134 706522
rect 329514 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 330134 706438
rect 318954 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 319574 680614
rect 318954 680294 319574 680378
rect 318954 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 319574 680294
rect 318954 644614 319574 680058
rect 318954 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 319574 644614
rect 318954 644294 319574 644378
rect 318954 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 319574 644294
rect 318954 608614 319574 644058
rect 318954 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 319574 608614
rect 318954 608294 319574 608378
rect 318954 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 319574 608294
rect 318954 572614 319574 608058
rect 318954 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 319574 572614
rect 318954 572294 319574 572378
rect 318954 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 319574 572294
rect 318954 537993 319574 572058
rect 325794 704838 326414 705830
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 543454 326414 578898
rect 325794 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 326414 543454
rect 325794 543134 326414 543218
rect 325794 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 326414 543134
rect 325794 537993 326414 542898
rect 329514 691174 330134 706202
rect 329514 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 330134 691174
rect 329514 690854 330134 690938
rect 329514 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 330134 690854
rect 329514 655174 330134 690618
rect 329514 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 330134 655174
rect 329514 654854 330134 654938
rect 329514 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 330134 654854
rect 329514 619174 330134 654618
rect 329514 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 330134 619174
rect 329514 618854 330134 618938
rect 329514 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 330134 618854
rect 329514 583174 330134 618618
rect 329514 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 330134 583174
rect 329514 582854 330134 582938
rect 329514 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 330134 582854
rect 329514 547174 330134 582618
rect 329514 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 330134 547174
rect 329514 546854 330134 546938
rect 329514 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 330134 546854
rect 329514 537993 330134 546618
rect 333234 694894 333854 708122
rect 333234 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 333854 694894
rect 333234 694574 333854 694658
rect 333234 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 333854 694574
rect 333234 658894 333854 694338
rect 333234 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 333854 658894
rect 333234 658574 333854 658658
rect 333234 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 333854 658574
rect 333234 622894 333854 658338
rect 333234 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 333854 622894
rect 333234 622574 333854 622658
rect 333234 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 333854 622574
rect 333234 586894 333854 622338
rect 333234 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 333854 586894
rect 333234 586574 333854 586658
rect 333234 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 333854 586574
rect 333234 550894 333854 586338
rect 333234 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 333854 550894
rect 333234 550574 333854 550658
rect 333234 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 333854 550574
rect 333234 537993 333854 550338
rect 336954 698614 337574 710042
rect 354954 711558 355574 711590
rect 354954 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 355574 711558
rect 354954 711238 355574 711322
rect 354954 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 355574 711238
rect 351234 709638 351854 709670
rect 351234 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 351854 709638
rect 351234 709318 351854 709402
rect 351234 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 351854 709318
rect 347514 707718 348134 707750
rect 347514 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 348134 707718
rect 347514 707398 348134 707482
rect 347514 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 348134 707398
rect 336954 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 337574 698614
rect 336954 698294 337574 698378
rect 336954 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 337574 698294
rect 336954 662614 337574 698058
rect 336954 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 337574 662614
rect 336954 662294 337574 662378
rect 336954 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 337574 662294
rect 336954 626614 337574 662058
rect 336954 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 337574 626614
rect 336954 626294 337574 626378
rect 336954 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 337574 626294
rect 336954 590614 337574 626058
rect 336954 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 337574 590614
rect 336954 590294 337574 590378
rect 336954 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 337574 590294
rect 336954 554614 337574 590058
rect 336954 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 337574 554614
rect 336954 554294 337574 554378
rect 336954 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 337574 554294
rect 336954 537993 337574 554058
rect 343794 705798 344414 705830
rect 343794 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 344414 705798
rect 343794 705478 344414 705562
rect 343794 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 344414 705478
rect 343794 669454 344414 705242
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 633454 344414 668898
rect 343794 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 344414 633454
rect 343794 633134 344414 633218
rect 343794 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 344414 633134
rect 343794 597454 344414 632898
rect 343794 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 344414 597454
rect 343794 597134 344414 597218
rect 343794 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 344414 597134
rect 343794 561454 344414 596898
rect 343794 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 344414 561454
rect 343794 561134 344414 561218
rect 343794 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 344414 561134
rect 343794 537993 344414 560898
rect 347514 673174 348134 707162
rect 347514 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 348134 673174
rect 347514 672854 348134 672938
rect 347514 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 348134 672854
rect 347514 637174 348134 672618
rect 347514 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 348134 637174
rect 347514 636854 348134 636938
rect 347514 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 348134 636854
rect 347514 601174 348134 636618
rect 347514 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 348134 601174
rect 347514 600854 348134 600938
rect 347514 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 348134 600854
rect 347514 565174 348134 600618
rect 347514 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 348134 565174
rect 347514 564854 348134 564938
rect 347514 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 348134 564854
rect 347514 537993 348134 564618
rect 351234 676894 351854 709082
rect 351234 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 351854 676894
rect 351234 676574 351854 676658
rect 351234 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 351854 676574
rect 351234 640894 351854 676338
rect 351234 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 351854 640894
rect 351234 640574 351854 640658
rect 351234 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 351854 640574
rect 351234 604894 351854 640338
rect 351234 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 351854 604894
rect 351234 604574 351854 604658
rect 351234 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 351854 604574
rect 351234 568894 351854 604338
rect 351234 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 351854 568894
rect 351234 568574 351854 568658
rect 351234 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 351854 568574
rect 351234 537993 351854 568338
rect 354954 680614 355574 711002
rect 372954 710598 373574 711590
rect 372954 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 373574 710598
rect 372954 710278 373574 710362
rect 372954 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 373574 710278
rect 369234 708678 369854 709670
rect 369234 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 369854 708678
rect 369234 708358 369854 708442
rect 369234 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 369854 708358
rect 365514 706758 366134 707750
rect 365514 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 366134 706758
rect 365514 706438 366134 706522
rect 365514 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 366134 706438
rect 354954 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 355574 680614
rect 354954 680294 355574 680378
rect 354954 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 355574 680294
rect 354954 644614 355574 680058
rect 354954 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 355574 644614
rect 354954 644294 355574 644378
rect 354954 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 355574 644294
rect 354954 608614 355574 644058
rect 354954 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 355574 608614
rect 354954 608294 355574 608378
rect 354954 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 355574 608294
rect 354954 572614 355574 608058
rect 354954 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 355574 572614
rect 354954 572294 355574 572378
rect 354954 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 355574 572294
rect 353339 545188 353405 545189
rect 353339 545124 353340 545188
rect 353404 545124 353405 545188
rect 353339 545123 353405 545124
rect 352051 538252 352117 538253
rect 352051 538188 352052 538252
rect 352116 538188 352117 538252
rect 352051 538187 352117 538188
rect 200132 533430 200682 533490
rect 200132 533428 200133 533430
rect 200067 533427 200133 533428
rect 219568 525454 219888 525486
rect 219568 525218 219610 525454
rect 219846 525218 219888 525454
rect 219568 525134 219888 525218
rect 219568 524898 219610 525134
rect 219846 524898 219888 525134
rect 219568 524866 219888 524898
rect 250288 525454 250608 525486
rect 250288 525218 250330 525454
rect 250566 525218 250608 525454
rect 250288 525134 250608 525218
rect 250288 524898 250330 525134
rect 250566 524898 250608 525134
rect 250288 524866 250608 524898
rect 281008 525454 281328 525486
rect 281008 525218 281050 525454
rect 281286 525218 281328 525454
rect 281008 525134 281328 525218
rect 281008 524898 281050 525134
rect 281286 524898 281328 525134
rect 281008 524866 281328 524898
rect 311728 525454 312048 525486
rect 311728 525218 311770 525454
rect 312006 525218 312048 525454
rect 311728 525134 312048 525218
rect 311728 524898 311770 525134
rect 312006 524898 312048 525134
rect 311728 524866 312048 524898
rect 342448 525454 342768 525486
rect 342448 525218 342490 525454
rect 342726 525218 342768 525454
rect 342448 525134 342768 525218
rect 342448 524898 342490 525134
rect 342726 524898 342768 525134
rect 342448 524866 342768 524898
rect 204208 507454 204528 507486
rect 204208 507218 204250 507454
rect 204486 507218 204528 507454
rect 204208 507134 204528 507218
rect 204208 506898 204250 507134
rect 204486 506898 204528 507134
rect 204208 506866 204528 506898
rect 234928 507454 235248 507486
rect 234928 507218 234970 507454
rect 235206 507218 235248 507454
rect 234928 507134 235248 507218
rect 234928 506898 234970 507134
rect 235206 506898 235248 507134
rect 234928 506866 235248 506898
rect 265648 507454 265968 507486
rect 265648 507218 265690 507454
rect 265926 507218 265968 507454
rect 265648 507134 265968 507218
rect 265648 506898 265690 507134
rect 265926 506898 265968 507134
rect 265648 506866 265968 506898
rect 296368 507454 296688 507486
rect 296368 507218 296410 507454
rect 296646 507218 296688 507454
rect 296368 507134 296688 507218
rect 296368 506898 296410 507134
rect 296646 506898 296688 507134
rect 296368 506866 296688 506898
rect 327088 507454 327408 507486
rect 327088 507218 327130 507454
rect 327366 507218 327408 507454
rect 327088 507134 327408 507218
rect 327088 506898 327130 507134
rect 327366 506898 327408 507134
rect 327088 506866 327408 506898
rect 219568 489454 219888 489486
rect 219568 489218 219610 489454
rect 219846 489218 219888 489454
rect 219568 489134 219888 489218
rect 219568 488898 219610 489134
rect 219846 488898 219888 489134
rect 219568 488866 219888 488898
rect 250288 489454 250608 489486
rect 250288 489218 250330 489454
rect 250566 489218 250608 489454
rect 250288 489134 250608 489218
rect 250288 488898 250330 489134
rect 250566 488898 250608 489134
rect 250288 488866 250608 488898
rect 281008 489454 281328 489486
rect 281008 489218 281050 489454
rect 281286 489218 281328 489454
rect 281008 489134 281328 489218
rect 281008 488898 281050 489134
rect 281286 488898 281328 489134
rect 281008 488866 281328 488898
rect 311728 489454 312048 489486
rect 311728 489218 311770 489454
rect 312006 489218 312048 489454
rect 311728 489134 312048 489218
rect 311728 488898 311770 489134
rect 312006 488898 312048 489134
rect 311728 488866 312048 488898
rect 342448 489454 342768 489486
rect 342448 489218 342490 489454
rect 342726 489218 342768 489454
rect 342448 489134 342768 489218
rect 342448 488898 342490 489134
rect 342726 488898 342768 489134
rect 342448 488866 342768 488898
rect 204208 471454 204528 471486
rect 204208 471218 204250 471454
rect 204486 471218 204528 471454
rect 204208 471134 204528 471218
rect 204208 470898 204250 471134
rect 204486 470898 204528 471134
rect 204208 470866 204528 470898
rect 234928 471454 235248 471486
rect 234928 471218 234970 471454
rect 235206 471218 235248 471454
rect 234928 471134 235248 471218
rect 234928 470898 234970 471134
rect 235206 470898 235248 471134
rect 234928 470866 235248 470898
rect 265648 471454 265968 471486
rect 265648 471218 265690 471454
rect 265926 471218 265968 471454
rect 265648 471134 265968 471218
rect 265648 470898 265690 471134
rect 265926 470898 265968 471134
rect 265648 470866 265968 470898
rect 296368 471454 296688 471486
rect 296368 471218 296410 471454
rect 296646 471218 296688 471454
rect 296368 471134 296688 471218
rect 296368 470898 296410 471134
rect 296646 470898 296688 471134
rect 296368 470866 296688 470898
rect 327088 471454 327408 471486
rect 327088 471218 327130 471454
rect 327366 471218 327408 471454
rect 327088 471134 327408 471218
rect 327088 470898 327130 471134
rect 327366 470898 327408 471134
rect 327088 470866 327408 470898
rect 219568 453454 219888 453486
rect 219568 453218 219610 453454
rect 219846 453218 219888 453454
rect 219568 453134 219888 453218
rect 219568 452898 219610 453134
rect 219846 452898 219888 453134
rect 219568 452866 219888 452898
rect 250288 453454 250608 453486
rect 250288 453218 250330 453454
rect 250566 453218 250608 453454
rect 250288 453134 250608 453218
rect 250288 452898 250330 453134
rect 250566 452898 250608 453134
rect 250288 452866 250608 452898
rect 281008 453454 281328 453486
rect 281008 453218 281050 453454
rect 281286 453218 281328 453454
rect 281008 453134 281328 453218
rect 281008 452898 281050 453134
rect 281286 452898 281328 453134
rect 281008 452866 281328 452898
rect 311728 453454 312048 453486
rect 311728 453218 311770 453454
rect 312006 453218 312048 453454
rect 311728 453134 312048 453218
rect 311728 452898 311770 453134
rect 312006 452898 312048 453134
rect 311728 452866 312048 452898
rect 342448 453454 342768 453486
rect 342448 453218 342490 453454
rect 342726 453218 342768 453454
rect 342448 453134 342768 453218
rect 342448 452898 342490 453134
rect 342726 452898 342768 453134
rect 342448 452866 342768 452898
rect 204208 435454 204528 435486
rect 204208 435218 204250 435454
rect 204486 435218 204528 435454
rect 204208 435134 204528 435218
rect 204208 434898 204250 435134
rect 204486 434898 204528 435134
rect 204208 434866 204528 434898
rect 234928 435454 235248 435486
rect 234928 435218 234970 435454
rect 235206 435218 235248 435454
rect 234928 435134 235248 435218
rect 234928 434898 234970 435134
rect 235206 434898 235248 435134
rect 234928 434866 235248 434898
rect 265648 435454 265968 435486
rect 265648 435218 265690 435454
rect 265926 435218 265968 435454
rect 265648 435134 265968 435218
rect 265648 434898 265690 435134
rect 265926 434898 265968 435134
rect 265648 434866 265968 434898
rect 296368 435454 296688 435486
rect 296368 435218 296410 435454
rect 296646 435218 296688 435454
rect 296368 435134 296688 435218
rect 296368 434898 296410 435134
rect 296646 434898 296688 435134
rect 296368 434866 296688 434898
rect 327088 435454 327408 435486
rect 327088 435218 327130 435454
rect 327366 435218 327408 435454
rect 327088 435134 327408 435218
rect 327088 434898 327130 435134
rect 327366 434898 327408 435134
rect 327088 434866 327408 434898
rect 219568 417454 219888 417486
rect 219568 417218 219610 417454
rect 219846 417218 219888 417454
rect 219568 417134 219888 417218
rect 219568 416898 219610 417134
rect 219846 416898 219888 417134
rect 219568 416866 219888 416898
rect 250288 417454 250608 417486
rect 250288 417218 250330 417454
rect 250566 417218 250608 417454
rect 250288 417134 250608 417218
rect 250288 416898 250330 417134
rect 250566 416898 250608 417134
rect 250288 416866 250608 416898
rect 281008 417454 281328 417486
rect 281008 417218 281050 417454
rect 281286 417218 281328 417454
rect 281008 417134 281328 417218
rect 281008 416898 281050 417134
rect 281286 416898 281328 417134
rect 281008 416866 281328 416898
rect 311728 417454 312048 417486
rect 311728 417218 311770 417454
rect 312006 417218 312048 417454
rect 311728 417134 312048 417218
rect 311728 416898 311770 417134
rect 312006 416898 312048 417134
rect 311728 416866 312048 416898
rect 342448 417454 342768 417486
rect 342448 417218 342490 417454
rect 342726 417218 342768 417454
rect 342448 417134 342768 417218
rect 342448 416898 342490 417134
rect 342726 416898 342768 417134
rect 342448 416866 342768 416898
rect 204208 399454 204528 399486
rect 204208 399218 204250 399454
rect 204486 399218 204528 399454
rect 204208 399134 204528 399218
rect 204208 398898 204250 399134
rect 204486 398898 204528 399134
rect 204208 398866 204528 398898
rect 234928 399454 235248 399486
rect 234928 399218 234970 399454
rect 235206 399218 235248 399454
rect 234928 399134 235248 399218
rect 234928 398898 234970 399134
rect 235206 398898 235248 399134
rect 234928 398866 235248 398898
rect 265648 399454 265968 399486
rect 265648 399218 265690 399454
rect 265926 399218 265968 399454
rect 265648 399134 265968 399218
rect 265648 398898 265690 399134
rect 265926 398898 265968 399134
rect 265648 398866 265968 398898
rect 296368 399454 296688 399486
rect 296368 399218 296410 399454
rect 296646 399218 296688 399454
rect 296368 399134 296688 399218
rect 296368 398898 296410 399134
rect 296646 398898 296688 399134
rect 296368 398866 296688 398898
rect 327088 399454 327408 399486
rect 327088 399218 327130 399454
rect 327366 399218 327408 399454
rect 327088 399134 327408 399218
rect 327088 398898 327130 399134
rect 327366 398898 327408 399134
rect 327088 398866 327408 398898
rect 219568 381454 219888 381486
rect 219568 381218 219610 381454
rect 219846 381218 219888 381454
rect 200067 381172 200133 381173
rect 200067 381108 200068 381172
rect 200132 381170 200133 381172
rect 200132 381110 200314 381170
rect 200132 381108 200133 381110
rect 200067 381107 200133 381108
rect 200254 380490 200314 381110
rect 219568 381134 219888 381218
rect 219568 380898 219610 381134
rect 219846 380898 219888 381134
rect 219568 380866 219888 380898
rect 250288 381454 250608 381486
rect 250288 381218 250330 381454
rect 250566 381218 250608 381454
rect 250288 381134 250608 381218
rect 250288 380898 250330 381134
rect 250566 380898 250608 381134
rect 250288 380866 250608 380898
rect 281008 381454 281328 381486
rect 281008 381218 281050 381454
rect 281286 381218 281328 381454
rect 281008 381134 281328 381218
rect 281008 380898 281050 381134
rect 281286 380898 281328 381134
rect 281008 380866 281328 380898
rect 311728 381454 312048 381486
rect 311728 381218 311770 381454
rect 312006 381218 312048 381454
rect 311728 381134 312048 381218
rect 311728 380898 311770 381134
rect 312006 380898 312048 381134
rect 311728 380866 312048 380898
rect 342448 381454 342768 381486
rect 342448 381218 342490 381454
rect 342726 381218 342768 381454
rect 342448 381134 342768 381218
rect 342448 380898 342490 381134
rect 342726 380898 342768 381134
rect 342448 380866 342768 380898
rect 200254 380430 200682 380490
rect 199515 353564 199581 353565
rect 199515 353500 199516 353564
rect 199580 353500 199581 353564
rect 199515 353499 199581 353500
rect 199794 345454 200414 375600
rect 199794 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 200414 345454
rect 199794 345134 200414 345218
rect 199794 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 200414 345134
rect 198595 314804 198661 314805
rect 198595 314740 198596 314804
rect 198660 314740 198661 314804
rect 198595 314739 198661 314740
rect 198598 278085 198658 314739
rect 199794 309454 200414 344898
rect 200622 312493 200682 380430
rect 203514 349174 204134 375600
rect 203514 348938 203546 349174
rect 203782 348938 203866 349174
rect 204102 348938 204134 349174
rect 203514 348854 204134 348938
rect 203514 348618 203546 348854
rect 203782 348618 203866 348854
rect 204102 348618 204134 348854
rect 202643 337652 202709 337653
rect 202643 337588 202644 337652
rect 202708 337588 202709 337652
rect 202643 337587 202709 337588
rect 200619 312492 200685 312493
rect 200619 312428 200620 312492
rect 200684 312428 200685 312492
rect 200619 312427 200685 312428
rect 199794 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 200414 309454
rect 199794 309134 200414 309218
rect 199794 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 200414 309134
rect 199331 287468 199397 287469
rect 199331 287404 199332 287468
rect 199396 287404 199397 287468
rect 199331 287403 199397 287404
rect 198779 284476 198845 284477
rect 198779 284412 198780 284476
rect 198844 284412 198845 284476
rect 198779 284411 198845 284412
rect 198782 279445 198842 284411
rect 198779 279444 198845 279445
rect 198779 279380 198780 279444
rect 198844 279380 198845 279444
rect 198779 279379 198845 279380
rect 198779 279308 198845 279309
rect 198779 279244 198780 279308
rect 198844 279244 198845 279308
rect 198779 279243 198845 279244
rect 198595 278084 198661 278085
rect 198595 278020 198596 278084
rect 198660 278020 198661 278084
rect 198595 278019 198661 278020
rect 198782 265573 198842 279243
rect 199334 271149 199394 287403
rect 199794 286182 200414 308898
rect 200619 294540 200685 294541
rect 200619 294476 200620 294540
rect 200684 294476 200685 294540
rect 200619 294475 200685 294476
rect 200622 285701 200682 294475
rect 200619 285700 200685 285701
rect 200619 285636 200620 285700
rect 200684 285636 200685 285700
rect 200619 285635 200685 285636
rect 201355 283932 201421 283933
rect 201355 283868 201356 283932
rect 201420 283868 201421 283932
rect 201355 283867 201421 283868
rect 199331 271148 199397 271149
rect 199331 271084 199332 271148
rect 199396 271084 199397 271148
rect 199331 271083 199397 271084
rect 198779 265572 198845 265573
rect 198779 265508 198780 265572
rect 198844 265508 198845 265572
rect 198779 265507 198845 265508
rect 199331 263124 199397 263125
rect 199331 263060 199332 263124
rect 199396 263060 199397 263124
rect 199331 263059 199397 263060
rect 197859 252652 197925 252653
rect 197859 252588 197860 252652
rect 197924 252588 197925 252652
rect 197859 252587 197925 252588
rect 197123 205596 197189 205597
rect 197123 205532 197124 205596
rect 197188 205532 197189 205596
rect 197123 205531 197189 205532
rect 199334 202333 199394 263059
rect 199794 237454 200414 238182
rect 199794 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 200414 237454
rect 199794 237134 200414 237218
rect 199794 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 200414 237134
rect 199331 202332 199397 202333
rect 199331 202268 199332 202332
rect 199396 202268 199397 202332
rect 199331 202267 199397 202268
rect 192954 194378 192986 194614
rect 193222 194378 193306 194614
rect 193542 194378 193574 194614
rect 192954 194294 193574 194378
rect 192954 194058 192986 194294
rect 193222 194058 193306 194294
rect 193542 194058 193574 194294
rect 192954 158614 193574 194058
rect 192954 158378 192986 158614
rect 193222 158378 193306 158614
rect 193542 158378 193574 158614
rect 192954 158294 193574 158378
rect 192954 158058 192986 158294
rect 193222 158058 193306 158294
rect 193542 158058 193574 158294
rect 192954 122614 193574 158058
rect 192954 122378 192986 122614
rect 193222 122378 193306 122614
rect 193542 122378 193574 122614
rect 192954 122294 193574 122378
rect 192954 122058 192986 122294
rect 193222 122058 193306 122294
rect 193542 122058 193574 122294
rect 192954 86614 193574 122058
rect 192954 86378 192986 86614
rect 193222 86378 193306 86614
rect 193542 86378 193574 86614
rect 192954 86294 193574 86378
rect 192954 86058 192986 86294
rect 193222 86058 193306 86294
rect 193542 86058 193574 86294
rect 192954 50614 193574 86058
rect 192954 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 193574 50614
rect 192954 50294 193574 50378
rect 192954 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 193574 50294
rect 189947 17372 190013 17373
rect 189947 17308 189948 17372
rect 190012 17308 190013 17372
rect 189947 17307 190013 17308
rect 189234 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 189854 10894
rect 189234 10574 189854 10658
rect 189234 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 189854 10574
rect 189234 -4186 189854 10338
rect 189234 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 189854 -4186
rect 189234 -4506 189854 -4422
rect 189234 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 189854 -4506
rect 189234 -5734 189854 -4742
rect 192954 14614 193574 50058
rect 192954 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 193574 14614
rect 192954 14294 193574 14378
rect 192954 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 193574 14294
rect 174954 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 175574 -7066
rect 174954 -7386 175574 -7302
rect 174954 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 175574 -7386
rect 174954 -7654 175574 -7622
rect 192954 -6106 193574 14058
rect 199794 201454 200414 236898
rect 199794 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 200414 201454
rect 199794 201134 200414 201218
rect 199794 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 200414 201134
rect 199794 165454 200414 200898
rect 199794 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 200414 165454
rect 199794 165134 200414 165218
rect 199794 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 200414 165134
rect 199794 129454 200414 164898
rect 199794 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 200414 129454
rect 199794 129134 200414 129218
rect 199794 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 200414 129134
rect 199794 93454 200414 128898
rect 201358 95165 201418 283867
rect 202646 240141 202706 337587
rect 203514 313174 204134 348618
rect 203514 312938 203546 313174
rect 203782 312938 203866 313174
rect 204102 312938 204134 313174
rect 203514 312854 204134 312938
rect 203514 312618 203546 312854
rect 203782 312618 203866 312854
rect 204102 312618 204134 312854
rect 203195 295356 203261 295357
rect 203195 295292 203196 295356
rect 203260 295292 203261 295356
rect 203195 295291 203261 295292
rect 203198 240141 203258 295291
rect 203514 286182 204134 312618
rect 207234 352894 207854 375600
rect 207234 352658 207266 352894
rect 207502 352658 207586 352894
rect 207822 352658 207854 352894
rect 207234 352574 207854 352658
rect 207234 352338 207266 352574
rect 207502 352338 207586 352574
rect 207822 352338 207854 352574
rect 207234 316894 207854 352338
rect 210954 356614 211574 375600
rect 210954 356378 210986 356614
rect 211222 356378 211306 356614
rect 211542 356378 211574 356614
rect 210954 356294 211574 356378
rect 210954 356058 210986 356294
rect 211222 356058 211306 356294
rect 211542 356058 211574 356294
rect 210739 338740 210805 338741
rect 210739 338676 210740 338740
rect 210804 338676 210805 338740
rect 210739 338675 210805 338676
rect 207234 316658 207266 316894
rect 207502 316658 207586 316894
rect 207822 316658 207854 316894
rect 207234 316574 207854 316658
rect 207234 316338 207266 316574
rect 207502 316338 207586 316574
rect 207822 316338 207854 316574
rect 206875 296308 206941 296309
rect 206875 296244 206876 296308
rect 206940 296244 206941 296308
rect 206875 296243 206941 296244
rect 204408 255454 204728 255486
rect 204408 255218 204450 255454
rect 204686 255218 204728 255454
rect 204408 255134 204728 255218
rect 204408 254898 204450 255134
rect 204686 254898 204728 255134
rect 204408 254866 204728 254898
rect 202643 240140 202709 240141
rect 202643 240076 202644 240140
rect 202708 240076 202709 240140
rect 202643 240075 202709 240076
rect 203195 240140 203261 240141
rect 203195 240076 203196 240140
rect 203260 240076 203261 240140
rect 203195 240075 203261 240076
rect 206878 238645 206938 296243
rect 207234 286182 207854 316338
rect 207979 305828 208045 305829
rect 207979 305764 207980 305828
rect 208044 305764 208045 305828
rect 207979 305763 208045 305764
rect 207982 240005 208042 305763
rect 209635 285700 209701 285701
rect 209635 285636 209636 285700
rect 209700 285636 209701 285700
rect 209635 285635 209701 285636
rect 208163 284204 208229 284205
rect 208163 284140 208164 284204
rect 208228 284140 208229 284204
rect 208163 284139 208229 284140
rect 208166 240141 208226 284139
rect 208163 240140 208229 240141
rect 208163 240076 208164 240140
rect 208228 240076 208229 240140
rect 208163 240075 208229 240076
rect 207979 240004 208045 240005
rect 207979 239940 207980 240004
rect 208044 239940 208045 240004
rect 207979 239939 208045 239940
rect 206875 238644 206941 238645
rect 206875 238580 206876 238644
rect 206940 238580 206941 238644
rect 206875 238579 206941 238580
rect 203514 205174 204134 238182
rect 203514 204938 203546 205174
rect 203782 204938 203866 205174
rect 204102 204938 204134 205174
rect 203514 204854 204134 204938
rect 203514 204618 203546 204854
rect 203782 204618 203866 204854
rect 204102 204618 204134 204854
rect 203514 169174 204134 204618
rect 203514 168938 203546 169174
rect 203782 168938 203866 169174
rect 204102 168938 204134 169174
rect 203514 168854 204134 168938
rect 203514 168618 203546 168854
rect 203782 168618 203866 168854
rect 204102 168618 204134 168854
rect 203514 133174 204134 168618
rect 203514 132938 203546 133174
rect 203782 132938 203866 133174
rect 204102 132938 204134 133174
rect 203514 132854 204134 132938
rect 203514 132618 203546 132854
rect 203782 132618 203866 132854
rect 204102 132618 204134 132854
rect 203514 97174 204134 132618
rect 203514 96938 203546 97174
rect 203782 96938 203866 97174
rect 204102 96938 204134 97174
rect 203514 96854 204134 96938
rect 203514 96618 203546 96854
rect 203782 96618 203866 96854
rect 204102 96618 204134 96854
rect 201355 95164 201421 95165
rect 201355 95100 201356 95164
rect 201420 95100 201421 95164
rect 201355 95099 201421 95100
rect 199794 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 200414 93454
rect 199794 93134 200414 93218
rect 199794 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 200414 93134
rect 199794 57454 200414 92898
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 199794 57134 200414 57218
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 199794 21454 200414 56898
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -1306 200414 20898
rect 199794 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 200414 -1306
rect 199794 -1626 200414 -1542
rect 199794 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 200414 -1626
rect 199794 -1894 200414 -1862
rect 203514 61174 204134 96618
rect 203514 60938 203546 61174
rect 203782 60938 203866 61174
rect 204102 60938 204134 61174
rect 203514 60854 204134 60938
rect 203514 60618 203546 60854
rect 203782 60618 203866 60854
rect 204102 60618 204134 60854
rect 203514 25174 204134 60618
rect 203514 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 204134 25174
rect 203514 24854 204134 24938
rect 203514 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 204134 24854
rect 203514 -3226 204134 24618
rect 203514 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 204134 -3226
rect 203514 -3546 204134 -3462
rect 203514 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 204134 -3546
rect 203514 -3814 204134 -3782
rect 207234 208894 207854 238182
rect 209638 211309 209698 285635
rect 210742 240141 210802 338675
rect 210954 320614 211574 356058
rect 217794 363454 218414 375600
rect 217794 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 218414 363454
rect 217794 363134 218414 363218
rect 217794 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 218414 363134
rect 211659 351388 211725 351389
rect 211659 351324 211660 351388
rect 211724 351324 211725 351388
rect 211659 351323 211725 351324
rect 210954 320378 210986 320614
rect 211222 320378 211306 320614
rect 211542 320378 211574 320614
rect 210954 320294 211574 320378
rect 210954 320058 210986 320294
rect 211222 320058 211306 320294
rect 211542 320058 211574 320294
rect 210954 286182 211574 320058
rect 210739 240140 210805 240141
rect 210739 240076 210740 240140
rect 210804 240076 210805 240140
rect 210739 240075 210805 240076
rect 210954 212614 211574 238182
rect 210954 212378 210986 212614
rect 211222 212378 211306 212614
rect 211542 212378 211574 212614
rect 210954 212294 211574 212378
rect 210954 212058 210986 212294
rect 211222 212058 211306 212294
rect 211542 212058 211574 212294
rect 209635 211308 209701 211309
rect 209635 211244 209636 211308
rect 209700 211244 209701 211308
rect 209635 211243 209701 211244
rect 207234 208658 207266 208894
rect 207502 208658 207586 208894
rect 207822 208658 207854 208894
rect 207234 208574 207854 208658
rect 207234 208338 207266 208574
rect 207502 208338 207586 208574
rect 207822 208338 207854 208574
rect 207234 172894 207854 208338
rect 207234 172658 207266 172894
rect 207502 172658 207586 172894
rect 207822 172658 207854 172894
rect 207234 172574 207854 172658
rect 207234 172338 207266 172574
rect 207502 172338 207586 172574
rect 207822 172338 207854 172574
rect 207234 136894 207854 172338
rect 207234 136658 207266 136894
rect 207502 136658 207586 136894
rect 207822 136658 207854 136894
rect 207234 136574 207854 136658
rect 207234 136338 207266 136574
rect 207502 136338 207586 136574
rect 207822 136338 207854 136574
rect 207234 100894 207854 136338
rect 207234 100658 207266 100894
rect 207502 100658 207586 100894
rect 207822 100658 207854 100894
rect 207234 100574 207854 100658
rect 207234 100338 207266 100574
rect 207502 100338 207586 100574
rect 207822 100338 207854 100574
rect 207234 64894 207854 100338
rect 207234 64658 207266 64894
rect 207502 64658 207586 64894
rect 207822 64658 207854 64894
rect 207234 64574 207854 64658
rect 207234 64338 207266 64574
rect 207502 64338 207586 64574
rect 207822 64338 207854 64574
rect 207234 28894 207854 64338
rect 207234 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 207854 28894
rect 207234 28574 207854 28658
rect 207234 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 207854 28574
rect 207234 -5146 207854 28338
rect 207234 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 207854 -5146
rect 207234 -5466 207854 -5382
rect 207234 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 207854 -5466
rect 207234 -5734 207854 -5702
rect 210954 176614 211574 212058
rect 211662 197301 211722 351323
rect 212579 339692 212645 339693
rect 212579 339628 212580 339692
rect 212644 339628 212645 339692
rect 212579 339627 212645 339628
rect 212582 238645 212642 339627
rect 214419 334660 214485 334661
rect 214419 334596 214420 334660
rect 214484 334596 214485 334660
rect 214419 334595 214485 334596
rect 213867 312492 213933 312493
rect 213867 312428 213868 312492
rect 213932 312428 213933 312492
rect 213867 312427 213933 312428
rect 213870 240141 213930 312427
rect 214422 240141 214482 334595
rect 217794 327454 218414 362898
rect 217794 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 218414 327454
rect 217794 327134 218414 327218
rect 217794 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 218414 327134
rect 215339 314124 215405 314125
rect 215339 314060 215340 314124
rect 215404 314060 215405 314124
rect 215339 314059 215405 314060
rect 215342 285701 215402 314059
rect 217547 291820 217613 291821
rect 217547 291756 217548 291820
rect 217612 291756 217613 291820
rect 217547 291755 217613 291756
rect 215339 285700 215405 285701
rect 215339 285636 215340 285700
rect 215404 285636 215405 285700
rect 215339 285635 215405 285636
rect 216443 284068 216509 284069
rect 216443 284004 216444 284068
rect 216508 284004 216509 284068
rect 216443 284003 216509 284004
rect 215523 283932 215589 283933
rect 215523 283868 215524 283932
rect 215588 283868 215589 283932
rect 215523 283867 215589 283868
rect 213867 240140 213933 240141
rect 213867 240076 213868 240140
rect 213932 240076 213933 240140
rect 213867 240075 213933 240076
rect 214419 240140 214485 240141
rect 214419 240076 214420 240140
rect 214484 240076 214485 240140
rect 214419 240075 214485 240076
rect 212579 238644 212645 238645
rect 212579 238580 212580 238644
rect 212644 238580 212645 238644
rect 212579 238579 212645 238580
rect 215155 222324 215221 222325
rect 215155 222260 215156 222324
rect 215220 222260 215221 222324
rect 215155 222259 215221 222260
rect 211659 197300 211725 197301
rect 211659 197236 211660 197300
rect 211724 197236 211725 197300
rect 211659 197235 211725 197236
rect 212395 197300 212461 197301
rect 212395 197236 212396 197300
rect 212460 197236 212461 197300
rect 212395 197235 212461 197236
rect 212398 196621 212458 197235
rect 212395 196620 212461 196621
rect 212395 196556 212396 196620
rect 212460 196556 212461 196620
rect 212395 196555 212461 196556
rect 210954 176378 210986 176614
rect 211222 176378 211306 176614
rect 211542 176378 211574 176614
rect 210954 176294 211574 176378
rect 210954 176058 210986 176294
rect 211222 176058 211306 176294
rect 211542 176058 211574 176294
rect 210954 140614 211574 176058
rect 210954 140378 210986 140614
rect 211222 140378 211306 140614
rect 211542 140378 211574 140614
rect 210954 140294 211574 140378
rect 210954 140058 210986 140294
rect 211222 140058 211306 140294
rect 211542 140058 211574 140294
rect 210954 104614 211574 140058
rect 210954 104378 210986 104614
rect 211222 104378 211306 104614
rect 211542 104378 211574 104614
rect 210954 104294 211574 104378
rect 210954 104058 210986 104294
rect 211222 104058 211306 104294
rect 211542 104058 211574 104294
rect 210954 68614 211574 104058
rect 215158 90405 215218 222259
rect 215526 214573 215586 283867
rect 215523 214572 215589 214573
rect 215523 214508 215524 214572
rect 215588 214508 215589 214572
rect 215523 214507 215589 214508
rect 216446 188461 216506 284003
rect 217550 240141 217610 291755
rect 217794 291454 218414 326898
rect 221514 367174 222134 375600
rect 225234 370894 225854 375600
rect 225234 370658 225266 370894
rect 225502 370658 225586 370894
rect 225822 370658 225854 370894
rect 225234 370574 225854 370658
rect 225234 370338 225266 370574
rect 225502 370338 225586 370574
rect 225822 370338 225854 370574
rect 224907 367844 224973 367845
rect 224907 367780 224908 367844
rect 224972 367780 224973 367844
rect 224907 367779 224973 367780
rect 221514 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 222134 367174
rect 221514 366854 222134 366938
rect 221514 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 222134 366854
rect 221514 331174 222134 366618
rect 222331 334252 222397 334253
rect 222331 334188 222332 334252
rect 222396 334188 222397 334252
rect 222331 334187 222397 334188
rect 221514 330938 221546 331174
rect 221782 330938 221866 331174
rect 222102 330938 222134 331174
rect 221514 330854 222134 330938
rect 221514 330618 221546 330854
rect 221782 330618 221866 330854
rect 222102 330618 222134 330854
rect 219203 296172 219269 296173
rect 219203 296108 219204 296172
rect 219268 296108 219269 296172
rect 219203 296107 219269 296108
rect 217794 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 218414 291454
rect 217794 291134 218414 291218
rect 217794 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 218414 291134
rect 217794 286182 218414 290898
rect 219206 240141 219266 296107
rect 221514 295174 222134 330618
rect 221514 294938 221546 295174
rect 221782 294938 221866 295174
rect 222102 294938 222134 295174
rect 221514 294854 222134 294938
rect 221514 294618 221546 294854
rect 221782 294618 221866 294854
rect 222102 294618 222134 294854
rect 221043 287332 221109 287333
rect 221043 287268 221044 287332
rect 221108 287268 221109 287332
rect 221043 287267 221109 287268
rect 220859 283932 220925 283933
rect 220859 283868 220860 283932
rect 220924 283868 220925 283932
rect 220859 283867 220925 283868
rect 219768 273454 220088 273486
rect 219768 273218 219810 273454
rect 220046 273218 220088 273454
rect 219768 273134 220088 273218
rect 219768 272898 219810 273134
rect 220046 272898 220088 273134
rect 219768 272866 220088 272898
rect 217547 240140 217613 240141
rect 217547 240076 217548 240140
rect 217612 240076 217613 240140
rect 217547 240075 217613 240076
rect 219203 240140 219269 240141
rect 219203 240076 219204 240140
rect 219268 240076 219269 240140
rect 219203 240075 219269 240076
rect 217794 219454 218414 238182
rect 217794 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 218414 219454
rect 217794 219134 218414 219218
rect 217794 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 218414 219134
rect 216443 188460 216509 188461
rect 216443 188396 216444 188460
rect 216508 188396 216509 188460
rect 216443 188395 216509 188396
rect 217794 183454 218414 218898
rect 220862 192541 220922 283867
rect 221046 240141 221106 287267
rect 221514 286182 222134 294618
rect 221043 240140 221109 240141
rect 221043 240076 221044 240140
rect 221108 240076 221109 240140
rect 221043 240075 221109 240076
rect 222334 238645 222394 334187
rect 224723 283932 224789 283933
rect 224723 283868 224724 283932
rect 224788 283868 224789 283932
rect 224723 283867 224789 283868
rect 222331 238644 222397 238645
rect 222331 238580 222332 238644
rect 222396 238580 222397 238644
rect 222331 238579 222397 238580
rect 221514 223174 222134 238182
rect 221514 222938 221546 223174
rect 221782 222938 221866 223174
rect 222102 222938 222134 223174
rect 221514 222854 222134 222938
rect 221514 222618 221546 222854
rect 221782 222618 221866 222854
rect 222102 222618 222134 222854
rect 220859 192540 220925 192541
rect 220859 192476 220860 192540
rect 220924 192476 220925 192540
rect 220859 192475 220925 192476
rect 217794 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 218414 183454
rect 217794 183134 218414 183218
rect 217794 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 218414 183134
rect 217794 178000 218414 182898
rect 221514 187174 222134 222618
rect 221514 186938 221546 187174
rect 221782 186938 221866 187174
rect 222102 186938 222134 187174
rect 221514 186854 222134 186938
rect 221514 186618 221546 186854
rect 221782 186618 221866 186854
rect 222102 186618 222134 186854
rect 221514 178000 222134 186618
rect 224726 180165 224786 283867
rect 224910 238509 224970 367779
rect 225234 334894 225854 370338
rect 225234 334658 225266 334894
rect 225502 334658 225586 334894
rect 225822 334658 225854 334894
rect 225234 334574 225854 334658
rect 225234 334338 225266 334574
rect 225502 334338 225586 334574
rect 225822 334338 225854 334574
rect 225234 298894 225854 334338
rect 228954 374614 229574 375600
rect 228954 374378 228986 374614
rect 229222 374378 229306 374614
rect 229542 374378 229574 374614
rect 228954 374294 229574 374378
rect 228954 374058 228986 374294
rect 229222 374058 229306 374294
rect 229542 374058 229574 374294
rect 228954 338614 229574 374058
rect 234475 352612 234541 352613
rect 234475 352548 234476 352612
rect 234540 352548 234541 352612
rect 234475 352547 234541 352548
rect 230427 339556 230493 339557
rect 230427 339492 230428 339556
rect 230492 339492 230493 339556
rect 230427 339491 230493 339492
rect 228954 338378 228986 338614
rect 229222 338378 229306 338614
rect 229542 338378 229574 338614
rect 228954 338294 229574 338378
rect 228954 338058 228986 338294
rect 229222 338058 229306 338294
rect 229542 338058 229574 338294
rect 227667 302836 227733 302837
rect 227667 302772 227668 302836
rect 227732 302772 227733 302836
rect 227667 302771 227733 302772
rect 225234 298658 225266 298894
rect 225502 298658 225586 298894
rect 225822 298658 225854 298894
rect 225234 298574 225854 298658
rect 225234 298338 225266 298574
rect 225502 298338 225586 298574
rect 225822 298338 225854 298574
rect 225234 286182 225854 298338
rect 226931 285836 226997 285837
rect 226931 285772 226932 285836
rect 226996 285772 226997 285836
rect 226931 285771 226997 285772
rect 226195 285700 226261 285701
rect 226195 285636 226196 285700
rect 226260 285636 226261 285700
rect 226195 285635 226261 285636
rect 226198 238509 226258 285635
rect 224907 238508 224973 238509
rect 224907 238444 224908 238508
rect 224972 238444 224973 238508
rect 224907 238443 224973 238444
rect 226195 238508 226261 238509
rect 226195 238444 226196 238508
rect 226260 238444 226261 238508
rect 226195 238443 226261 238444
rect 225234 226894 225854 238182
rect 225234 226658 225266 226894
rect 225502 226658 225586 226894
rect 225822 226658 225854 226894
rect 225234 226574 225854 226658
rect 225234 226338 225266 226574
rect 225502 226338 225586 226574
rect 225822 226338 225854 226574
rect 224907 199612 224973 199613
rect 224907 199548 224908 199612
rect 224972 199548 224973 199612
rect 224907 199547 224973 199548
rect 224910 181253 224970 199547
rect 225234 190894 225854 226338
rect 225234 190658 225266 190894
rect 225502 190658 225586 190894
rect 225822 190658 225854 190894
rect 225234 190574 225854 190658
rect 225234 190338 225266 190574
rect 225502 190338 225586 190574
rect 225822 190338 225854 190574
rect 224907 181252 224973 181253
rect 224907 181188 224908 181252
rect 224972 181188 224973 181252
rect 224907 181187 224973 181188
rect 224723 180164 224789 180165
rect 224723 180100 224724 180164
rect 224788 180100 224789 180164
rect 224723 180099 224789 180100
rect 225234 178000 225854 190338
rect 226934 180301 226994 285771
rect 227670 283933 227730 302771
rect 228954 302614 229574 338058
rect 228954 302378 228986 302614
rect 229222 302378 229306 302614
rect 229542 302378 229574 302614
rect 228954 302294 229574 302378
rect 228954 302058 228986 302294
rect 229222 302058 229306 302294
rect 229542 302058 229574 302294
rect 228219 287196 228285 287197
rect 228219 287132 228220 287196
rect 228284 287132 228285 287196
rect 228219 287131 228285 287132
rect 227667 283932 227733 283933
rect 227667 283868 227668 283932
rect 227732 283868 227733 283932
rect 227667 283867 227733 283868
rect 228222 219605 228282 287131
rect 228954 286182 229574 302058
rect 228771 283932 228837 283933
rect 228771 283868 228772 283932
rect 228836 283868 228837 283932
rect 228771 283867 228837 283868
rect 229691 283932 229757 283933
rect 229691 283868 229692 283932
rect 229756 283868 229757 283932
rect 229691 283867 229757 283868
rect 228219 219604 228285 219605
rect 228219 219540 228220 219604
rect 228284 219540 228285 219604
rect 228219 219539 228285 219540
rect 226931 180300 226997 180301
rect 226931 180236 226932 180300
rect 226996 180236 226997 180300
rect 226931 180235 226997 180236
rect 228774 178669 228834 283867
rect 228954 230614 229574 238182
rect 228954 230378 228986 230614
rect 229222 230378 229306 230614
rect 229542 230378 229574 230614
rect 228954 230294 229574 230378
rect 228954 230058 228986 230294
rect 229222 230058 229306 230294
rect 229542 230058 229574 230294
rect 228954 194614 229574 230058
rect 228954 194378 228986 194614
rect 229222 194378 229306 194614
rect 229542 194378 229574 194614
rect 228954 194294 229574 194378
rect 228954 194058 228986 194294
rect 229222 194058 229306 194294
rect 229542 194058 229574 194294
rect 228771 178668 228837 178669
rect 228771 178604 228772 178668
rect 228836 178604 228837 178668
rect 228771 178603 228837 178604
rect 228954 178000 229574 194058
rect 229139 177036 229205 177037
rect 229139 176972 229140 177036
rect 229204 176972 229205 177036
rect 229139 176971 229205 176972
rect 221207 165454 221527 165486
rect 221207 165218 221249 165454
rect 221485 165218 221527 165454
rect 221207 165134 221527 165218
rect 221207 164898 221249 165134
rect 221485 164898 221527 165134
rect 221207 164866 221527 164898
rect 224471 165454 224791 165486
rect 224471 165218 224513 165454
rect 224749 165218 224791 165454
rect 224471 165134 224791 165218
rect 224471 164898 224513 165134
rect 224749 164898 224791 165134
rect 224471 164866 224791 164898
rect 229142 149701 229202 176971
rect 229139 149700 229205 149701
rect 229139 149636 229140 149700
rect 229204 149636 229205 149700
rect 229139 149635 229205 149636
rect 229139 148068 229205 148069
rect 229139 148004 229140 148068
rect 229204 148004 229205 148068
rect 229139 148003 229205 148004
rect 219575 147454 219895 147486
rect 219575 147218 219617 147454
rect 219853 147218 219895 147454
rect 219575 147134 219895 147218
rect 219575 146898 219617 147134
rect 219853 146898 219895 147134
rect 219575 146866 219895 146898
rect 222839 147454 223159 147486
rect 222839 147218 222881 147454
rect 223117 147218 223159 147454
rect 222839 147134 223159 147218
rect 222839 146898 222881 147134
rect 223117 146898 223159 147134
rect 222839 146866 223159 146898
rect 226103 147454 226423 147486
rect 226103 147218 226145 147454
rect 226381 147218 226423 147454
rect 226103 147134 226423 147218
rect 226103 146898 226145 147134
rect 226381 146898 226423 147134
rect 226103 146866 226423 146898
rect 229142 141133 229202 148003
rect 229139 141132 229205 141133
rect 229139 141068 229140 141132
rect 229204 141068 229205 141132
rect 229139 141067 229205 141068
rect 229694 137325 229754 283867
rect 230430 240141 230490 339491
rect 232083 331804 232149 331805
rect 232083 331740 232084 331804
rect 232148 331740 232149 331804
rect 232083 331739 232149 331740
rect 231899 287332 231965 287333
rect 231899 287268 231900 287332
rect 231964 287268 231965 287332
rect 231899 287267 231965 287268
rect 230979 283932 231045 283933
rect 230979 283868 230980 283932
rect 231044 283868 231045 283932
rect 230979 283867 231045 283868
rect 230982 240141 231042 283867
rect 230427 240140 230493 240141
rect 230427 240076 230428 240140
rect 230492 240076 230493 240140
rect 230427 240075 230493 240076
rect 230979 240140 231045 240141
rect 230979 240076 230980 240140
rect 231044 240076 231045 240140
rect 230979 240075 231045 240076
rect 230430 147933 230490 240075
rect 230611 176900 230677 176901
rect 230611 176836 230612 176900
rect 230676 176836 230677 176900
rect 230611 176835 230677 176836
rect 230614 169557 230674 176835
rect 230611 169556 230677 169557
rect 230611 169492 230612 169556
rect 230676 169492 230677 169556
rect 230611 169491 230677 169492
rect 231902 167653 231962 287267
rect 232086 240141 232146 331739
rect 234478 240141 234538 352547
rect 235794 345454 236414 375600
rect 235794 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 236414 345454
rect 235794 345134 236414 345218
rect 235794 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 236414 345134
rect 235794 309454 236414 344898
rect 235794 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 236414 309454
rect 235794 309134 236414 309218
rect 235794 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 236414 309134
rect 235794 286182 236414 308898
rect 239514 349174 240134 375600
rect 241651 375324 241717 375325
rect 241651 375260 241652 375324
rect 241716 375260 241717 375324
rect 241651 375259 241717 375260
rect 240731 351252 240797 351253
rect 240731 351188 240732 351252
rect 240796 351188 240797 351252
rect 240731 351187 240797 351188
rect 239514 348938 239546 349174
rect 239782 348938 239866 349174
rect 240102 348938 240134 349174
rect 239514 348854 240134 348938
rect 239514 348618 239546 348854
rect 239782 348618 239866 348854
rect 240102 348618 240134 348854
rect 239514 313174 240134 348618
rect 239514 312938 239546 313174
rect 239782 312938 239866 313174
rect 240102 312938 240134 313174
rect 239514 312854 240134 312938
rect 239514 312618 239546 312854
rect 239782 312618 239866 312854
rect 240102 312618 240134 312854
rect 238707 287196 238773 287197
rect 238707 287132 238708 287196
rect 238772 287132 238773 287196
rect 238707 287131 238773 287132
rect 238710 287070 238770 287131
rect 238526 287010 238770 287070
rect 234659 285972 234725 285973
rect 234659 285908 234660 285972
rect 234724 285908 234725 285972
rect 234659 285907 234725 285908
rect 232083 240140 232149 240141
rect 232083 240076 232084 240140
rect 232148 240076 232149 240140
rect 232083 240075 232149 240076
rect 234475 240140 234541 240141
rect 234475 240076 234476 240140
rect 234540 240076 234541 240140
rect 234475 240075 234541 240076
rect 233187 223548 233253 223549
rect 233187 223484 233188 223548
rect 233252 223484 233253 223548
rect 233187 223483 233253 223484
rect 232083 185740 232149 185741
rect 232083 185676 232084 185740
rect 232148 185676 232149 185740
rect 232083 185675 232149 185676
rect 231899 167652 231965 167653
rect 231899 167588 231900 167652
rect 231964 167588 231965 167652
rect 231899 167587 231965 167588
rect 230979 167244 231045 167245
rect 230979 167180 230980 167244
rect 231044 167180 231045 167244
rect 230979 167179 231045 167180
rect 230982 159629 231042 167179
rect 230979 159628 231045 159629
rect 230979 159564 230980 159628
rect 231044 159564 231045 159628
rect 230979 159563 231045 159564
rect 230427 147932 230493 147933
rect 230427 147868 230428 147932
rect 230492 147868 230493 147932
rect 230427 147867 230493 147868
rect 232086 147253 232146 185675
rect 233190 153101 233250 223483
rect 233371 185876 233437 185877
rect 233371 185812 233372 185876
rect 233436 185812 233437 185876
rect 233371 185811 233437 185812
rect 233374 171189 233434 185811
rect 233371 171188 233437 171189
rect 233371 171124 233372 171188
rect 233436 171124 233437 171188
rect 233371 171123 233437 171124
rect 234662 154869 234722 285907
rect 236499 283932 236565 283933
rect 236499 283868 236500 283932
rect 236564 283868 236565 283932
rect 236499 283867 236565 283868
rect 237971 283932 238037 283933
rect 237971 283868 237972 283932
rect 238036 283868 238037 283932
rect 237971 283867 238037 283868
rect 235128 255454 235448 255486
rect 235128 255218 235170 255454
rect 235406 255218 235448 255454
rect 235128 255134 235448 255218
rect 235128 254898 235170 255134
rect 235406 254898 235448 255134
rect 235128 254866 235448 254898
rect 235794 237454 236414 238182
rect 235794 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 236414 237454
rect 235794 237134 236414 237218
rect 235794 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 236414 237134
rect 235794 201454 236414 236898
rect 235794 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 236414 201454
rect 235794 201134 236414 201218
rect 235794 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 236414 201134
rect 235794 165454 236414 200898
rect 236502 175133 236562 283867
rect 237974 212533 238034 283867
rect 238526 244290 238586 287010
rect 239514 286182 240134 312618
rect 240363 298484 240429 298485
rect 240363 298420 240364 298484
rect 240428 298420 240429 298484
rect 240363 298419 240429 298420
rect 238526 244230 238770 244290
rect 238710 240141 238770 244230
rect 238707 240140 238773 240141
rect 238707 240076 238708 240140
rect 238772 240076 238773 240140
rect 238707 240075 238773 240076
rect 239259 235652 239325 235653
rect 239259 235588 239260 235652
rect 239324 235588 239325 235652
rect 239259 235587 239325 235588
rect 237971 212532 238037 212533
rect 237971 212468 237972 212532
rect 238036 212468 238037 212532
rect 237971 212467 238037 212468
rect 237419 188596 237485 188597
rect 237419 188532 237420 188596
rect 237484 188532 237485 188596
rect 237419 188531 237485 188532
rect 236683 175268 236749 175269
rect 236683 175204 236684 175268
rect 236748 175204 236749 175268
rect 236683 175203 236749 175204
rect 236499 175132 236565 175133
rect 236499 175068 236500 175132
rect 236564 175068 236565 175132
rect 236499 175067 236565 175068
rect 235794 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 236414 165454
rect 235794 165134 236414 165218
rect 235794 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 236414 165134
rect 234659 154868 234725 154869
rect 234659 154804 234660 154868
rect 234724 154804 234725 154868
rect 234659 154803 234725 154804
rect 233187 153100 233253 153101
rect 233187 153036 233188 153100
rect 233252 153036 233253 153100
rect 233187 153035 233253 153036
rect 232083 147252 232149 147253
rect 232083 147188 232084 147252
rect 232148 147188 232149 147252
rect 232083 147187 232149 147188
rect 231715 146980 231781 146981
rect 231715 146916 231716 146980
rect 231780 146916 231781 146980
rect 231715 146915 231781 146916
rect 231718 145893 231778 146915
rect 231715 145892 231781 145893
rect 231715 145828 231716 145892
rect 231780 145828 231781 145892
rect 231715 145827 231781 145828
rect 230427 144124 230493 144125
rect 230427 144060 230428 144124
rect 230492 144060 230493 144124
rect 230427 144059 230493 144060
rect 230430 141677 230490 144059
rect 230427 141676 230493 141677
rect 230427 141612 230428 141676
rect 230492 141612 230493 141676
rect 230427 141611 230493 141612
rect 232451 141676 232517 141677
rect 232451 141612 232452 141676
rect 232516 141612 232517 141676
rect 232451 141611 232517 141612
rect 230979 141540 231045 141541
rect 230979 141476 230980 141540
rect 231044 141476 231045 141540
rect 230979 141475 231045 141476
rect 229691 137324 229757 137325
rect 229691 137260 229692 137324
rect 229756 137260 229757 137324
rect 229691 137259 229757 137260
rect 230982 132157 231042 141475
rect 231715 141404 231781 141405
rect 231715 141340 231716 141404
rect 231780 141340 231781 141404
rect 231715 141339 231781 141340
rect 231718 135013 231778 141339
rect 231715 135012 231781 135013
rect 231715 134948 231716 135012
rect 231780 134948 231781 135012
rect 231715 134947 231781 134948
rect 230979 132156 231045 132157
rect 230979 132092 230980 132156
rect 231044 132092 231045 132156
rect 230979 132091 231045 132092
rect 221207 129454 221527 129486
rect 221207 129218 221249 129454
rect 221485 129218 221527 129454
rect 221207 129134 221527 129218
rect 221207 128898 221249 129134
rect 221485 128898 221527 129134
rect 221207 128866 221527 128898
rect 224471 129454 224791 129486
rect 224471 129218 224513 129454
rect 224749 129218 224791 129454
rect 224471 129134 224791 129218
rect 224471 128898 224513 129134
rect 224749 128898 224791 129134
rect 231163 129028 231229 129029
rect 231163 128964 231164 129028
rect 231228 128964 231229 129028
rect 231163 128963 231229 128964
rect 224471 128866 224791 128898
rect 230979 126036 231045 126037
rect 230979 125972 230980 126036
rect 231044 125972 231045 126036
rect 230979 125971 231045 125972
rect 229691 114884 229757 114885
rect 229691 114820 229692 114884
rect 229756 114820 229757 114884
rect 229691 114819 229757 114820
rect 219575 111454 219895 111486
rect 219575 111218 219617 111454
rect 219853 111218 219895 111454
rect 219575 111134 219895 111218
rect 219575 110898 219617 111134
rect 219853 110898 219895 111134
rect 219575 110866 219895 110898
rect 222839 111454 223159 111486
rect 222839 111218 222881 111454
rect 223117 111218 223159 111454
rect 222839 111134 223159 111218
rect 222839 110898 222881 111134
rect 223117 110898 223159 111134
rect 222839 110866 223159 110898
rect 226103 111454 226423 111486
rect 226103 111218 226145 111454
rect 226381 111218 226423 111454
rect 226103 111134 226423 111218
rect 226103 110898 226145 111134
rect 226381 110898 226423 111134
rect 226103 110866 226423 110898
rect 229139 97884 229205 97885
rect 229139 97820 229140 97884
rect 229204 97820 229205 97884
rect 229139 97819 229205 97820
rect 229142 97610 229202 97819
rect 228774 97550 229202 97610
rect 223619 95572 223685 95573
rect 223619 95508 223620 95572
rect 223684 95508 223685 95572
rect 223619 95507 223685 95508
rect 223435 95436 223501 95437
rect 223435 95372 223436 95436
rect 223500 95372 223501 95436
rect 223435 95371 223501 95372
rect 219387 94076 219453 94077
rect 219387 94012 219388 94076
rect 219452 94012 219453 94076
rect 219387 94011 219453 94012
rect 215155 90404 215221 90405
rect 215155 90340 215156 90404
rect 215220 90340 215221 90404
rect 215155 90339 215221 90340
rect 210954 68378 210986 68614
rect 211222 68378 211306 68614
rect 211542 68378 211574 68614
rect 210954 68294 211574 68378
rect 210954 68058 210986 68294
rect 211222 68058 211306 68294
rect 211542 68058 211574 68294
rect 210954 32614 211574 68058
rect 210954 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 211574 32614
rect 210954 32294 211574 32378
rect 210954 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 211574 32294
rect 192954 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 193574 -6106
rect 192954 -6426 193574 -6342
rect 192954 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 193574 -6426
rect 192954 -7654 193574 -6662
rect 210954 -7066 211574 32058
rect 217794 75454 218414 94000
rect 219390 93530 219450 94011
rect 217794 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 218414 75454
rect 217794 75134 218414 75218
rect 217794 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 218414 75134
rect 217794 39454 218414 74898
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 219206 93470 219450 93530
rect 219206 33829 219266 93470
rect 221514 79174 222134 94000
rect 223438 88229 223498 95371
rect 223435 88228 223501 88229
rect 223435 88164 223436 88228
rect 223500 88164 223501 88228
rect 223435 88163 223501 88164
rect 221514 78938 221546 79174
rect 221782 78938 221866 79174
rect 222102 78938 222134 79174
rect 221514 78854 222134 78938
rect 221514 78618 221546 78854
rect 221782 78618 221866 78854
rect 222102 78618 222134 78854
rect 221514 43174 222134 78618
rect 221514 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 222134 43174
rect 221514 42854 222134 42938
rect 221514 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 222134 42854
rect 219203 33828 219269 33829
rect 219203 33764 219204 33828
rect 219268 33764 219269 33828
rect 219203 33763 219269 33764
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -1894 218414 -902
rect 221514 7174 222134 42618
rect 223622 17237 223682 95507
rect 228774 95437 228834 97550
rect 229139 97204 229205 97205
rect 229139 97140 229140 97204
rect 229204 97140 229205 97204
rect 229139 97139 229205 97140
rect 229142 96930 229202 97139
rect 228958 96870 229202 96930
rect 228958 95573 229018 96870
rect 228955 95572 229021 95573
rect 228955 95508 228956 95572
rect 229020 95508 229021 95572
rect 228955 95507 229021 95508
rect 228771 95436 228837 95437
rect 228771 95372 228772 95436
rect 228836 95372 228837 95436
rect 228771 95371 228837 95372
rect 225234 82894 225854 94000
rect 227667 90404 227733 90405
rect 227667 90340 227668 90404
rect 227732 90340 227733 90404
rect 227667 90339 227733 90340
rect 225234 82658 225266 82894
rect 225502 82658 225586 82894
rect 225822 82658 225854 82894
rect 225234 82574 225854 82658
rect 225234 82338 225266 82574
rect 225502 82338 225586 82574
rect 225822 82338 225854 82574
rect 225234 46894 225854 82338
rect 225234 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 225854 46894
rect 225234 46574 225854 46658
rect 225234 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 225854 46574
rect 223619 17236 223685 17237
rect 223619 17172 223620 17236
rect 223684 17172 223685 17236
rect 223619 17171 223685 17172
rect 221514 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 222134 7174
rect 221514 6854 222134 6938
rect 221514 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 222134 6854
rect 221514 -2266 222134 6618
rect 221514 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 222134 -2266
rect 221514 -2586 222134 -2502
rect 221514 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 222134 -2586
rect 221514 -3814 222134 -2822
rect 225234 10894 225854 46338
rect 225234 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 225854 10894
rect 225234 10574 225854 10658
rect 225234 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 225854 10574
rect 225234 -4186 225854 10338
rect 227670 8941 227730 90339
rect 228954 86614 229574 94000
rect 228954 86378 228986 86614
rect 229222 86378 229306 86614
rect 229542 86378 229574 86614
rect 228954 86294 229574 86378
rect 228954 86058 228986 86294
rect 229222 86058 229306 86294
rect 229542 86058 229574 86294
rect 228954 50614 229574 86058
rect 229694 57221 229754 114819
rect 229691 57220 229757 57221
rect 229691 57156 229692 57220
rect 229756 57156 229757 57220
rect 229691 57155 229757 57156
rect 228954 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 229574 50614
rect 228954 50294 229574 50378
rect 228954 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 229574 50294
rect 228954 14614 229574 50058
rect 230982 42125 231042 125971
rect 231166 119781 231226 128963
rect 231163 119780 231229 119781
rect 231163 119716 231164 119780
rect 231228 119716 231229 119780
rect 231163 119715 231229 119716
rect 232454 98565 232514 141611
rect 233739 134196 233805 134197
rect 233739 134132 233740 134196
rect 233804 134132 233805 134196
rect 233739 134131 233805 134132
rect 232451 98564 232517 98565
rect 232451 98500 232452 98564
rect 232516 98500 232517 98564
rect 232451 98499 232517 98500
rect 230979 42124 231045 42125
rect 230979 42060 230980 42124
rect 231044 42060 231045 42124
rect 230979 42059 231045 42060
rect 233742 26893 233802 134131
rect 235794 129454 236414 164898
rect 236686 145349 236746 175203
rect 237422 161533 237482 188531
rect 237971 180164 238037 180165
rect 237971 180100 237972 180164
rect 238036 180100 238037 180164
rect 237971 180099 238037 180100
rect 237419 161532 237485 161533
rect 237419 161468 237420 161532
rect 237484 161468 237485 161532
rect 237419 161467 237485 161468
rect 236683 145348 236749 145349
rect 236683 145284 236684 145348
rect 236748 145284 236749 145348
rect 236683 145283 236749 145284
rect 237974 142493 238034 180099
rect 239262 156637 239322 235587
rect 239514 205174 240134 238182
rect 239514 204938 239546 205174
rect 239782 204938 239866 205174
rect 240102 204938 240134 205174
rect 239514 204854 240134 204938
rect 239514 204618 239546 204854
rect 239782 204618 239866 204854
rect 240102 204618 240134 204854
rect 239514 169174 240134 204618
rect 240366 174317 240426 298419
rect 240734 288421 240794 351187
rect 240731 288420 240797 288421
rect 240731 288356 240732 288420
rect 240796 288356 240797 288420
rect 240731 288355 240797 288356
rect 241654 215933 241714 375259
rect 243234 352894 243854 375600
rect 244779 374644 244845 374645
rect 244779 374580 244780 374644
rect 244844 374580 244845 374644
rect 244779 374579 244845 374580
rect 243234 352658 243266 352894
rect 243502 352658 243586 352894
rect 243822 352658 243854 352894
rect 243234 352574 243854 352658
rect 243234 352338 243266 352574
rect 243502 352338 243586 352574
rect 243822 352338 243854 352574
rect 243234 316894 243854 352338
rect 243234 316658 243266 316894
rect 243502 316658 243586 316894
rect 243822 316658 243854 316894
rect 243234 316574 243854 316658
rect 243234 316338 243266 316574
rect 243502 316338 243586 316574
rect 243822 316338 243854 316574
rect 242939 298756 243005 298757
rect 242939 298692 242940 298756
rect 243004 298692 243005 298756
rect 242939 298691 243005 298692
rect 242942 277410 243002 298691
rect 243234 286182 243854 316338
rect 244411 298212 244477 298213
rect 244411 298148 244412 298212
rect 244476 298148 244477 298212
rect 244411 298147 244477 298148
rect 244043 285972 244109 285973
rect 244043 285908 244044 285972
rect 244108 285908 244109 285972
rect 244043 285907 244109 285908
rect 242942 277350 243554 277410
rect 243494 269109 243554 277350
rect 243491 269108 243557 269109
rect 243491 269044 243492 269108
rect 243556 269044 243557 269108
rect 243491 269043 243557 269044
rect 244046 244290 244106 285907
rect 244227 269924 244293 269925
rect 244227 269860 244228 269924
rect 244292 269860 244293 269924
rect 244227 269859 244293 269860
rect 243862 244230 244106 244290
rect 243491 241364 243557 241365
rect 243491 241300 243492 241364
rect 243556 241300 243557 241364
rect 243491 241299 243557 241300
rect 243494 238370 243554 241299
rect 243862 238645 243922 244230
rect 244230 243810 244290 269859
rect 244414 259589 244474 298147
rect 244782 280125 244842 374579
rect 246954 356614 247574 375600
rect 246954 356378 246986 356614
rect 247222 356378 247306 356614
rect 247542 356378 247574 356614
rect 246954 356294 247574 356378
rect 246954 356058 246986 356294
rect 247222 356058 247306 356294
rect 247542 356058 247574 356294
rect 245699 345812 245765 345813
rect 245699 345748 245700 345812
rect 245764 345748 245765 345812
rect 245699 345747 245765 345748
rect 244779 280124 244845 280125
rect 244779 280060 244780 280124
rect 244844 280060 244845 280124
rect 244779 280059 244845 280060
rect 245702 275365 245762 345747
rect 246954 320614 247574 356058
rect 253794 363454 254414 375600
rect 253794 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 254414 363454
rect 253794 363134 254414 363218
rect 253794 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 254414 363134
rect 248459 347172 248525 347173
rect 248459 347108 248460 347172
rect 248524 347108 248525 347172
rect 248459 347107 248525 347108
rect 246954 320378 246986 320614
rect 247222 320378 247306 320614
rect 247542 320378 247574 320614
rect 246954 320294 247574 320378
rect 246954 320058 246986 320294
rect 247222 320058 247306 320294
rect 247542 320058 247574 320294
rect 246954 284614 247574 320058
rect 247723 303652 247789 303653
rect 247723 303588 247724 303652
rect 247788 303588 247789 303652
rect 247723 303587 247789 303588
rect 246954 284378 246986 284614
rect 247222 284378 247306 284614
rect 247542 284378 247574 284614
rect 246954 284294 247574 284378
rect 246954 284058 246986 284294
rect 247222 284058 247306 284294
rect 247542 284058 247574 284294
rect 245699 275364 245765 275365
rect 245699 275300 245700 275364
rect 245764 275300 245765 275364
rect 245699 275299 245765 275300
rect 244411 259588 244477 259589
rect 244411 259524 244412 259588
rect 244476 259524 244477 259588
rect 244411 259523 244477 259524
rect 244046 243750 244290 243810
rect 246954 248614 247574 284058
rect 247726 256053 247786 303587
rect 247723 256052 247789 256053
rect 247723 255988 247724 256052
rect 247788 255988 247789 256052
rect 247723 255987 247789 255988
rect 248462 252245 248522 347107
rect 251771 341460 251837 341461
rect 251771 341396 251772 341460
rect 251836 341396 251837 341460
rect 251771 341395 251837 341396
rect 249747 315348 249813 315349
rect 249747 315284 249748 315348
rect 249812 315284 249813 315348
rect 249747 315283 249813 315284
rect 249011 285836 249077 285837
rect 249011 285772 249012 285836
rect 249076 285772 249077 285836
rect 249011 285771 249077 285772
rect 249014 261493 249074 285771
rect 249011 261492 249077 261493
rect 249011 261428 249012 261492
rect 249076 261428 249077 261492
rect 249011 261427 249077 261428
rect 248459 252244 248525 252245
rect 248459 252180 248460 252244
rect 248524 252180 248525 252244
rect 248459 252179 248525 252180
rect 248459 249932 248525 249933
rect 248459 249868 248460 249932
rect 248524 249868 248525 249932
rect 248459 249867 248525 249868
rect 246954 248378 246986 248614
rect 247222 248378 247306 248614
rect 247542 248378 247574 248614
rect 246954 248294 247574 248378
rect 246954 248058 246986 248294
rect 247222 248058 247306 248294
rect 247542 248058 247574 248294
rect 243859 238644 243925 238645
rect 243859 238580 243860 238644
rect 243924 238580 243925 238644
rect 243859 238579 243925 238580
rect 242942 238310 243554 238370
rect 242942 226133 243002 238310
rect 242939 226132 243005 226133
rect 242939 226068 242940 226132
rect 243004 226068 243005 226132
rect 242939 226067 243005 226068
rect 241651 215932 241717 215933
rect 241651 215868 241652 215932
rect 241716 215868 241717 215932
rect 241651 215867 241717 215868
rect 243234 208894 243854 238182
rect 244046 234630 244106 243750
rect 245699 242996 245765 242997
rect 245699 242932 245700 242996
rect 245764 242932 245765 242996
rect 245699 242931 245765 242932
rect 244046 234570 244290 234630
rect 243234 208658 243266 208894
rect 243502 208658 243586 208894
rect 243822 208658 243854 208894
rect 243234 208574 243854 208658
rect 243234 208338 243266 208574
rect 243502 208338 243586 208574
rect 243822 208338 243854 208574
rect 242939 189140 243005 189141
rect 242939 189076 242940 189140
rect 243004 189076 243005 189140
rect 242939 189075 243005 189076
rect 241651 178804 241717 178805
rect 241651 178740 241652 178804
rect 241716 178740 241717 178804
rect 241651 178739 241717 178740
rect 240547 177308 240613 177309
rect 240547 177244 240548 177308
rect 240612 177244 240613 177308
rect 240547 177243 240613 177244
rect 240363 174316 240429 174317
rect 240363 174252 240364 174316
rect 240428 174252 240429 174316
rect 240363 174251 240429 174252
rect 239514 168938 239546 169174
rect 239782 168938 239866 169174
rect 240102 168938 240134 169174
rect 239514 168854 240134 168938
rect 239514 168618 239546 168854
rect 239782 168618 239866 168854
rect 240102 168618 240134 168854
rect 239259 156636 239325 156637
rect 239259 156572 239260 156636
rect 239324 156572 239325 156636
rect 239259 156571 239325 156572
rect 237971 142492 238037 142493
rect 237971 142428 237972 142492
rect 238036 142428 238037 142492
rect 237971 142427 238037 142428
rect 237971 138684 238037 138685
rect 237971 138620 237972 138684
rect 238036 138620 238037 138684
rect 237971 138619 238037 138620
rect 235794 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 236414 129454
rect 235794 129134 236414 129218
rect 235794 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 236414 129134
rect 235794 93454 236414 128898
rect 237974 98021 238034 138619
rect 239514 133174 240134 168618
rect 240550 152557 240610 177243
rect 241283 175268 241349 175269
rect 241283 175204 241284 175268
rect 241348 175204 241349 175268
rect 241283 175203 241349 175204
rect 240547 152556 240613 152557
rect 240547 152492 240548 152556
rect 240612 152492 240613 152556
rect 240547 152491 240613 152492
rect 239514 132938 239546 133174
rect 239782 132938 239866 133174
rect 240102 132938 240134 133174
rect 239514 132854 240134 132938
rect 239514 132618 239546 132854
rect 239782 132618 239866 132854
rect 240102 132618 240134 132854
rect 237971 98020 238037 98021
rect 237971 97956 237972 98020
rect 238036 97956 238037 98020
rect 237971 97955 238037 97956
rect 235794 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 236414 93454
rect 235794 93134 236414 93218
rect 235794 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 236414 93134
rect 235794 57454 236414 92898
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 233739 26892 233805 26893
rect 233739 26828 233740 26892
rect 233804 26828 233805 26892
rect 233739 26827 233805 26828
rect 228954 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 229574 14614
rect 228954 14294 229574 14378
rect 228954 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 229574 14294
rect 227667 8940 227733 8941
rect 227667 8876 227668 8940
rect 227732 8876 227733 8940
rect 227667 8875 227733 8876
rect 225234 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 225854 -4186
rect 225234 -4506 225854 -4422
rect 225234 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 225854 -4506
rect 225234 -5734 225854 -4742
rect 210954 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 211574 -7066
rect 210954 -7386 211574 -7302
rect 210954 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 211574 -7386
rect 210954 -7654 211574 -7622
rect 228954 -6106 229574 14058
rect 235794 21454 236414 56898
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -1306 236414 20898
rect 235794 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 236414 -1306
rect 235794 -1626 236414 -1542
rect 235794 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 236414 -1626
rect 235794 -1894 236414 -1862
rect 239514 97174 240134 132618
rect 239514 96938 239546 97174
rect 239782 96938 239866 97174
rect 240102 96938 240134 97174
rect 239514 96854 240134 96938
rect 239514 96618 239546 96854
rect 239782 96618 239866 96854
rect 240102 96618 240134 96854
rect 239514 61174 240134 96618
rect 239514 60938 239546 61174
rect 239782 60938 239866 61174
rect 240102 60938 240134 61174
rect 239514 60854 240134 60938
rect 239514 60618 239546 60854
rect 239782 60618 239866 60854
rect 240102 60618 240134 60854
rect 239514 25174 240134 60618
rect 239514 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 240134 25174
rect 239514 24854 240134 24938
rect 239514 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 240134 24854
rect 239514 -3226 240134 24618
rect 241286 3365 241346 175203
rect 241654 138821 241714 178739
rect 242942 149157 243002 189075
rect 243234 172894 243854 208338
rect 243234 172658 243266 172894
rect 243502 172658 243586 172894
rect 243822 172658 243854 172894
rect 244230 172821 244290 234570
rect 245702 231437 245762 242931
rect 245699 231436 245765 231437
rect 245699 231372 245700 231436
rect 245764 231372 245765 231436
rect 245699 231371 245765 231372
rect 246954 212614 247574 248058
rect 248462 239597 248522 249867
rect 248459 239596 248525 239597
rect 248459 239532 248460 239596
rect 248524 239532 248525 239596
rect 248459 239531 248525 239532
rect 246954 212378 246986 212614
rect 247222 212378 247306 212614
rect 247542 212378 247574 212614
rect 246954 212294 247574 212378
rect 246954 212058 246986 212294
rect 247222 212058 247306 212294
rect 247542 212058 247574 212294
rect 246251 199340 246317 199341
rect 246251 199276 246252 199340
rect 246316 199276 246317 199340
rect 246251 199275 246317 199276
rect 244411 175948 244477 175949
rect 244411 175884 244412 175948
rect 244476 175884 244477 175948
rect 244411 175883 244477 175884
rect 244227 172820 244293 172821
rect 244227 172756 244228 172820
rect 244292 172756 244293 172820
rect 244227 172755 244293 172756
rect 243234 172574 243854 172658
rect 243234 172338 243266 172574
rect 243502 172338 243586 172574
rect 243822 172338 243854 172574
rect 242939 149156 243005 149157
rect 242939 149092 242940 149156
rect 243004 149092 243005 149156
rect 242939 149091 243005 149092
rect 241651 138820 241717 138821
rect 241651 138756 241652 138820
rect 241716 138756 241717 138820
rect 241651 138755 241717 138756
rect 243234 136894 243854 172338
rect 244414 151061 244474 175883
rect 244411 151060 244477 151061
rect 244411 150996 244412 151060
rect 244476 150996 244477 151060
rect 244411 150995 244477 150996
rect 244779 140044 244845 140045
rect 244779 139980 244780 140044
rect 244844 139980 244845 140044
rect 244779 139979 244845 139980
rect 243234 136658 243266 136894
rect 243502 136658 243586 136894
rect 243822 136658 243854 136894
rect 243234 136574 243854 136658
rect 243234 136338 243266 136574
rect 243502 136338 243586 136574
rect 243822 136338 243854 136574
rect 242019 127124 242085 127125
rect 242019 127060 242020 127124
rect 242084 127060 242085 127124
rect 242019 127059 242085 127060
rect 242022 61437 242082 127059
rect 243234 100894 243854 136338
rect 243234 100658 243266 100894
rect 243502 100658 243586 100894
rect 243822 100658 243854 100894
rect 244782 100741 244842 139979
rect 244963 126308 245029 126309
rect 244963 126244 244964 126308
rect 245028 126244 245029 126308
rect 244963 126243 245029 126244
rect 244966 105501 245026 126243
rect 244963 105500 245029 105501
rect 244963 105436 244964 105500
rect 245028 105436 245029 105500
rect 244963 105435 245029 105436
rect 244779 100740 244845 100741
rect 244779 100676 244780 100740
rect 244844 100676 244845 100740
rect 244779 100675 244845 100676
rect 243234 100574 243854 100658
rect 243234 100338 243266 100574
rect 243502 100338 243586 100574
rect 243822 100338 243854 100574
rect 243234 64894 243854 100338
rect 243234 64658 243266 64894
rect 243502 64658 243586 64894
rect 243822 64658 243854 64894
rect 243234 64574 243854 64658
rect 243234 64338 243266 64574
rect 243502 64338 243586 64574
rect 243822 64338 243854 64574
rect 242019 61436 242085 61437
rect 242019 61372 242020 61436
rect 242084 61372 242085 61436
rect 242019 61371 242085 61372
rect 243234 28894 243854 64338
rect 243234 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 243854 28894
rect 243234 28574 243854 28658
rect 243234 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 243854 28574
rect 241283 3364 241349 3365
rect 241283 3300 241284 3364
rect 241348 3300 241349 3364
rect 241283 3299 241349 3300
rect 239514 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 240134 -3226
rect 239514 -3546 240134 -3462
rect 239514 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 240134 -3546
rect 239514 -3814 240134 -3782
rect 243234 -5146 243854 28338
rect 246254 3501 246314 199275
rect 246954 176614 247574 212058
rect 248459 197980 248525 197981
rect 248459 197916 248460 197980
rect 248524 197916 248525 197980
rect 248459 197915 248525 197916
rect 246954 176378 246986 176614
rect 247222 176378 247306 176614
rect 247542 176378 247574 176614
rect 246954 176294 247574 176378
rect 246954 176058 246986 176294
rect 247222 176058 247306 176294
rect 247542 176058 247574 176294
rect 246954 140614 247574 176058
rect 247723 173908 247789 173909
rect 247723 173844 247724 173908
rect 247788 173844 247789 173908
rect 247723 173843 247789 173844
rect 247726 150109 247786 173843
rect 247723 150108 247789 150109
rect 247723 150044 247724 150108
rect 247788 150044 247789 150108
rect 247723 150043 247789 150044
rect 248462 144125 248522 197915
rect 249750 150517 249810 315283
rect 249931 292772 249997 292773
rect 249931 292708 249932 292772
rect 249996 292708 249997 292772
rect 249931 292707 249997 292708
rect 249934 278765 249994 292707
rect 249931 278764 249997 278765
rect 249931 278700 249932 278764
rect 249996 278700 249997 278764
rect 249931 278699 249997 278700
rect 249931 215116 249997 215117
rect 249931 215052 249932 215116
rect 249996 215052 249997 215116
rect 249931 215051 249997 215052
rect 249747 150516 249813 150517
rect 249747 150452 249748 150516
rect 249812 150452 249813 150516
rect 249747 150451 249813 150452
rect 249934 147117 249994 215051
rect 249931 147116 249997 147117
rect 249931 147052 249932 147116
rect 249996 147052 249997 147116
rect 249931 147051 249997 147052
rect 248459 144124 248525 144125
rect 248459 144060 248460 144124
rect 248524 144060 248525 144124
rect 248459 144059 248525 144060
rect 246954 140378 246986 140614
rect 247222 140378 247306 140614
rect 247542 140378 247574 140614
rect 246954 140294 247574 140378
rect 246954 140058 246986 140294
rect 247222 140058 247306 140294
rect 247542 140058 247574 140294
rect 246954 104614 247574 140058
rect 250299 129980 250365 129981
rect 250299 129916 250300 129980
rect 250364 129916 250365 129980
rect 250299 129915 250365 129916
rect 246954 104378 246986 104614
rect 247222 104378 247306 104614
rect 247542 104378 247574 104614
rect 246954 104294 247574 104378
rect 246954 104058 246986 104294
rect 247222 104058 247306 104294
rect 247542 104058 247574 104294
rect 246954 68614 247574 104058
rect 246954 68378 246986 68614
rect 247222 68378 247306 68614
rect 247542 68378 247574 68614
rect 246954 68294 247574 68378
rect 246954 68058 246986 68294
rect 247222 68058 247306 68294
rect 247542 68058 247574 68294
rect 246954 32614 247574 68058
rect 250302 50285 250362 129915
rect 250299 50284 250365 50285
rect 250299 50220 250300 50284
rect 250364 50220 250365 50284
rect 250299 50219 250365 50220
rect 246954 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 247574 32614
rect 246954 32294 247574 32378
rect 246954 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 247574 32294
rect 246251 3500 246317 3501
rect 246251 3436 246252 3500
rect 246316 3436 246317 3500
rect 246251 3435 246317 3436
rect 243234 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 243854 -5146
rect 243234 -5466 243854 -5382
rect 243234 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 243854 -5466
rect 243234 -5734 243854 -5702
rect 228954 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 229574 -6106
rect 228954 -6426 229574 -6342
rect 228954 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 229574 -6426
rect 228954 -7654 229574 -6662
rect 246954 -7066 247574 32058
rect 251774 3501 251834 341395
rect 253794 327454 254414 362898
rect 257514 367174 258134 375600
rect 257514 366938 257546 367174
rect 257782 366938 257866 367174
rect 258102 366938 258134 367174
rect 257514 366854 258134 366938
rect 257514 366618 257546 366854
rect 257782 366618 257866 366854
rect 258102 366618 258134 366854
rect 257514 331174 258134 366618
rect 257514 330938 257546 331174
rect 257782 330938 257866 331174
rect 258102 330938 258134 331174
rect 257514 330854 258134 330938
rect 257514 330618 257546 330854
rect 257782 330618 257866 330854
rect 258102 330618 258134 330854
rect 255267 328540 255333 328541
rect 255267 328476 255268 328540
rect 255332 328476 255333 328540
rect 255267 328475 255333 328476
rect 253794 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 254414 327454
rect 253794 327134 254414 327218
rect 253794 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 254414 327134
rect 253059 322148 253125 322149
rect 253059 322084 253060 322148
rect 253124 322084 253125 322148
rect 253059 322083 253125 322084
rect 253062 22133 253122 322083
rect 253794 291454 254414 326898
rect 253794 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 254414 291454
rect 253794 291134 254414 291218
rect 253794 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 254414 291134
rect 253794 255454 254414 290898
rect 255270 280125 255330 328475
rect 257514 295174 258134 330618
rect 257514 294938 257546 295174
rect 257782 294938 257866 295174
rect 258102 294938 258134 295174
rect 257514 294854 258134 294938
rect 257514 294618 257546 294854
rect 257782 294618 257866 294854
rect 258102 294618 258134 294854
rect 255267 280124 255333 280125
rect 255267 280060 255268 280124
rect 255332 280060 255333 280124
rect 255267 280059 255333 280060
rect 253794 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 254414 255454
rect 253794 255134 254414 255218
rect 253794 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 254414 255134
rect 253794 219454 254414 254898
rect 253794 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 254414 219454
rect 253794 219134 254414 219218
rect 253794 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 254414 219134
rect 253794 183454 254414 218898
rect 253794 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 254414 183454
rect 253794 183134 254414 183218
rect 253794 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 254414 183134
rect 253794 147454 254414 182898
rect 257514 259174 258134 294618
rect 257514 258938 257546 259174
rect 257782 258938 257866 259174
rect 258102 258938 258134 259174
rect 257514 258854 258134 258938
rect 257514 258618 257546 258854
rect 257782 258618 257866 258854
rect 258102 258618 258134 258854
rect 257514 223174 258134 258618
rect 257514 222938 257546 223174
rect 257782 222938 257866 223174
rect 258102 222938 258134 223174
rect 257514 222854 258134 222938
rect 257514 222618 257546 222854
rect 257782 222618 257866 222854
rect 258102 222618 258134 222854
rect 257514 187174 258134 222618
rect 261234 370894 261854 375600
rect 261234 370658 261266 370894
rect 261502 370658 261586 370894
rect 261822 370658 261854 370894
rect 261234 370574 261854 370658
rect 261234 370338 261266 370574
rect 261502 370338 261586 370574
rect 261822 370338 261854 370574
rect 261234 334894 261854 370338
rect 261234 334658 261266 334894
rect 261502 334658 261586 334894
rect 261822 334658 261854 334894
rect 261234 334574 261854 334658
rect 261234 334338 261266 334574
rect 261502 334338 261586 334574
rect 261822 334338 261854 334574
rect 261234 298894 261854 334338
rect 264954 374614 265574 375600
rect 264954 374378 264986 374614
rect 265222 374378 265306 374614
rect 265542 374378 265574 374614
rect 264954 374294 265574 374378
rect 264954 374058 264986 374294
rect 265222 374058 265306 374294
rect 265542 374058 265574 374294
rect 264954 338614 265574 374058
rect 264954 338378 264986 338614
rect 265222 338378 265306 338614
rect 265542 338378 265574 338614
rect 264954 338294 265574 338378
rect 264954 338058 264986 338294
rect 265222 338058 265306 338294
rect 265542 338058 265574 338294
rect 263547 306508 263613 306509
rect 263547 306444 263548 306508
rect 263612 306444 263613 306508
rect 263547 306443 263613 306444
rect 261234 298658 261266 298894
rect 261502 298658 261586 298894
rect 261822 298658 261854 298894
rect 261234 298574 261854 298658
rect 261234 298338 261266 298574
rect 261502 298338 261586 298574
rect 261822 298338 261854 298574
rect 261234 262894 261854 298338
rect 261234 262658 261266 262894
rect 261502 262658 261586 262894
rect 261822 262658 261854 262894
rect 261234 262574 261854 262658
rect 261234 262338 261266 262574
rect 261502 262338 261586 262574
rect 261822 262338 261854 262574
rect 261234 226894 261854 262338
rect 261234 226658 261266 226894
rect 261502 226658 261586 226894
rect 261822 226658 261854 226894
rect 261234 226574 261854 226658
rect 261234 226338 261266 226574
rect 261502 226338 261586 226574
rect 261822 226338 261854 226574
rect 258579 196620 258645 196621
rect 258579 196556 258580 196620
rect 258644 196556 258645 196620
rect 258579 196555 258645 196556
rect 257514 186938 257546 187174
rect 257782 186938 257866 187174
rect 258102 186938 258134 187174
rect 257514 186854 258134 186938
rect 257514 186618 257546 186854
rect 257782 186618 257866 186854
rect 258102 186618 258134 186854
rect 255819 177308 255885 177309
rect 255819 177244 255820 177308
rect 255884 177244 255885 177308
rect 255819 177243 255885 177244
rect 253794 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 254414 147454
rect 253794 147134 254414 147218
rect 253794 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 254414 147134
rect 253794 111454 254414 146898
rect 253794 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 254414 111454
rect 253794 111134 254414 111218
rect 253794 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 254414 111134
rect 253794 75454 254414 110898
rect 255822 91901 255882 177243
rect 257514 151174 258134 186618
rect 257514 150938 257546 151174
rect 257782 150938 257866 151174
rect 258102 150938 258134 151174
rect 257514 150854 258134 150938
rect 257514 150618 257546 150854
rect 257782 150618 257866 150854
rect 258102 150618 258134 150854
rect 257514 115174 258134 150618
rect 257514 114938 257546 115174
rect 257782 114938 257866 115174
rect 258102 114938 258134 115174
rect 257514 114854 258134 114938
rect 257514 114618 257546 114854
rect 257782 114618 257866 114854
rect 258102 114618 258134 114854
rect 255819 91900 255885 91901
rect 255819 91836 255820 91900
rect 255884 91836 255885 91900
rect 255819 91835 255885 91836
rect 253794 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 254414 75454
rect 253794 75134 254414 75218
rect 253794 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 254414 75134
rect 253794 39454 254414 74898
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253059 22132 253125 22133
rect 253059 22068 253060 22132
rect 253124 22068 253125 22132
rect 253059 22067 253125 22068
rect 251771 3500 251837 3501
rect 251771 3436 251772 3500
rect 251836 3436 251837 3500
rect 251771 3435 251837 3436
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -1894 254414 -902
rect 257514 79174 258134 114618
rect 257514 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 258134 79174
rect 257514 78854 258134 78938
rect 257514 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 258134 78854
rect 257514 43174 258134 78618
rect 257514 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 258134 43174
rect 257514 42854 258134 42938
rect 257514 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 258134 42854
rect 257514 7174 258134 42618
rect 258582 37229 258642 196555
rect 261234 190894 261854 226338
rect 261234 190658 261266 190894
rect 261502 190658 261586 190894
rect 261822 190658 261854 190894
rect 261234 190574 261854 190658
rect 261234 190338 261266 190574
rect 261502 190338 261586 190574
rect 261822 190338 261854 190574
rect 261234 154894 261854 190338
rect 261234 154658 261266 154894
rect 261502 154658 261586 154894
rect 261822 154658 261854 154894
rect 261234 154574 261854 154658
rect 261234 154338 261266 154574
rect 261502 154338 261586 154574
rect 261822 154338 261854 154574
rect 261234 118894 261854 154338
rect 262811 131476 262877 131477
rect 262811 131412 262812 131476
rect 262876 131412 262877 131476
rect 262811 131411 262877 131412
rect 261234 118658 261266 118894
rect 261502 118658 261586 118894
rect 261822 118658 261854 118894
rect 261234 118574 261854 118658
rect 261234 118338 261266 118574
rect 261502 118338 261586 118574
rect 261822 118338 261854 118574
rect 260051 103868 260117 103869
rect 260051 103804 260052 103868
rect 260116 103804 260117 103868
rect 260051 103803 260117 103804
rect 260054 93261 260114 103803
rect 260051 93260 260117 93261
rect 260051 93196 260052 93260
rect 260116 93196 260117 93260
rect 260051 93195 260117 93196
rect 261234 82894 261854 118338
rect 261234 82658 261266 82894
rect 261502 82658 261586 82894
rect 261822 82658 261854 82894
rect 261234 82574 261854 82658
rect 261234 82338 261266 82574
rect 261502 82338 261586 82574
rect 261822 82338 261854 82574
rect 261234 46894 261854 82338
rect 262814 71093 262874 131411
rect 263550 109173 263610 306443
rect 264954 302614 265574 338058
rect 264954 302378 264986 302614
rect 265222 302378 265306 302614
rect 265542 302378 265574 302614
rect 264954 302294 265574 302378
rect 264954 302058 264986 302294
rect 265222 302058 265306 302294
rect 265542 302058 265574 302294
rect 264954 266614 265574 302058
rect 264954 266378 264986 266614
rect 265222 266378 265306 266614
rect 265542 266378 265574 266614
rect 264954 266294 265574 266378
rect 264954 266058 264986 266294
rect 265222 266058 265306 266294
rect 265542 266058 265574 266294
rect 264954 230614 265574 266058
rect 264954 230378 264986 230614
rect 265222 230378 265306 230614
rect 265542 230378 265574 230614
rect 264954 230294 265574 230378
rect 264954 230058 264986 230294
rect 265222 230058 265306 230294
rect 265542 230058 265574 230294
rect 264954 194614 265574 230058
rect 264954 194378 264986 194614
rect 265222 194378 265306 194614
rect 265542 194378 265574 194614
rect 264954 194294 265574 194378
rect 264954 194058 264986 194294
rect 265222 194058 265306 194294
rect 265542 194058 265574 194294
rect 264954 158614 265574 194058
rect 271794 345454 272414 375600
rect 271794 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 272414 345454
rect 271794 345134 272414 345218
rect 271794 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 272414 345134
rect 271794 309454 272414 344898
rect 271794 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 272414 309454
rect 271794 309134 272414 309218
rect 271794 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 272414 309134
rect 271794 273454 272414 308898
rect 271794 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 272414 273454
rect 271794 273134 272414 273218
rect 271794 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 272414 273134
rect 271794 237454 272414 272898
rect 271794 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 272414 237454
rect 271794 237134 272414 237218
rect 271794 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 272414 237134
rect 271794 201454 272414 236898
rect 271794 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 272414 201454
rect 271794 201134 272414 201218
rect 271794 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 272414 201134
rect 271794 178000 272414 200898
rect 275514 349174 276134 375600
rect 275514 348938 275546 349174
rect 275782 348938 275866 349174
rect 276102 348938 276134 349174
rect 275514 348854 276134 348938
rect 275514 348618 275546 348854
rect 275782 348618 275866 348854
rect 276102 348618 276134 348854
rect 275514 313174 276134 348618
rect 279234 352894 279854 375600
rect 279234 352658 279266 352894
rect 279502 352658 279586 352894
rect 279822 352658 279854 352894
rect 279234 352574 279854 352658
rect 279234 352338 279266 352574
rect 279502 352338 279586 352574
rect 279822 352338 279854 352574
rect 279234 316894 279854 352338
rect 279234 316658 279266 316894
rect 279502 316658 279586 316894
rect 279822 316658 279854 316894
rect 279234 316574 279854 316658
rect 279234 316338 279266 316574
rect 279502 316338 279586 316574
rect 279822 316338 279854 316574
rect 277899 314804 277965 314805
rect 277899 314740 277900 314804
rect 277964 314740 277965 314804
rect 277899 314739 277965 314740
rect 275514 312938 275546 313174
rect 275782 312938 275866 313174
rect 276102 312938 276134 313174
rect 275514 312854 276134 312938
rect 275514 312618 275546 312854
rect 275782 312618 275866 312854
rect 276102 312618 276134 312854
rect 275514 277174 276134 312618
rect 275514 276938 275546 277174
rect 275782 276938 275866 277174
rect 276102 276938 276134 277174
rect 275514 276854 276134 276938
rect 275514 276618 275546 276854
rect 275782 276618 275866 276854
rect 276102 276618 276134 276854
rect 275514 241174 276134 276618
rect 275514 240938 275546 241174
rect 275782 240938 275866 241174
rect 276102 240938 276134 241174
rect 275514 240854 276134 240938
rect 275514 240618 275546 240854
rect 275782 240618 275866 240854
rect 276102 240618 276134 240854
rect 275514 205174 276134 240618
rect 275514 204938 275546 205174
rect 275782 204938 275866 205174
rect 276102 204938 276134 205174
rect 275514 204854 276134 204938
rect 275514 204618 275546 204854
rect 275782 204618 275866 204854
rect 276102 204618 276134 204854
rect 275514 178000 276134 204618
rect 277902 175130 277962 314739
rect 279234 280894 279854 316338
rect 282954 356614 283574 375600
rect 288387 375324 288453 375325
rect 288387 375260 288388 375324
rect 288452 375260 288453 375324
rect 288387 375259 288453 375260
rect 285627 365804 285693 365805
rect 285627 365740 285628 365804
rect 285692 365740 285693 365804
rect 285627 365739 285693 365740
rect 282954 356378 282986 356614
rect 283222 356378 283306 356614
rect 283542 356378 283574 356614
rect 282954 356294 283574 356378
rect 282954 356058 282986 356294
rect 283222 356058 283306 356294
rect 283542 356058 283574 356294
rect 282954 320614 283574 356058
rect 282954 320378 282986 320614
rect 283222 320378 283306 320614
rect 283542 320378 283574 320614
rect 282954 320294 283574 320378
rect 282954 320058 282986 320294
rect 283222 320058 283306 320294
rect 283542 320058 283574 320294
rect 281579 307732 281645 307733
rect 281579 307668 281580 307732
rect 281644 307668 281645 307732
rect 281579 307667 281645 307668
rect 279234 280658 279266 280894
rect 279502 280658 279586 280894
rect 279822 280658 279854 280894
rect 279234 280574 279854 280658
rect 279234 280338 279266 280574
rect 279502 280338 279586 280574
rect 279822 280338 279854 280574
rect 279234 244894 279854 280338
rect 279234 244658 279266 244894
rect 279502 244658 279586 244894
rect 279822 244658 279854 244894
rect 279234 244574 279854 244658
rect 279234 244338 279266 244574
rect 279502 244338 279586 244574
rect 279822 244338 279854 244574
rect 279234 208894 279854 244338
rect 279234 208658 279266 208894
rect 279502 208658 279586 208894
rect 279822 208658 279854 208894
rect 279234 208574 279854 208658
rect 279234 208338 279266 208574
rect 279502 208338 279586 208574
rect 279822 208338 279854 208574
rect 279003 178668 279069 178669
rect 279003 178604 279004 178668
rect 279068 178604 279069 178668
rect 279003 178603 279069 178604
rect 279006 177850 279066 178603
rect 279234 178000 279854 208338
rect 280475 183156 280541 183157
rect 280475 183092 280476 183156
rect 280540 183092 280541 183156
rect 280475 183091 280541 183092
rect 280291 181524 280357 181525
rect 280291 181460 280292 181524
rect 280356 181460 280357 181524
rect 280291 181459 280357 181460
rect 279006 177790 279618 177850
rect 279371 177308 279437 177309
rect 279371 177244 279372 177308
rect 279436 177244 279437 177308
rect 279371 177243 279437 177244
rect 279374 175269 279434 177243
rect 279371 175268 279437 175269
rect 279371 175204 279372 175268
rect 279436 175204 279437 175268
rect 279371 175203 279437 175204
rect 277902 175070 278882 175130
rect 278822 173770 278882 175070
rect 279371 173772 279437 173773
rect 279371 173770 279372 173772
rect 278822 173710 279372 173770
rect 279371 173708 279372 173710
rect 279436 173708 279437 173772
rect 279371 173707 279437 173708
rect 279558 170645 279618 177790
rect 280107 172412 280173 172413
rect 280107 172348 280108 172412
rect 280172 172348 280173 172412
rect 280107 172347 280173 172348
rect 279555 170644 279621 170645
rect 279555 170580 279556 170644
rect 279620 170580 279621 170644
rect 279555 170579 279621 170580
rect 272207 165454 272527 165486
rect 272207 165218 272249 165454
rect 272485 165218 272527 165454
rect 272207 165134 272527 165218
rect 272207 164898 272249 165134
rect 272485 164898 272527 165134
rect 272207 164866 272527 164898
rect 275471 165454 275791 165486
rect 275471 165218 275513 165454
rect 275749 165218 275791 165454
rect 275471 165134 275791 165218
rect 275471 164898 275513 165134
rect 275749 164898 275791 165134
rect 275471 164866 275791 164898
rect 280110 161490 280170 172347
rect 264954 158378 264986 158614
rect 265222 158378 265306 158614
rect 265542 158378 265574 158614
rect 264954 158294 265574 158378
rect 264954 158058 264986 158294
rect 265222 158058 265306 158294
rect 265542 158058 265574 158294
rect 264099 133108 264165 133109
rect 264099 133044 264100 133108
rect 264164 133044 264165 133108
rect 264099 133043 264165 133044
rect 263547 109172 263613 109173
rect 263547 109108 263548 109172
rect 263612 109108 263613 109172
rect 263547 109107 263613 109108
rect 263547 103052 263613 103053
rect 263547 102988 263548 103052
rect 263612 102988 263613 103052
rect 263547 102987 263613 102988
rect 263550 95845 263610 102987
rect 263547 95844 263613 95845
rect 263547 95780 263548 95844
rect 263612 95780 263613 95844
rect 263547 95779 263613 95780
rect 262811 71092 262877 71093
rect 262811 71028 262812 71092
rect 262876 71028 262877 71092
rect 262811 71027 262877 71028
rect 261234 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 261854 46894
rect 261234 46574 261854 46658
rect 261234 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 261854 46574
rect 258579 37228 258645 37229
rect 258579 37164 258580 37228
rect 258644 37164 258645 37228
rect 258579 37163 258645 37164
rect 257514 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 258134 7174
rect 257514 6854 258134 6938
rect 257514 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 258134 6854
rect 257514 -2266 258134 6618
rect 257514 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 258134 -2266
rect 257514 -2586 258134 -2502
rect 257514 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 258134 -2586
rect 257514 -3814 258134 -2822
rect 261234 10894 261854 46338
rect 264102 44845 264162 133043
rect 264954 122614 265574 158058
rect 278822 161430 280170 161490
rect 278822 157350 278882 161430
rect 278822 157290 279434 157350
rect 270575 147454 270895 147486
rect 270575 147218 270617 147454
rect 270853 147218 270895 147454
rect 270575 147134 270895 147218
rect 270575 146898 270617 147134
rect 270853 146898 270895 147134
rect 270575 146866 270895 146898
rect 273839 147454 274159 147486
rect 273839 147218 273881 147454
rect 274117 147218 274159 147454
rect 273839 147134 274159 147218
rect 273839 146898 273881 147134
rect 274117 146898 274159 147134
rect 273839 146866 274159 146898
rect 277103 147454 277423 147486
rect 277103 147218 277145 147454
rect 277381 147218 277423 147454
rect 277103 147134 277423 147218
rect 277103 146898 277145 147134
rect 277381 146898 277423 147134
rect 277103 146866 277423 146898
rect 266859 140452 266925 140453
rect 266859 140388 266860 140452
rect 266924 140388 266925 140452
rect 266859 140387 266925 140388
rect 264954 122378 264986 122614
rect 265222 122378 265306 122614
rect 265542 122378 265574 122614
rect 264954 122294 265574 122378
rect 264954 122058 264986 122294
rect 265222 122058 265306 122294
rect 265542 122058 265574 122294
rect 264954 86614 265574 122058
rect 264954 86378 264986 86614
rect 265222 86378 265306 86614
rect 265542 86378 265574 86614
rect 264954 86294 265574 86378
rect 264954 86058 264986 86294
rect 265222 86058 265306 86294
rect 265542 86058 265574 86294
rect 264954 50614 265574 86058
rect 264954 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 265574 50614
rect 264954 50294 265574 50378
rect 264954 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 265574 50294
rect 264099 44844 264165 44845
rect 264099 44780 264100 44844
rect 264164 44780 264165 44844
rect 264099 44779 264165 44780
rect 261234 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 261854 10894
rect 261234 10574 261854 10658
rect 261234 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 261854 10574
rect 261234 -4186 261854 10338
rect 261234 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 261854 -4186
rect 261234 -4506 261854 -4422
rect 261234 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 261854 -4506
rect 261234 -5734 261854 -4742
rect 264954 14614 265574 50058
rect 266862 35189 266922 140387
rect 267779 138684 267845 138685
rect 267779 138620 267780 138684
rect 267844 138620 267845 138684
rect 267779 138619 267845 138620
rect 267595 128484 267661 128485
rect 267595 128420 267596 128484
rect 267660 128420 267661 128484
rect 267595 128419 267661 128420
rect 267598 93261 267658 128419
rect 267595 93260 267661 93261
rect 267595 93196 267596 93260
rect 267660 93196 267661 93260
rect 267595 93195 267661 93196
rect 267782 92581 267842 138619
rect 279374 135285 279434 157290
rect 279371 135284 279437 135285
rect 279371 135220 279372 135284
rect 279436 135220 279437 135284
rect 279371 135219 279437 135220
rect 272207 129454 272527 129486
rect 272207 129218 272249 129454
rect 272485 129218 272527 129454
rect 272207 129134 272527 129218
rect 272207 128898 272249 129134
rect 272485 128898 272527 129134
rect 272207 128866 272527 128898
rect 275471 129454 275791 129486
rect 275471 129218 275513 129454
rect 275749 129218 275791 129454
rect 275471 129134 275791 129218
rect 275471 128898 275513 129134
rect 275749 128898 275791 129134
rect 275471 128866 275791 128898
rect 280294 126853 280354 181459
rect 280478 172413 280538 183091
rect 280475 172412 280541 172413
rect 280475 172348 280476 172412
rect 280540 172348 280541 172412
rect 280475 172347 280541 172348
rect 281582 156501 281642 307667
rect 282954 284614 283574 320058
rect 282954 284378 282986 284614
rect 283222 284378 283306 284614
rect 283542 284378 283574 284614
rect 282954 284294 283574 284378
rect 282954 284058 282986 284294
rect 283222 284058 283306 284294
rect 283542 284058 283574 284294
rect 281763 268428 281829 268429
rect 281763 268364 281764 268428
rect 281828 268364 281829 268428
rect 281763 268363 281829 268364
rect 281766 157317 281826 268363
rect 282954 248614 283574 284058
rect 282954 248378 282986 248614
rect 283222 248378 283306 248614
rect 283542 248378 283574 248614
rect 282954 248294 283574 248378
rect 282954 248058 282986 248294
rect 283222 248058 283306 248294
rect 283542 248058 283574 248294
rect 282954 212614 283574 248058
rect 282954 212378 282986 212614
rect 283222 212378 283306 212614
rect 283542 212378 283574 212614
rect 282954 212294 283574 212378
rect 282954 212058 282986 212294
rect 283222 212058 283306 212294
rect 283542 212058 283574 212294
rect 282954 176614 283574 212058
rect 284523 188460 284589 188461
rect 284523 188396 284524 188460
rect 284588 188396 284589 188460
rect 284523 188395 284589 188396
rect 284339 178804 284405 178805
rect 284339 178740 284340 178804
rect 284404 178740 284405 178804
rect 284339 178739 284405 178740
rect 283787 177444 283853 177445
rect 283787 177380 283788 177444
rect 283852 177380 283853 177444
rect 283787 177379 283853 177380
rect 282954 176378 282986 176614
rect 283222 176378 283306 176614
rect 283542 176378 283574 176614
rect 282954 176294 283574 176378
rect 282954 176058 282986 176294
rect 283222 176058 283306 176294
rect 283542 176058 283574 176294
rect 281763 157316 281829 157317
rect 281763 157252 281764 157316
rect 281828 157252 281829 157316
rect 281763 157251 281829 157252
rect 281579 156500 281645 156501
rect 281579 156436 281580 156500
rect 281644 156436 281645 156500
rect 281579 156435 281645 156436
rect 282954 140614 283574 176058
rect 283790 146573 283850 177379
rect 283787 146572 283853 146573
rect 283787 146508 283788 146572
rect 283852 146508 283853 146572
rect 283787 146507 283853 146508
rect 282954 140378 282986 140614
rect 283222 140378 283306 140614
rect 283542 140378 283574 140614
rect 282954 140294 283574 140378
rect 282954 140058 282986 140294
rect 283222 140058 283306 140294
rect 283542 140058 283574 140294
rect 280291 126852 280357 126853
rect 280291 126788 280292 126852
rect 280356 126788 280357 126852
rect 280291 126787 280357 126788
rect 270575 111454 270895 111486
rect 270575 111218 270617 111454
rect 270853 111218 270895 111454
rect 270575 111134 270895 111218
rect 270575 110898 270617 111134
rect 270853 110898 270895 111134
rect 270575 110866 270895 110898
rect 273839 111454 274159 111486
rect 273839 111218 273881 111454
rect 274117 111218 274159 111454
rect 273839 111134 274159 111218
rect 273839 110898 273881 111134
rect 274117 110898 274159 111134
rect 273839 110866 274159 110898
rect 277103 111454 277423 111486
rect 277103 111218 277145 111454
rect 277381 111218 277423 111454
rect 277103 111134 277423 111218
rect 277103 110898 277145 111134
rect 277381 110898 277423 111134
rect 277103 110866 277423 110898
rect 282954 104614 283574 140058
rect 282954 104378 282986 104614
rect 283222 104378 283306 104614
rect 283542 104378 283574 104614
rect 282954 104294 283574 104378
rect 282954 104058 282986 104294
rect 283222 104058 283306 104294
rect 283542 104058 283574 104294
rect 268515 96796 268581 96797
rect 268515 96732 268516 96796
rect 268580 96732 268581 96796
rect 268515 96731 268581 96732
rect 268518 95029 268578 96731
rect 268515 95028 268581 95029
rect 268515 94964 268516 95028
rect 268580 94964 268581 95028
rect 268515 94963 268581 94964
rect 271794 93454 272414 94000
rect 271794 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 272414 93454
rect 271794 93134 272414 93218
rect 271794 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 272414 93134
rect 267779 92580 267845 92581
rect 267779 92516 267780 92580
rect 267844 92516 267845 92580
rect 267779 92515 267845 92516
rect 271794 57454 272414 92898
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 266859 35188 266925 35189
rect 266859 35124 266860 35188
rect 266924 35124 266925 35188
rect 266859 35123 266925 35124
rect 264954 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 265574 14614
rect 264954 14294 265574 14378
rect 264954 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 265574 14294
rect 246954 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 247574 -7066
rect 246954 -7386 247574 -7302
rect 246954 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 247574 -7386
rect 246954 -7654 247574 -7622
rect 264954 -6106 265574 14058
rect 271794 21454 272414 56898
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -1306 272414 20898
rect 271794 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 272414 -1306
rect 271794 -1626 272414 -1542
rect 271794 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 272414 -1626
rect 271794 -1894 272414 -1862
rect 275514 61174 276134 94000
rect 275514 60938 275546 61174
rect 275782 60938 275866 61174
rect 276102 60938 276134 61174
rect 275514 60854 276134 60938
rect 275514 60618 275546 60854
rect 275782 60618 275866 60854
rect 276102 60618 276134 60854
rect 275514 25174 276134 60618
rect 275514 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 276134 25174
rect 275514 24854 276134 24938
rect 275514 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 276134 24854
rect 275514 -3226 276134 24618
rect 275514 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 276134 -3226
rect 275514 -3546 276134 -3462
rect 275514 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 276134 -3546
rect 275514 -3814 276134 -3782
rect 279234 64894 279854 94000
rect 279234 64658 279266 64894
rect 279502 64658 279586 64894
rect 279822 64658 279854 64894
rect 279234 64574 279854 64658
rect 279234 64338 279266 64574
rect 279502 64338 279586 64574
rect 279822 64338 279854 64574
rect 279234 28894 279854 64338
rect 279234 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 279854 28894
rect 279234 28574 279854 28658
rect 279234 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 279854 28574
rect 279234 -5146 279854 28338
rect 279234 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 279854 -5146
rect 279234 -5466 279854 -5382
rect 279234 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 279854 -5466
rect 279234 -5734 279854 -5702
rect 282954 68614 283574 104058
rect 284342 97069 284402 178739
rect 284526 140453 284586 188395
rect 284523 140452 284589 140453
rect 284523 140388 284524 140452
rect 284588 140388 284589 140452
rect 284523 140387 284589 140388
rect 284339 97068 284405 97069
rect 284339 97004 284340 97068
rect 284404 97004 284405 97068
rect 284339 97003 284405 97004
rect 282954 68378 282986 68614
rect 283222 68378 283306 68614
rect 283542 68378 283574 68614
rect 282954 68294 283574 68378
rect 282954 68058 282986 68294
rect 283222 68058 283306 68294
rect 283542 68058 283574 68294
rect 282954 32614 283574 68058
rect 282954 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 283574 32614
rect 282954 32294 283574 32378
rect 282954 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 283574 32294
rect 264954 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 265574 -6106
rect 264954 -6426 265574 -6342
rect 264954 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 265574 -6426
rect 264954 -7654 265574 -6662
rect 282954 -7066 283574 32058
rect 285630 3501 285690 365739
rect 288390 189685 288450 375259
rect 289794 363454 290414 375600
rect 289794 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 290414 363454
rect 289794 363134 290414 363218
rect 289794 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 290414 363134
rect 289794 327454 290414 362898
rect 289794 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 290414 327454
rect 289794 327134 290414 327218
rect 289794 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 290414 327134
rect 289794 291454 290414 326898
rect 293514 367174 294134 375600
rect 293514 366938 293546 367174
rect 293782 366938 293866 367174
rect 294102 366938 294134 367174
rect 293514 366854 294134 366938
rect 293514 366618 293546 366854
rect 293782 366618 293866 366854
rect 294102 366618 294134 366854
rect 293514 331174 294134 366618
rect 297234 370894 297854 375600
rect 297234 370658 297266 370894
rect 297502 370658 297586 370894
rect 297822 370658 297854 370894
rect 297234 370574 297854 370658
rect 297234 370338 297266 370574
rect 297502 370338 297586 370574
rect 297822 370338 297854 370574
rect 295379 343772 295445 343773
rect 295379 343708 295380 343772
rect 295444 343708 295445 343772
rect 295379 343707 295445 343708
rect 293514 330938 293546 331174
rect 293782 330938 293866 331174
rect 294102 330938 294134 331174
rect 293514 330854 294134 330938
rect 293514 330618 293546 330854
rect 293782 330618 293866 330854
rect 294102 330618 294134 330854
rect 291147 323644 291213 323645
rect 291147 323580 291148 323644
rect 291212 323580 291213 323644
rect 291147 323579 291213 323580
rect 289794 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 290414 291454
rect 289794 291134 290414 291218
rect 289794 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 290414 291134
rect 289794 255454 290414 290898
rect 289794 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 290414 255454
rect 289794 255134 290414 255218
rect 289794 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 290414 255134
rect 289794 219454 290414 254898
rect 289794 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 290414 219454
rect 289794 219134 290414 219218
rect 289794 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 290414 219134
rect 287651 189684 287717 189685
rect 287651 189620 287652 189684
rect 287716 189620 287717 189684
rect 287651 189619 287717 189620
rect 288387 189684 288453 189685
rect 288387 189620 288388 189684
rect 288452 189620 288453 189684
rect 288387 189619 288453 189620
rect 287099 180300 287165 180301
rect 287099 180236 287100 180300
rect 287164 180236 287165 180300
rect 287099 180235 287165 180236
rect 285811 176900 285877 176901
rect 285811 176836 285812 176900
rect 285876 176836 285877 176900
rect 285811 176835 285877 176836
rect 285814 102373 285874 176835
rect 287102 167109 287162 180235
rect 287099 167108 287165 167109
rect 287099 167044 287100 167108
rect 287164 167044 287165 167108
rect 287099 167043 287165 167044
rect 285811 102372 285877 102373
rect 285811 102308 285812 102372
rect 285876 102308 285877 102372
rect 285811 102307 285877 102308
rect 287654 3501 287714 189619
rect 289794 183454 290414 218898
rect 289794 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 290414 183454
rect 289794 183134 290414 183218
rect 288571 183020 288637 183021
rect 288571 182956 288572 183020
rect 288636 182956 288637 183020
rect 288571 182955 288637 182956
rect 288574 143581 288634 182955
rect 289794 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 290414 183134
rect 289794 147454 290414 182898
rect 290595 180164 290661 180165
rect 290595 180100 290596 180164
rect 290660 180100 290661 180164
rect 290595 180099 290661 180100
rect 289794 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 290414 147454
rect 289794 147134 290414 147218
rect 289794 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 290414 147134
rect 288571 143580 288637 143581
rect 288571 143516 288572 143580
rect 288636 143516 288637 143580
rect 288571 143515 288637 143516
rect 289794 111454 290414 146898
rect 290598 117333 290658 180099
rect 290595 117332 290661 117333
rect 290595 117268 290596 117332
rect 290660 117268 290661 117332
rect 290595 117267 290661 117268
rect 289794 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 290414 111454
rect 289794 111134 290414 111218
rect 289794 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 290414 111134
rect 289794 75454 290414 110898
rect 289794 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 290414 75454
rect 289794 75134 290414 75218
rect 289794 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 290414 75134
rect 289794 39454 290414 74898
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 285627 3500 285693 3501
rect 285627 3436 285628 3500
rect 285692 3436 285693 3500
rect 285627 3435 285693 3436
rect 287651 3500 287717 3501
rect 287651 3436 287652 3500
rect 287716 3436 287717 3500
rect 287651 3435 287717 3436
rect 289794 3454 290414 38898
rect 291150 3501 291210 323579
rect 293514 295174 294134 330618
rect 293514 294938 293546 295174
rect 293782 294938 293866 295174
rect 294102 294938 294134 295174
rect 293514 294854 294134 294938
rect 293514 294618 293546 294854
rect 293782 294618 293866 294854
rect 294102 294618 294134 294854
rect 293514 259174 294134 294618
rect 293514 258938 293546 259174
rect 293782 258938 293866 259174
rect 294102 258938 294134 259174
rect 293514 258854 294134 258938
rect 293514 258618 293546 258854
rect 293782 258618 293866 258854
rect 294102 258618 294134 258854
rect 293514 223174 294134 258618
rect 293514 222938 293546 223174
rect 293782 222938 293866 223174
rect 294102 222938 294134 223174
rect 293514 222854 294134 222938
rect 293514 222618 293546 222854
rect 293782 222618 293866 222854
rect 294102 222618 294134 222854
rect 293171 207636 293237 207637
rect 293171 207572 293172 207636
rect 293236 207572 293237 207636
rect 293171 207571 293237 207572
rect 293174 3501 293234 207571
rect 293514 187174 294134 222618
rect 293514 186938 293546 187174
rect 293782 186938 293866 187174
rect 294102 186938 294134 187174
rect 293514 186854 294134 186938
rect 293514 186618 293546 186854
rect 293782 186618 293866 186854
rect 294102 186618 294134 186854
rect 293514 151174 294134 186618
rect 293514 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 294134 151174
rect 293514 150854 294134 150938
rect 293514 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 294134 150854
rect 293514 115174 294134 150618
rect 293514 114938 293546 115174
rect 293782 114938 293866 115174
rect 294102 114938 294134 115174
rect 293514 114854 294134 114938
rect 293514 114618 293546 114854
rect 293782 114618 293866 114854
rect 294102 114618 294134 114854
rect 293514 79174 294134 114618
rect 293514 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 294134 79174
rect 293514 78854 294134 78938
rect 293514 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 294134 78854
rect 293514 43174 294134 78618
rect 293514 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 294134 43174
rect 293514 42854 294134 42938
rect 293514 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 294134 42854
rect 293514 7174 294134 42618
rect 295382 22677 295442 343707
rect 297234 334894 297854 370338
rect 297234 334658 297266 334894
rect 297502 334658 297586 334894
rect 297822 334658 297854 334894
rect 297234 334574 297854 334658
rect 297234 334338 297266 334574
rect 297502 334338 297586 334574
rect 297822 334338 297854 334574
rect 297234 298894 297854 334338
rect 297234 298658 297266 298894
rect 297502 298658 297586 298894
rect 297822 298658 297854 298894
rect 297234 298574 297854 298658
rect 297234 298338 297266 298574
rect 297502 298338 297586 298574
rect 297822 298338 297854 298574
rect 297234 262894 297854 298338
rect 297234 262658 297266 262894
rect 297502 262658 297586 262894
rect 297822 262658 297854 262894
rect 297234 262574 297854 262658
rect 297234 262338 297266 262574
rect 297502 262338 297586 262574
rect 297822 262338 297854 262574
rect 297234 226894 297854 262338
rect 297234 226658 297266 226894
rect 297502 226658 297586 226894
rect 297822 226658 297854 226894
rect 297234 226574 297854 226658
rect 297234 226338 297266 226574
rect 297502 226338 297586 226574
rect 297822 226338 297854 226574
rect 297234 190894 297854 226338
rect 300954 374614 301574 375600
rect 300954 374378 300986 374614
rect 301222 374378 301306 374614
rect 301542 374378 301574 374614
rect 300954 374294 301574 374378
rect 300954 374058 300986 374294
rect 301222 374058 301306 374294
rect 301542 374058 301574 374294
rect 300954 338614 301574 374058
rect 303659 374100 303725 374101
rect 303659 374036 303660 374100
rect 303724 374036 303725 374100
rect 303659 374035 303725 374036
rect 300954 338378 300986 338614
rect 301222 338378 301306 338614
rect 301542 338378 301574 338614
rect 300954 338294 301574 338378
rect 300954 338058 300986 338294
rect 301222 338058 301306 338294
rect 301542 338058 301574 338294
rect 300954 302614 301574 338058
rect 300954 302378 300986 302614
rect 301222 302378 301306 302614
rect 301542 302378 301574 302614
rect 300954 302294 301574 302378
rect 300954 302058 300986 302294
rect 301222 302058 301306 302294
rect 301542 302058 301574 302294
rect 300954 266614 301574 302058
rect 300954 266378 300986 266614
rect 301222 266378 301306 266614
rect 301542 266378 301574 266614
rect 300954 266294 301574 266378
rect 300954 266058 300986 266294
rect 301222 266058 301306 266294
rect 301542 266058 301574 266294
rect 300954 230614 301574 266058
rect 300954 230378 300986 230614
rect 301222 230378 301306 230614
rect 301542 230378 301574 230614
rect 300954 230294 301574 230378
rect 300954 230058 300986 230294
rect 301222 230058 301306 230294
rect 301542 230058 301574 230294
rect 298139 217292 298205 217293
rect 298139 217228 298140 217292
rect 298204 217228 298205 217292
rect 298139 217227 298205 217228
rect 297234 190658 297266 190894
rect 297502 190658 297586 190894
rect 297822 190658 297854 190894
rect 297234 190574 297854 190658
rect 297234 190338 297266 190574
rect 297502 190338 297586 190574
rect 297822 190338 297854 190574
rect 297234 154894 297854 190338
rect 297234 154658 297266 154894
rect 297502 154658 297586 154894
rect 297822 154658 297854 154894
rect 297234 154574 297854 154658
rect 297234 154338 297266 154574
rect 297502 154338 297586 154574
rect 297822 154338 297854 154574
rect 297234 118894 297854 154338
rect 297234 118658 297266 118894
rect 297502 118658 297586 118894
rect 297822 118658 297854 118894
rect 297234 118574 297854 118658
rect 297234 118338 297266 118574
rect 297502 118338 297586 118574
rect 297822 118338 297854 118574
rect 297234 82894 297854 118338
rect 297234 82658 297266 82894
rect 297502 82658 297586 82894
rect 297822 82658 297854 82894
rect 297234 82574 297854 82658
rect 297234 82338 297266 82574
rect 297502 82338 297586 82574
rect 297822 82338 297854 82574
rect 297234 46894 297854 82338
rect 297234 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 297854 46894
rect 297234 46574 297854 46658
rect 297234 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 297854 46574
rect 295379 22676 295445 22677
rect 295379 22612 295380 22676
rect 295444 22612 295445 22676
rect 295379 22611 295445 22612
rect 293514 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 294134 7174
rect 293514 6854 294134 6938
rect 293514 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 294134 6854
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 291147 3500 291213 3501
rect 291147 3436 291148 3500
rect 291212 3436 291213 3500
rect 291147 3435 291213 3436
rect 293171 3500 293237 3501
rect 293171 3436 293172 3500
rect 293236 3436 293237 3500
rect 293171 3435 293237 3436
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -1894 290414 -902
rect 293514 -2266 294134 6618
rect 293514 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 294134 -2266
rect 293514 -2586 294134 -2502
rect 293514 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 294134 -2586
rect 293514 -3814 294134 -2822
rect 297234 10894 297854 46338
rect 297234 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 297854 10894
rect 297234 10574 297854 10658
rect 297234 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 297854 10574
rect 297234 -4186 297854 10338
rect 298142 3365 298202 217227
rect 300954 194614 301574 230058
rect 302739 214708 302805 214709
rect 302739 214644 302740 214708
rect 302804 214644 302805 214708
rect 302739 214643 302805 214644
rect 300954 194378 300986 194614
rect 301222 194378 301306 194614
rect 301542 194378 301574 194614
rect 300954 194294 301574 194378
rect 300954 194058 300986 194294
rect 301222 194058 301306 194294
rect 301542 194058 301574 194294
rect 299611 185060 299677 185061
rect 299611 184996 299612 185060
rect 299676 184996 299677 185060
rect 299611 184995 299677 184996
rect 299614 3501 299674 184995
rect 300954 158614 301574 194058
rect 300954 158378 300986 158614
rect 301222 158378 301306 158614
rect 301542 158378 301574 158614
rect 300954 158294 301574 158378
rect 300954 158058 300986 158294
rect 301222 158058 301306 158294
rect 301542 158058 301574 158294
rect 300954 122614 301574 158058
rect 300954 122378 300986 122614
rect 301222 122378 301306 122614
rect 301542 122378 301574 122614
rect 300954 122294 301574 122378
rect 300954 122058 300986 122294
rect 301222 122058 301306 122294
rect 301542 122058 301574 122294
rect 300954 86614 301574 122058
rect 300954 86378 300986 86614
rect 301222 86378 301306 86614
rect 301542 86378 301574 86614
rect 300954 86294 301574 86378
rect 300954 86058 300986 86294
rect 301222 86058 301306 86294
rect 301542 86058 301574 86294
rect 300954 50614 301574 86058
rect 300954 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 301574 50614
rect 300954 50294 301574 50378
rect 300954 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 301574 50294
rect 300954 14614 301574 50058
rect 300954 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 301574 14614
rect 300954 14294 301574 14378
rect 300954 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 301574 14294
rect 299611 3500 299677 3501
rect 299611 3436 299612 3500
rect 299676 3436 299677 3500
rect 299611 3435 299677 3436
rect 298139 3364 298205 3365
rect 298139 3300 298140 3364
rect 298204 3300 298205 3364
rect 298139 3299 298205 3300
rect 297234 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 297854 -4186
rect 297234 -4506 297854 -4422
rect 297234 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 297854 -4506
rect 297234 -5734 297854 -4742
rect 282954 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 283574 -7066
rect 282954 -7386 283574 -7302
rect 282954 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 283574 -7386
rect 282954 -7654 283574 -7622
rect 300954 -6106 301574 14058
rect 302742 3365 302802 214643
rect 303662 19957 303722 374035
rect 307794 345454 308414 375600
rect 307794 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 308414 345454
rect 307794 345134 308414 345218
rect 307794 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 308414 345134
rect 307794 309454 308414 344898
rect 307794 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 308414 309454
rect 307794 309134 308414 309218
rect 307794 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 308414 309134
rect 307794 273454 308414 308898
rect 307794 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 308414 273454
rect 307794 273134 308414 273218
rect 307794 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 308414 273134
rect 307794 237454 308414 272898
rect 307794 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 308414 237454
rect 307794 237134 308414 237218
rect 307794 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 308414 237134
rect 307794 201454 308414 236898
rect 307794 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 308414 201454
rect 307794 201134 308414 201218
rect 307794 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 308414 201134
rect 307794 165454 308414 200898
rect 307794 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 308414 165454
rect 307794 165134 308414 165218
rect 307794 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 308414 165134
rect 307794 129454 308414 164898
rect 307794 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 308414 129454
rect 307794 129134 308414 129218
rect 307794 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 308414 129134
rect 307794 93454 308414 128898
rect 307794 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 308414 93454
rect 307794 93134 308414 93218
rect 307794 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 308414 93134
rect 307794 57454 308414 92898
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 303659 19956 303725 19957
rect 303659 19892 303660 19956
rect 303724 19892 303725 19956
rect 303659 19891 303725 19892
rect 302739 3364 302805 3365
rect 302739 3300 302740 3364
rect 302804 3300 302805 3364
rect 302739 3299 302805 3300
rect 307794 -1306 308414 20898
rect 307794 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 308414 -1306
rect 307794 -1626 308414 -1542
rect 307794 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 308414 -1626
rect 307794 -1894 308414 -1862
rect 311514 349174 312134 375600
rect 311514 348938 311546 349174
rect 311782 348938 311866 349174
rect 312102 348938 312134 349174
rect 311514 348854 312134 348938
rect 311514 348618 311546 348854
rect 311782 348618 311866 348854
rect 312102 348618 312134 348854
rect 311514 313174 312134 348618
rect 311514 312938 311546 313174
rect 311782 312938 311866 313174
rect 312102 312938 312134 313174
rect 311514 312854 312134 312938
rect 311514 312618 311546 312854
rect 311782 312618 311866 312854
rect 312102 312618 312134 312854
rect 311514 277174 312134 312618
rect 311514 276938 311546 277174
rect 311782 276938 311866 277174
rect 312102 276938 312134 277174
rect 311514 276854 312134 276938
rect 311514 276618 311546 276854
rect 311782 276618 311866 276854
rect 312102 276618 312134 276854
rect 311514 241174 312134 276618
rect 311514 240938 311546 241174
rect 311782 240938 311866 241174
rect 312102 240938 312134 241174
rect 311514 240854 312134 240938
rect 311514 240618 311546 240854
rect 311782 240618 311866 240854
rect 312102 240618 312134 240854
rect 311514 205174 312134 240618
rect 311514 204938 311546 205174
rect 311782 204938 311866 205174
rect 312102 204938 312134 205174
rect 311514 204854 312134 204938
rect 311514 204618 311546 204854
rect 311782 204618 311866 204854
rect 312102 204618 312134 204854
rect 311514 169174 312134 204618
rect 311514 168938 311546 169174
rect 311782 168938 311866 169174
rect 312102 168938 312134 169174
rect 311514 168854 312134 168938
rect 311514 168618 311546 168854
rect 311782 168618 311866 168854
rect 312102 168618 312134 168854
rect 311514 133174 312134 168618
rect 311514 132938 311546 133174
rect 311782 132938 311866 133174
rect 312102 132938 312134 133174
rect 311514 132854 312134 132938
rect 311514 132618 311546 132854
rect 311782 132618 311866 132854
rect 312102 132618 312134 132854
rect 311514 97174 312134 132618
rect 311514 96938 311546 97174
rect 311782 96938 311866 97174
rect 312102 96938 312134 97174
rect 311514 96854 312134 96938
rect 311514 96618 311546 96854
rect 311782 96618 311866 96854
rect 312102 96618 312134 96854
rect 311514 61174 312134 96618
rect 311514 60938 311546 61174
rect 311782 60938 311866 61174
rect 312102 60938 312134 61174
rect 311514 60854 312134 60938
rect 311514 60618 311546 60854
rect 311782 60618 311866 60854
rect 312102 60618 312134 60854
rect 311514 25174 312134 60618
rect 311514 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 312134 25174
rect 311514 24854 312134 24938
rect 311514 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 312134 24854
rect 311514 -3226 312134 24618
rect 311514 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 312134 -3226
rect 311514 -3546 312134 -3462
rect 311514 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 312134 -3546
rect 311514 -3814 312134 -3782
rect 315234 352894 315854 375600
rect 315234 352658 315266 352894
rect 315502 352658 315586 352894
rect 315822 352658 315854 352894
rect 315234 352574 315854 352658
rect 315234 352338 315266 352574
rect 315502 352338 315586 352574
rect 315822 352338 315854 352574
rect 315234 316894 315854 352338
rect 315234 316658 315266 316894
rect 315502 316658 315586 316894
rect 315822 316658 315854 316894
rect 315234 316574 315854 316658
rect 315234 316338 315266 316574
rect 315502 316338 315586 316574
rect 315822 316338 315854 316574
rect 315234 280894 315854 316338
rect 315234 280658 315266 280894
rect 315502 280658 315586 280894
rect 315822 280658 315854 280894
rect 315234 280574 315854 280658
rect 315234 280338 315266 280574
rect 315502 280338 315586 280574
rect 315822 280338 315854 280574
rect 315234 244894 315854 280338
rect 315234 244658 315266 244894
rect 315502 244658 315586 244894
rect 315822 244658 315854 244894
rect 315234 244574 315854 244658
rect 315234 244338 315266 244574
rect 315502 244338 315586 244574
rect 315822 244338 315854 244574
rect 315234 208894 315854 244338
rect 315234 208658 315266 208894
rect 315502 208658 315586 208894
rect 315822 208658 315854 208894
rect 315234 208574 315854 208658
rect 315234 208338 315266 208574
rect 315502 208338 315586 208574
rect 315822 208338 315854 208574
rect 315234 172894 315854 208338
rect 315234 172658 315266 172894
rect 315502 172658 315586 172894
rect 315822 172658 315854 172894
rect 315234 172574 315854 172658
rect 315234 172338 315266 172574
rect 315502 172338 315586 172574
rect 315822 172338 315854 172574
rect 315234 136894 315854 172338
rect 315234 136658 315266 136894
rect 315502 136658 315586 136894
rect 315822 136658 315854 136894
rect 315234 136574 315854 136658
rect 315234 136338 315266 136574
rect 315502 136338 315586 136574
rect 315822 136338 315854 136574
rect 315234 100894 315854 136338
rect 315234 100658 315266 100894
rect 315502 100658 315586 100894
rect 315822 100658 315854 100894
rect 315234 100574 315854 100658
rect 315234 100338 315266 100574
rect 315502 100338 315586 100574
rect 315822 100338 315854 100574
rect 315234 64894 315854 100338
rect 315234 64658 315266 64894
rect 315502 64658 315586 64894
rect 315822 64658 315854 64894
rect 315234 64574 315854 64658
rect 315234 64338 315266 64574
rect 315502 64338 315586 64574
rect 315822 64338 315854 64574
rect 315234 28894 315854 64338
rect 315234 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 315854 28894
rect 315234 28574 315854 28658
rect 315234 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 315854 28574
rect 315234 -5146 315854 28338
rect 315234 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 315854 -5146
rect 315234 -5466 315854 -5382
rect 315234 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 315854 -5466
rect 315234 -5734 315854 -5702
rect 318954 356614 319574 375600
rect 318954 356378 318986 356614
rect 319222 356378 319306 356614
rect 319542 356378 319574 356614
rect 318954 356294 319574 356378
rect 318954 356058 318986 356294
rect 319222 356058 319306 356294
rect 319542 356058 319574 356294
rect 318954 320614 319574 356058
rect 318954 320378 318986 320614
rect 319222 320378 319306 320614
rect 319542 320378 319574 320614
rect 318954 320294 319574 320378
rect 318954 320058 318986 320294
rect 319222 320058 319306 320294
rect 319542 320058 319574 320294
rect 318954 284614 319574 320058
rect 318954 284378 318986 284614
rect 319222 284378 319306 284614
rect 319542 284378 319574 284614
rect 318954 284294 319574 284378
rect 318954 284058 318986 284294
rect 319222 284058 319306 284294
rect 319542 284058 319574 284294
rect 318954 248614 319574 284058
rect 318954 248378 318986 248614
rect 319222 248378 319306 248614
rect 319542 248378 319574 248614
rect 318954 248294 319574 248378
rect 318954 248058 318986 248294
rect 319222 248058 319306 248294
rect 319542 248058 319574 248294
rect 318954 212614 319574 248058
rect 318954 212378 318986 212614
rect 319222 212378 319306 212614
rect 319542 212378 319574 212614
rect 318954 212294 319574 212378
rect 318954 212058 318986 212294
rect 319222 212058 319306 212294
rect 319542 212058 319574 212294
rect 318954 176614 319574 212058
rect 318954 176378 318986 176614
rect 319222 176378 319306 176614
rect 319542 176378 319574 176614
rect 318954 176294 319574 176378
rect 318954 176058 318986 176294
rect 319222 176058 319306 176294
rect 319542 176058 319574 176294
rect 318954 140614 319574 176058
rect 318954 140378 318986 140614
rect 319222 140378 319306 140614
rect 319542 140378 319574 140614
rect 318954 140294 319574 140378
rect 318954 140058 318986 140294
rect 319222 140058 319306 140294
rect 319542 140058 319574 140294
rect 318954 104614 319574 140058
rect 318954 104378 318986 104614
rect 319222 104378 319306 104614
rect 319542 104378 319574 104614
rect 318954 104294 319574 104378
rect 318954 104058 318986 104294
rect 319222 104058 319306 104294
rect 319542 104058 319574 104294
rect 318954 68614 319574 104058
rect 318954 68378 318986 68614
rect 319222 68378 319306 68614
rect 319542 68378 319574 68614
rect 318954 68294 319574 68378
rect 318954 68058 318986 68294
rect 319222 68058 319306 68294
rect 319542 68058 319574 68294
rect 318954 32614 319574 68058
rect 318954 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 319574 32614
rect 318954 32294 319574 32378
rect 318954 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 319574 32294
rect 300954 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 301574 -6106
rect 300954 -6426 301574 -6342
rect 300954 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 301574 -6426
rect 300954 -7654 301574 -6662
rect 318954 -7066 319574 32058
rect 325794 363454 326414 375600
rect 325794 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 326414 363454
rect 325794 363134 326414 363218
rect 325794 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 326414 363134
rect 325794 327454 326414 362898
rect 325794 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 326414 327454
rect 325794 327134 326414 327218
rect 325794 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 326414 327134
rect 325794 291454 326414 326898
rect 325794 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 326414 291454
rect 325794 291134 326414 291218
rect 325794 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 326414 291134
rect 325794 255454 326414 290898
rect 325794 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 326414 255454
rect 325794 255134 326414 255218
rect 325794 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 326414 255134
rect 325794 219454 326414 254898
rect 325794 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 326414 219454
rect 325794 219134 326414 219218
rect 325794 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 326414 219134
rect 325794 183454 326414 218898
rect 325794 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 326414 183454
rect 325794 183134 326414 183218
rect 325794 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 326414 183134
rect 325794 147454 326414 182898
rect 325794 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 326414 147454
rect 325794 147134 326414 147218
rect 325794 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 326414 147134
rect 325794 111454 326414 146898
rect 325794 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 326414 111454
rect 325794 111134 326414 111218
rect 325794 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 326414 111134
rect 325794 75454 326414 110898
rect 325794 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 326414 75454
rect 325794 75134 326414 75218
rect 325794 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 326414 75134
rect 325794 39454 326414 74898
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -1894 326414 -902
rect 329514 367174 330134 375600
rect 329514 366938 329546 367174
rect 329782 366938 329866 367174
rect 330102 366938 330134 367174
rect 329514 366854 330134 366938
rect 329514 366618 329546 366854
rect 329782 366618 329866 366854
rect 330102 366618 330134 366854
rect 329514 331174 330134 366618
rect 329514 330938 329546 331174
rect 329782 330938 329866 331174
rect 330102 330938 330134 331174
rect 329514 330854 330134 330938
rect 329514 330618 329546 330854
rect 329782 330618 329866 330854
rect 330102 330618 330134 330854
rect 329514 295174 330134 330618
rect 329514 294938 329546 295174
rect 329782 294938 329866 295174
rect 330102 294938 330134 295174
rect 329514 294854 330134 294938
rect 329514 294618 329546 294854
rect 329782 294618 329866 294854
rect 330102 294618 330134 294854
rect 329514 259174 330134 294618
rect 329514 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 330134 259174
rect 329514 258854 330134 258938
rect 329514 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 330134 258854
rect 329514 223174 330134 258618
rect 329514 222938 329546 223174
rect 329782 222938 329866 223174
rect 330102 222938 330134 223174
rect 329514 222854 330134 222938
rect 329514 222618 329546 222854
rect 329782 222618 329866 222854
rect 330102 222618 330134 222854
rect 329514 187174 330134 222618
rect 329514 186938 329546 187174
rect 329782 186938 329866 187174
rect 330102 186938 330134 187174
rect 329514 186854 330134 186938
rect 329514 186618 329546 186854
rect 329782 186618 329866 186854
rect 330102 186618 330134 186854
rect 329514 151174 330134 186618
rect 329514 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 330134 151174
rect 329514 150854 330134 150938
rect 329514 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 330134 150854
rect 329514 115174 330134 150618
rect 329514 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 330134 115174
rect 329514 114854 330134 114938
rect 329514 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 330134 114854
rect 329514 79174 330134 114618
rect 329514 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 330134 79174
rect 329514 78854 330134 78938
rect 329514 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 330134 78854
rect 329514 43174 330134 78618
rect 329514 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 330134 43174
rect 329514 42854 330134 42938
rect 329514 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 330134 42854
rect 329514 7174 330134 42618
rect 329514 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 330134 7174
rect 329514 6854 330134 6938
rect 329514 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 330134 6854
rect 329514 -2266 330134 6618
rect 329514 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 330134 -2266
rect 329514 -2586 330134 -2502
rect 329514 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 330134 -2586
rect 329514 -3814 330134 -2822
rect 333234 370894 333854 375600
rect 333234 370658 333266 370894
rect 333502 370658 333586 370894
rect 333822 370658 333854 370894
rect 333234 370574 333854 370658
rect 333234 370338 333266 370574
rect 333502 370338 333586 370574
rect 333822 370338 333854 370574
rect 333234 334894 333854 370338
rect 333234 334658 333266 334894
rect 333502 334658 333586 334894
rect 333822 334658 333854 334894
rect 333234 334574 333854 334658
rect 333234 334338 333266 334574
rect 333502 334338 333586 334574
rect 333822 334338 333854 334574
rect 333234 298894 333854 334338
rect 333234 298658 333266 298894
rect 333502 298658 333586 298894
rect 333822 298658 333854 298894
rect 333234 298574 333854 298658
rect 333234 298338 333266 298574
rect 333502 298338 333586 298574
rect 333822 298338 333854 298574
rect 333234 262894 333854 298338
rect 333234 262658 333266 262894
rect 333502 262658 333586 262894
rect 333822 262658 333854 262894
rect 333234 262574 333854 262658
rect 333234 262338 333266 262574
rect 333502 262338 333586 262574
rect 333822 262338 333854 262574
rect 333234 226894 333854 262338
rect 333234 226658 333266 226894
rect 333502 226658 333586 226894
rect 333822 226658 333854 226894
rect 333234 226574 333854 226658
rect 333234 226338 333266 226574
rect 333502 226338 333586 226574
rect 333822 226338 333854 226574
rect 333234 190894 333854 226338
rect 333234 190658 333266 190894
rect 333502 190658 333586 190894
rect 333822 190658 333854 190894
rect 333234 190574 333854 190658
rect 333234 190338 333266 190574
rect 333502 190338 333586 190574
rect 333822 190338 333854 190574
rect 333234 154894 333854 190338
rect 333234 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 333854 154894
rect 333234 154574 333854 154658
rect 333234 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 333854 154574
rect 333234 118894 333854 154338
rect 333234 118658 333266 118894
rect 333502 118658 333586 118894
rect 333822 118658 333854 118894
rect 333234 118574 333854 118658
rect 333234 118338 333266 118574
rect 333502 118338 333586 118574
rect 333822 118338 333854 118574
rect 333234 82894 333854 118338
rect 333234 82658 333266 82894
rect 333502 82658 333586 82894
rect 333822 82658 333854 82894
rect 333234 82574 333854 82658
rect 333234 82338 333266 82574
rect 333502 82338 333586 82574
rect 333822 82338 333854 82574
rect 333234 46894 333854 82338
rect 333234 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 333854 46894
rect 333234 46574 333854 46658
rect 333234 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 333854 46574
rect 333234 10894 333854 46338
rect 333234 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 333854 10894
rect 333234 10574 333854 10658
rect 333234 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 333854 10574
rect 333234 -4186 333854 10338
rect 333234 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 333854 -4186
rect 333234 -4506 333854 -4422
rect 333234 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 333854 -4506
rect 333234 -5734 333854 -4742
rect 336954 374614 337574 375600
rect 336954 374378 336986 374614
rect 337222 374378 337306 374614
rect 337542 374378 337574 374614
rect 336954 374294 337574 374378
rect 336954 374058 336986 374294
rect 337222 374058 337306 374294
rect 337542 374058 337574 374294
rect 336954 338614 337574 374058
rect 336954 338378 336986 338614
rect 337222 338378 337306 338614
rect 337542 338378 337574 338614
rect 336954 338294 337574 338378
rect 336954 338058 336986 338294
rect 337222 338058 337306 338294
rect 337542 338058 337574 338294
rect 336954 302614 337574 338058
rect 336954 302378 336986 302614
rect 337222 302378 337306 302614
rect 337542 302378 337574 302614
rect 336954 302294 337574 302378
rect 336954 302058 336986 302294
rect 337222 302058 337306 302294
rect 337542 302058 337574 302294
rect 336954 266614 337574 302058
rect 336954 266378 336986 266614
rect 337222 266378 337306 266614
rect 337542 266378 337574 266614
rect 336954 266294 337574 266378
rect 336954 266058 336986 266294
rect 337222 266058 337306 266294
rect 337542 266058 337574 266294
rect 336954 230614 337574 266058
rect 336954 230378 336986 230614
rect 337222 230378 337306 230614
rect 337542 230378 337574 230614
rect 336954 230294 337574 230378
rect 336954 230058 336986 230294
rect 337222 230058 337306 230294
rect 337542 230058 337574 230294
rect 336954 194614 337574 230058
rect 336954 194378 336986 194614
rect 337222 194378 337306 194614
rect 337542 194378 337574 194614
rect 336954 194294 337574 194378
rect 336954 194058 336986 194294
rect 337222 194058 337306 194294
rect 337542 194058 337574 194294
rect 336954 158614 337574 194058
rect 336954 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 337574 158614
rect 336954 158294 337574 158378
rect 336954 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 337574 158294
rect 336954 122614 337574 158058
rect 336954 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 337574 122614
rect 336954 122294 337574 122378
rect 336954 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 337574 122294
rect 336954 86614 337574 122058
rect 336954 86378 336986 86614
rect 337222 86378 337306 86614
rect 337542 86378 337574 86614
rect 336954 86294 337574 86378
rect 336954 86058 336986 86294
rect 337222 86058 337306 86294
rect 337542 86058 337574 86294
rect 336954 50614 337574 86058
rect 336954 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 337574 50614
rect 336954 50294 337574 50378
rect 336954 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 337574 50294
rect 336954 14614 337574 50058
rect 336954 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 337574 14614
rect 336954 14294 337574 14378
rect 336954 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 337574 14294
rect 318954 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 319574 -7066
rect 318954 -7386 319574 -7302
rect 318954 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 319574 -7386
rect 318954 -7654 319574 -7622
rect 336954 -6106 337574 14058
rect 343794 345454 344414 375600
rect 343794 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 344414 345454
rect 343794 345134 344414 345218
rect 343794 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 344414 345134
rect 343794 309454 344414 344898
rect 343794 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 344414 309454
rect 343794 309134 344414 309218
rect 343794 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 344414 309134
rect 343794 273454 344414 308898
rect 343794 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 344414 273454
rect 343794 273134 344414 273218
rect 343794 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 344414 273134
rect 343794 237454 344414 272898
rect 343794 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 344414 237454
rect 343794 237134 344414 237218
rect 343794 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 344414 237134
rect 343794 201454 344414 236898
rect 343794 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 344414 201454
rect 343794 201134 344414 201218
rect 343794 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 344414 201134
rect 343794 165454 344414 200898
rect 343794 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 344414 165454
rect 343794 165134 344414 165218
rect 343794 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 344414 165134
rect 343794 129454 344414 164898
rect 343794 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 344414 129454
rect 343794 129134 344414 129218
rect 343794 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 344414 129134
rect 343794 93454 344414 128898
rect 343794 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 344414 93454
rect 343794 93134 344414 93218
rect 343794 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 344414 93134
rect 343794 57454 344414 92898
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -1306 344414 20898
rect 343794 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 344414 -1306
rect 343794 -1626 344414 -1542
rect 343794 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 344414 -1626
rect 343794 -1894 344414 -1862
rect 347514 349174 348134 375600
rect 347514 348938 347546 349174
rect 347782 348938 347866 349174
rect 348102 348938 348134 349174
rect 347514 348854 348134 348938
rect 347514 348618 347546 348854
rect 347782 348618 347866 348854
rect 348102 348618 348134 348854
rect 347514 313174 348134 348618
rect 347514 312938 347546 313174
rect 347782 312938 347866 313174
rect 348102 312938 348134 313174
rect 347514 312854 348134 312938
rect 347514 312618 347546 312854
rect 347782 312618 347866 312854
rect 348102 312618 348134 312854
rect 347514 277174 348134 312618
rect 347514 276938 347546 277174
rect 347782 276938 347866 277174
rect 348102 276938 348134 277174
rect 347514 276854 348134 276938
rect 347514 276618 347546 276854
rect 347782 276618 347866 276854
rect 348102 276618 348134 276854
rect 347514 241174 348134 276618
rect 347514 240938 347546 241174
rect 347782 240938 347866 241174
rect 348102 240938 348134 241174
rect 347514 240854 348134 240938
rect 347514 240618 347546 240854
rect 347782 240618 347866 240854
rect 348102 240618 348134 240854
rect 347514 205174 348134 240618
rect 347514 204938 347546 205174
rect 347782 204938 347866 205174
rect 348102 204938 348134 205174
rect 347514 204854 348134 204938
rect 347514 204618 347546 204854
rect 347782 204618 347866 204854
rect 348102 204618 348134 204854
rect 347514 169174 348134 204618
rect 347514 168938 347546 169174
rect 347782 168938 347866 169174
rect 348102 168938 348134 169174
rect 347514 168854 348134 168938
rect 347514 168618 347546 168854
rect 347782 168618 347866 168854
rect 348102 168618 348134 168854
rect 347514 133174 348134 168618
rect 347514 132938 347546 133174
rect 347782 132938 347866 133174
rect 348102 132938 348134 133174
rect 347514 132854 348134 132938
rect 347514 132618 347546 132854
rect 347782 132618 347866 132854
rect 348102 132618 348134 132854
rect 347514 97174 348134 132618
rect 347514 96938 347546 97174
rect 347782 96938 347866 97174
rect 348102 96938 348134 97174
rect 347514 96854 348134 96938
rect 347514 96618 347546 96854
rect 347782 96618 347866 96854
rect 348102 96618 348134 96854
rect 347514 61174 348134 96618
rect 347514 60938 347546 61174
rect 347782 60938 347866 61174
rect 348102 60938 348134 61174
rect 347514 60854 348134 60938
rect 347514 60618 347546 60854
rect 347782 60618 347866 60854
rect 348102 60618 348134 60854
rect 347514 25174 348134 60618
rect 347514 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 348134 25174
rect 347514 24854 348134 24938
rect 347514 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 348134 24854
rect 347514 -3226 348134 24618
rect 347514 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 348134 -3226
rect 347514 -3546 348134 -3462
rect 347514 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 348134 -3546
rect 347514 -3814 348134 -3782
rect 351234 352894 351854 375600
rect 352054 355469 352114 538187
rect 353342 376005 353402 545123
rect 354954 537993 355574 572058
rect 361794 704838 362414 705830
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 361794 543454 362414 578898
rect 361794 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 362414 543454
rect 361794 543134 362414 543218
rect 361794 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 362414 543134
rect 357571 537164 357637 537165
rect 357571 537100 357572 537164
rect 357636 537100 357637 537164
rect 357571 537099 357637 537100
rect 356283 507108 356349 507109
rect 356283 507044 356284 507108
rect 356348 507044 356349 507108
rect 356283 507043 356349 507044
rect 356099 389332 356165 389333
rect 356099 389330 356100 389332
rect 354446 389270 356100 389330
rect 354446 389190 354506 389270
rect 356099 389268 356100 389270
rect 356164 389268 356165 389332
rect 356099 389267 356165 389268
rect 354446 389130 354690 389190
rect 354630 379530 354690 389130
rect 356099 386612 356165 386613
rect 356099 386610 356100 386612
rect 354446 379470 354690 379530
rect 354814 386550 356100 386610
rect 353339 376004 353405 376005
rect 353339 375940 353340 376004
rect 353404 375940 353405 376004
rect 353339 375939 353405 375940
rect 354446 375325 354506 379470
rect 354814 376413 354874 386550
rect 356099 386548 356100 386550
rect 356164 386548 356165 386612
rect 356099 386547 356165 386548
rect 356286 384029 356346 507043
rect 356467 394500 356533 394501
rect 356467 394436 356468 394500
rect 356532 394436 356533 394500
rect 356467 394435 356533 394436
rect 356283 384028 356349 384029
rect 356283 383964 356284 384028
rect 356348 383964 356349 384028
rect 356283 383963 356349 383964
rect 356283 383756 356349 383757
rect 356283 383692 356284 383756
rect 356348 383692 356349 383756
rect 356283 383691 356349 383692
rect 356099 381580 356165 381581
rect 356099 381516 356100 381580
rect 356164 381516 356165 381580
rect 356099 381515 356165 381516
rect 354811 376412 354877 376413
rect 354811 376348 354812 376412
rect 354876 376348 354877 376412
rect 354811 376347 354877 376348
rect 354443 375324 354509 375325
rect 354443 375260 354444 375324
rect 354508 375260 354509 375324
rect 354443 375259 354509 375260
rect 354954 356614 355574 375600
rect 356102 371381 356162 381515
rect 356099 371380 356165 371381
rect 356099 371316 356100 371380
rect 356164 371316 356165 371380
rect 356099 371315 356165 371316
rect 354954 356378 354986 356614
rect 355222 356378 355306 356614
rect 355542 356378 355574 356614
rect 354954 356294 355574 356378
rect 354954 356058 354986 356294
rect 355222 356058 355306 356294
rect 355542 356058 355574 356294
rect 352051 355468 352117 355469
rect 352051 355404 352052 355468
rect 352116 355404 352117 355468
rect 352051 355403 352117 355404
rect 351234 352658 351266 352894
rect 351502 352658 351586 352894
rect 351822 352658 351854 352894
rect 351234 352574 351854 352658
rect 351234 352338 351266 352574
rect 351502 352338 351586 352574
rect 351822 352338 351854 352574
rect 351234 316894 351854 352338
rect 351234 316658 351266 316894
rect 351502 316658 351586 316894
rect 351822 316658 351854 316894
rect 351234 316574 351854 316658
rect 351234 316338 351266 316574
rect 351502 316338 351586 316574
rect 351822 316338 351854 316574
rect 351234 280894 351854 316338
rect 351234 280658 351266 280894
rect 351502 280658 351586 280894
rect 351822 280658 351854 280894
rect 351234 280574 351854 280658
rect 351234 280338 351266 280574
rect 351502 280338 351586 280574
rect 351822 280338 351854 280574
rect 351234 244894 351854 280338
rect 351234 244658 351266 244894
rect 351502 244658 351586 244894
rect 351822 244658 351854 244894
rect 351234 244574 351854 244658
rect 351234 244338 351266 244574
rect 351502 244338 351586 244574
rect 351822 244338 351854 244574
rect 351234 208894 351854 244338
rect 351234 208658 351266 208894
rect 351502 208658 351586 208894
rect 351822 208658 351854 208894
rect 351234 208574 351854 208658
rect 351234 208338 351266 208574
rect 351502 208338 351586 208574
rect 351822 208338 351854 208574
rect 351234 172894 351854 208338
rect 351234 172658 351266 172894
rect 351502 172658 351586 172894
rect 351822 172658 351854 172894
rect 351234 172574 351854 172658
rect 351234 172338 351266 172574
rect 351502 172338 351586 172574
rect 351822 172338 351854 172574
rect 351234 136894 351854 172338
rect 351234 136658 351266 136894
rect 351502 136658 351586 136894
rect 351822 136658 351854 136894
rect 351234 136574 351854 136658
rect 351234 136338 351266 136574
rect 351502 136338 351586 136574
rect 351822 136338 351854 136574
rect 351234 100894 351854 136338
rect 351234 100658 351266 100894
rect 351502 100658 351586 100894
rect 351822 100658 351854 100894
rect 351234 100574 351854 100658
rect 351234 100338 351266 100574
rect 351502 100338 351586 100574
rect 351822 100338 351854 100574
rect 351234 64894 351854 100338
rect 351234 64658 351266 64894
rect 351502 64658 351586 64894
rect 351822 64658 351854 64894
rect 351234 64574 351854 64658
rect 351234 64338 351266 64574
rect 351502 64338 351586 64574
rect 351822 64338 351854 64574
rect 351234 28894 351854 64338
rect 351234 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 351854 28894
rect 351234 28574 351854 28658
rect 351234 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 351854 28574
rect 351234 -5146 351854 28338
rect 351234 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 351854 -5146
rect 351234 -5466 351854 -5382
rect 351234 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 351854 -5466
rect 351234 -5734 351854 -5702
rect 354954 320614 355574 356058
rect 354954 320378 354986 320614
rect 355222 320378 355306 320614
rect 355542 320378 355574 320614
rect 354954 320294 355574 320378
rect 354954 320058 354986 320294
rect 355222 320058 355306 320294
rect 355542 320058 355574 320294
rect 354954 284614 355574 320058
rect 354954 284378 354986 284614
rect 355222 284378 355306 284614
rect 355542 284378 355574 284614
rect 354954 284294 355574 284378
rect 354954 284058 354986 284294
rect 355222 284058 355306 284294
rect 355542 284058 355574 284294
rect 354954 248614 355574 284058
rect 354954 248378 354986 248614
rect 355222 248378 355306 248614
rect 355542 248378 355574 248614
rect 354954 248294 355574 248378
rect 354954 248058 354986 248294
rect 355222 248058 355306 248294
rect 355542 248058 355574 248294
rect 354954 212614 355574 248058
rect 354954 212378 354986 212614
rect 355222 212378 355306 212614
rect 355542 212378 355574 212614
rect 354954 212294 355574 212378
rect 354954 212058 354986 212294
rect 355222 212058 355306 212294
rect 355542 212058 355574 212294
rect 354954 176614 355574 212058
rect 354954 176378 354986 176614
rect 355222 176378 355306 176614
rect 355542 176378 355574 176614
rect 354954 176294 355574 176378
rect 354954 176058 354986 176294
rect 355222 176058 355306 176294
rect 355542 176058 355574 176294
rect 354954 140614 355574 176058
rect 354954 140378 354986 140614
rect 355222 140378 355306 140614
rect 355542 140378 355574 140614
rect 354954 140294 355574 140378
rect 354954 140058 354986 140294
rect 355222 140058 355306 140294
rect 355542 140058 355574 140294
rect 354954 104614 355574 140058
rect 354954 104378 354986 104614
rect 355222 104378 355306 104614
rect 355542 104378 355574 104614
rect 354954 104294 355574 104378
rect 354954 104058 354986 104294
rect 355222 104058 355306 104294
rect 355542 104058 355574 104294
rect 354954 68614 355574 104058
rect 354954 68378 354986 68614
rect 355222 68378 355306 68614
rect 355542 68378 355574 68614
rect 354954 68294 355574 68378
rect 354954 68058 354986 68294
rect 355222 68058 355306 68294
rect 355542 68058 355574 68294
rect 354954 32614 355574 68058
rect 354954 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 355574 32614
rect 354954 32294 355574 32378
rect 354954 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 355574 32294
rect 336954 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 337574 -6106
rect 336954 -6426 337574 -6342
rect 336954 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 337574 -6426
rect 336954 -7654 337574 -6662
rect 354954 -7066 355574 32058
rect 356102 4861 356162 371315
rect 356286 359413 356346 383691
rect 356470 381581 356530 394435
rect 356467 381580 356533 381581
rect 356467 381516 356468 381580
rect 356532 381516 356533 381580
rect 356467 381515 356533 381516
rect 357574 379530 357634 537099
rect 361794 507454 362414 542898
rect 365514 691174 366134 706202
rect 365514 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 366134 691174
rect 365514 690854 366134 690938
rect 365514 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 366134 690854
rect 365514 655174 366134 690618
rect 365514 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 366134 655174
rect 365514 654854 366134 654938
rect 365514 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 366134 654854
rect 365514 619174 366134 654618
rect 365514 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 366134 619174
rect 365514 618854 366134 618938
rect 365514 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 366134 618854
rect 365514 583174 366134 618618
rect 365514 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 366134 583174
rect 365514 582854 366134 582938
rect 365514 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 366134 582854
rect 365514 547174 366134 582618
rect 365514 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 366134 547174
rect 365514 546854 366134 546938
rect 365514 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 366134 546854
rect 362907 539748 362973 539749
rect 362907 539684 362908 539748
rect 362972 539684 362973 539748
rect 362907 539683 362973 539684
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 360147 480452 360213 480453
rect 360147 480388 360148 480452
rect 360212 480388 360213 480452
rect 360147 480387 360213 480388
rect 358859 458420 358925 458421
rect 358859 458356 358860 458420
rect 358924 458356 358925 458420
rect 358859 458355 358925 458356
rect 357390 379470 357634 379530
rect 356283 359412 356349 359413
rect 356283 359348 356284 359412
rect 356348 359348 356349 359412
rect 356283 359347 356349 359348
rect 357390 354690 357450 379470
rect 357571 378044 357637 378045
rect 357571 377980 357572 378044
rect 357636 377980 357637 378044
rect 357571 377979 357637 377980
rect 357574 362269 357634 377979
rect 357571 362268 357637 362269
rect 357571 362204 357572 362268
rect 357636 362204 357637 362268
rect 357571 362203 357637 362204
rect 358862 356693 358922 458355
rect 360150 389190 360210 480387
rect 359966 389130 360210 389190
rect 361794 471454 362414 506898
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 361794 435454 362414 470898
rect 361794 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 362414 435454
rect 361794 435134 362414 435218
rect 361794 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 362414 435134
rect 361794 399454 362414 434898
rect 361794 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 362414 399454
rect 361794 399134 362414 399218
rect 361794 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 362414 399134
rect 359966 379530 360026 389130
rect 359966 379470 360210 379530
rect 358859 356692 358925 356693
rect 358859 356628 358860 356692
rect 358924 356628 358925 356692
rect 358859 356627 358925 356628
rect 357390 354630 357634 354690
rect 357574 296717 357634 354630
rect 360150 344317 360210 379470
rect 361794 363454 362414 398898
rect 361794 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 362414 363454
rect 361794 363134 362414 363218
rect 361794 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 362414 363134
rect 360147 344316 360213 344317
rect 360147 344252 360148 344316
rect 360212 344252 360213 344316
rect 360147 344251 360213 344252
rect 361794 327454 362414 362898
rect 361794 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 362414 327454
rect 361794 327134 362414 327218
rect 361794 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 362414 327134
rect 357571 296716 357637 296717
rect 357571 296652 357572 296716
rect 357636 296652 357637 296716
rect 357571 296651 357637 296652
rect 357574 296037 357634 296651
rect 357571 296036 357637 296037
rect 357571 295972 357572 296036
rect 357636 295972 357637 296036
rect 357571 295971 357637 295972
rect 361794 291454 362414 326898
rect 361794 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 362414 291454
rect 361794 291134 362414 291218
rect 361794 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 362414 291134
rect 361794 255454 362414 290898
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 361794 219454 362414 254898
rect 361794 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 362414 219454
rect 361794 219134 362414 219218
rect 361794 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 362414 219134
rect 361794 183454 362414 218898
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 361794 147454 362414 182898
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 361794 39454 362414 74898
rect 362910 67557 362970 539683
rect 365514 511174 366134 546618
rect 365514 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 366134 511174
rect 365514 510854 366134 510938
rect 365514 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 366134 510854
rect 365514 475174 366134 510618
rect 365514 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 366134 475174
rect 365514 474854 366134 474938
rect 365514 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 366134 474854
rect 365514 439174 366134 474618
rect 365514 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 366134 439174
rect 365514 438854 366134 438938
rect 365514 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 366134 438854
rect 365514 403174 366134 438618
rect 365514 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 366134 403174
rect 365514 402854 366134 402938
rect 365514 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 366134 402854
rect 363091 384708 363157 384709
rect 363091 384644 363092 384708
rect 363156 384644 363157 384708
rect 363091 384643 363157 384644
rect 362907 67556 362973 67557
rect 362907 67492 362908 67556
rect 362972 67492 362973 67556
rect 362907 67491 362973 67492
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 356099 4860 356165 4861
rect 356099 4796 356100 4860
rect 356164 4796 356165 4860
rect 356099 4795 356165 4796
rect 361794 3454 362414 38898
rect 363094 10301 363154 384643
rect 365514 367174 366134 402618
rect 365514 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 366134 367174
rect 365514 366854 366134 366938
rect 365514 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 366134 366854
rect 365514 331174 366134 366618
rect 365514 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 366134 331174
rect 365514 330854 366134 330938
rect 365514 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 366134 330854
rect 365514 295174 366134 330618
rect 365514 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 366134 295174
rect 365514 294854 366134 294938
rect 365514 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 366134 294854
rect 365514 259174 366134 294618
rect 365514 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 366134 259174
rect 365514 258854 366134 258938
rect 365514 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 366134 258854
rect 365514 223174 366134 258618
rect 365514 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 366134 223174
rect 365514 222854 366134 222938
rect 365514 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 366134 222854
rect 365514 187174 366134 222618
rect 365514 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 366134 187174
rect 365514 186854 366134 186938
rect 365514 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 366134 186854
rect 365514 151174 366134 186618
rect 365514 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 366134 151174
rect 365514 150854 366134 150938
rect 365514 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 366134 150854
rect 365514 115174 366134 150618
rect 365514 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 366134 115174
rect 365514 114854 366134 114938
rect 365514 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 366134 114854
rect 365514 79174 366134 114618
rect 365514 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 366134 79174
rect 365514 78854 366134 78938
rect 365514 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 366134 78854
rect 365514 43174 366134 78618
rect 365514 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 366134 43174
rect 365514 42854 366134 42938
rect 365514 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 366134 42854
rect 363091 10300 363157 10301
rect 363091 10236 363092 10300
rect 363156 10236 363157 10300
rect 363091 10235 363157 10236
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -1894 362414 -902
rect 365514 7174 366134 42618
rect 365514 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 366134 7174
rect 365514 6854 366134 6938
rect 365514 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 366134 6854
rect 365514 -2266 366134 6618
rect 365514 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 366134 -2266
rect 365514 -2586 366134 -2502
rect 365514 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 366134 -2586
rect 365514 -3814 366134 -2822
rect 369234 694894 369854 708122
rect 369234 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 369854 694894
rect 369234 694574 369854 694658
rect 369234 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 369854 694574
rect 369234 658894 369854 694338
rect 369234 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 369854 658894
rect 369234 658574 369854 658658
rect 369234 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 369854 658574
rect 369234 622894 369854 658338
rect 369234 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 369854 622894
rect 369234 622574 369854 622658
rect 369234 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 369854 622574
rect 369234 586894 369854 622338
rect 369234 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 369854 586894
rect 369234 586574 369854 586658
rect 369234 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 369854 586574
rect 369234 550894 369854 586338
rect 369234 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 369854 550894
rect 369234 550574 369854 550658
rect 369234 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 369854 550574
rect 369234 514894 369854 550338
rect 369234 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 369854 514894
rect 369234 514574 369854 514658
rect 369234 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 369854 514574
rect 369234 478894 369854 514338
rect 369234 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 369854 478894
rect 369234 478574 369854 478658
rect 369234 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 369854 478574
rect 369234 442894 369854 478338
rect 369234 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 369854 442894
rect 369234 442574 369854 442658
rect 369234 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 369854 442574
rect 369234 406894 369854 442338
rect 369234 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 369854 406894
rect 369234 406574 369854 406658
rect 369234 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 369854 406574
rect 369234 370894 369854 406338
rect 369234 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 369854 370894
rect 369234 370574 369854 370658
rect 369234 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 369854 370574
rect 369234 334894 369854 370338
rect 369234 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 369854 334894
rect 369234 334574 369854 334658
rect 369234 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 369854 334574
rect 369234 298894 369854 334338
rect 369234 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 369854 298894
rect 369234 298574 369854 298658
rect 369234 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 369854 298574
rect 369234 262894 369854 298338
rect 369234 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 369854 262894
rect 369234 262574 369854 262658
rect 369234 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 369854 262574
rect 369234 226894 369854 262338
rect 369234 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 369854 226894
rect 369234 226574 369854 226658
rect 369234 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 369854 226574
rect 369234 190894 369854 226338
rect 369234 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 369854 190894
rect 369234 190574 369854 190658
rect 369234 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 369854 190574
rect 369234 154894 369854 190338
rect 369234 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 369854 154894
rect 369234 154574 369854 154658
rect 369234 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 369854 154574
rect 369234 118894 369854 154338
rect 369234 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 369854 118894
rect 369234 118574 369854 118658
rect 369234 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 369854 118574
rect 369234 82894 369854 118338
rect 369234 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 369854 82894
rect 369234 82574 369854 82658
rect 369234 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 369854 82574
rect 369234 46894 369854 82338
rect 369234 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 369854 46894
rect 369234 46574 369854 46658
rect 369234 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 369854 46574
rect 369234 10894 369854 46338
rect 369234 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 369854 10894
rect 369234 10574 369854 10658
rect 369234 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 369854 10574
rect 369234 -4186 369854 10338
rect 369234 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 369854 -4186
rect 369234 -4506 369854 -4422
rect 369234 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 369854 -4506
rect 369234 -5734 369854 -4742
rect 372954 698614 373574 710042
rect 390954 711558 391574 711590
rect 390954 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 391574 711558
rect 390954 711238 391574 711322
rect 390954 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 391574 711238
rect 387234 709638 387854 709670
rect 387234 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 387854 709638
rect 387234 709318 387854 709402
rect 387234 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 387854 709318
rect 383514 707718 384134 707750
rect 383514 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 384134 707718
rect 383514 707398 384134 707482
rect 383514 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 384134 707398
rect 372954 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 373574 698614
rect 372954 698294 373574 698378
rect 372954 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 373574 698294
rect 372954 662614 373574 698058
rect 372954 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 373574 662614
rect 372954 662294 373574 662378
rect 372954 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 373574 662294
rect 372954 626614 373574 662058
rect 372954 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 373574 626614
rect 372954 626294 373574 626378
rect 372954 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 373574 626294
rect 372954 590614 373574 626058
rect 372954 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 373574 590614
rect 372954 590294 373574 590378
rect 372954 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 373574 590294
rect 372954 554614 373574 590058
rect 372954 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 373574 554614
rect 372954 554294 373574 554378
rect 372954 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 373574 554294
rect 372954 518614 373574 554058
rect 372954 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 373574 518614
rect 372954 518294 373574 518378
rect 372954 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 373574 518294
rect 372954 482614 373574 518058
rect 372954 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 373574 482614
rect 372954 482294 373574 482378
rect 372954 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 373574 482294
rect 372954 446614 373574 482058
rect 372954 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 373574 446614
rect 372954 446294 373574 446378
rect 372954 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 373574 446294
rect 372954 410614 373574 446058
rect 372954 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 373574 410614
rect 372954 410294 373574 410378
rect 372954 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 373574 410294
rect 372954 374614 373574 410058
rect 372954 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 373574 374614
rect 372954 374294 373574 374378
rect 372954 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 373574 374294
rect 372954 338614 373574 374058
rect 372954 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 373574 338614
rect 372954 338294 373574 338378
rect 372954 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 373574 338294
rect 372954 302614 373574 338058
rect 372954 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 373574 302614
rect 372954 302294 373574 302378
rect 372954 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 373574 302294
rect 372954 266614 373574 302058
rect 372954 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 373574 266614
rect 372954 266294 373574 266378
rect 372954 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 373574 266294
rect 372954 230614 373574 266058
rect 372954 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 373574 230614
rect 372954 230294 373574 230378
rect 372954 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 373574 230294
rect 372954 194614 373574 230058
rect 372954 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 373574 194614
rect 372954 194294 373574 194378
rect 372954 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 373574 194294
rect 372954 158614 373574 194058
rect 372954 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 373574 158614
rect 372954 158294 373574 158378
rect 372954 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 373574 158294
rect 372954 122614 373574 158058
rect 372954 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 373574 122614
rect 372954 122294 373574 122378
rect 372954 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 373574 122294
rect 372954 86614 373574 122058
rect 372954 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 373574 86614
rect 372954 86294 373574 86378
rect 372954 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 373574 86294
rect 372954 50614 373574 86058
rect 372954 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 373574 50614
rect 372954 50294 373574 50378
rect 372954 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 373574 50294
rect 372954 14614 373574 50058
rect 372954 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 373574 14614
rect 372954 14294 373574 14378
rect 372954 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 373574 14294
rect 354954 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 355574 -7066
rect 354954 -7386 355574 -7302
rect 354954 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 355574 -7386
rect 354954 -7654 355574 -7622
rect 372954 -6106 373574 14058
rect 379794 705798 380414 705830
rect 379794 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 380414 705798
rect 379794 705478 380414 705562
rect 379794 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 380414 705478
rect 379794 669454 380414 705242
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 633454 380414 668898
rect 379794 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 380414 633454
rect 379794 633134 380414 633218
rect 379794 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 380414 633134
rect 379794 597454 380414 632898
rect 379794 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 380414 597454
rect 379794 597134 380414 597218
rect 379794 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 380414 597134
rect 379794 561454 380414 596898
rect 379794 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 380414 561454
rect 379794 561134 380414 561218
rect 379794 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 380414 561134
rect 379794 525454 380414 560898
rect 379794 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 380414 525454
rect 379794 525134 380414 525218
rect 379794 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 380414 525134
rect 379794 489454 380414 524898
rect 379794 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 380414 489454
rect 379794 489134 380414 489218
rect 379794 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 380414 489134
rect 379794 453454 380414 488898
rect 379794 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 380414 453454
rect 379794 453134 380414 453218
rect 379794 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 380414 453134
rect 379794 417454 380414 452898
rect 379794 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 380414 417454
rect 379794 417134 380414 417218
rect 379794 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 380414 417134
rect 379794 381454 380414 416898
rect 379794 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 380414 381454
rect 379794 381134 380414 381218
rect 379794 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 380414 381134
rect 379794 345454 380414 380898
rect 379794 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 380414 345454
rect 379794 345134 380414 345218
rect 379794 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 380414 345134
rect 379794 309454 380414 344898
rect 379794 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 380414 309454
rect 379794 309134 380414 309218
rect 379794 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 380414 309134
rect 379794 273454 380414 308898
rect 379794 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 380414 273454
rect 379794 273134 380414 273218
rect 379794 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 380414 273134
rect 379794 237454 380414 272898
rect 379794 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 380414 237454
rect 379794 237134 380414 237218
rect 379794 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 380414 237134
rect 379794 201454 380414 236898
rect 379794 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 380414 201454
rect 379794 201134 380414 201218
rect 379794 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 380414 201134
rect 379794 165454 380414 200898
rect 379794 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 380414 165454
rect 379794 165134 380414 165218
rect 379794 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 380414 165134
rect 379794 129454 380414 164898
rect 379794 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 380414 129454
rect 379794 129134 380414 129218
rect 379794 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 380414 129134
rect 379794 93454 380414 128898
rect 379794 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 380414 93454
rect 379794 93134 380414 93218
rect 379794 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 380414 93134
rect 379794 57454 380414 92898
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -1306 380414 20898
rect 379794 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 380414 -1306
rect 379794 -1626 380414 -1542
rect 379794 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 380414 -1626
rect 379794 -1894 380414 -1862
rect 383514 673174 384134 707162
rect 383514 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 384134 673174
rect 383514 672854 384134 672938
rect 383514 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 384134 672854
rect 383514 637174 384134 672618
rect 383514 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 384134 637174
rect 383514 636854 384134 636938
rect 383514 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 384134 636854
rect 383514 601174 384134 636618
rect 383514 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 384134 601174
rect 383514 600854 384134 600938
rect 383514 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 384134 600854
rect 383514 565174 384134 600618
rect 383514 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 384134 565174
rect 383514 564854 384134 564938
rect 383514 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 384134 564854
rect 383514 529174 384134 564618
rect 383514 528938 383546 529174
rect 383782 528938 383866 529174
rect 384102 528938 384134 529174
rect 383514 528854 384134 528938
rect 383514 528618 383546 528854
rect 383782 528618 383866 528854
rect 384102 528618 384134 528854
rect 383514 493174 384134 528618
rect 383514 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 384134 493174
rect 383514 492854 384134 492938
rect 383514 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 384134 492854
rect 383514 457174 384134 492618
rect 383514 456938 383546 457174
rect 383782 456938 383866 457174
rect 384102 456938 384134 457174
rect 383514 456854 384134 456938
rect 383514 456618 383546 456854
rect 383782 456618 383866 456854
rect 384102 456618 384134 456854
rect 383514 421174 384134 456618
rect 383514 420938 383546 421174
rect 383782 420938 383866 421174
rect 384102 420938 384134 421174
rect 383514 420854 384134 420938
rect 383514 420618 383546 420854
rect 383782 420618 383866 420854
rect 384102 420618 384134 420854
rect 383514 385174 384134 420618
rect 383514 384938 383546 385174
rect 383782 384938 383866 385174
rect 384102 384938 384134 385174
rect 383514 384854 384134 384938
rect 383514 384618 383546 384854
rect 383782 384618 383866 384854
rect 384102 384618 384134 384854
rect 383514 349174 384134 384618
rect 383514 348938 383546 349174
rect 383782 348938 383866 349174
rect 384102 348938 384134 349174
rect 383514 348854 384134 348938
rect 383514 348618 383546 348854
rect 383782 348618 383866 348854
rect 384102 348618 384134 348854
rect 383514 313174 384134 348618
rect 383514 312938 383546 313174
rect 383782 312938 383866 313174
rect 384102 312938 384134 313174
rect 383514 312854 384134 312938
rect 383514 312618 383546 312854
rect 383782 312618 383866 312854
rect 384102 312618 384134 312854
rect 383514 277174 384134 312618
rect 383514 276938 383546 277174
rect 383782 276938 383866 277174
rect 384102 276938 384134 277174
rect 383514 276854 384134 276938
rect 383514 276618 383546 276854
rect 383782 276618 383866 276854
rect 384102 276618 384134 276854
rect 383514 241174 384134 276618
rect 383514 240938 383546 241174
rect 383782 240938 383866 241174
rect 384102 240938 384134 241174
rect 383514 240854 384134 240938
rect 383514 240618 383546 240854
rect 383782 240618 383866 240854
rect 384102 240618 384134 240854
rect 383514 205174 384134 240618
rect 383514 204938 383546 205174
rect 383782 204938 383866 205174
rect 384102 204938 384134 205174
rect 383514 204854 384134 204938
rect 383514 204618 383546 204854
rect 383782 204618 383866 204854
rect 384102 204618 384134 204854
rect 383514 169174 384134 204618
rect 383514 168938 383546 169174
rect 383782 168938 383866 169174
rect 384102 168938 384134 169174
rect 383514 168854 384134 168938
rect 383514 168618 383546 168854
rect 383782 168618 383866 168854
rect 384102 168618 384134 168854
rect 383514 133174 384134 168618
rect 383514 132938 383546 133174
rect 383782 132938 383866 133174
rect 384102 132938 384134 133174
rect 383514 132854 384134 132938
rect 383514 132618 383546 132854
rect 383782 132618 383866 132854
rect 384102 132618 384134 132854
rect 383514 97174 384134 132618
rect 383514 96938 383546 97174
rect 383782 96938 383866 97174
rect 384102 96938 384134 97174
rect 383514 96854 384134 96938
rect 383514 96618 383546 96854
rect 383782 96618 383866 96854
rect 384102 96618 384134 96854
rect 383514 61174 384134 96618
rect 383514 60938 383546 61174
rect 383782 60938 383866 61174
rect 384102 60938 384134 61174
rect 383514 60854 384134 60938
rect 383514 60618 383546 60854
rect 383782 60618 383866 60854
rect 384102 60618 384134 60854
rect 383514 25174 384134 60618
rect 383514 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 384134 25174
rect 383514 24854 384134 24938
rect 383514 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 384134 24854
rect 383514 -3226 384134 24618
rect 383514 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 384134 -3226
rect 383514 -3546 384134 -3462
rect 383514 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 384134 -3546
rect 383514 -3814 384134 -3782
rect 387234 676894 387854 709082
rect 387234 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 387854 676894
rect 387234 676574 387854 676658
rect 387234 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 387854 676574
rect 387234 640894 387854 676338
rect 387234 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 387854 640894
rect 387234 640574 387854 640658
rect 387234 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 387854 640574
rect 387234 604894 387854 640338
rect 387234 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 387854 604894
rect 387234 604574 387854 604658
rect 387234 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 387854 604574
rect 387234 568894 387854 604338
rect 387234 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 387854 568894
rect 387234 568574 387854 568658
rect 387234 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 387854 568574
rect 387234 532894 387854 568338
rect 387234 532658 387266 532894
rect 387502 532658 387586 532894
rect 387822 532658 387854 532894
rect 387234 532574 387854 532658
rect 387234 532338 387266 532574
rect 387502 532338 387586 532574
rect 387822 532338 387854 532574
rect 387234 496894 387854 532338
rect 387234 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 387854 496894
rect 387234 496574 387854 496658
rect 387234 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 387854 496574
rect 387234 460894 387854 496338
rect 387234 460658 387266 460894
rect 387502 460658 387586 460894
rect 387822 460658 387854 460894
rect 387234 460574 387854 460658
rect 387234 460338 387266 460574
rect 387502 460338 387586 460574
rect 387822 460338 387854 460574
rect 387234 424894 387854 460338
rect 387234 424658 387266 424894
rect 387502 424658 387586 424894
rect 387822 424658 387854 424894
rect 387234 424574 387854 424658
rect 387234 424338 387266 424574
rect 387502 424338 387586 424574
rect 387822 424338 387854 424574
rect 387234 388894 387854 424338
rect 387234 388658 387266 388894
rect 387502 388658 387586 388894
rect 387822 388658 387854 388894
rect 387234 388574 387854 388658
rect 387234 388338 387266 388574
rect 387502 388338 387586 388574
rect 387822 388338 387854 388574
rect 387234 352894 387854 388338
rect 387234 352658 387266 352894
rect 387502 352658 387586 352894
rect 387822 352658 387854 352894
rect 387234 352574 387854 352658
rect 387234 352338 387266 352574
rect 387502 352338 387586 352574
rect 387822 352338 387854 352574
rect 387234 316894 387854 352338
rect 387234 316658 387266 316894
rect 387502 316658 387586 316894
rect 387822 316658 387854 316894
rect 387234 316574 387854 316658
rect 387234 316338 387266 316574
rect 387502 316338 387586 316574
rect 387822 316338 387854 316574
rect 387234 280894 387854 316338
rect 387234 280658 387266 280894
rect 387502 280658 387586 280894
rect 387822 280658 387854 280894
rect 387234 280574 387854 280658
rect 387234 280338 387266 280574
rect 387502 280338 387586 280574
rect 387822 280338 387854 280574
rect 387234 244894 387854 280338
rect 387234 244658 387266 244894
rect 387502 244658 387586 244894
rect 387822 244658 387854 244894
rect 387234 244574 387854 244658
rect 387234 244338 387266 244574
rect 387502 244338 387586 244574
rect 387822 244338 387854 244574
rect 387234 208894 387854 244338
rect 387234 208658 387266 208894
rect 387502 208658 387586 208894
rect 387822 208658 387854 208894
rect 387234 208574 387854 208658
rect 387234 208338 387266 208574
rect 387502 208338 387586 208574
rect 387822 208338 387854 208574
rect 387234 172894 387854 208338
rect 387234 172658 387266 172894
rect 387502 172658 387586 172894
rect 387822 172658 387854 172894
rect 387234 172574 387854 172658
rect 387234 172338 387266 172574
rect 387502 172338 387586 172574
rect 387822 172338 387854 172574
rect 387234 136894 387854 172338
rect 387234 136658 387266 136894
rect 387502 136658 387586 136894
rect 387822 136658 387854 136894
rect 387234 136574 387854 136658
rect 387234 136338 387266 136574
rect 387502 136338 387586 136574
rect 387822 136338 387854 136574
rect 387234 100894 387854 136338
rect 387234 100658 387266 100894
rect 387502 100658 387586 100894
rect 387822 100658 387854 100894
rect 387234 100574 387854 100658
rect 387234 100338 387266 100574
rect 387502 100338 387586 100574
rect 387822 100338 387854 100574
rect 387234 64894 387854 100338
rect 387234 64658 387266 64894
rect 387502 64658 387586 64894
rect 387822 64658 387854 64894
rect 387234 64574 387854 64658
rect 387234 64338 387266 64574
rect 387502 64338 387586 64574
rect 387822 64338 387854 64574
rect 387234 28894 387854 64338
rect 387234 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 387854 28894
rect 387234 28574 387854 28658
rect 387234 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 387854 28574
rect 387234 -5146 387854 28338
rect 387234 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 387854 -5146
rect 387234 -5466 387854 -5382
rect 387234 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 387854 -5466
rect 387234 -5734 387854 -5702
rect 390954 680614 391574 711002
rect 408954 710598 409574 711590
rect 408954 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 409574 710598
rect 408954 710278 409574 710362
rect 408954 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 409574 710278
rect 405234 708678 405854 709670
rect 405234 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 405854 708678
rect 405234 708358 405854 708442
rect 405234 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 405854 708358
rect 401514 706758 402134 707750
rect 401514 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 402134 706758
rect 401514 706438 402134 706522
rect 401514 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 402134 706438
rect 390954 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 391574 680614
rect 390954 680294 391574 680378
rect 390954 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 391574 680294
rect 390954 644614 391574 680058
rect 390954 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 391574 644614
rect 390954 644294 391574 644378
rect 390954 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 391574 644294
rect 390954 608614 391574 644058
rect 390954 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 391574 608614
rect 390954 608294 391574 608378
rect 390954 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 391574 608294
rect 390954 572614 391574 608058
rect 390954 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 391574 572614
rect 390954 572294 391574 572378
rect 390954 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 391574 572294
rect 390954 536614 391574 572058
rect 390954 536378 390986 536614
rect 391222 536378 391306 536614
rect 391542 536378 391574 536614
rect 390954 536294 391574 536378
rect 390954 536058 390986 536294
rect 391222 536058 391306 536294
rect 391542 536058 391574 536294
rect 390954 500614 391574 536058
rect 390954 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 391574 500614
rect 390954 500294 391574 500378
rect 390954 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 391574 500294
rect 390954 464614 391574 500058
rect 390954 464378 390986 464614
rect 391222 464378 391306 464614
rect 391542 464378 391574 464614
rect 390954 464294 391574 464378
rect 390954 464058 390986 464294
rect 391222 464058 391306 464294
rect 391542 464058 391574 464294
rect 390954 428614 391574 464058
rect 390954 428378 390986 428614
rect 391222 428378 391306 428614
rect 391542 428378 391574 428614
rect 390954 428294 391574 428378
rect 390954 428058 390986 428294
rect 391222 428058 391306 428294
rect 391542 428058 391574 428294
rect 390954 392614 391574 428058
rect 390954 392378 390986 392614
rect 391222 392378 391306 392614
rect 391542 392378 391574 392614
rect 390954 392294 391574 392378
rect 390954 392058 390986 392294
rect 391222 392058 391306 392294
rect 391542 392058 391574 392294
rect 390954 356614 391574 392058
rect 390954 356378 390986 356614
rect 391222 356378 391306 356614
rect 391542 356378 391574 356614
rect 390954 356294 391574 356378
rect 390954 356058 390986 356294
rect 391222 356058 391306 356294
rect 391542 356058 391574 356294
rect 390954 320614 391574 356058
rect 390954 320378 390986 320614
rect 391222 320378 391306 320614
rect 391542 320378 391574 320614
rect 390954 320294 391574 320378
rect 390954 320058 390986 320294
rect 391222 320058 391306 320294
rect 391542 320058 391574 320294
rect 390954 284614 391574 320058
rect 390954 284378 390986 284614
rect 391222 284378 391306 284614
rect 391542 284378 391574 284614
rect 390954 284294 391574 284378
rect 390954 284058 390986 284294
rect 391222 284058 391306 284294
rect 391542 284058 391574 284294
rect 390954 248614 391574 284058
rect 390954 248378 390986 248614
rect 391222 248378 391306 248614
rect 391542 248378 391574 248614
rect 390954 248294 391574 248378
rect 390954 248058 390986 248294
rect 391222 248058 391306 248294
rect 391542 248058 391574 248294
rect 390954 212614 391574 248058
rect 390954 212378 390986 212614
rect 391222 212378 391306 212614
rect 391542 212378 391574 212614
rect 390954 212294 391574 212378
rect 390954 212058 390986 212294
rect 391222 212058 391306 212294
rect 391542 212058 391574 212294
rect 390954 176614 391574 212058
rect 390954 176378 390986 176614
rect 391222 176378 391306 176614
rect 391542 176378 391574 176614
rect 390954 176294 391574 176378
rect 390954 176058 390986 176294
rect 391222 176058 391306 176294
rect 391542 176058 391574 176294
rect 390954 140614 391574 176058
rect 390954 140378 390986 140614
rect 391222 140378 391306 140614
rect 391542 140378 391574 140614
rect 390954 140294 391574 140378
rect 390954 140058 390986 140294
rect 391222 140058 391306 140294
rect 391542 140058 391574 140294
rect 390954 104614 391574 140058
rect 390954 104378 390986 104614
rect 391222 104378 391306 104614
rect 391542 104378 391574 104614
rect 390954 104294 391574 104378
rect 390954 104058 390986 104294
rect 391222 104058 391306 104294
rect 391542 104058 391574 104294
rect 390954 68614 391574 104058
rect 390954 68378 390986 68614
rect 391222 68378 391306 68614
rect 391542 68378 391574 68614
rect 390954 68294 391574 68378
rect 390954 68058 390986 68294
rect 391222 68058 391306 68294
rect 391542 68058 391574 68294
rect 390954 32614 391574 68058
rect 390954 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 391574 32614
rect 390954 32294 391574 32378
rect 390954 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 391574 32294
rect 372954 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 373574 -6106
rect 372954 -6426 373574 -6342
rect 372954 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 373574 -6426
rect 372954 -7654 373574 -6662
rect 390954 -7066 391574 32058
rect 397794 704838 398414 705830
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 543454 398414 578898
rect 397794 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 398414 543454
rect 397794 543134 398414 543218
rect 397794 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 398414 543134
rect 397794 507454 398414 542898
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 435454 398414 470898
rect 397794 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 398414 435454
rect 397794 435134 398414 435218
rect 397794 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 398414 435134
rect 397794 399454 398414 434898
rect 397794 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 398414 399454
rect 397794 399134 398414 399218
rect 397794 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 398414 399134
rect 397794 363454 398414 398898
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 397794 327454 398414 362898
rect 397794 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 398414 327454
rect 397794 327134 398414 327218
rect 397794 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 398414 327134
rect 397794 291454 398414 326898
rect 397794 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 398414 291454
rect 397794 291134 398414 291218
rect 397794 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 398414 291134
rect 397794 255454 398414 290898
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 219454 398414 254898
rect 397794 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 398414 219454
rect 397794 219134 398414 219218
rect 397794 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 398414 219134
rect 397794 183454 398414 218898
rect 397794 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 398414 183454
rect 397794 183134 398414 183218
rect 397794 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 398414 183134
rect 397794 147454 398414 182898
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 111454 398414 146898
rect 397794 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 398414 111454
rect 397794 111134 398414 111218
rect 397794 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 398414 111134
rect 397794 75454 398414 110898
rect 397794 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 398414 75454
rect 397794 75134 398414 75218
rect 397794 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 398414 75134
rect 397794 39454 398414 74898
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -1894 398414 -902
rect 401514 691174 402134 706202
rect 401514 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 402134 691174
rect 401514 690854 402134 690938
rect 401514 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 402134 690854
rect 401514 655174 402134 690618
rect 401514 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 402134 655174
rect 401514 654854 402134 654938
rect 401514 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 402134 654854
rect 401514 619174 402134 654618
rect 401514 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 402134 619174
rect 401514 618854 402134 618938
rect 401514 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 402134 618854
rect 401514 583174 402134 618618
rect 401514 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 402134 583174
rect 401514 582854 402134 582938
rect 401514 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 402134 582854
rect 401514 547174 402134 582618
rect 401514 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 402134 547174
rect 401514 546854 402134 546938
rect 401514 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 402134 546854
rect 401514 511174 402134 546618
rect 401514 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 402134 511174
rect 401514 510854 402134 510938
rect 401514 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 402134 510854
rect 401514 475174 402134 510618
rect 401514 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 402134 475174
rect 401514 474854 402134 474938
rect 401514 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 402134 474854
rect 401514 439174 402134 474618
rect 401514 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 402134 439174
rect 401514 438854 402134 438938
rect 401514 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 402134 438854
rect 401514 403174 402134 438618
rect 401514 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 402134 403174
rect 401514 402854 402134 402938
rect 401514 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 402134 402854
rect 401514 367174 402134 402618
rect 401514 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 402134 367174
rect 401514 366854 402134 366938
rect 401514 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 402134 366854
rect 401514 331174 402134 366618
rect 401514 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 402134 331174
rect 401514 330854 402134 330938
rect 401514 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 402134 330854
rect 401514 295174 402134 330618
rect 401514 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 402134 295174
rect 401514 294854 402134 294938
rect 401514 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 402134 294854
rect 401514 259174 402134 294618
rect 401514 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 402134 259174
rect 401514 258854 402134 258938
rect 401514 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 402134 258854
rect 401514 223174 402134 258618
rect 401514 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 402134 223174
rect 401514 222854 402134 222938
rect 401514 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 402134 222854
rect 401514 187174 402134 222618
rect 401514 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 402134 187174
rect 401514 186854 402134 186938
rect 401514 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 402134 186854
rect 401514 151174 402134 186618
rect 401514 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 402134 151174
rect 401514 150854 402134 150938
rect 401514 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 402134 150854
rect 401514 115174 402134 150618
rect 401514 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 402134 115174
rect 401514 114854 402134 114938
rect 401514 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 402134 114854
rect 401514 79174 402134 114618
rect 401514 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 402134 79174
rect 401514 78854 402134 78938
rect 401514 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 402134 78854
rect 401514 43174 402134 78618
rect 401514 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 402134 43174
rect 401514 42854 402134 42938
rect 401514 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 402134 42854
rect 401514 7174 402134 42618
rect 401514 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 402134 7174
rect 401514 6854 402134 6938
rect 401514 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 402134 6854
rect 401514 -2266 402134 6618
rect 401514 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 402134 -2266
rect 401514 -2586 402134 -2502
rect 401514 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 402134 -2586
rect 401514 -3814 402134 -2822
rect 405234 694894 405854 708122
rect 405234 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 405854 694894
rect 405234 694574 405854 694658
rect 405234 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 405854 694574
rect 405234 658894 405854 694338
rect 405234 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 405854 658894
rect 405234 658574 405854 658658
rect 405234 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 405854 658574
rect 405234 622894 405854 658338
rect 405234 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 405854 622894
rect 405234 622574 405854 622658
rect 405234 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 405854 622574
rect 405234 586894 405854 622338
rect 405234 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 405854 586894
rect 405234 586574 405854 586658
rect 405234 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 405854 586574
rect 405234 550894 405854 586338
rect 405234 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 405854 550894
rect 405234 550574 405854 550658
rect 405234 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 405854 550574
rect 405234 514894 405854 550338
rect 405234 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 405854 514894
rect 405234 514574 405854 514658
rect 405234 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 405854 514574
rect 405234 478894 405854 514338
rect 405234 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 405854 478894
rect 405234 478574 405854 478658
rect 405234 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 405854 478574
rect 405234 442894 405854 478338
rect 405234 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 405854 442894
rect 405234 442574 405854 442658
rect 405234 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 405854 442574
rect 405234 406894 405854 442338
rect 405234 406658 405266 406894
rect 405502 406658 405586 406894
rect 405822 406658 405854 406894
rect 405234 406574 405854 406658
rect 405234 406338 405266 406574
rect 405502 406338 405586 406574
rect 405822 406338 405854 406574
rect 405234 370894 405854 406338
rect 405234 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 405854 370894
rect 405234 370574 405854 370658
rect 405234 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 405854 370574
rect 405234 334894 405854 370338
rect 405234 334658 405266 334894
rect 405502 334658 405586 334894
rect 405822 334658 405854 334894
rect 405234 334574 405854 334658
rect 405234 334338 405266 334574
rect 405502 334338 405586 334574
rect 405822 334338 405854 334574
rect 405234 298894 405854 334338
rect 405234 298658 405266 298894
rect 405502 298658 405586 298894
rect 405822 298658 405854 298894
rect 405234 298574 405854 298658
rect 405234 298338 405266 298574
rect 405502 298338 405586 298574
rect 405822 298338 405854 298574
rect 405234 262894 405854 298338
rect 405234 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 405854 262894
rect 405234 262574 405854 262658
rect 405234 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 405854 262574
rect 405234 226894 405854 262338
rect 405234 226658 405266 226894
rect 405502 226658 405586 226894
rect 405822 226658 405854 226894
rect 405234 226574 405854 226658
rect 405234 226338 405266 226574
rect 405502 226338 405586 226574
rect 405822 226338 405854 226574
rect 405234 190894 405854 226338
rect 405234 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 405854 190894
rect 405234 190574 405854 190658
rect 405234 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 405854 190574
rect 405234 154894 405854 190338
rect 405234 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 405854 154894
rect 405234 154574 405854 154658
rect 405234 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 405854 154574
rect 405234 118894 405854 154338
rect 405234 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 405854 118894
rect 405234 118574 405854 118658
rect 405234 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 405854 118574
rect 405234 82894 405854 118338
rect 405234 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 405854 82894
rect 405234 82574 405854 82658
rect 405234 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 405854 82574
rect 405234 46894 405854 82338
rect 405234 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 405854 46894
rect 405234 46574 405854 46658
rect 405234 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 405854 46574
rect 405234 10894 405854 46338
rect 405234 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 405854 10894
rect 405234 10574 405854 10658
rect 405234 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 405854 10574
rect 405234 -4186 405854 10338
rect 405234 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 405854 -4186
rect 405234 -4506 405854 -4422
rect 405234 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 405854 -4506
rect 405234 -5734 405854 -4742
rect 408954 698614 409574 710042
rect 426954 711558 427574 711590
rect 426954 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 427574 711558
rect 426954 711238 427574 711322
rect 426954 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 427574 711238
rect 423234 709638 423854 709670
rect 423234 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 423854 709638
rect 423234 709318 423854 709402
rect 423234 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 423854 709318
rect 419514 707718 420134 707750
rect 419514 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 420134 707718
rect 419514 707398 420134 707482
rect 419514 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 420134 707398
rect 408954 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 409574 698614
rect 408954 698294 409574 698378
rect 408954 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 409574 698294
rect 408954 662614 409574 698058
rect 408954 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 409574 662614
rect 408954 662294 409574 662378
rect 408954 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 409574 662294
rect 408954 626614 409574 662058
rect 408954 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 409574 626614
rect 408954 626294 409574 626378
rect 408954 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 409574 626294
rect 408954 590614 409574 626058
rect 408954 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 409574 590614
rect 408954 590294 409574 590378
rect 408954 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 409574 590294
rect 408954 554614 409574 590058
rect 408954 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 409574 554614
rect 408954 554294 409574 554378
rect 408954 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 409574 554294
rect 408954 518614 409574 554058
rect 408954 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 409574 518614
rect 408954 518294 409574 518378
rect 408954 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 409574 518294
rect 408954 482614 409574 518058
rect 408954 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 409574 482614
rect 408954 482294 409574 482378
rect 408954 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 409574 482294
rect 408954 446614 409574 482058
rect 408954 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 409574 446614
rect 408954 446294 409574 446378
rect 408954 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 409574 446294
rect 408954 410614 409574 446058
rect 408954 410378 408986 410614
rect 409222 410378 409306 410614
rect 409542 410378 409574 410614
rect 408954 410294 409574 410378
rect 408954 410058 408986 410294
rect 409222 410058 409306 410294
rect 409542 410058 409574 410294
rect 408954 374614 409574 410058
rect 408954 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 409574 374614
rect 408954 374294 409574 374378
rect 408954 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 409574 374294
rect 408954 338614 409574 374058
rect 408954 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 409574 338614
rect 408954 338294 409574 338378
rect 408954 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 409574 338294
rect 408954 302614 409574 338058
rect 408954 302378 408986 302614
rect 409222 302378 409306 302614
rect 409542 302378 409574 302614
rect 408954 302294 409574 302378
rect 408954 302058 408986 302294
rect 409222 302058 409306 302294
rect 409542 302058 409574 302294
rect 408954 266614 409574 302058
rect 408954 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 409574 266614
rect 408954 266294 409574 266378
rect 408954 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 409574 266294
rect 408954 230614 409574 266058
rect 408954 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 409574 230614
rect 408954 230294 409574 230378
rect 408954 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 409574 230294
rect 408954 194614 409574 230058
rect 408954 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 409574 194614
rect 408954 194294 409574 194378
rect 408954 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 409574 194294
rect 408954 158614 409574 194058
rect 408954 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 409574 158614
rect 408954 158294 409574 158378
rect 408954 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 409574 158294
rect 408954 122614 409574 158058
rect 408954 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 409574 122614
rect 408954 122294 409574 122378
rect 408954 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 409574 122294
rect 408954 86614 409574 122058
rect 408954 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 409574 86614
rect 408954 86294 409574 86378
rect 408954 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 409574 86294
rect 408954 50614 409574 86058
rect 408954 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 409574 50614
rect 408954 50294 409574 50378
rect 408954 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 409574 50294
rect 408954 14614 409574 50058
rect 408954 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 409574 14614
rect 408954 14294 409574 14378
rect 408954 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 409574 14294
rect 390954 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 391574 -7066
rect 390954 -7386 391574 -7302
rect 390954 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 391574 -7386
rect 390954 -7654 391574 -7622
rect 408954 -6106 409574 14058
rect 415794 705798 416414 705830
rect 415794 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 416414 705798
rect 415794 705478 416414 705562
rect 415794 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 416414 705478
rect 415794 669454 416414 705242
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 633454 416414 668898
rect 415794 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 416414 633454
rect 415794 633134 416414 633218
rect 415794 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 416414 633134
rect 415794 597454 416414 632898
rect 415794 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 416414 597454
rect 415794 597134 416414 597218
rect 415794 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 416414 597134
rect 415794 561454 416414 596898
rect 415794 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 416414 561454
rect 415794 561134 416414 561218
rect 415794 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 416414 561134
rect 415794 525454 416414 560898
rect 415794 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 416414 525454
rect 415794 525134 416414 525218
rect 415794 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 416414 525134
rect 415794 489454 416414 524898
rect 415794 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 416414 489454
rect 415794 489134 416414 489218
rect 415794 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 416414 489134
rect 415794 453454 416414 488898
rect 415794 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 416414 453454
rect 415794 453134 416414 453218
rect 415794 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 416414 453134
rect 415794 417454 416414 452898
rect 415794 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 416414 417454
rect 415794 417134 416414 417218
rect 415794 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 416414 417134
rect 415794 381454 416414 416898
rect 415794 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 416414 381454
rect 415794 381134 416414 381218
rect 415794 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 416414 381134
rect 415794 345454 416414 380898
rect 415794 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 416414 345454
rect 415794 345134 416414 345218
rect 415794 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 416414 345134
rect 415794 309454 416414 344898
rect 415794 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 416414 309454
rect 415794 309134 416414 309218
rect 415794 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 416414 309134
rect 415794 273454 416414 308898
rect 415794 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 416414 273454
rect 415794 273134 416414 273218
rect 415794 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 416414 273134
rect 415794 237454 416414 272898
rect 415794 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 416414 237454
rect 415794 237134 416414 237218
rect 415794 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 416414 237134
rect 415794 201454 416414 236898
rect 415794 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 416414 201454
rect 415794 201134 416414 201218
rect 415794 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 416414 201134
rect 415794 165454 416414 200898
rect 415794 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 416414 165454
rect 415794 165134 416414 165218
rect 415794 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 416414 165134
rect 415794 129454 416414 164898
rect 415794 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 416414 129454
rect 415794 129134 416414 129218
rect 415794 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 416414 129134
rect 415794 93454 416414 128898
rect 415794 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 416414 93454
rect 415794 93134 416414 93218
rect 415794 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 416414 93134
rect 415794 57454 416414 92898
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -1306 416414 20898
rect 415794 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 416414 -1306
rect 415794 -1626 416414 -1542
rect 415794 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 416414 -1626
rect 415794 -1894 416414 -1862
rect 419514 673174 420134 707162
rect 419514 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 420134 673174
rect 419514 672854 420134 672938
rect 419514 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 420134 672854
rect 419514 637174 420134 672618
rect 419514 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 420134 637174
rect 419514 636854 420134 636938
rect 419514 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 420134 636854
rect 419514 601174 420134 636618
rect 419514 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 420134 601174
rect 419514 600854 420134 600938
rect 419514 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 420134 600854
rect 419514 565174 420134 600618
rect 419514 564938 419546 565174
rect 419782 564938 419866 565174
rect 420102 564938 420134 565174
rect 419514 564854 420134 564938
rect 419514 564618 419546 564854
rect 419782 564618 419866 564854
rect 420102 564618 420134 564854
rect 419514 529174 420134 564618
rect 419514 528938 419546 529174
rect 419782 528938 419866 529174
rect 420102 528938 420134 529174
rect 419514 528854 420134 528938
rect 419514 528618 419546 528854
rect 419782 528618 419866 528854
rect 420102 528618 420134 528854
rect 419514 493174 420134 528618
rect 419514 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 420134 493174
rect 419514 492854 420134 492938
rect 419514 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 420134 492854
rect 419514 457174 420134 492618
rect 419514 456938 419546 457174
rect 419782 456938 419866 457174
rect 420102 456938 420134 457174
rect 419514 456854 420134 456938
rect 419514 456618 419546 456854
rect 419782 456618 419866 456854
rect 420102 456618 420134 456854
rect 419514 421174 420134 456618
rect 419514 420938 419546 421174
rect 419782 420938 419866 421174
rect 420102 420938 420134 421174
rect 419514 420854 420134 420938
rect 419514 420618 419546 420854
rect 419782 420618 419866 420854
rect 420102 420618 420134 420854
rect 419514 385174 420134 420618
rect 419514 384938 419546 385174
rect 419782 384938 419866 385174
rect 420102 384938 420134 385174
rect 419514 384854 420134 384938
rect 419514 384618 419546 384854
rect 419782 384618 419866 384854
rect 420102 384618 420134 384854
rect 419514 349174 420134 384618
rect 419514 348938 419546 349174
rect 419782 348938 419866 349174
rect 420102 348938 420134 349174
rect 419514 348854 420134 348938
rect 419514 348618 419546 348854
rect 419782 348618 419866 348854
rect 420102 348618 420134 348854
rect 419514 313174 420134 348618
rect 419514 312938 419546 313174
rect 419782 312938 419866 313174
rect 420102 312938 420134 313174
rect 419514 312854 420134 312938
rect 419514 312618 419546 312854
rect 419782 312618 419866 312854
rect 420102 312618 420134 312854
rect 419514 277174 420134 312618
rect 419514 276938 419546 277174
rect 419782 276938 419866 277174
rect 420102 276938 420134 277174
rect 419514 276854 420134 276938
rect 419514 276618 419546 276854
rect 419782 276618 419866 276854
rect 420102 276618 420134 276854
rect 419514 241174 420134 276618
rect 419514 240938 419546 241174
rect 419782 240938 419866 241174
rect 420102 240938 420134 241174
rect 419514 240854 420134 240938
rect 419514 240618 419546 240854
rect 419782 240618 419866 240854
rect 420102 240618 420134 240854
rect 419514 205174 420134 240618
rect 419514 204938 419546 205174
rect 419782 204938 419866 205174
rect 420102 204938 420134 205174
rect 419514 204854 420134 204938
rect 419514 204618 419546 204854
rect 419782 204618 419866 204854
rect 420102 204618 420134 204854
rect 419514 169174 420134 204618
rect 419514 168938 419546 169174
rect 419782 168938 419866 169174
rect 420102 168938 420134 169174
rect 419514 168854 420134 168938
rect 419514 168618 419546 168854
rect 419782 168618 419866 168854
rect 420102 168618 420134 168854
rect 419514 133174 420134 168618
rect 419514 132938 419546 133174
rect 419782 132938 419866 133174
rect 420102 132938 420134 133174
rect 419514 132854 420134 132938
rect 419514 132618 419546 132854
rect 419782 132618 419866 132854
rect 420102 132618 420134 132854
rect 419514 97174 420134 132618
rect 419514 96938 419546 97174
rect 419782 96938 419866 97174
rect 420102 96938 420134 97174
rect 419514 96854 420134 96938
rect 419514 96618 419546 96854
rect 419782 96618 419866 96854
rect 420102 96618 420134 96854
rect 419514 61174 420134 96618
rect 419514 60938 419546 61174
rect 419782 60938 419866 61174
rect 420102 60938 420134 61174
rect 419514 60854 420134 60938
rect 419514 60618 419546 60854
rect 419782 60618 419866 60854
rect 420102 60618 420134 60854
rect 419514 25174 420134 60618
rect 419514 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 420134 25174
rect 419514 24854 420134 24938
rect 419514 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 420134 24854
rect 419514 -3226 420134 24618
rect 419514 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 420134 -3226
rect 419514 -3546 420134 -3462
rect 419514 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 420134 -3546
rect 419514 -3814 420134 -3782
rect 423234 676894 423854 709082
rect 423234 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 423854 676894
rect 423234 676574 423854 676658
rect 423234 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 423854 676574
rect 423234 640894 423854 676338
rect 423234 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 423854 640894
rect 423234 640574 423854 640658
rect 423234 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 423854 640574
rect 423234 604894 423854 640338
rect 423234 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 423854 604894
rect 423234 604574 423854 604658
rect 423234 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 423854 604574
rect 423234 568894 423854 604338
rect 423234 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 423854 568894
rect 423234 568574 423854 568658
rect 423234 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 423854 568574
rect 423234 532894 423854 568338
rect 423234 532658 423266 532894
rect 423502 532658 423586 532894
rect 423822 532658 423854 532894
rect 423234 532574 423854 532658
rect 423234 532338 423266 532574
rect 423502 532338 423586 532574
rect 423822 532338 423854 532574
rect 423234 496894 423854 532338
rect 423234 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 423854 496894
rect 423234 496574 423854 496658
rect 423234 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 423854 496574
rect 423234 460894 423854 496338
rect 423234 460658 423266 460894
rect 423502 460658 423586 460894
rect 423822 460658 423854 460894
rect 423234 460574 423854 460658
rect 423234 460338 423266 460574
rect 423502 460338 423586 460574
rect 423822 460338 423854 460574
rect 423234 424894 423854 460338
rect 423234 424658 423266 424894
rect 423502 424658 423586 424894
rect 423822 424658 423854 424894
rect 423234 424574 423854 424658
rect 423234 424338 423266 424574
rect 423502 424338 423586 424574
rect 423822 424338 423854 424574
rect 423234 388894 423854 424338
rect 423234 388658 423266 388894
rect 423502 388658 423586 388894
rect 423822 388658 423854 388894
rect 423234 388574 423854 388658
rect 423234 388338 423266 388574
rect 423502 388338 423586 388574
rect 423822 388338 423854 388574
rect 423234 352894 423854 388338
rect 423234 352658 423266 352894
rect 423502 352658 423586 352894
rect 423822 352658 423854 352894
rect 423234 352574 423854 352658
rect 423234 352338 423266 352574
rect 423502 352338 423586 352574
rect 423822 352338 423854 352574
rect 423234 316894 423854 352338
rect 423234 316658 423266 316894
rect 423502 316658 423586 316894
rect 423822 316658 423854 316894
rect 423234 316574 423854 316658
rect 423234 316338 423266 316574
rect 423502 316338 423586 316574
rect 423822 316338 423854 316574
rect 423234 280894 423854 316338
rect 423234 280658 423266 280894
rect 423502 280658 423586 280894
rect 423822 280658 423854 280894
rect 423234 280574 423854 280658
rect 423234 280338 423266 280574
rect 423502 280338 423586 280574
rect 423822 280338 423854 280574
rect 423234 244894 423854 280338
rect 423234 244658 423266 244894
rect 423502 244658 423586 244894
rect 423822 244658 423854 244894
rect 423234 244574 423854 244658
rect 423234 244338 423266 244574
rect 423502 244338 423586 244574
rect 423822 244338 423854 244574
rect 423234 208894 423854 244338
rect 423234 208658 423266 208894
rect 423502 208658 423586 208894
rect 423822 208658 423854 208894
rect 423234 208574 423854 208658
rect 423234 208338 423266 208574
rect 423502 208338 423586 208574
rect 423822 208338 423854 208574
rect 423234 172894 423854 208338
rect 423234 172658 423266 172894
rect 423502 172658 423586 172894
rect 423822 172658 423854 172894
rect 423234 172574 423854 172658
rect 423234 172338 423266 172574
rect 423502 172338 423586 172574
rect 423822 172338 423854 172574
rect 423234 136894 423854 172338
rect 423234 136658 423266 136894
rect 423502 136658 423586 136894
rect 423822 136658 423854 136894
rect 423234 136574 423854 136658
rect 423234 136338 423266 136574
rect 423502 136338 423586 136574
rect 423822 136338 423854 136574
rect 423234 100894 423854 136338
rect 423234 100658 423266 100894
rect 423502 100658 423586 100894
rect 423822 100658 423854 100894
rect 423234 100574 423854 100658
rect 423234 100338 423266 100574
rect 423502 100338 423586 100574
rect 423822 100338 423854 100574
rect 423234 64894 423854 100338
rect 423234 64658 423266 64894
rect 423502 64658 423586 64894
rect 423822 64658 423854 64894
rect 423234 64574 423854 64658
rect 423234 64338 423266 64574
rect 423502 64338 423586 64574
rect 423822 64338 423854 64574
rect 423234 28894 423854 64338
rect 423234 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 423854 28894
rect 423234 28574 423854 28658
rect 423234 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 423854 28574
rect 423234 -5146 423854 28338
rect 423234 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 423854 -5146
rect 423234 -5466 423854 -5382
rect 423234 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 423854 -5466
rect 423234 -5734 423854 -5702
rect 426954 680614 427574 711002
rect 444954 710598 445574 711590
rect 444954 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 445574 710598
rect 444954 710278 445574 710362
rect 444954 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 445574 710278
rect 441234 708678 441854 709670
rect 441234 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 441854 708678
rect 441234 708358 441854 708442
rect 441234 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 441854 708358
rect 437514 706758 438134 707750
rect 437514 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 438134 706758
rect 437514 706438 438134 706522
rect 437514 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 438134 706438
rect 426954 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 427574 680614
rect 426954 680294 427574 680378
rect 426954 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 427574 680294
rect 426954 644614 427574 680058
rect 426954 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 427574 644614
rect 426954 644294 427574 644378
rect 426954 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 427574 644294
rect 426954 608614 427574 644058
rect 426954 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 427574 608614
rect 426954 608294 427574 608378
rect 426954 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 427574 608294
rect 426954 572614 427574 608058
rect 426954 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 427574 572614
rect 426954 572294 427574 572378
rect 426954 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 427574 572294
rect 426954 536614 427574 572058
rect 426954 536378 426986 536614
rect 427222 536378 427306 536614
rect 427542 536378 427574 536614
rect 426954 536294 427574 536378
rect 426954 536058 426986 536294
rect 427222 536058 427306 536294
rect 427542 536058 427574 536294
rect 426954 500614 427574 536058
rect 426954 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 427574 500614
rect 426954 500294 427574 500378
rect 426954 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 427574 500294
rect 426954 464614 427574 500058
rect 426954 464378 426986 464614
rect 427222 464378 427306 464614
rect 427542 464378 427574 464614
rect 426954 464294 427574 464378
rect 426954 464058 426986 464294
rect 427222 464058 427306 464294
rect 427542 464058 427574 464294
rect 426954 428614 427574 464058
rect 426954 428378 426986 428614
rect 427222 428378 427306 428614
rect 427542 428378 427574 428614
rect 426954 428294 427574 428378
rect 426954 428058 426986 428294
rect 427222 428058 427306 428294
rect 427542 428058 427574 428294
rect 426954 392614 427574 428058
rect 426954 392378 426986 392614
rect 427222 392378 427306 392614
rect 427542 392378 427574 392614
rect 426954 392294 427574 392378
rect 426954 392058 426986 392294
rect 427222 392058 427306 392294
rect 427542 392058 427574 392294
rect 426954 356614 427574 392058
rect 426954 356378 426986 356614
rect 427222 356378 427306 356614
rect 427542 356378 427574 356614
rect 426954 356294 427574 356378
rect 426954 356058 426986 356294
rect 427222 356058 427306 356294
rect 427542 356058 427574 356294
rect 426954 320614 427574 356058
rect 426954 320378 426986 320614
rect 427222 320378 427306 320614
rect 427542 320378 427574 320614
rect 426954 320294 427574 320378
rect 426954 320058 426986 320294
rect 427222 320058 427306 320294
rect 427542 320058 427574 320294
rect 426954 284614 427574 320058
rect 426954 284378 426986 284614
rect 427222 284378 427306 284614
rect 427542 284378 427574 284614
rect 426954 284294 427574 284378
rect 426954 284058 426986 284294
rect 427222 284058 427306 284294
rect 427542 284058 427574 284294
rect 426954 248614 427574 284058
rect 426954 248378 426986 248614
rect 427222 248378 427306 248614
rect 427542 248378 427574 248614
rect 426954 248294 427574 248378
rect 426954 248058 426986 248294
rect 427222 248058 427306 248294
rect 427542 248058 427574 248294
rect 426954 212614 427574 248058
rect 426954 212378 426986 212614
rect 427222 212378 427306 212614
rect 427542 212378 427574 212614
rect 426954 212294 427574 212378
rect 426954 212058 426986 212294
rect 427222 212058 427306 212294
rect 427542 212058 427574 212294
rect 426954 176614 427574 212058
rect 426954 176378 426986 176614
rect 427222 176378 427306 176614
rect 427542 176378 427574 176614
rect 426954 176294 427574 176378
rect 426954 176058 426986 176294
rect 427222 176058 427306 176294
rect 427542 176058 427574 176294
rect 426954 140614 427574 176058
rect 426954 140378 426986 140614
rect 427222 140378 427306 140614
rect 427542 140378 427574 140614
rect 426954 140294 427574 140378
rect 426954 140058 426986 140294
rect 427222 140058 427306 140294
rect 427542 140058 427574 140294
rect 426954 104614 427574 140058
rect 426954 104378 426986 104614
rect 427222 104378 427306 104614
rect 427542 104378 427574 104614
rect 426954 104294 427574 104378
rect 426954 104058 426986 104294
rect 427222 104058 427306 104294
rect 427542 104058 427574 104294
rect 426954 68614 427574 104058
rect 426954 68378 426986 68614
rect 427222 68378 427306 68614
rect 427542 68378 427574 68614
rect 426954 68294 427574 68378
rect 426954 68058 426986 68294
rect 427222 68058 427306 68294
rect 427542 68058 427574 68294
rect 426954 32614 427574 68058
rect 426954 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 427574 32614
rect 426954 32294 427574 32378
rect 426954 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 427574 32294
rect 408954 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 409574 -6106
rect 408954 -6426 409574 -6342
rect 408954 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 409574 -6426
rect 408954 -7654 409574 -6662
rect 426954 -7066 427574 32058
rect 433794 704838 434414 705830
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 433794 507454 434414 542898
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 471454 434414 506898
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 435454 434414 470898
rect 433794 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 434414 435454
rect 433794 435134 434414 435218
rect 433794 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 434414 435134
rect 433794 399454 434414 434898
rect 433794 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 434414 399454
rect 433794 399134 434414 399218
rect 433794 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 434414 399134
rect 433794 363454 434414 398898
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 433794 327454 434414 362898
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 433794 291454 434414 326898
rect 433794 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 434414 291454
rect 433794 291134 434414 291218
rect 433794 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 434414 291134
rect 433794 255454 434414 290898
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 219454 434414 254898
rect 433794 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 434414 219454
rect 433794 219134 434414 219218
rect 433794 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 434414 219134
rect 433794 183454 434414 218898
rect 433794 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 434414 183454
rect 433794 183134 434414 183218
rect 433794 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 434414 183134
rect 433794 147454 434414 182898
rect 433794 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 434414 147454
rect 433794 147134 434414 147218
rect 433794 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 434414 147134
rect 433794 111454 434414 146898
rect 433794 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 434414 111454
rect 433794 111134 434414 111218
rect 433794 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 434414 111134
rect 433794 75454 434414 110898
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 433794 39454 434414 74898
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -1894 434414 -902
rect 437514 691174 438134 706202
rect 437514 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 438134 691174
rect 437514 690854 438134 690938
rect 437514 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 438134 690854
rect 437514 655174 438134 690618
rect 437514 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 438134 655174
rect 437514 654854 438134 654938
rect 437514 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 438134 654854
rect 437514 619174 438134 654618
rect 437514 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 438134 619174
rect 437514 618854 438134 618938
rect 437514 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 438134 618854
rect 437514 583174 438134 618618
rect 437514 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 438134 583174
rect 437514 582854 438134 582938
rect 437514 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 438134 582854
rect 437514 547174 438134 582618
rect 437514 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 438134 547174
rect 437514 546854 438134 546938
rect 437514 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 438134 546854
rect 437514 511174 438134 546618
rect 437514 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 438134 511174
rect 437514 510854 438134 510938
rect 437514 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 438134 510854
rect 437514 475174 438134 510618
rect 437514 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 438134 475174
rect 437514 474854 438134 474938
rect 437514 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 438134 474854
rect 437514 439174 438134 474618
rect 437514 438938 437546 439174
rect 437782 438938 437866 439174
rect 438102 438938 438134 439174
rect 437514 438854 438134 438938
rect 437514 438618 437546 438854
rect 437782 438618 437866 438854
rect 438102 438618 438134 438854
rect 437514 403174 438134 438618
rect 437514 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 438134 403174
rect 437514 402854 438134 402938
rect 437514 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 438134 402854
rect 437514 367174 438134 402618
rect 437514 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 438134 367174
rect 437514 366854 438134 366938
rect 437514 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 438134 366854
rect 437514 331174 438134 366618
rect 437514 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 438134 331174
rect 437514 330854 438134 330938
rect 437514 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 438134 330854
rect 437514 295174 438134 330618
rect 437514 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 438134 295174
rect 437514 294854 438134 294938
rect 437514 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 438134 294854
rect 437514 259174 438134 294618
rect 437514 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 438134 259174
rect 437514 258854 438134 258938
rect 437514 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 438134 258854
rect 437514 223174 438134 258618
rect 437514 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 438134 223174
rect 437514 222854 438134 222938
rect 437514 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 438134 222854
rect 437514 187174 438134 222618
rect 437514 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 438134 187174
rect 437514 186854 438134 186938
rect 437514 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 438134 186854
rect 437514 151174 438134 186618
rect 437514 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 438134 151174
rect 437514 150854 438134 150938
rect 437514 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 438134 150854
rect 437514 115174 438134 150618
rect 437514 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 438134 115174
rect 437514 114854 438134 114938
rect 437514 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 438134 114854
rect 437514 79174 438134 114618
rect 437514 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 438134 79174
rect 437514 78854 438134 78938
rect 437514 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 438134 78854
rect 437514 43174 438134 78618
rect 437514 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 438134 43174
rect 437514 42854 438134 42938
rect 437514 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 438134 42854
rect 437514 7174 438134 42618
rect 437514 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 438134 7174
rect 437514 6854 438134 6938
rect 437514 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 438134 6854
rect 437514 -2266 438134 6618
rect 437514 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 438134 -2266
rect 437514 -2586 438134 -2502
rect 437514 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 438134 -2586
rect 437514 -3814 438134 -2822
rect 441234 694894 441854 708122
rect 441234 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 441854 694894
rect 441234 694574 441854 694658
rect 441234 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 441854 694574
rect 441234 658894 441854 694338
rect 441234 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 441854 658894
rect 441234 658574 441854 658658
rect 441234 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 441854 658574
rect 441234 622894 441854 658338
rect 441234 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 441854 622894
rect 441234 622574 441854 622658
rect 441234 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 441854 622574
rect 441234 586894 441854 622338
rect 441234 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 441854 586894
rect 441234 586574 441854 586658
rect 441234 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 441854 586574
rect 441234 550894 441854 586338
rect 441234 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 441854 550894
rect 441234 550574 441854 550658
rect 441234 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 441854 550574
rect 441234 514894 441854 550338
rect 441234 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 441854 514894
rect 441234 514574 441854 514658
rect 441234 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 441854 514574
rect 441234 478894 441854 514338
rect 441234 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 441854 478894
rect 441234 478574 441854 478658
rect 441234 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 441854 478574
rect 441234 442894 441854 478338
rect 441234 442658 441266 442894
rect 441502 442658 441586 442894
rect 441822 442658 441854 442894
rect 441234 442574 441854 442658
rect 441234 442338 441266 442574
rect 441502 442338 441586 442574
rect 441822 442338 441854 442574
rect 441234 406894 441854 442338
rect 441234 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 441854 406894
rect 441234 406574 441854 406658
rect 441234 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 441854 406574
rect 441234 370894 441854 406338
rect 441234 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 441854 370894
rect 441234 370574 441854 370658
rect 441234 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 441854 370574
rect 441234 334894 441854 370338
rect 441234 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 441854 334894
rect 441234 334574 441854 334658
rect 441234 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 441854 334574
rect 441234 298894 441854 334338
rect 441234 298658 441266 298894
rect 441502 298658 441586 298894
rect 441822 298658 441854 298894
rect 441234 298574 441854 298658
rect 441234 298338 441266 298574
rect 441502 298338 441586 298574
rect 441822 298338 441854 298574
rect 441234 262894 441854 298338
rect 441234 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 441854 262894
rect 441234 262574 441854 262658
rect 441234 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 441854 262574
rect 441234 226894 441854 262338
rect 441234 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 441854 226894
rect 441234 226574 441854 226658
rect 441234 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 441854 226574
rect 441234 190894 441854 226338
rect 441234 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 441854 190894
rect 441234 190574 441854 190658
rect 441234 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 441854 190574
rect 441234 154894 441854 190338
rect 441234 154658 441266 154894
rect 441502 154658 441586 154894
rect 441822 154658 441854 154894
rect 441234 154574 441854 154658
rect 441234 154338 441266 154574
rect 441502 154338 441586 154574
rect 441822 154338 441854 154574
rect 441234 118894 441854 154338
rect 441234 118658 441266 118894
rect 441502 118658 441586 118894
rect 441822 118658 441854 118894
rect 441234 118574 441854 118658
rect 441234 118338 441266 118574
rect 441502 118338 441586 118574
rect 441822 118338 441854 118574
rect 441234 82894 441854 118338
rect 441234 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 441854 82894
rect 441234 82574 441854 82658
rect 441234 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 441854 82574
rect 441234 46894 441854 82338
rect 441234 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 441854 46894
rect 441234 46574 441854 46658
rect 441234 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 441854 46574
rect 441234 10894 441854 46338
rect 441234 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 441854 10894
rect 441234 10574 441854 10658
rect 441234 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 441854 10574
rect 441234 -4186 441854 10338
rect 441234 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 441854 -4186
rect 441234 -4506 441854 -4422
rect 441234 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 441854 -4506
rect 441234 -5734 441854 -4742
rect 444954 698614 445574 710042
rect 462954 711558 463574 711590
rect 462954 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 463574 711558
rect 462954 711238 463574 711322
rect 462954 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 463574 711238
rect 459234 709638 459854 709670
rect 459234 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 459854 709638
rect 459234 709318 459854 709402
rect 459234 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 459854 709318
rect 455514 707718 456134 707750
rect 455514 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 456134 707718
rect 455514 707398 456134 707482
rect 455514 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 456134 707398
rect 444954 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 445574 698614
rect 444954 698294 445574 698378
rect 444954 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 445574 698294
rect 444954 662614 445574 698058
rect 444954 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 445574 662614
rect 444954 662294 445574 662378
rect 444954 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 445574 662294
rect 444954 626614 445574 662058
rect 444954 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 445574 626614
rect 444954 626294 445574 626378
rect 444954 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 445574 626294
rect 444954 590614 445574 626058
rect 444954 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 445574 590614
rect 444954 590294 445574 590378
rect 444954 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 445574 590294
rect 444954 554614 445574 590058
rect 444954 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 445574 554614
rect 444954 554294 445574 554378
rect 444954 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 445574 554294
rect 444954 518614 445574 554058
rect 444954 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 445574 518614
rect 444954 518294 445574 518378
rect 444954 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 445574 518294
rect 444954 482614 445574 518058
rect 444954 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 445574 482614
rect 444954 482294 445574 482378
rect 444954 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 445574 482294
rect 444954 446614 445574 482058
rect 444954 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 445574 446614
rect 444954 446294 445574 446378
rect 444954 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 445574 446294
rect 444954 410614 445574 446058
rect 444954 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 445574 410614
rect 444954 410294 445574 410378
rect 444954 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 445574 410294
rect 444954 374614 445574 410058
rect 444954 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 445574 374614
rect 444954 374294 445574 374378
rect 444954 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 445574 374294
rect 444954 338614 445574 374058
rect 444954 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 445574 338614
rect 444954 338294 445574 338378
rect 444954 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 445574 338294
rect 444954 302614 445574 338058
rect 444954 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 445574 302614
rect 444954 302294 445574 302378
rect 444954 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 445574 302294
rect 444954 266614 445574 302058
rect 444954 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 445574 266614
rect 444954 266294 445574 266378
rect 444954 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 445574 266294
rect 444954 230614 445574 266058
rect 444954 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 445574 230614
rect 444954 230294 445574 230378
rect 444954 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 445574 230294
rect 444954 194614 445574 230058
rect 444954 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 445574 194614
rect 444954 194294 445574 194378
rect 444954 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 445574 194294
rect 444954 158614 445574 194058
rect 444954 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 445574 158614
rect 444954 158294 445574 158378
rect 444954 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 445574 158294
rect 444954 122614 445574 158058
rect 444954 122378 444986 122614
rect 445222 122378 445306 122614
rect 445542 122378 445574 122614
rect 444954 122294 445574 122378
rect 444954 122058 444986 122294
rect 445222 122058 445306 122294
rect 445542 122058 445574 122294
rect 444954 86614 445574 122058
rect 444954 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 445574 86614
rect 444954 86294 445574 86378
rect 444954 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 445574 86294
rect 444954 50614 445574 86058
rect 444954 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 445574 50614
rect 444954 50294 445574 50378
rect 444954 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 445574 50294
rect 444954 14614 445574 50058
rect 444954 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 445574 14614
rect 444954 14294 445574 14378
rect 444954 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 445574 14294
rect 426954 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 427574 -7066
rect 426954 -7386 427574 -7302
rect 426954 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 427574 -7386
rect 426954 -7654 427574 -7622
rect 444954 -6106 445574 14058
rect 451794 705798 452414 705830
rect 451794 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 452414 705798
rect 451794 705478 452414 705562
rect 451794 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 452414 705478
rect 451794 669454 452414 705242
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597454 452414 632898
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 561454 452414 596898
rect 451794 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 452414 561454
rect 451794 561134 452414 561218
rect 451794 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 452414 561134
rect 451794 525454 452414 560898
rect 451794 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 452414 525454
rect 451794 525134 452414 525218
rect 451794 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 452414 525134
rect 451794 489454 452414 524898
rect 451794 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 452414 489454
rect 451794 489134 452414 489218
rect 451794 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 452414 489134
rect 451794 453454 452414 488898
rect 451794 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 452414 453454
rect 451794 453134 452414 453218
rect 451794 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 452414 453134
rect 451794 417454 452414 452898
rect 451794 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 452414 417454
rect 451794 417134 452414 417218
rect 451794 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 452414 417134
rect 451794 381454 452414 416898
rect 451794 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 452414 381454
rect 451794 381134 452414 381218
rect 451794 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 452414 381134
rect 451794 345454 452414 380898
rect 451794 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 452414 345454
rect 451794 345134 452414 345218
rect 451794 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 452414 345134
rect 451794 309454 452414 344898
rect 451794 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 452414 309454
rect 451794 309134 452414 309218
rect 451794 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 452414 309134
rect 451794 273454 452414 308898
rect 451794 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 452414 273454
rect 451794 273134 452414 273218
rect 451794 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 452414 273134
rect 451794 237454 452414 272898
rect 451794 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 452414 237454
rect 451794 237134 452414 237218
rect 451794 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 452414 237134
rect 451794 201454 452414 236898
rect 451794 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 452414 201454
rect 451794 201134 452414 201218
rect 451794 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 452414 201134
rect 451794 165454 452414 200898
rect 451794 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 452414 165454
rect 451794 165134 452414 165218
rect 451794 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 452414 165134
rect 451794 129454 452414 164898
rect 451794 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 452414 129454
rect 451794 129134 452414 129218
rect 451794 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 452414 129134
rect 451794 93454 452414 128898
rect 451794 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 452414 93454
rect 451794 93134 452414 93218
rect 451794 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 452414 93134
rect 451794 57454 452414 92898
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -1306 452414 20898
rect 451794 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 452414 -1306
rect 451794 -1626 452414 -1542
rect 451794 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 452414 -1626
rect 451794 -1894 452414 -1862
rect 455514 673174 456134 707162
rect 455514 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 456134 673174
rect 455514 672854 456134 672938
rect 455514 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 456134 672854
rect 455514 637174 456134 672618
rect 455514 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 456134 637174
rect 455514 636854 456134 636938
rect 455514 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 456134 636854
rect 455514 601174 456134 636618
rect 455514 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 456134 601174
rect 455514 600854 456134 600938
rect 455514 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 456134 600854
rect 455514 565174 456134 600618
rect 455514 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 456134 565174
rect 455514 564854 456134 564938
rect 455514 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 456134 564854
rect 455514 529174 456134 564618
rect 455514 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 456134 529174
rect 455514 528854 456134 528938
rect 455514 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 456134 528854
rect 455514 493174 456134 528618
rect 455514 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 456134 493174
rect 455514 492854 456134 492938
rect 455514 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 456134 492854
rect 455514 457174 456134 492618
rect 455514 456938 455546 457174
rect 455782 456938 455866 457174
rect 456102 456938 456134 457174
rect 455514 456854 456134 456938
rect 455514 456618 455546 456854
rect 455782 456618 455866 456854
rect 456102 456618 456134 456854
rect 455514 421174 456134 456618
rect 455514 420938 455546 421174
rect 455782 420938 455866 421174
rect 456102 420938 456134 421174
rect 455514 420854 456134 420938
rect 455514 420618 455546 420854
rect 455782 420618 455866 420854
rect 456102 420618 456134 420854
rect 455514 385174 456134 420618
rect 455514 384938 455546 385174
rect 455782 384938 455866 385174
rect 456102 384938 456134 385174
rect 455514 384854 456134 384938
rect 455514 384618 455546 384854
rect 455782 384618 455866 384854
rect 456102 384618 456134 384854
rect 455514 349174 456134 384618
rect 455514 348938 455546 349174
rect 455782 348938 455866 349174
rect 456102 348938 456134 349174
rect 455514 348854 456134 348938
rect 455514 348618 455546 348854
rect 455782 348618 455866 348854
rect 456102 348618 456134 348854
rect 455514 313174 456134 348618
rect 455514 312938 455546 313174
rect 455782 312938 455866 313174
rect 456102 312938 456134 313174
rect 455514 312854 456134 312938
rect 455514 312618 455546 312854
rect 455782 312618 455866 312854
rect 456102 312618 456134 312854
rect 455514 277174 456134 312618
rect 455514 276938 455546 277174
rect 455782 276938 455866 277174
rect 456102 276938 456134 277174
rect 455514 276854 456134 276938
rect 455514 276618 455546 276854
rect 455782 276618 455866 276854
rect 456102 276618 456134 276854
rect 455514 241174 456134 276618
rect 455514 240938 455546 241174
rect 455782 240938 455866 241174
rect 456102 240938 456134 241174
rect 455514 240854 456134 240938
rect 455514 240618 455546 240854
rect 455782 240618 455866 240854
rect 456102 240618 456134 240854
rect 455514 205174 456134 240618
rect 455514 204938 455546 205174
rect 455782 204938 455866 205174
rect 456102 204938 456134 205174
rect 455514 204854 456134 204938
rect 455514 204618 455546 204854
rect 455782 204618 455866 204854
rect 456102 204618 456134 204854
rect 455514 169174 456134 204618
rect 455514 168938 455546 169174
rect 455782 168938 455866 169174
rect 456102 168938 456134 169174
rect 455514 168854 456134 168938
rect 455514 168618 455546 168854
rect 455782 168618 455866 168854
rect 456102 168618 456134 168854
rect 455514 133174 456134 168618
rect 455514 132938 455546 133174
rect 455782 132938 455866 133174
rect 456102 132938 456134 133174
rect 455514 132854 456134 132938
rect 455514 132618 455546 132854
rect 455782 132618 455866 132854
rect 456102 132618 456134 132854
rect 455514 97174 456134 132618
rect 455514 96938 455546 97174
rect 455782 96938 455866 97174
rect 456102 96938 456134 97174
rect 455514 96854 456134 96938
rect 455514 96618 455546 96854
rect 455782 96618 455866 96854
rect 456102 96618 456134 96854
rect 455514 61174 456134 96618
rect 455514 60938 455546 61174
rect 455782 60938 455866 61174
rect 456102 60938 456134 61174
rect 455514 60854 456134 60938
rect 455514 60618 455546 60854
rect 455782 60618 455866 60854
rect 456102 60618 456134 60854
rect 455514 25174 456134 60618
rect 455514 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 456134 25174
rect 455514 24854 456134 24938
rect 455514 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 456134 24854
rect 455514 -3226 456134 24618
rect 455514 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 456134 -3226
rect 455514 -3546 456134 -3462
rect 455514 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 456134 -3546
rect 455514 -3814 456134 -3782
rect 459234 676894 459854 709082
rect 459234 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 459854 676894
rect 459234 676574 459854 676658
rect 459234 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 459854 676574
rect 459234 640894 459854 676338
rect 459234 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 459854 640894
rect 459234 640574 459854 640658
rect 459234 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 459854 640574
rect 459234 604894 459854 640338
rect 459234 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 459854 604894
rect 459234 604574 459854 604658
rect 459234 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 459854 604574
rect 459234 568894 459854 604338
rect 459234 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 459854 568894
rect 459234 568574 459854 568658
rect 459234 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 459854 568574
rect 459234 532894 459854 568338
rect 459234 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 459854 532894
rect 459234 532574 459854 532658
rect 459234 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 459854 532574
rect 459234 496894 459854 532338
rect 459234 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 459854 496894
rect 459234 496574 459854 496658
rect 459234 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 459854 496574
rect 459234 460894 459854 496338
rect 459234 460658 459266 460894
rect 459502 460658 459586 460894
rect 459822 460658 459854 460894
rect 459234 460574 459854 460658
rect 459234 460338 459266 460574
rect 459502 460338 459586 460574
rect 459822 460338 459854 460574
rect 459234 424894 459854 460338
rect 459234 424658 459266 424894
rect 459502 424658 459586 424894
rect 459822 424658 459854 424894
rect 459234 424574 459854 424658
rect 459234 424338 459266 424574
rect 459502 424338 459586 424574
rect 459822 424338 459854 424574
rect 459234 388894 459854 424338
rect 459234 388658 459266 388894
rect 459502 388658 459586 388894
rect 459822 388658 459854 388894
rect 459234 388574 459854 388658
rect 459234 388338 459266 388574
rect 459502 388338 459586 388574
rect 459822 388338 459854 388574
rect 459234 352894 459854 388338
rect 459234 352658 459266 352894
rect 459502 352658 459586 352894
rect 459822 352658 459854 352894
rect 459234 352574 459854 352658
rect 459234 352338 459266 352574
rect 459502 352338 459586 352574
rect 459822 352338 459854 352574
rect 459234 316894 459854 352338
rect 459234 316658 459266 316894
rect 459502 316658 459586 316894
rect 459822 316658 459854 316894
rect 459234 316574 459854 316658
rect 459234 316338 459266 316574
rect 459502 316338 459586 316574
rect 459822 316338 459854 316574
rect 459234 280894 459854 316338
rect 459234 280658 459266 280894
rect 459502 280658 459586 280894
rect 459822 280658 459854 280894
rect 459234 280574 459854 280658
rect 459234 280338 459266 280574
rect 459502 280338 459586 280574
rect 459822 280338 459854 280574
rect 459234 244894 459854 280338
rect 459234 244658 459266 244894
rect 459502 244658 459586 244894
rect 459822 244658 459854 244894
rect 459234 244574 459854 244658
rect 459234 244338 459266 244574
rect 459502 244338 459586 244574
rect 459822 244338 459854 244574
rect 459234 208894 459854 244338
rect 459234 208658 459266 208894
rect 459502 208658 459586 208894
rect 459822 208658 459854 208894
rect 459234 208574 459854 208658
rect 459234 208338 459266 208574
rect 459502 208338 459586 208574
rect 459822 208338 459854 208574
rect 459234 172894 459854 208338
rect 459234 172658 459266 172894
rect 459502 172658 459586 172894
rect 459822 172658 459854 172894
rect 459234 172574 459854 172658
rect 459234 172338 459266 172574
rect 459502 172338 459586 172574
rect 459822 172338 459854 172574
rect 459234 136894 459854 172338
rect 459234 136658 459266 136894
rect 459502 136658 459586 136894
rect 459822 136658 459854 136894
rect 459234 136574 459854 136658
rect 459234 136338 459266 136574
rect 459502 136338 459586 136574
rect 459822 136338 459854 136574
rect 459234 100894 459854 136338
rect 459234 100658 459266 100894
rect 459502 100658 459586 100894
rect 459822 100658 459854 100894
rect 459234 100574 459854 100658
rect 459234 100338 459266 100574
rect 459502 100338 459586 100574
rect 459822 100338 459854 100574
rect 459234 64894 459854 100338
rect 459234 64658 459266 64894
rect 459502 64658 459586 64894
rect 459822 64658 459854 64894
rect 459234 64574 459854 64658
rect 459234 64338 459266 64574
rect 459502 64338 459586 64574
rect 459822 64338 459854 64574
rect 459234 28894 459854 64338
rect 459234 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 459854 28894
rect 459234 28574 459854 28658
rect 459234 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 459854 28574
rect 459234 -5146 459854 28338
rect 459234 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 459854 -5146
rect 459234 -5466 459854 -5382
rect 459234 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 459854 -5466
rect 459234 -5734 459854 -5702
rect 462954 680614 463574 711002
rect 480954 710598 481574 711590
rect 480954 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 481574 710598
rect 480954 710278 481574 710362
rect 480954 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 481574 710278
rect 477234 708678 477854 709670
rect 477234 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 477854 708678
rect 477234 708358 477854 708442
rect 477234 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 477854 708358
rect 473514 706758 474134 707750
rect 473514 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 474134 706758
rect 473514 706438 474134 706522
rect 473514 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 474134 706438
rect 462954 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 463574 680614
rect 462954 680294 463574 680378
rect 462954 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 463574 680294
rect 462954 644614 463574 680058
rect 462954 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 463574 644614
rect 462954 644294 463574 644378
rect 462954 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 463574 644294
rect 462954 608614 463574 644058
rect 462954 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 463574 608614
rect 462954 608294 463574 608378
rect 462954 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 463574 608294
rect 462954 572614 463574 608058
rect 462954 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 463574 572614
rect 462954 572294 463574 572378
rect 462954 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 463574 572294
rect 462954 536614 463574 572058
rect 462954 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 463574 536614
rect 462954 536294 463574 536378
rect 462954 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 463574 536294
rect 462954 500614 463574 536058
rect 462954 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 463574 500614
rect 462954 500294 463574 500378
rect 462954 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 463574 500294
rect 462954 464614 463574 500058
rect 462954 464378 462986 464614
rect 463222 464378 463306 464614
rect 463542 464378 463574 464614
rect 462954 464294 463574 464378
rect 462954 464058 462986 464294
rect 463222 464058 463306 464294
rect 463542 464058 463574 464294
rect 462954 428614 463574 464058
rect 462954 428378 462986 428614
rect 463222 428378 463306 428614
rect 463542 428378 463574 428614
rect 462954 428294 463574 428378
rect 462954 428058 462986 428294
rect 463222 428058 463306 428294
rect 463542 428058 463574 428294
rect 462954 392614 463574 428058
rect 462954 392378 462986 392614
rect 463222 392378 463306 392614
rect 463542 392378 463574 392614
rect 462954 392294 463574 392378
rect 462954 392058 462986 392294
rect 463222 392058 463306 392294
rect 463542 392058 463574 392294
rect 462954 356614 463574 392058
rect 462954 356378 462986 356614
rect 463222 356378 463306 356614
rect 463542 356378 463574 356614
rect 462954 356294 463574 356378
rect 462954 356058 462986 356294
rect 463222 356058 463306 356294
rect 463542 356058 463574 356294
rect 462954 320614 463574 356058
rect 462954 320378 462986 320614
rect 463222 320378 463306 320614
rect 463542 320378 463574 320614
rect 462954 320294 463574 320378
rect 462954 320058 462986 320294
rect 463222 320058 463306 320294
rect 463542 320058 463574 320294
rect 462954 284614 463574 320058
rect 462954 284378 462986 284614
rect 463222 284378 463306 284614
rect 463542 284378 463574 284614
rect 462954 284294 463574 284378
rect 462954 284058 462986 284294
rect 463222 284058 463306 284294
rect 463542 284058 463574 284294
rect 462954 248614 463574 284058
rect 462954 248378 462986 248614
rect 463222 248378 463306 248614
rect 463542 248378 463574 248614
rect 462954 248294 463574 248378
rect 462954 248058 462986 248294
rect 463222 248058 463306 248294
rect 463542 248058 463574 248294
rect 462954 212614 463574 248058
rect 462954 212378 462986 212614
rect 463222 212378 463306 212614
rect 463542 212378 463574 212614
rect 462954 212294 463574 212378
rect 462954 212058 462986 212294
rect 463222 212058 463306 212294
rect 463542 212058 463574 212294
rect 462954 176614 463574 212058
rect 462954 176378 462986 176614
rect 463222 176378 463306 176614
rect 463542 176378 463574 176614
rect 462954 176294 463574 176378
rect 462954 176058 462986 176294
rect 463222 176058 463306 176294
rect 463542 176058 463574 176294
rect 462954 140614 463574 176058
rect 462954 140378 462986 140614
rect 463222 140378 463306 140614
rect 463542 140378 463574 140614
rect 462954 140294 463574 140378
rect 462954 140058 462986 140294
rect 463222 140058 463306 140294
rect 463542 140058 463574 140294
rect 462954 104614 463574 140058
rect 462954 104378 462986 104614
rect 463222 104378 463306 104614
rect 463542 104378 463574 104614
rect 462954 104294 463574 104378
rect 462954 104058 462986 104294
rect 463222 104058 463306 104294
rect 463542 104058 463574 104294
rect 462954 68614 463574 104058
rect 462954 68378 462986 68614
rect 463222 68378 463306 68614
rect 463542 68378 463574 68614
rect 462954 68294 463574 68378
rect 462954 68058 462986 68294
rect 463222 68058 463306 68294
rect 463542 68058 463574 68294
rect 462954 32614 463574 68058
rect 462954 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 463574 32614
rect 462954 32294 463574 32378
rect 462954 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 463574 32294
rect 444954 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 445574 -6106
rect 444954 -6426 445574 -6342
rect 444954 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 445574 -6426
rect 444954 -7654 445574 -6662
rect 462954 -7066 463574 32058
rect 469794 704838 470414 705830
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 579454 470414 614898
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 399454 470414 434898
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 469794 363454 470414 398898
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 469794 327454 470414 362898
rect 469794 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 470414 327454
rect 469794 327134 470414 327218
rect 469794 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 470414 327134
rect 469794 291454 470414 326898
rect 469794 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 470414 291454
rect 469794 291134 470414 291218
rect 469794 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 470414 291134
rect 469794 255454 470414 290898
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 219454 470414 254898
rect 469794 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 470414 219454
rect 469794 219134 470414 219218
rect 469794 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 470414 219134
rect 469794 183454 470414 218898
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 147454 470414 182898
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 111454 470414 146898
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -1894 470414 -902
rect 473514 691174 474134 706202
rect 473514 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 474134 691174
rect 473514 690854 474134 690938
rect 473514 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 474134 690854
rect 473514 655174 474134 690618
rect 473514 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 474134 655174
rect 473514 654854 474134 654938
rect 473514 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 474134 654854
rect 473514 619174 474134 654618
rect 473514 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 474134 619174
rect 473514 618854 474134 618938
rect 473514 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 474134 618854
rect 473514 583174 474134 618618
rect 473514 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 474134 583174
rect 473514 582854 474134 582938
rect 473514 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 474134 582854
rect 473514 547174 474134 582618
rect 473514 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 474134 547174
rect 473514 546854 474134 546938
rect 473514 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 474134 546854
rect 473514 511174 474134 546618
rect 473514 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 474134 511174
rect 473514 510854 474134 510938
rect 473514 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 474134 510854
rect 473514 475174 474134 510618
rect 473514 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 474134 475174
rect 473514 474854 474134 474938
rect 473514 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 474134 474854
rect 473514 439174 474134 474618
rect 473514 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 474134 439174
rect 473514 438854 474134 438938
rect 473514 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 474134 438854
rect 473514 403174 474134 438618
rect 473514 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 474134 403174
rect 473514 402854 474134 402938
rect 473514 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 474134 402854
rect 473514 367174 474134 402618
rect 473514 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 474134 367174
rect 473514 366854 474134 366938
rect 473514 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 474134 366854
rect 473514 331174 474134 366618
rect 473514 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 474134 331174
rect 473514 330854 474134 330938
rect 473514 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 474134 330854
rect 473514 295174 474134 330618
rect 473514 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 474134 295174
rect 473514 294854 474134 294938
rect 473514 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 474134 294854
rect 473514 259174 474134 294618
rect 473514 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 474134 259174
rect 473514 258854 474134 258938
rect 473514 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 474134 258854
rect 473514 223174 474134 258618
rect 473514 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 474134 223174
rect 473514 222854 474134 222938
rect 473514 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 474134 222854
rect 473514 187174 474134 222618
rect 473514 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 474134 187174
rect 473514 186854 474134 186938
rect 473514 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 474134 186854
rect 473514 151174 474134 186618
rect 473514 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 474134 151174
rect 473514 150854 474134 150938
rect 473514 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 474134 150854
rect 473514 115174 474134 150618
rect 473514 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 474134 115174
rect 473514 114854 474134 114938
rect 473514 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 474134 114854
rect 473514 79174 474134 114618
rect 473514 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 474134 79174
rect 473514 78854 474134 78938
rect 473514 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 474134 78854
rect 473514 43174 474134 78618
rect 473514 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 474134 43174
rect 473514 42854 474134 42938
rect 473514 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 474134 42854
rect 473514 7174 474134 42618
rect 473514 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 474134 7174
rect 473514 6854 474134 6938
rect 473514 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 474134 6854
rect 473514 -2266 474134 6618
rect 473514 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 474134 -2266
rect 473514 -2586 474134 -2502
rect 473514 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 474134 -2586
rect 473514 -3814 474134 -2822
rect 477234 694894 477854 708122
rect 477234 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 477854 694894
rect 477234 694574 477854 694658
rect 477234 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 477854 694574
rect 477234 658894 477854 694338
rect 477234 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 477854 658894
rect 477234 658574 477854 658658
rect 477234 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 477854 658574
rect 477234 622894 477854 658338
rect 477234 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 477854 622894
rect 477234 622574 477854 622658
rect 477234 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 477854 622574
rect 477234 586894 477854 622338
rect 477234 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 477854 586894
rect 477234 586574 477854 586658
rect 477234 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 477854 586574
rect 477234 550894 477854 586338
rect 477234 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 477854 550894
rect 477234 550574 477854 550658
rect 477234 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 477854 550574
rect 477234 514894 477854 550338
rect 477234 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 477854 514894
rect 477234 514574 477854 514658
rect 477234 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 477854 514574
rect 477234 478894 477854 514338
rect 477234 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 477854 478894
rect 477234 478574 477854 478658
rect 477234 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 477854 478574
rect 477234 442894 477854 478338
rect 477234 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 477854 442894
rect 477234 442574 477854 442658
rect 477234 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 477854 442574
rect 477234 406894 477854 442338
rect 477234 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 477854 406894
rect 477234 406574 477854 406658
rect 477234 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 477854 406574
rect 477234 370894 477854 406338
rect 477234 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 477854 370894
rect 477234 370574 477854 370658
rect 477234 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 477854 370574
rect 477234 334894 477854 370338
rect 477234 334658 477266 334894
rect 477502 334658 477586 334894
rect 477822 334658 477854 334894
rect 477234 334574 477854 334658
rect 477234 334338 477266 334574
rect 477502 334338 477586 334574
rect 477822 334338 477854 334574
rect 477234 298894 477854 334338
rect 477234 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 477854 298894
rect 477234 298574 477854 298658
rect 477234 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 477854 298574
rect 477234 262894 477854 298338
rect 477234 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 477854 262894
rect 477234 262574 477854 262658
rect 477234 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 477854 262574
rect 477234 226894 477854 262338
rect 477234 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 477854 226894
rect 477234 226574 477854 226658
rect 477234 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 477854 226574
rect 477234 190894 477854 226338
rect 477234 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 477854 190894
rect 477234 190574 477854 190658
rect 477234 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 477854 190574
rect 477234 154894 477854 190338
rect 477234 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 477854 154894
rect 477234 154574 477854 154658
rect 477234 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 477854 154574
rect 477234 118894 477854 154338
rect 477234 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 477854 118894
rect 477234 118574 477854 118658
rect 477234 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 477854 118574
rect 477234 82894 477854 118338
rect 477234 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 477854 82894
rect 477234 82574 477854 82658
rect 477234 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 477854 82574
rect 477234 46894 477854 82338
rect 477234 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 477854 46894
rect 477234 46574 477854 46658
rect 477234 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 477854 46574
rect 477234 10894 477854 46338
rect 477234 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 477854 10894
rect 477234 10574 477854 10658
rect 477234 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 477854 10574
rect 477234 -4186 477854 10338
rect 477234 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 477854 -4186
rect 477234 -4506 477854 -4422
rect 477234 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 477854 -4506
rect 477234 -5734 477854 -4742
rect 480954 698614 481574 710042
rect 498954 711558 499574 711590
rect 498954 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 499574 711558
rect 498954 711238 499574 711322
rect 498954 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 499574 711238
rect 495234 709638 495854 709670
rect 495234 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 495854 709638
rect 495234 709318 495854 709402
rect 495234 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 495854 709318
rect 491514 707718 492134 707750
rect 491514 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 492134 707718
rect 491514 707398 492134 707482
rect 491514 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 492134 707398
rect 480954 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 481574 698614
rect 480954 698294 481574 698378
rect 480954 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 481574 698294
rect 480954 662614 481574 698058
rect 480954 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 481574 662614
rect 480954 662294 481574 662378
rect 480954 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 481574 662294
rect 480954 626614 481574 662058
rect 480954 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 481574 626614
rect 480954 626294 481574 626378
rect 480954 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 481574 626294
rect 480954 590614 481574 626058
rect 480954 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 481574 590614
rect 480954 590294 481574 590378
rect 480954 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 481574 590294
rect 480954 554614 481574 590058
rect 480954 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 481574 554614
rect 480954 554294 481574 554378
rect 480954 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 481574 554294
rect 480954 518614 481574 554058
rect 480954 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 481574 518614
rect 480954 518294 481574 518378
rect 480954 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 481574 518294
rect 480954 482614 481574 518058
rect 480954 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 481574 482614
rect 480954 482294 481574 482378
rect 480954 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 481574 482294
rect 480954 446614 481574 482058
rect 480954 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 481574 446614
rect 480954 446294 481574 446378
rect 480954 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 481574 446294
rect 480954 410614 481574 446058
rect 480954 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 481574 410614
rect 480954 410294 481574 410378
rect 480954 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 481574 410294
rect 480954 374614 481574 410058
rect 480954 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 481574 374614
rect 480954 374294 481574 374378
rect 480954 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 481574 374294
rect 480954 338614 481574 374058
rect 480954 338378 480986 338614
rect 481222 338378 481306 338614
rect 481542 338378 481574 338614
rect 480954 338294 481574 338378
rect 480954 338058 480986 338294
rect 481222 338058 481306 338294
rect 481542 338058 481574 338294
rect 480954 302614 481574 338058
rect 480954 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 481574 302614
rect 480954 302294 481574 302378
rect 480954 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 481574 302294
rect 480954 266614 481574 302058
rect 480954 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 481574 266614
rect 480954 266294 481574 266378
rect 480954 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 481574 266294
rect 480954 230614 481574 266058
rect 480954 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 481574 230614
rect 480954 230294 481574 230378
rect 480954 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 481574 230294
rect 480954 194614 481574 230058
rect 480954 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 481574 194614
rect 480954 194294 481574 194378
rect 480954 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 481574 194294
rect 480954 158614 481574 194058
rect 480954 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 481574 158614
rect 480954 158294 481574 158378
rect 480954 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 481574 158294
rect 480954 122614 481574 158058
rect 480954 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 481574 122614
rect 480954 122294 481574 122378
rect 480954 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 481574 122294
rect 480954 86614 481574 122058
rect 480954 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 481574 86614
rect 480954 86294 481574 86378
rect 480954 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 481574 86294
rect 480954 50614 481574 86058
rect 480954 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 481574 50614
rect 480954 50294 481574 50378
rect 480954 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 481574 50294
rect 480954 14614 481574 50058
rect 480954 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 481574 14614
rect 480954 14294 481574 14378
rect 480954 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 481574 14294
rect 462954 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 463574 -7066
rect 462954 -7386 463574 -7302
rect 462954 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 463574 -7386
rect 462954 -7654 463574 -7622
rect 480954 -6106 481574 14058
rect 487794 705798 488414 705830
rect 487794 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 488414 705798
rect 487794 705478 488414 705562
rect 487794 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 488414 705478
rect 487794 669454 488414 705242
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 633454 488414 668898
rect 487794 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 488414 633454
rect 487794 633134 488414 633218
rect 487794 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 488414 633134
rect 487794 597454 488414 632898
rect 487794 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 488414 597454
rect 487794 597134 488414 597218
rect 487794 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 488414 597134
rect 487794 561454 488414 596898
rect 487794 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 488414 561454
rect 487794 561134 488414 561218
rect 487794 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 488414 561134
rect 487794 525454 488414 560898
rect 487794 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 488414 525454
rect 487794 525134 488414 525218
rect 487794 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 488414 525134
rect 487794 489454 488414 524898
rect 487794 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 488414 489454
rect 487794 489134 488414 489218
rect 487794 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 488414 489134
rect 487794 453454 488414 488898
rect 487794 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 488414 453454
rect 487794 453134 488414 453218
rect 487794 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 488414 453134
rect 487794 417454 488414 452898
rect 487794 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 488414 417454
rect 487794 417134 488414 417218
rect 487794 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 488414 417134
rect 487794 381454 488414 416898
rect 487794 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 488414 381454
rect 487794 381134 488414 381218
rect 487794 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 488414 381134
rect 487794 345454 488414 380898
rect 487794 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 488414 345454
rect 487794 345134 488414 345218
rect 487794 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 488414 345134
rect 487794 309454 488414 344898
rect 487794 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 488414 309454
rect 487794 309134 488414 309218
rect 487794 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 488414 309134
rect 487794 273454 488414 308898
rect 487794 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 488414 273454
rect 487794 273134 488414 273218
rect 487794 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 488414 273134
rect 487794 237454 488414 272898
rect 487794 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 488414 237454
rect 487794 237134 488414 237218
rect 487794 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 488414 237134
rect 487794 201454 488414 236898
rect 487794 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 488414 201454
rect 487794 201134 488414 201218
rect 487794 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 488414 201134
rect 487794 165454 488414 200898
rect 487794 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 488414 165454
rect 487794 165134 488414 165218
rect 487794 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 488414 165134
rect 487794 129454 488414 164898
rect 487794 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 488414 129454
rect 487794 129134 488414 129218
rect 487794 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 488414 129134
rect 487794 93454 488414 128898
rect 487794 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 488414 93454
rect 487794 93134 488414 93218
rect 487794 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 488414 93134
rect 487794 57454 488414 92898
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -1306 488414 20898
rect 487794 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 488414 -1306
rect 487794 -1626 488414 -1542
rect 487794 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 488414 -1626
rect 487794 -1894 488414 -1862
rect 491514 673174 492134 707162
rect 491514 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 492134 673174
rect 491514 672854 492134 672938
rect 491514 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 492134 672854
rect 491514 637174 492134 672618
rect 491514 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 492134 637174
rect 491514 636854 492134 636938
rect 491514 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 492134 636854
rect 491514 601174 492134 636618
rect 491514 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 492134 601174
rect 491514 600854 492134 600938
rect 491514 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 492134 600854
rect 491514 565174 492134 600618
rect 491514 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 492134 565174
rect 491514 564854 492134 564938
rect 491514 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 492134 564854
rect 491514 529174 492134 564618
rect 491514 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 492134 529174
rect 491514 528854 492134 528938
rect 491514 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 492134 528854
rect 491514 493174 492134 528618
rect 491514 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 492134 493174
rect 491514 492854 492134 492938
rect 491514 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 492134 492854
rect 491514 457174 492134 492618
rect 491514 456938 491546 457174
rect 491782 456938 491866 457174
rect 492102 456938 492134 457174
rect 491514 456854 492134 456938
rect 491514 456618 491546 456854
rect 491782 456618 491866 456854
rect 492102 456618 492134 456854
rect 491514 421174 492134 456618
rect 491514 420938 491546 421174
rect 491782 420938 491866 421174
rect 492102 420938 492134 421174
rect 491514 420854 492134 420938
rect 491514 420618 491546 420854
rect 491782 420618 491866 420854
rect 492102 420618 492134 420854
rect 491514 385174 492134 420618
rect 491514 384938 491546 385174
rect 491782 384938 491866 385174
rect 492102 384938 492134 385174
rect 491514 384854 492134 384938
rect 491514 384618 491546 384854
rect 491782 384618 491866 384854
rect 492102 384618 492134 384854
rect 491514 349174 492134 384618
rect 491514 348938 491546 349174
rect 491782 348938 491866 349174
rect 492102 348938 492134 349174
rect 491514 348854 492134 348938
rect 491514 348618 491546 348854
rect 491782 348618 491866 348854
rect 492102 348618 492134 348854
rect 491514 313174 492134 348618
rect 491514 312938 491546 313174
rect 491782 312938 491866 313174
rect 492102 312938 492134 313174
rect 491514 312854 492134 312938
rect 491514 312618 491546 312854
rect 491782 312618 491866 312854
rect 492102 312618 492134 312854
rect 491514 277174 492134 312618
rect 491514 276938 491546 277174
rect 491782 276938 491866 277174
rect 492102 276938 492134 277174
rect 491514 276854 492134 276938
rect 491514 276618 491546 276854
rect 491782 276618 491866 276854
rect 492102 276618 492134 276854
rect 491514 241174 492134 276618
rect 491514 240938 491546 241174
rect 491782 240938 491866 241174
rect 492102 240938 492134 241174
rect 491514 240854 492134 240938
rect 491514 240618 491546 240854
rect 491782 240618 491866 240854
rect 492102 240618 492134 240854
rect 491514 205174 492134 240618
rect 491514 204938 491546 205174
rect 491782 204938 491866 205174
rect 492102 204938 492134 205174
rect 491514 204854 492134 204938
rect 491514 204618 491546 204854
rect 491782 204618 491866 204854
rect 492102 204618 492134 204854
rect 491514 169174 492134 204618
rect 491514 168938 491546 169174
rect 491782 168938 491866 169174
rect 492102 168938 492134 169174
rect 491514 168854 492134 168938
rect 491514 168618 491546 168854
rect 491782 168618 491866 168854
rect 492102 168618 492134 168854
rect 491514 133174 492134 168618
rect 491514 132938 491546 133174
rect 491782 132938 491866 133174
rect 492102 132938 492134 133174
rect 491514 132854 492134 132938
rect 491514 132618 491546 132854
rect 491782 132618 491866 132854
rect 492102 132618 492134 132854
rect 491514 97174 492134 132618
rect 491514 96938 491546 97174
rect 491782 96938 491866 97174
rect 492102 96938 492134 97174
rect 491514 96854 492134 96938
rect 491514 96618 491546 96854
rect 491782 96618 491866 96854
rect 492102 96618 492134 96854
rect 491514 61174 492134 96618
rect 491514 60938 491546 61174
rect 491782 60938 491866 61174
rect 492102 60938 492134 61174
rect 491514 60854 492134 60938
rect 491514 60618 491546 60854
rect 491782 60618 491866 60854
rect 492102 60618 492134 60854
rect 491514 25174 492134 60618
rect 491514 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 492134 25174
rect 491514 24854 492134 24938
rect 491514 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 492134 24854
rect 491514 -3226 492134 24618
rect 491514 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 492134 -3226
rect 491514 -3546 492134 -3462
rect 491514 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 492134 -3546
rect 491514 -3814 492134 -3782
rect 495234 676894 495854 709082
rect 495234 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 495854 676894
rect 495234 676574 495854 676658
rect 495234 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 495854 676574
rect 495234 640894 495854 676338
rect 495234 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 495854 640894
rect 495234 640574 495854 640658
rect 495234 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 495854 640574
rect 495234 604894 495854 640338
rect 495234 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 495854 604894
rect 495234 604574 495854 604658
rect 495234 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 495854 604574
rect 495234 568894 495854 604338
rect 495234 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 495854 568894
rect 495234 568574 495854 568658
rect 495234 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 495854 568574
rect 495234 532894 495854 568338
rect 495234 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 495854 532894
rect 495234 532574 495854 532658
rect 495234 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 495854 532574
rect 495234 496894 495854 532338
rect 495234 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 495854 496894
rect 495234 496574 495854 496658
rect 495234 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 495854 496574
rect 495234 460894 495854 496338
rect 495234 460658 495266 460894
rect 495502 460658 495586 460894
rect 495822 460658 495854 460894
rect 495234 460574 495854 460658
rect 495234 460338 495266 460574
rect 495502 460338 495586 460574
rect 495822 460338 495854 460574
rect 495234 424894 495854 460338
rect 495234 424658 495266 424894
rect 495502 424658 495586 424894
rect 495822 424658 495854 424894
rect 495234 424574 495854 424658
rect 495234 424338 495266 424574
rect 495502 424338 495586 424574
rect 495822 424338 495854 424574
rect 495234 388894 495854 424338
rect 495234 388658 495266 388894
rect 495502 388658 495586 388894
rect 495822 388658 495854 388894
rect 495234 388574 495854 388658
rect 495234 388338 495266 388574
rect 495502 388338 495586 388574
rect 495822 388338 495854 388574
rect 495234 352894 495854 388338
rect 495234 352658 495266 352894
rect 495502 352658 495586 352894
rect 495822 352658 495854 352894
rect 495234 352574 495854 352658
rect 495234 352338 495266 352574
rect 495502 352338 495586 352574
rect 495822 352338 495854 352574
rect 495234 316894 495854 352338
rect 495234 316658 495266 316894
rect 495502 316658 495586 316894
rect 495822 316658 495854 316894
rect 495234 316574 495854 316658
rect 495234 316338 495266 316574
rect 495502 316338 495586 316574
rect 495822 316338 495854 316574
rect 495234 280894 495854 316338
rect 495234 280658 495266 280894
rect 495502 280658 495586 280894
rect 495822 280658 495854 280894
rect 495234 280574 495854 280658
rect 495234 280338 495266 280574
rect 495502 280338 495586 280574
rect 495822 280338 495854 280574
rect 495234 244894 495854 280338
rect 495234 244658 495266 244894
rect 495502 244658 495586 244894
rect 495822 244658 495854 244894
rect 495234 244574 495854 244658
rect 495234 244338 495266 244574
rect 495502 244338 495586 244574
rect 495822 244338 495854 244574
rect 495234 208894 495854 244338
rect 495234 208658 495266 208894
rect 495502 208658 495586 208894
rect 495822 208658 495854 208894
rect 495234 208574 495854 208658
rect 495234 208338 495266 208574
rect 495502 208338 495586 208574
rect 495822 208338 495854 208574
rect 495234 172894 495854 208338
rect 495234 172658 495266 172894
rect 495502 172658 495586 172894
rect 495822 172658 495854 172894
rect 495234 172574 495854 172658
rect 495234 172338 495266 172574
rect 495502 172338 495586 172574
rect 495822 172338 495854 172574
rect 495234 136894 495854 172338
rect 495234 136658 495266 136894
rect 495502 136658 495586 136894
rect 495822 136658 495854 136894
rect 495234 136574 495854 136658
rect 495234 136338 495266 136574
rect 495502 136338 495586 136574
rect 495822 136338 495854 136574
rect 495234 100894 495854 136338
rect 495234 100658 495266 100894
rect 495502 100658 495586 100894
rect 495822 100658 495854 100894
rect 495234 100574 495854 100658
rect 495234 100338 495266 100574
rect 495502 100338 495586 100574
rect 495822 100338 495854 100574
rect 495234 64894 495854 100338
rect 495234 64658 495266 64894
rect 495502 64658 495586 64894
rect 495822 64658 495854 64894
rect 495234 64574 495854 64658
rect 495234 64338 495266 64574
rect 495502 64338 495586 64574
rect 495822 64338 495854 64574
rect 495234 28894 495854 64338
rect 495234 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 495854 28894
rect 495234 28574 495854 28658
rect 495234 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 495854 28574
rect 495234 -5146 495854 28338
rect 495234 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 495854 -5146
rect 495234 -5466 495854 -5382
rect 495234 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 495854 -5466
rect 495234 -5734 495854 -5702
rect 498954 680614 499574 711002
rect 516954 710598 517574 711590
rect 516954 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 517574 710598
rect 516954 710278 517574 710362
rect 516954 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 517574 710278
rect 513234 708678 513854 709670
rect 513234 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 513854 708678
rect 513234 708358 513854 708442
rect 513234 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 513854 708358
rect 509514 706758 510134 707750
rect 509514 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 510134 706758
rect 509514 706438 510134 706522
rect 509514 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 510134 706438
rect 498954 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 499574 680614
rect 498954 680294 499574 680378
rect 498954 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 499574 680294
rect 498954 644614 499574 680058
rect 498954 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 499574 644614
rect 498954 644294 499574 644378
rect 498954 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 499574 644294
rect 498954 608614 499574 644058
rect 498954 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 499574 608614
rect 498954 608294 499574 608378
rect 498954 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 499574 608294
rect 498954 572614 499574 608058
rect 498954 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 499574 572614
rect 498954 572294 499574 572378
rect 498954 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 499574 572294
rect 498954 536614 499574 572058
rect 498954 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 499574 536614
rect 498954 536294 499574 536378
rect 498954 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 499574 536294
rect 498954 500614 499574 536058
rect 498954 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 499574 500614
rect 498954 500294 499574 500378
rect 498954 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 499574 500294
rect 498954 464614 499574 500058
rect 498954 464378 498986 464614
rect 499222 464378 499306 464614
rect 499542 464378 499574 464614
rect 498954 464294 499574 464378
rect 498954 464058 498986 464294
rect 499222 464058 499306 464294
rect 499542 464058 499574 464294
rect 498954 428614 499574 464058
rect 498954 428378 498986 428614
rect 499222 428378 499306 428614
rect 499542 428378 499574 428614
rect 498954 428294 499574 428378
rect 498954 428058 498986 428294
rect 499222 428058 499306 428294
rect 499542 428058 499574 428294
rect 498954 392614 499574 428058
rect 498954 392378 498986 392614
rect 499222 392378 499306 392614
rect 499542 392378 499574 392614
rect 498954 392294 499574 392378
rect 498954 392058 498986 392294
rect 499222 392058 499306 392294
rect 499542 392058 499574 392294
rect 498954 356614 499574 392058
rect 498954 356378 498986 356614
rect 499222 356378 499306 356614
rect 499542 356378 499574 356614
rect 498954 356294 499574 356378
rect 498954 356058 498986 356294
rect 499222 356058 499306 356294
rect 499542 356058 499574 356294
rect 498954 320614 499574 356058
rect 498954 320378 498986 320614
rect 499222 320378 499306 320614
rect 499542 320378 499574 320614
rect 498954 320294 499574 320378
rect 498954 320058 498986 320294
rect 499222 320058 499306 320294
rect 499542 320058 499574 320294
rect 498954 284614 499574 320058
rect 498954 284378 498986 284614
rect 499222 284378 499306 284614
rect 499542 284378 499574 284614
rect 498954 284294 499574 284378
rect 498954 284058 498986 284294
rect 499222 284058 499306 284294
rect 499542 284058 499574 284294
rect 498954 248614 499574 284058
rect 498954 248378 498986 248614
rect 499222 248378 499306 248614
rect 499542 248378 499574 248614
rect 498954 248294 499574 248378
rect 498954 248058 498986 248294
rect 499222 248058 499306 248294
rect 499542 248058 499574 248294
rect 498954 212614 499574 248058
rect 498954 212378 498986 212614
rect 499222 212378 499306 212614
rect 499542 212378 499574 212614
rect 498954 212294 499574 212378
rect 498954 212058 498986 212294
rect 499222 212058 499306 212294
rect 499542 212058 499574 212294
rect 498954 176614 499574 212058
rect 498954 176378 498986 176614
rect 499222 176378 499306 176614
rect 499542 176378 499574 176614
rect 498954 176294 499574 176378
rect 498954 176058 498986 176294
rect 499222 176058 499306 176294
rect 499542 176058 499574 176294
rect 498954 140614 499574 176058
rect 498954 140378 498986 140614
rect 499222 140378 499306 140614
rect 499542 140378 499574 140614
rect 498954 140294 499574 140378
rect 498954 140058 498986 140294
rect 499222 140058 499306 140294
rect 499542 140058 499574 140294
rect 498954 104614 499574 140058
rect 498954 104378 498986 104614
rect 499222 104378 499306 104614
rect 499542 104378 499574 104614
rect 498954 104294 499574 104378
rect 498954 104058 498986 104294
rect 499222 104058 499306 104294
rect 499542 104058 499574 104294
rect 498954 68614 499574 104058
rect 498954 68378 498986 68614
rect 499222 68378 499306 68614
rect 499542 68378 499574 68614
rect 498954 68294 499574 68378
rect 498954 68058 498986 68294
rect 499222 68058 499306 68294
rect 499542 68058 499574 68294
rect 498954 32614 499574 68058
rect 498954 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 499574 32614
rect 498954 32294 499574 32378
rect 498954 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 499574 32294
rect 480954 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 481574 -6106
rect 480954 -6426 481574 -6342
rect 480954 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 481574 -6426
rect 480954 -7654 481574 -6662
rect 498954 -7066 499574 32058
rect 505794 704838 506414 705830
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 505794 579454 506414 614898
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 291454 506414 326898
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 255454 506414 290898
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 219454 506414 254898
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 111454 506414 146898
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -1894 506414 -902
rect 509514 691174 510134 706202
rect 509514 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 510134 691174
rect 509514 690854 510134 690938
rect 509514 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 510134 690854
rect 509514 655174 510134 690618
rect 509514 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 510134 655174
rect 509514 654854 510134 654938
rect 509514 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 510134 654854
rect 509514 619174 510134 654618
rect 509514 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 510134 619174
rect 509514 618854 510134 618938
rect 509514 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 510134 618854
rect 509514 583174 510134 618618
rect 509514 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 510134 583174
rect 509514 582854 510134 582938
rect 509514 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 510134 582854
rect 509514 547174 510134 582618
rect 509514 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 510134 547174
rect 509514 546854 510134 546938
rect 509514 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 510134 546854
rect 509514 511174 510134 546618
rect 509514 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 510134 511174
rect 509514 510854 510134 510938
rect 509514 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 510134 510854
rect 509514 475174 510134 510618
rect 509514 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 510134 475174
rect 509514 474854 510134 474938
rect 509514 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 510134 474854
rect 509514 439174 510134 474618
rect 509514 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 510134 439174
rect 509514 438854 510134 438938
rect 509514 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 510134 438854
rect 509514 403174 510134 438618
rect 509514 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 510134 403174
rect 509514 402854 510134 402938
rect 509514 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 510134 402854
rect 509514 367174 510134 402618
rect 509514 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 510134 367174
rect 509514 366854 510134 366938
rect 509514 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 510134 366854
rect 509514 331174 510134 366618
rect 509514 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 510134 331174
rect 509514 330854 510134 330938
rect 509514 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 510134 330854
rect 509514 295174 510134 330618
rect 509514 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 510134 295174
rect 509514 294854 510134 294938
rect 509514 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 510134 294854
rect 509514 259174 510134 294618
rect 509514 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 510134 259174
rect 509514 258854 510134 258938
rect 509514 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 510134 258854
rect 509514 223174 510134 258618
rect 509514 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 510134 223174
rect 509514 222854 510134 222938
rect 509514 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 510134 222854
rect 509514 187174 510134 222618
rect 509514 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 510134 187174
rect 509514 186854 510134 186938
rect 509514 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 510134 186854
rect 509514 151174 510134 186618
rect 509514 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 510134 151174
rect 509514 150854 510134 150938
rect 509514 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 510134 150854
rect 509514 115174 510134 150618
rect 509514 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 510134 115174
rect 509514 114854 510134 114938
rect 509514 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 510134 114854
rect 509514 79174 510134 114618
rect 509514 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 510134 79174
rect 509514 78854 510134 78938
rect 509514 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 510134 78854
rect 509514 43174 510134 78618
rect 509514 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 510134 43174
rect 509514 42854 510134 42938
rect 509514 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 510134 42854
rect 509514 7174 510134 42618
rect 509514 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 510134 7174
rect 509514 6854 510134 6938
rect 509514 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 510134 6854
rect 509514 -2266 510134 6618
rect 509514 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 510134 -2266
rect 509514 -2586 510134 -2502
rect 509514 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 510134 -2586
rect 509514 -3814 510134 -2822
rect 513234 694894 513854 708122
rect 513234 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 513854 694894
rect 513234 694574 513854 694658
rect 513234 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 513854 694574
rect 513234 658894 513854 694338
rect 513234 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 513854 658894
rect 513234 658574 513854 658658
rect 513234 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 513854 658574
rect 513234 622894 513854 658338
rect 513234 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 513854 622894
rect 513234 622574 513854 622658
rect 513234 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 513854 622574
rect 513234 586894 513854 622338
rect 513234 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 513854 586894
rect 513234 586574 513854 586658
rect 513234 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 513854 586574
rect 513234 550894 513854 586338
rect 513234 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 513854 550894
rect 513234 550574 513854 550658
rect 513234 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 513854 550574
rect 513234 514894 513854 550338
rect 513234 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 513854 514894
rect 513234 514574 513854 514658
rect 513234 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 513854 514574
rect 513234 478894 513854 514338
rect 513234 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 513854 478894
rect 513234 478574 513854 478658
rect 513234 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 513854 478574
rect 513234 442894 513854 478338
rect 513234 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 513854 442894
rect 513234 442574 513854 442658
rect 513234 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 513854 442574
rect 513234 406894 513854 442338
rect 513234 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 513854 406894
rect 513234 406574 513854 406658
rect 513234 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 513854 406574
rect 513234 370894 513854 406338
rect 513234 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 513854 370894
rect 513234 370574 513854 370658
rect 513234 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 513854 370574
rect 513234 334894 513854 370338
rect 513234 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 513854 334894
rect 513234 334574 513854 334658
rect 513234 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 513854 334574
rect 513234 298894 513854 334338
rect 513234 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 513854 298894
rect 513234 298574 513854 298658
rect 513234 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 513854 298574
rect 513234 262894 513854 298338
rect 513234 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 513854 262894
rect 513234 262574 513854 262658
rect 513234 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 513854 262574
rect 513234 226894 513854 262338
rect 513234 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 513854 226894
rect 513234 226574 513854 226658
rect 513234 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 513854 226574
rect 513234 190894 513854 226338
rect 513234 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 513854 190894
rect 513234 190574 513854 190658
rect 513234 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 513854 190574
rect 513234 154894 513854 190338
rect 513234 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 513854 154894
rect 513234 154574 513854 154658
rect 513234 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 513854 154574
rect 513234 118894 513854 154338
rect 513234 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 513854 118894
rect 513234 118574 513854 118658
rect 513234 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 513854 118574
rect 513234 82894 513854 118338
rect 513234 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 513854 82894
rect 513234 82574 513854 82658
rect 513234 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 513854 82574
rect 513234 46894 513854 82338
rect 513234 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 513854 46894
rect 513234 46574 513854 46658
rect 513234 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 513854 46574
rect 513234 10894 513854 46338
rect 513234 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 513854 10894
rect 513234 10574 513854 10658
rect 513234 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 513854 10574
rect 513234 -4186 513854 10338
rect 513234 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 513854 -4186
rect 513234 -4506 513854 -4422
rect 513234 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 513854 -4506
rect 513234 -5734 513854 -4742
rect 516954 698614 517574 710042
rect 534954 711558 535574 711590
rect 534954 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 535574 711558
rect 534954 711238 535574 711322
rect 534954 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 535574 711238
rect 531234 709638 531854 709670
rect 531234 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 531854 709638
rect 531234 709318 531854 709402
rect 531234 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 531854 709318
rect 527514 707718 528134 707750
rect 527514 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 528134 707718
rect 527514 707398 528134 707482
rect 527514 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 528134 707398
rect 516954 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 517574 698614
rect 516954 698294 517574 698378
rect 516954 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 517574 698294
rect 516954 662614 517574 698058
rect 516954 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 517574 662614
rect 516954 662294 517574 662378
rect 516954 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 517574 662294
rect 516954 626614 517574 662058
rect 516954 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 517574 626614
rect 516954 626294 517574 626378
rect 516954 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 517574 626294
rect 516954 590614 517574 626058
rect 516954 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 517574 590614
rect 516954 590294 517574 590378
rect 516954 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 517574 590294
rect 516954 554614 517574 590058
rect 516954 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 517574 554614
rect 516954 554294 517574 554378
rect 516954 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 517574 554294
rect 516954 518614 517574 554058
rect 516954 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 517574 518614
rect 516954 518294 517574 518378
rect 516954 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 517574 518294
rect 516954 482614 517574 518058
rect 516954 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 517574 482614
rect 516954 482294 517574 482378
rect 516954 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 517574 482294
rect 516954 446614 517574 482058
rect 516954 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 517574 446614
rect 516954 446294 517574 446378
rect 516954 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 517574 446294
rect 516954 410614 517574 446058
rect 516954 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 517574 410614
rect 516954 410294 517574 410378
rect 516954 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 517574 410294
rect 516954 374614 517574 410058
rect 516954 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 517574 374614
rect 516954 374294 517574 374378
rect 516954 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 517574 374294
rect 516954 338614 517574 374058
rect 516954 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 517574 338614
rect 516954 338294 517574 338378
rect 516954 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 517574 338294
rect 516954 302614 517574 338058
rect 516954 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 517574 302614
rect 516954 302294 517574 302378
rect 516954 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 517574 302294
rect 516954 266614 517574 302058
rect 516954 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 517574 266614
rect 516954 266294 517574 266378
rect 516954 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 517574 266294
rect 516954 230614 517574 266058
rect 516954 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 517574 230614
rect 516954 230294 517574 230378
rect 516954 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 517574 230294
rect 516954 194614 517574 230058
rect 516954 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 517574 194614
rect 516954 194294 517574 194378
rect 516954 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 517574 194294
rect 516954 158614 517574 194058
rect 516954 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 517574 158614
rect 516954 158294 517574 158378
rect 516954 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 517574 158294
rect 516954 122614 517574 158058
rect 516954 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 517574 122614
rect 516954 122294 517574 122378
rect 516954 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 517574 122294
rect 516954 86614 517574 122058
rect 516954 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 517574 86614
rect 516954 86294 517574 86378
rect 516954 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 517574 86294
rect 516954 50614 517574 86058
rect 516954 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 517574 50614
rect 516954 50294 517574 50378
rect 516954 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 517574 50294
rect 516954 14614 517574 50058
rect 516954 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 517574 14614
rect 516954 14294 517574 14378
rect 516954 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 517574 14294
rect 498954 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 499574 -7066
rect 498954 -7386 499574 -7302
rect 498954 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 499574 -7386
rect 498954 -7654 499574 -7622
rect 516954 -6106 517574 14058
rect 523794 705798 524414 705830
rect 523794 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 524414 705798
rect 523794 705478 524414 705562
rect 523794 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 524414 705478
rect 523794 669454 524414 705242
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 523794 309454 524414 344898
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 523794 273454 524414 308898
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -1306 524414 20898
rect 523794 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 524414 -1306
rect 523794 -1626 524414 -1542
rect 523794 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 524414 -1626
rect 523794 -1894 524414 -1862
rect 527514 673174 528134 707162
rect 527514 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 528134 673174
rect 527514 672854 528134 672938
rect 527514 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 528134 672854
rect 527514 637174 528134 672618
rect 527514 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 528134 637174
rect 527514 636854 528134 636938
rect 527514 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 528134 636854
rect 527514 601174 528134 636618
rect 527514 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 528134 601174
rect 527514 600854 528134 600938
rect 527514 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 528134 600854
rect 527514 565174 528134 600618
rect 527514 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 528134 565174
rect 527514 564854 528134 564938
rect 527514 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 528134 564854
rect 527514 529174 528134 564618
rect 527514 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 528134 529174
rect 527514 528854 528134 528938
rect 527514 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 528134 528854
rect 527514 493174 528134 528618
rect 527514 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 528134 493174
rect 527514 492854 528134 492938
rect 527514 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 528134 492854
rect 527514 457174 528134 492618
rect 527514 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 528134 457174
rect 527514 456854 528134 456938
rect 527514 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 528134 456854
rect 527514 421174 528134 456618
rect 527514 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 528134 421174
rect 527514 420854 528134 420938
rect 527514 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 528134 420854
rect 527514 385174 528134 420618
rect 527514 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 528134 385174
rect 527514 384854 528134 384938
rect 527514 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 528134 384854
rect 527514 349174 528134 384618
rect 527514 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 528134 349174
rect 527514 348854 528134 348938
rect 527514 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 528134 348854
rect 527514 313174 528134 348618
rect 527514 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 528134 313174
rect 527514 312854 528134 312938
rect 527514 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 528134 312854
rect 527514 277174 528134 312618
rect 527514 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 528134 277174
rect 527514 276854 528134 276938
rect 527514 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 528134 276854
rect 527514 241174 528134 276618
rect 527514 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 528134 241174
rect 527514 240854 528134 240938
rect 527514 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 528134 240854
rect 527514 205174 528134 240618
rect 527514 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 528134 205174
rect 527514 204854 528134 204938
rect 527514 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 528134 204854
rect 527514 169174 528134 204618
rect 527514 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 528134 169174
rect 527514 168854 528134 168938
rect 527514 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 528134 168854
rect 527514 133174 528134 168618
rect 527514 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 528134 133174
rect 527514 132854 528134 132938
rect 527514 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 528134 132854
rect 527514 97174 528134 132618
rect 527514 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 528134 97174
rect 527514 96854 528134 96938
rect 527514 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 528134 96854
rect 527514 61174 528134 96618
rect 527514 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 528134 61174
rect 527514 60854 528134 60938
rect 527514 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 528134 60854
rect 527514 25174 528134 60618
rect 527514 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 528134 25174
rect 527514 24854 528134 24938
rect 527514 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 528134 24854
rect 527514 -3226 528134 24618
rect 527514 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 528134 -3226
rect 527514 -3546 528134 -3462
rect 527514 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 528134 -3546
rect 527514 -3814 528134 -3782
rect 531234 676894 531854 709082
rect 531234 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 531854 676894
rect 531234 676574 531854 676658
rect 531234 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 531854 676574
rect 531234 640894 531854 676338
rect 531234 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 531854 640894
rect 531234 640574 531854 640658
rect 531234 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 531854 640574
rect 531234 604894 531854 640338
rect 531234 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 531854 604894
rect 531234 604574 531854 604658
rect 531234 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 531854 604574
rect 531234 568894 531854 604338
rect 531234 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 531854 568894
rect 531234 568574 531854 568658
rect 531234 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 531854 568574
rect 531234 532894 531854 568338
rect 531234 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 531854 532894
rect 531234 532574 531854 532658
rect 531234 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 531854 532574
rect 531234 496894 531854 532338
rect 531234 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 531854 496894
rect 531234 496574 531854 496658
rect 531234 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 531854 496574
rect 531234 460894 531854 496338
rect 531234 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 531854 460894
rect 531234 460574 531854 460658
rect 531234 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 531854 460574
rect 531234 424894 531854 460338
rect 531234 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 531854 424894
rect 531234 424574 531854 424658
rect 531234 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 531854 424574
rect 531234 388894 531854 424338
rect 531234 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 531854 388894
rect 531234 388574 531854 388658
rect 531234 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 531854 388574
rect 531234 352894 531854 388338
rect 531234 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 531854 352894
rect 531234 352574 531854 352658
rect 531234 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 531854 352574
rect 531234 316894 531854 352338
rect 531234 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 531854 316894
rect 531234 316574 531854 316658
rect 531234 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 531854 316574
rect 531234 280894 531854 316338
rect 531234 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 531854 280894
rect 531234 280574 531854 280658
rect 531234 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 531854 280574
rect 531234 244894 531854 280338
rect 531234 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 531854 244894
rect 531234 244574 531854 244658
rect 531234 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 531854 244574
rect 531234 208894 531854 244338
rect 531234 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 531854 208894
rect 531234 208574 531854 208658
rect 531234 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 531854 208574
rect 531234 172894 531854 208338
rect 531234 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 531854 172894
rect 531234 172574 531854 172658
rect 531234 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 531854 172574
rect 531234 136894 531854 172338
rect 531234 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 531854 136894
rect 531234 136574 531854 136658
rect 531234 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 531854 136574
rect 531234 100894 531854 136338
rect 531234 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 531854 100894
rect 531234 100574 531854 100658
rect 531234 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 531854 100574
rect 531234 64894 531854 100338
rect 531234 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 531854 64894
rect 531234 64574 531854 64658
rect 531234 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 531854 64574
rect 531234 28894 531854 64338
rect 531234 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 531854 28894
rect 531234 28574 531854 28658
rect 531234 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 531854 28574
rect 531234 -5146 531854 28338
rect 531234 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 531854 -5146
rect 531234 -5466 531854 -5382
rect 531234 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 531854 -5466
rect 531234 -5734 531854 -5702
rect 534954 680614 535574 711002
rect 552954 710598 553574 711590
rect 552954 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 553574 710598
rect 552954 710278 553574 710362
rect 552954 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 553574 710278
rect 549234 708678 549854 709670
rect 549234 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 549854 708678
rect 549234 708358 549854 708442
rect 549234 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 549854 708358
rect 545514 706758 546134 707750
rect 545514 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 546134 706758
rect 545514 706438 546134 706522
rect 545514 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 546134 706438
rect 534954 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 535574 680614
rect 534954 680294 535574 680378
rect 534954 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 535574 680294
rect 534954 644614 535574 680058
rect 534954 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 535574 644614
rect 534954 644294 535574 644378
rect 534954 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 535574 644294
rect 534954 608614 535574 644058
rect 534954 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 535574 608614
rect 534954 608294 535574 608378
rect 534954 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 535574 608294
rect 534954 572614 535574 608058
rect 534954 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 535574 572614
rect 534954 572294 535574 572378
rect 534954 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 535574 572294
rect 534954 536614 535574 572058
rect 534954 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 535574 536614
rect 534954 536294 535574 536378
rect 534954 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 535574 536294
rect 534954 500614 535574 536058
rect 534954 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 535574 500614
rect 534954 500294 535574 500378
rect 534954 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 535574 500294
rect 534954 464614 535574 500058
rect 534954 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 535574 464614
rect 534954 464294 535574 464378
rect 534954 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 535574 464294
rect 534954 428614 535574 464058
rect 534954 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 535574 428614
rect 534954 428294 535574 428378
rect 534954 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 535574 428294
rect 534954 392614 535574 428058
rect 534954 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 535574 392614
rect 534954 392294 535574 392378
rect 534954 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 535574 392294
rect 534954 356614 535574 392058
rect 534954 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 535574 356614
rect 534954 356294 535574 356378
rect 534954 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 535574 356294
rect 534954 320614 535574 356058
rect 534954 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 535574 320614
rect 534954 320294 535574 320378
rect 534954 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 535574 320294
rect 534954 284614 535574 320058
rect 534954 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 535574 284614
rect 534954 284294 535574 284378
rect 534954 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 535574 284294
rect 534954 248614 535574 284058
rect 534954 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 535574 248614
rect 534954 248294 535574 248378
rect 534954 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 535574 248294
rect 534954 212614 535574 248058
rect 534954 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 535574 212614
rect 534954 212294 535574 212378
rect 534954 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 535574 212294
rect 534954 176614 535574 212058
rect 534954 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 535574 176614
rect 534954 176294 535574 176378
rect 534954 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 535574 176294
rect 534954 140614 535574 176058
rect 534954 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 535574 140614
rect 534954 140294 535574 140378
rect 534954 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 535574 140294
rect 534954 104614 535574 140058
rect 534954 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 535574 104614
rect 534954 104294 535574 104378
rect 534954 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 535574 104294
rect 534954 68614 535574 104058
rect 534954 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 535574 68614
rect 534954 68294 535574 68378
rect 534954 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 535574 68294
rect 534954 32614 535574 68058
rect 534954 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 535574 32614
rect 534954 32294 535574 32378
rect 534954 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 535574 32294
rect 516954 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 517574 -6106
rect 516954 -6426 517574 -6342
rect 516954 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 517574 -6426
rect 516954 -7654 517574 -6662
rect 534954 -7066 535574 32058
rect 541794 704838 542414 705830
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -1894 542414 -902
rect 545514 691174 546134 706202
rect 545514 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 546134 691174
rect 545514 690854 546134 690938
rect 545514 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 546134 690854
rect 545514 655174 546134 690618
rect 545514 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 546134 655174
rect 545514 654854 546134 654938
rect 545514 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 546134 654854
rect 545514 619174 546134 654618
rect 545514 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 546134 619174
rect 545514 618854 546134 618938
rect 545514 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 546134 618854
rect 545514 583174 546134 618618
rect 545514 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 546134 583174
rect 545514 582854 546134 582938
rect 545514 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 546134 582854
rect 545514 547174 546134 582618
rect 545514 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 546134 547174
rect 545514 546854 546134 546938
rect 545514 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 546134 546854
rect 545514 511174 546134 546618
rect 545514 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 546134 511174
rect 545514 510854 546134 510938
rect 545514 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 546134 510854
rect 545514 475174 546134 510618
rect 545514 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 546134 475174
rect 545514 474854 546134 474938
rect 545514 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 546134 474854
rect 545514 439174 546134 474618
rect 545514 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 546134 439174
rect 545514 438854 546134 438938
rect 545514 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 546134 438854
rect 545514 403174 546134 438618
rect 545514 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 546134 403174
rect 545514 402854 546134 402938
rect 545514 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 546134 402854
rect 545514 367174 546134 402618
rect 545514 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 546134 367174
rect 545514 366854 546134 366938
rect 545514 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 546134 366854
rect 545514 331174 546134 366618
rect 545514 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 546134 331174
rect 545514 330854 546134 330938
rect 545514 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 546134 330854
rect 545514 295174 546134 330618
rect 545514 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 546134 295174
rect 545514 294854 546134 294938
rect 545514 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 546134 294854
rect 545514 259174 546134 294618
rect 545514 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 546134 259174
rect 545514 258854 546134 258938
rect 545514 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 546134 258854
rect 545514 223174 546134 258618
rect 545514 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 546134 223174
rect 545514 222854 546134 222938
rect 545514 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 546134 222854
rect 545514 187174 546134 222618
rect 545514 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 546134 187174
rect 545514 186854 546134 186938
rect 545514 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 546134 186854
rect 545514 151174 546134 186618
rect 545514 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 546134 151174
rect 545514 150854 546134 150938
rect 545514 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 546134 150854
rect 545514 115174 546134 150618
rect 545514 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 546134 115174
rect 545514 114854 546134 114938
rect 545514 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 546134 114854
rect 545514 79174 546134 114618
rect 545514 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 546134 79174
rect 545514 78854 546134 78938
rect 545514 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 546134 78854
rect 545514 43174 546134 78618
rect 545514 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 546134 43174
rect 545514 42854 546134 42938
rect 545514 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 546134 42854
rect 545514 7174 546134 42618
rect 545514 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 546134 7174
rect 545514 6854 546134 6938
rect 545514 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 546134 6854
rect 545514 -2266 546134 6618
rect 545514 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 546134 -2266
rect 545514 -2586 546134 -2502
rect 545514 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 546134 -2586
rect 545514 -3814 546134 -2822
rect 549234 694894 549854 708122
rect 549234 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 549854 694894
rect 549234 694574 549854 694658
rect 549234 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 549854 694574
rect 549234 658894 549854 694338
rect 549234 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 549854 658894
rect 549234 658574 549854 658658
rect 549234 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 549854 658574
rect 549234 622894 549854 658338
rect 549234 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 549854 622894
rect 549234 622574 549854 622658
rect 549234 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 549854 622574
rect 549234 586894 549854 622338
rect 549234 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 549854 586894
rect 549234 586574 549854 586658
rect 549234 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 549854 586574
rect 549234 550894 549854 586338
rect 549234 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 549854 550894
rect 549234 550574 549854 550658
rect 549234 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 549854 550574
rect 549234 514894 549854 550338
rect 549234 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 549854 514894
rect 549234 514574 549854 514658
rect 549234 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 549854 514574
rect 549234 478894 549854 514338
rect 549234 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 549854 478894
rect 549234 478574 549854 478658
rect 549234 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 549854 478574
rect 549234 442894 549854 478338
rect 549234 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 549854 442894
rect 549234 442574 549854 442658
rect 549234 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 549854 442574
rect 549234 406894 549854 442338
rect 549234 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 549854 406894
rect 549234 406574 549854 406658
rect 549234 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 549854 406574
rect 549234 370894 549854 406338
rect 549234 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 549854 370894
rect 549234 370574 549854 370658
rect 549234 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 549854 370574
rect 549234 334894 549854 370338
rect 549234 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 549854 334894
rect 549234 334574 549854 334658
rect 549234 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 549854 334574
rect 549234 298894 549854 334338
rect 549234 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 549854 298894
rect 549234 298574 549854 298658
rect 549234 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 549854 298574
rect 549234 262894 549854 298338
rect 549234 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 549854 262894
rect 549234 262574 549854 262658
rect 549234 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 549854 262574
rect 549234 226894 549854 262338
rect 549234 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 549854 226894
rect 549234 226574 549854 226658
rect 549234 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 549854 226574
rect 549234 190894 549854 226338
rect 549234 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 549854 190894
rect 549234 190574 549854 190658
rect 549234 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 549854 190574
rect 549234 154894 549854 190338
rect 549234 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 549854 154894
rect 549234 154574 549854 154658
rect 549234 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 549854 154574
rect 549234 118894 549854 154338
rect 549234 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 549854 118894
rect 549234 118574 549854 118658
rect 549234 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 549854 118574
rect 549234 82894 549854 118338
rect 549234 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 549854 82894
rect 549234 82574 549854 82658
rect 549234 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 549854 82574
rect 549234 46894 549854 82338
rect 549234 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 549854 46894
rect 549234 46574 549854 46658
rect 549234 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 549854 46574
rect 549234 10894 549854 46338
rect 549234 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 549854 10894
rect 549234 10574 549854 10658
rect 549234 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 549854 10574
rect 549234 -4186 549854 10338
rect 549234 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 549854 -4186
rect 549234 -4506 549854 -4422
rect 549234 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 549854 -4506
rect 549234 -5734 549854 -4742
rect 552954 698614 553574 710042
rect 570954 711558 571574 711590
rect 570954 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 571574 711558
rect 570954 711238 571574 711322
rect 570954 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 571574 711238
rect 567234 709638 567854 709670
rect 567234 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 567854 709638
rect 567234 709318 567854 709402
rect 567234 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 567854 709318
rect 563514 707718 564134 707750
rect 563514 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 564134 707718
rect 563514 707398 564134 707482
rect 563514 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 564134 707398
rect 552954 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 553574 698614
rect 552954 698294 553574 698378
rect 552954 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 553574 698294
rect 552954 662614 553574 698058
rect 552954 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 553574 662614
rect 552954 662294 553574 662378
rect 552954 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 553574 662294
rect 552954 626614 553574 662058
rect 552954 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 553574 626614
rect 552954 626294 553574 626378
rect 552954 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 553574 626294
rect 552954 590614 553574 626058
rect 552954 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 553574 590614
rect 552954 590294 553574 590378
rect 552954 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 553574 590294
rect 552954 554614 553574 590058
rect 552954 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 553574 554614
rect 552954 554294 553574 554378
rect 552954 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 553574 554294
rect 552954 518614 553574 554058
rect 552954 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 553574 518614
rect 552954 518294 553574 518378
rect 552954 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 553574 518294
rect 552954 482614 553574 518058
rect 552954 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 553574 482614
rect 552954 482294 553574 482378
rect 552954 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 553574 482294
rect 552954 446614 553574 482058
rect 552954 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 553574 446614
rect 552954 446294 553574 446378
rect 552954 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 553574 446294
rect 552954 410614 553574 446058
rect 552954 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 553574 410614
rect 552954 410294 553574 410378
rect 552954 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 553574 410294
rect 552954 374614 553574 410058
rect 552954 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 553574 374614
rect 552954 374294 553574 374378
rect 552954 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 553574 374294
rect 552954 338614 553574 374058
rect 552954 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 553574 338614
rect 552954 338294 553574 338378
rect 552954 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 553574 338294
rect 552954 302614 553574 338058
rect 552954 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 553574 302614
rect 552954 302294 553574 302378
rect 552954 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 553574 302294
rect 552954 266614 553574 302058
rect 552954 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 553574 266614
rect 552954 266294 553574 266378
rect 552954 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 553574 266294
rect 552954 230614 553574 266058
rect 552954 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 553574 230614
rect 552954 230294 553574 230378
rect 552954 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 553574 230294
rect 552954 194614 553574 230058
rect 552954 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 553574 194614
rect 552954 194294 553574 194378
rect 552954 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 553574 194294
rect 552954 158614 553574 194058
rect 552954 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 553574 158614
rect 552954 158294 553574 158378
rect 552954 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 553574 158294
rect 552954 122614 553574 158058
rect 552954 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 553574 122614
rect 552954 122294 553574 122378
rect 552954 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 553574 122294
rect 552954 86614 553574 122058
rect 552954 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 553574 86614
rect 552954 86294 553574 86378
rect 552954 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 553574 86294
rect 552954 50614 553574 86058
rect 552954 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 553574 50614
rect 552954 50294 553574 50378
rect 552954 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 553574 50294
rect 552954 14614 553574 50058
rect 552954 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 553574 14614
rect 552954 14294 553574 14378
rect 552954 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 553574 14294
rect 534954 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 535574 -7066
rect 534954 -7386 535574 -7302
rect 534954 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 535574 -7386
rect 534954 -7654 535574 -7622
rect 552954 -6106 553574 14058
rect 559794 705798 560414 705830
rect 559794 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 560414 705798
rect 559794 705478 560414 705562
rect 559794 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 560414 705478
rect 559794 669454 560414 705242
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -1306 560414 20898
rect 559794 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 560414 -1306
rect 559794 -1626 560414 -1542
rect 559794 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 560414 -1626
rect 559794 -1894 560414 -1862
rect 563514 673174 564134 707162
rect 563514 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 564134 673174
rect 563514 672854 564134 672938
rect 563514 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 564134 672854
rect 563514 637174 564134 672618
rect 563514 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 564134 637174
rect 563514 636854 564134 636938
rect 563514 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 564134 636854
rect 563514 601174 564134 636618
rect 563514 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 564134 601174
rect 563514 600854 564134 600938
rect 563514 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 564134 600854
rect 563514 565174 564134 600618
rect 563514 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 564134 565174
rect 563514 564854 564134 564938
rect 563514 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 564134 564854
rect 563514 529174 564134 564618
rect 563514 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 564134 529174
rect 563514 528854 564134 528938
rect 563514 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 564134 528854
rect 563514 493174 564134 528618
rect 563514 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 564134 493174
rect 563514 492854 564134 492938
rect 563514 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 564134 492854
rect 563514 457174 564134 492618
rect 563514 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 564134 457174
rect 563514 456854 564134 456938
rect 563514 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 564134 456854
rect 563514 421174 564134 456618
rect 563514 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 564134 421174
rect 563514 420854 564134 420938
rect 563514 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 564134 420854
rect 563514 385174 564134 420618
rect 563514 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 564134 385174
rect 563514 384854 564134 384938
rect 563514 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 564134 384854
rect 563514 349174 564134 384618
rect 563514 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 564134 349174
rect 563514 348854 564134 348938
rect 563514 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 564134 348854
rect 563514 313174 564134 348618
rect 563514 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 564134 313174
rect 563514 312854 564134 312938
rect 563514 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 564134 312854
rect 563514 277174 564134 312618
rect 563514 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 564134 277174
rect 563514 276854 564134 276938
rect 563514 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 564134 276854
rect 563514 241174 564134 276618
rect 563514 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 564134 241174
rect 563514 240854 564134 240938
rect 563514 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 564134 240854
rect 563514 205174 564134 240618
rect 563514 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 564134 205174
rect 563514 204854 564134 204938
rect 563514 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 564134 204854
rect 563514 169174 564134 204618
rect 563514 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 564134 169174
rect 563514 168854 564134 168938
rect 563514 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 564134 168854
rect 563514 133174 564134 168618
rect 563514 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 564134 133174
rect 563514 132854 564134 132938
rect 563514 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 564134 132854
rect 563514 97174 564134 132618
rect 563514 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 564134 97174
rect 563514 96854 564134 96938
rect 563514 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 564134 96854
rect 563514 61174 564134 96618
rect 563514 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 564134 61174
rect 563514 60854 564134 60938
rect 563514 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 564134 60854
rect 563514 25174 564134 60618
rect 563514 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 564134 25174
rect 563514 24854 564134 24938
rect 563514 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 564134 24854
rect 563514 -3226 564134 24618
rect 563514 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 564134 -3226
rect 563514 -3546 564134 -3462
rect 563514 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 564134 -3546
rect 563514 -3814 564134 -3782
rect 567234 676894 567854 709082
rect 567234 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 567854 676894
rect 567234 676574 567854 676658
rect 567234 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 567854 676574
rect 567234 640894 567854 676338
rect 567234 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 567854 640894
rect 567234 640574 567854 640658
rect 567234 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 567854 640574
rect 567234 604894 567854 640338
rect 567234 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 567854 604894
rect 567234 604574 567854 604658
rect 567234 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 567854 604574
rect 567234 568894 567854 604338
rect 567234 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 567854 568894
rect 567234 568574 567854 568658
rect 567234 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 567854 568574
rect 567234 532894 567854 568338
rect 567234 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 567854 532894
rect 567234 532574 567854 532658
rect 567234 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 567854 532574
rect 567234 496894 567854 532338
rect 567234 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 567854 496894
rect 567234 496574 567854 496658
rect 567234 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 567854 496574
rect 567234 460894 567854 496338
rect 567234 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 567854 460894
rect 567234 460574 567854 460658
rect 567234 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 567854 460574
rect 567234 424894 567854 460338
rect 567234 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 567854 424894
rect 567234 424574 567854 424658
rect 567234 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 567854 424574
rect 567234 388894 567854 424338
rect 567234 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 567854 388894
rect 567234 388574 567854 388658
rect 567234 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 567854 388574
rect 567234 352894 567854 388338
rect 567234 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 567854 352894
rect 567234 352574 567854 352658
rect 567234 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 567854 352574
rect 567234 316894 567854 352338
rect 567234 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 567854 316894
rect 567234 316574 567854 316658
rect 567234 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 567854 316574
rect 567234 280894 567854 316338
rect 567234 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 567854 280894
rect 567234 280574 567854 280658
rect 567234 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 567854 280574
rect 567234 244894 567854 280338
rect 567234 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 567854 244894
rect 567234 244574 567854 244658
rect 567234 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 567854 244574
rect 567234 208894 567854 244338
rect 567234 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 567854 208894
rect 567234 208574 567854 208658
rect 567234 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 567854 208574
rect 567234 172894 567854 208338
rect 567234 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 567854 172894
rect 567234 172574 567854 172658
rect 567234 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 567854 172574
rect 567234 136894 567854 172338
rect 567234 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 567854 136894
rect 567234 136574 567854 136658
rect 567234 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 567854 136574
rect 567234 100894 567854 136338
rect 567234 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 567854 100894
rect 567234 100574 567854 100658
rect 567234 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 567854 100574
rect 567234 64894 567854 100338
rect 567234 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 567854 64894
rect 567234 64574 567854 64658
rect 567234 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 567854 64574
rect 567234 28894 567854 64338
rect 567234 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 567854 28894
rect 567234 28574 567854 28658
rect 567234 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 567854 28574
rect 567234 -5146 567854 28338
rect 567234 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 567854 -5146
rect 567234 -5466 567854 -5382
rect 567234 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 567854 -5466
rect 567234 -5734 567854 -5702
rect 570954 680614 571574 711002
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 581514 706758 582134 707750
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 581514 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 582134 706758
rect 581514 706438 582134 706522
rect 581514 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 582134 706438
rect 570954 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 571574 680614
rect 570954 680294 571574 680378
rect 570954 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 571574 680294
rect 570954 644614 571574 680058
rect 570954 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 571574 644614
rect 570954 644294 571574 644378
rect 570954 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 571574 644294
rect 570954 608614 571574 644058
rect 570954 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 571574 608614
rect 570954 608294 571574 608378
rect 570954 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 571574 608294
rect 570954 572614 571574 608058
rect 570954 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 571574 572614
rect 570954 572294 571574 572378
rect 570954 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 571574 572294
rect 570954 536614 571574 572058
rect 570954 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 571574 536614
rect 570954 536294 571574 536378
rect 570954 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 571574 536294
rect 570954 500614 571574 536058
rect 570954 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 571574 500614
rect 570954 500294 571574 500378
rect 570954 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 571574 500294
rect 570954 464614 571574 500058
rect 570954 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 571574 464614
rect 570954 464294 571574 464378
rect 570954 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 571574 464294
rect 570954 428614 571574 464058
rect 570954 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 571574 428614
rect 570954 428294 571574 428378
rect 570954 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 571574 428294
rect 570954 392614 571574 428058
rect 570954 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 571574 392614
rect 570954 392294 571574 392378
rect 570954 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 571574 392294
rect 570954 356614 571574 392058
rect 570954 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 571574 356614
rect 570954 356294 571574 356378
rect 570954 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 571574 356294
rect 570954 320614 571574 356058
rect 570954 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 571574 320614
rect 570954 320294 571574 320378
rect 570954 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 571574 320294
rect 570954 284614 571574 320058
rect 570954 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 571574 284614
rect 570954 284294 571574 284378
rect 570954 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 571574 284294
rect 570954 248614 571574 284058
rect 570954 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 571574 248614
rect 570954 248294 571574 248378
rect 570954 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 571574 248294
rect 570954 212614 571574 248058
rect 570954 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 571574 212614
rect 570954 212294 571574 212378
rect 570954 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 571574 212294
rect 570954 176614 571574 212058
rect 570954 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 571574 176614
rect 570954 176294 571574 176378
rect 570954 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 571574 176294
rect 570954 140614 571574 176058
rect 570954 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 571574 140614
rect 570954 140294 571574 140378
rect 570954 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 571574 140294
rect 570954 104614 571574 140058
rect 570954 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 571574 104614
rect 570954 104294 571574 104378
rect 570954 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 571574 104294
rect 570954 68614 571574 104058
rect 570954 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 571574 68614
rect 570954 68294 571574 68378
rect 570954 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 571574 68294
rect 570954 32614 571574 68058
rect 570954 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 571574 32614
rect 570954 32294 571574 32378
rect 570954 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 571574 32294
rect 552954 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 553574 -6106
rect 552954 -6426 553574 -6342
rect 552954 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 553574 -6426
rect 552954 -7654 553574 -6662
rect 570954 -7066 571574 32058
rect 577794 704838 578414 705830
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -1894 578414 -902
rect 581514 691174 582134 706202
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581514 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 582134 691174
rect 581514 690854 582134 690938
rect 581514 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 582134 690854
rect 581514 655174 582134 690618
rect 581514 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 582134 655174
rect 581514 654854 582134 654938
rect 581514 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 582134 654854
rect 581514 619174 582134 654618
rect 581514 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 582134 619174
rect 581514 618854 582134 618938
rect 581514 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 582134 618854
rect 581514 583174 582134 618618
rect 581514 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 582134 583174
rect 581514 582854 582134 582938
rect 581514 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 582134 582854
rect 581514 547174 582134 582618
rect 581514 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 582134 547174
rect 581514 546854 582134 546938
rect 581514 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 582134 546854
rect 581514 511174 582134 546618
rect 581514 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 582134 511174
rect 581514 510854 582134 510938
rect 581514 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 582134 510854
rect 581514 475174 582134 510618
rect 581514 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 582134 475174
rect 581514 474854 582134 474938
rect 581514 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 582134 474854
rect 581514 439174 582134 474618
rect 581514 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 582134 439174
rect 581514 438854 582134 438938
rect 581514 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 582134 438854
rect 581514 403174 582134 438618
rect 581514 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 582134 403174
rect 581514 402854 582134 402938
rect 581514 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 582134 402854
rect 581514 367174 582134 402618
rect 581514 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 582134 367174
rect 581514 366854 582134 366938
rect 581514 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 582134 366854
rect 581514 331174 582134 366618
rect 581514 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 582134 331174
rect 581514 330854 582134 330938
rect 581514 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 582134 330854
rect 581514 295174 582134 330618
rect 581514 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 582134 295174
rect 581514 294854 582134 294938
rect 581514 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 582134 294854
rect 581514 259174 582134 294618
rect 581514 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 582134 259174
rect 581514 258854 582134 258938
rect 581514 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 582134 258854
rect 581514 223174 582134 258618
rect 581514 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 582134 223174
rect 581514 222854 582134 222938
rect 581514 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 582134 222854
rect 581514 187174 582134 222618
rect 581514 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 582134 187174
rect 581514 186854 582134 186938
rect 581514 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 582134 186854
rect 581514 151174 582134 186618
rect 581514 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 582134 151174
rect 581514 150854 582134 150938
rect 581514 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 582134 150854
rect 581514 115174 582134 150618
rect 581514 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 582134 115174
rect 581514 114854 582134 114938
rect 581514 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 582134 114854
rect 581514 79174 582134 114618
rect 581514 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 582134 79174
rect 581514 78854 582134 78938
rect 581514 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 582134 78854
rect 581514 43174 582134 78618
rect 581514 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 582134 43174
rect 581514 42854 582134 42938
rect 581514 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 582134 42854
rect 581514 7174 582134 42618
rect 581514 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 582134 7174
rect 581514 6854 582134 6938
rect 581514 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 582134 6854
rect 581514 -2266 582134 6618
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 669454 586890 705242
rect 586270 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect 586270 669134 586890 669218
rect 586270 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect 586270 633454 586890 668898
rect 586270 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect 586270 633134 586890 633218
rect 586270 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect 586270 597454 586890 632898
rect 586270 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect 586270 597134 586890 597218
rect 586270 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect 586270 561454 586890 596898
rect 586270 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect 586270 561134 586890 561218
rect 586270 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect 586270 525454 586890 560898
rect 586270 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect 586270 525134 586890 525218
rect 586270 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect 586270 489454 586890 524898
rect 586270 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect 586270 489134 586890 489218
rect 586270 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect 586270 453454 586890 488898
rect 586270 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect 586270 453134 586890 453218
rect 586270 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect 586270 417454 586890 452898
rect 586270 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect 586270 417134 586890 417218
rect 586270 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect 586270 381454 586890 416898
rect 586270 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect 586270 381134 586890 381218
rect 586270 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect 586270 345454 586890 380898
rect 586270 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect 586270 345134 586890 345218
rect 586270 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect 586270 309454 586890 344898
rect 586270 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect 586270 309134 586890 309218
rect 586270 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect 586270 273454 586890 308898
rect 586270 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect 586270 273134 586890 273218
rect 586270 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect 586270 237454 586890 272898
rect 586270 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect 586270 237134 586890 237218
rect 586270 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect 586270 201454 586890 236898
rect 586270 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect 586270 201134 586890 201218
rect 586270 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect 586270 165454 586890 200898
rect 586270 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect 586270 165134 586890 165218
rect 586270 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect 586270 129454 586890 164898
rect 586270 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect 586270 129134 586890 129218
rect 586270 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect 586270 93454 586890 128898
rect 586270 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect 586270 93134 586890 93218
rect 586270 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect 586270 57454 586890 92898
rect 586270 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect 586270 57134 586890 57218
rect 586270 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect 586270 21454 586890 56898
rect 586270 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect 586270 21134 586890 21218
rect 586270 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect 586270 -1306 586890 20898
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 691174 587850 706202
rect 587230 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 587850 691174
rect 587230 690854 587850 690938
rect 587230 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 587850 690854
rect 587230 655174 587850 690618
rect 587230 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 587850 655174
rect 587230 654854 587850 654938
rect 587230 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 587850 654854
rect 587230 619174 587850 654618
rect 587230 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 587850 619174
rect 587230 618854 587850 618938
rect 587230 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 587850 618854
rect 587230 583174 587850 618618
rect 587230 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 587850 583174
rect 587230 582854 587850 582938
rect 587230 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 587850 582854
rect 587230 547174 587850 582618
rect 587230 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 587850 547174
rect 587230 546854 587850 546938
rect 587230 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 587850 546854
rect 587230 511174 587850 546618
rect 587230 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 587850 511174
rect 587230 510854 587850 510938
rect 587230 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 587850 510854
rect 587230 475174 587850 510618
rect 587230 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 587850 475174
rect 587230 474854 587850 474938
rect 587230 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 587850 474854
rect 587230 439174 587850 474618
rect 587230 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 587850 439174
rect 587230 438854 587850 438938
rect 587230 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 587850 438854
rect 587230 403174 587850 438618
rect 587230 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 587850 403174
rect 587230 402854 587850 402938
rect 587230 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 587850 402854
rect 587230 367174 587850 402618
rect 587230 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 587850 367174
rect 587230 366854 587850 366938
rect 587230 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 587850 366854
rect 587230 331174 587850 366618
rect 587230 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 587850 331174
rect 587230 330854 587850 330938
rect 587230 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 587850 330854
rect 587230 295174 587850 330618
rect 587230 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 587850 295174
rect 587230 294854 587850 294938
rect 587230 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 587850 294854
rect 587230 259174 587850 294618
rect 587230 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 587850 259174
rect 587230 258854 587850 258938
rect 587230 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 587850 258854
rect 587230 223174 587850 258618
rect 587230 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 587850 223174
rect 587230 222854 587850 222938
rect 587230 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 587850 222854
rect 587230 187174 587850 222618
rect 587230 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 587850 187174
rect 587230 186854 587850 186938
rect 587230 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 587850 186854
rect 587230 151174 587850 186618
rect 587230 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 587850 151174
rect 587230 150854 587850 150938
rect 587230 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 587850 150854
rect 587230 115174 587850 150618
rect 587230 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 587850 115174
rect 587230 114854 587850 114938
rect 587230 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 587850 114854
rect 587230 79174 587850 114618
rect 587230 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 587850 79174
rect 587230 78854 587850 78938
rect 587230 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 587850 78854
rect 587230 43174 587850 78618
rect 587230 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 587850 43174
rect 587230 42854 587850 42938
rect 587230 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 587850 42854
rect 587230 7174 587850 42618
rect 587230 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 587850 7174
rect 587230 6854 587850 6938
rect 587230 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 587850 6854
rect 581514 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 582134 -2266
rect 581514 -2586 582134 -2502
rect 581514 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 582134 -2586
rect 581514 -3814 582134 -2822
rect 587230 -2266 587850 6618
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 673174 588810 707162
rect 588190 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect 588190 672854 588810 672938
rect 588190 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect 588190 637174 588810 672618
rect 588190 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect 588190 636854 588810 636938
rect 588190 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect 588190 601174 588810 636618
rect 588190 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect 588190 600854 588810 600938
rect 588190 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect 588190 565174 588810 600618
rect 588190 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect 588190 564854 588810 564938
rect 588190 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect 588190 529174 588810 564618
rect 588190 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect 588190 528854 588810 528938
rect 588190 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect 588190 493174 588810 528618
rect 588190 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect 588190 492854 588810 492938
rect 588190 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect 588190 457174 588810 492618
rect 588190 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect 588190 456854 588810 456938
rect 588190 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect 588190 421174 588810 456618
rect 588190 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect 588190 420854 588810 420938
rect 588190 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect 588190 385174 588810 420618
rect 588190 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect 588190 384854 588810 384938
rect 588190 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect 588190 349174 588810 384618
rect 588190 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect 588190 348854 588810 348938
rect 588190 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect 588190 313174 588810 348618
rect 588190 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect 588190 312854 588810 312938
rect 588190 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect 588190 277174 588810 312618
rect 588190 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect 588190 276854 588810 276938
rect 588190 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect 588190 241174 588810 276618
rect 588190 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect 588190 240854 588810 240938
rect 588190 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect 588190 205174 588810 240618
rect 588190 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect 588190 204854 588810 204938
rect 588190 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect 588190 169174 588810 204618
rect 588190 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect 588190 168854 588810 168938
rect 588190 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect 588190 133174 588810 168618
rect 588190 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect 588190 132854 588810 132938
rect 588190 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect 588190 97174 588810 132618
rect 588190 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect 588190 96854 588810 96938
rect 588190 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect 588190 61174 588810 96618
rect 588190 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect 588190 60854 588810 60938
rect 588190 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect 588190 25174 588810 60618
rect 588190 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect 588190 24854 588810 24938
rect 588190 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect 588190 -3226 588810 24618
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 694894 589770 708122
rect 589150 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 589770 694894
rect 589150 694574 589770 694658
rect 589150 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 589770 694574
rect 589150 658894 589770 694338
rect 589150 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 589770 658894
rect 589150 658574 589770 658658
rect 589150 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 589770 658574
rect 589150 622894 589770 658338
rect 589150 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 589770 622894
rect 589150 622574 589770 622658
rect 589150 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 589770 622574
rect 589150 586894 589770 622338
rect 589150 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 589770 586894
rect 589150 586574 589770 586658
rect 589150 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 589770 586574
rect 589150 550894 589770 586338
rect 589150 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 589770 550894
rect 589150 550574 589770 550658
rect 589150 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 589770 550574
rect 589150 514894 589770 550338
rect 589150 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 589770 514894
rect 589150 514574 589770 514658
rect 589150 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 589770 514574
rect 589150 478894 589770 514338
rect 589150 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 589770 478894
rect 589150 478574 589770 478658
rect 589150 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 589770 478574
rect 589150 442894 589770 478338
rect 589150 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 589770 442894
rect 589150 442574 589770 442658
rect 589150 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 589770 442574
rect 589150 406894 589770 442338
rect 589150 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 589770 406894
rect 589150 406574 589770 406658
rect 589150 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 589770 406574
rect 589150 370894 589770 406338
rect 589150 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 589770 370894
rect 589150 370574 589770 370658
rect 589150 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 589770 370574
rect 589150 334894 589770 370338
rect 589150 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 589770 334894
rect 589150 334574 589770 334658
rect 589150 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 589770 334574
rect 589150 298894 589770 334338
rect 589150 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 589770 298894
rect 589150 298574 589770 298658
rect 589150 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 589770 298574
rect 589150 262894 589770 298338
rect 589150 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 589770 262894
rect 589150 262574 589770 262658
rect 589150 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 589770 262574
rect 589150 226894 589770 262338
rect 589150 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 589770 226894
rect 589150 226574 589770 226658
rect 589150 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 589770 226574
rect 589150 190894 589770 226338
rect 589150 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 589770 190894
rect 589150 190574 589770 190658
rect 589150 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 589770 190574
rect 589150 154894 589770 190338
rect 589150 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 589770 154894
rect 589150 154574 589770 154658
rect 589150 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 589770 154574
rect 589150 118894 589770 154338
rect 589150 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 589770 118894
rect 589150 118574 589770 118658
rect 589150 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 589770 118574
rect 589150 82894 589770 118338
rect 589150 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 589770 82894
rect 589150 82574 589770 82658
rect 589150 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 589770 82574
rect 589150 46894 589770 82338
rect 589150 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 589770 46894
rect 589150 46574 589770 46658
rect 589150 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 589770 46574
rect 589150 10894 589770 46338
rect 589150 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 589770 10894
rect 589150 10574 589770 10658
rect 589150 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 589770 10574
rect 589150 -4186 589770 10338
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 676894 590730 709082
rect 590110 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect 590110 676574 590730 676658
rect 590110 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect 590110 640894 590730 676338
rect 590110 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect 590110 640574 590730 640658
rect 590110 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect 590110 604894 590730 640338
rect 590110 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect 590110 604574 590730 604658
rect 590110 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect 590110 568894 590730 604338
rect 590110 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect 590110 568574 590730 568658
rect 590110 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect 590110 532894 590730 568338
rect 590110 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect 590110 532574 590730 532658
rect 590110 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect 590110 496894 590730 532338
rect 590110 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect 590110 496574 590730 496658
rect 590110 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect 590110 460894 590730 496338
rect 590110 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect 590110 460574 590730 460658
rect 590110 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect 590110 424894 590730 460338
rect 590110 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect 590110 424574 590730 424658
rect 590110 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect 590110 388894 590730 424338
rect 590110 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect 590110 388574 590730 388658
rect 590110 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect 590110 352894 590730 388338
rect 590110 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect 590110 352574 590730 352658
rect 590110 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect 590110 316894 590730 352338
rect 590110 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect 590110 316574 590730 316658
rect 590110 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect 590110 280894 590730 316338
rect 590110 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect 590110 280574 590730 280658
rect 590110 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect 590110 244894 590730 280338
rect 590110 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect 590110 244574 590730 244658
rect 590110 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect 590110 208894 590730 244338
rect 590110 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect 590110 208574 590730 208658
rect 590110 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect 590110 172894 590730 208338
rect 590110 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect 590110 172574 590730 172658
rect 590110 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect 590110 136894 590730 172338
rect 590110 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect 590110 136574 590730 136658
rect 590110 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect 590110 100894 590730 136338
rect 590110 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect 590110 100574 590730 100658
rect 590110 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect 590110 64894 590730 100338
rect 590110 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect 590110 64574 590730 64658
rect 590110 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect 590110 28894 590730 64338
rect 590110 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect 590110 28574 590730 28658
rect 590110 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect 590110 -5146 590730 28338
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 698614 591690 710042
rect 591070 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 591690 698614
rect 591070 698294 591690 698378
rect 591070 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 591690 698294
rect 591070 662614 591690 698058
rect 591070 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 591690 662614
rect 591070 662294 591690 662378
rect 591070 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 591690 662294
rect 591070 626614 591690 662058
rect 591070 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 591690 626614
rect 591070 626294 591690 626378
rect 591070 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 591690 626294
rect 591070 590614 591690 626058
rect 591070 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 591690 590614
rect 591070 590294 591690 590378
rect 591070 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 591690 590294
rect 591070 554614 591690 590058
rect 591070 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 591690 554614
rect 591070 554294 591690 554378
rect 591070 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 591690 554294
rect 591070 518614 591690 554058
rect 591070 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 591690 518614
rect 591070 518294 591690 518378
rect 591070 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 591690 518294
rect 591070 482614 591690 518058
rect 591070 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 591690 482614
rect 591070 482294 591690 482378
rect 591070 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 591690 482294
rect 591070 446614 591690 482058
rect 591070 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 591690 446614
rect 591070 446294 591690 446378
rect 591070 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 591690 446294
rect 591070 410614 591690 446058
rect 591070 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 591690 410614
rect 591070 410294 591690 410378
rect 591070 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 591690 410294
rect 591070 374614 591690 410058
rect 591070 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 591690 374614
rect 591070 374294 591690 374378
rect 591070 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 591690 374294
rect 591070 338614 591690 374058
rect 591070 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 591690 338614
rect 591070 338294 591690 338378
rect 591070 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 591690 338294
rect 591070 302614 591690 338058
rect 591070 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 591690 302614
rect 591070 302294 591690 302378
rect 591070 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 591690 302294
rect 591070 266614 591690 302058
rect 591070 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 591690 266614
rect 591070 266294 591690 266378
rect 591070 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 591690 266294
rect 591070 230614 591690 266058
rect 591070 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 591690 230614
rect 591070 230294 591690 230378
rect 591070 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 591690 230294
rect 591070 194614 591690 230058
rect 591070 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 591690 194614
rect 591070 194294 591690 194378
rect 591070 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 591690 194294
rect 591070 158614 591690 194058
rect 591070 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 591690 158614
rect 591070 158294 591690 158378
rect 591070 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 591690 158294
rect 591070 122614 591690 158058
rect 591070 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 591690 122614
rect 591070 122294 591690 122378
rect 591070 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 591690 122294
rect 591070 86614 591690 122058
rect 591070 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 591690 86614
rect 591070 86294 591690 86378
rect 591070 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 591690 86294
rect 591070 50614 591690 86058
rect 591070 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 591690 50614
rect 591070 50294 591690 50378
rect 591070 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 591690 50294
rect 591070 14614 591690 50058
rect 591070 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 591690 14614
rect 591070 14294 591690 14378
rect 591070 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 591690 14294
rect 591070 -6106 591690 14058
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 680614 592650 711002
rect 592030 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect 592030 680294 592650 680378
rect 592030 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect 592030 644614 592650 680058
rect 592030 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect 592030 644294 592650 644378
rect 592030 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect 592030 608614 592650 644058
rect 592030 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect 592030 608294 592650 608378
rect 592030 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect 592030 572614 592650 608058
rect 592030 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect 592030 572294 592650 572378
rect 592030 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect 592030 536614 592650 572058
rect 592030 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect 592030 536294 592650 536378
rect 592030 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect 592030 500614 592650 536058
rect 592030 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect 592030 500294 592650 500378
rect 592030 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect 592030 464614 592650 500058
rect 592030 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect 592030 464294 592650 464378
rect 592030 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect 592030 428614 592650 464058
rect 592030 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect 592030 428294 592650 428378
rect 592030 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect 592030 392614 592650 428058
rect 592030 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect 592030 392294 592650 392378
rect 592030 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect 592030 356614 592650 392058
rect 592030 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect 592030 356294 592650 356378
rect 592030 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect 592030 320614 592650 356058
rect 592030 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect 592030 320294 592650 320378
rect 592030 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect 592030 284614 592650 320058
rect 592030 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect 592030 284294 592650 284378
rect 592030 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect 592030 248614 592650 284058
rect 592030 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect 592030 248294 592650 248378
rect 592030 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect 592030 212614 592650 248058
rect 592030 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect 592030 212294 592650 212378
rect 592030 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect 592030 176614 592650 212058
rect 592030 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect 592030 176294 592650 176378
rect 592030 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect 592030 140614 592650 176058
rect 592030 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect 592030 140294 592650 140378
rect 592030 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect 592030 104614 592650 140058
rect 592030 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect 592030 104294 592650 104378
rect 592030 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect 592030 68614 592650 104058
rect 592030 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect 592030 68294 592650 68378
rect 592030 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect 592030 32614 592650 68058
rect 592030 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect 592030 32294 592650 32378
rect 592030 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect 570954 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 571574 -7066
rect 570954 -7386 571574 -7302
rect 570954 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 571574 -7386
rect 570954 -7654 571574 -7622
rect 592030 -7066 592650 32058
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 680378 -8458 680614
rect -8374 680378 -8138 680614
rect -8694 680058 -8458 680294
rect -8374 680058 -8138 680294
rect -8694 644378 -8458 644614
rect -8374 644378 -8138 644614
rect -8694 644058 -8458 644294
rect -8374 644058 -8138 644294
rect -8694 608378 -8458 608614
rect -8374 608378 -8138 608614
rect -8694 608058 -8458 608294
rect -8374 608058 -8138 608294
rect -8694 572378 -8458 572614
rect -8374 572378 -8138 572614
rect -8694 572058 -8458 572294
rect -8374 572058 -8138 572294
rect -8694 536378 -8458 536614
rect -8374 536378 -8138 536614
rect -8694 536058 -8458 536294
rect -8374 536058 -8138 536294
rect -8694 500378 -8458 500614
rect -8374 500378 -8138 500614
rect -8694 500058 -8458 500294
rect -8374 500058 -8138 500294
rect -8694 464378 -8458 464614
rect -8374 464378 -8138 464614
rect -8694 464058 -8458 464294
rect -8374 464058 -8138 464294
rect -8694 428378 -8458 428614
rect -8374 428378 -8138 428614
rect -8694 428058 -8458 428294
rect -8374 428058 -8138 428294
rect -8694 392378 -8458 392614
rect -8374 392378 -8138 392614
rect -8694 392058 -8458 392294
rect -8374 392058 -8138 392294
rect -8694 356378 -8458 356614
rect -8374 356378 -8138 356614
rect -8694 356058 -8458 356294
rect -8374 356058 -8138 356294
rect -8694 320378 -8458 320614
rect -8374 320378 -8138 320614
rect -8694 320058 -8458 320294
rect -8374 320058 -8138 320294
rect -8694 284378 -8458 284614
rect -8374 284378 -8138 284614
rect -8694 284058 -8458 284294
rect -8374 284058 -8138 284294
rect -8694 248378 -8458 248614
rect -8374 248378 -8138 248614
rect -8694 248058 -8458 248294
rect -8374 248058 -8138 248294
rect -8694 212378 -8458 212614
rect -8374 212378 -8138 212614
rect -8694 212058 -8458 212294
rect -8374 212058 -8138 212294
rect -8694 176378 -8458 176614
rect -8374 176378 -8138 176614
rect -8694 176058 -8458 176294
rect -8374 176058 -8138 176294
rect -8694 140378 -8458 140614
rect -8374 140378 -8138 140614
rect -8694 140058 -8458 140294
rect -8374 140058 -8138 140294
rect -8694 104378 -8458 104614
rect -8374 104378 -8138 104614
rect -8694 104058 -8458 104294
rect -8374 104058 -8138 104294
rect -8694 68378 -8458 68614
rect -8374 68378 -8138 68614
rect -8694 68058 -8458 68294
rect -8374 68058 -8138 68294
rect -8694 32378 -8458 32614
rect -8374 32378 -8138 32614
rect -8694 32058 -8458 32294
rect -8374 32058 -8138 32294
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect 12986 710362 13222 710598
rect 13306 710362 13542 710598
rect 12986 710042 13222 710278
rect 13306 710042 13542 710278
rect -7734 698378 -7498 698614
rect -7414 698378 -7178 698614
rect -7734 698058 -7498 698294
rect -7414 698058 -7178 698294
rect -7734 662378 -7498 662614
rect -7414 662378 -7178 662614
rect -7734 662058 -7498 662294
rect -7414 662058 -7178 662294
rect -7734 626378 -7498 626614
rect -7414 626378 -7178 626614
rect -7734 626058 -7498 626294
rect -7414 626058 -7178 626294
rect -7734 590378 -7498 590614
rect -7414 590378 -7178 590614
rect -7734 590058 -7498 590294
rect -7414 590058 -7178 590294
rect -7734 554378 -7498 554614
rect -7414 554378 -7178 554614
rect -7734 554058 -7498 554294
rect -7414 554058 -7178 554294
rect -7734 518378 -7498 518614
rect -7414 518378 -7178 518614
rect -7734 518058 -7498 518294
rect -7414 518058 -7178 518294
rect -7734 482378 -7498 482614
rect -7414 482378 -7178 482614
rect -7734 482058 -7498 482294
rect -7414 482058 -7178 482294
rect -7734 446378 -7498 446614
rect -7414 446378 -7178 446614
rect -7734 446058 -7498 446294
rect -7414 446058 -7178 446294
rect -7734 410378 -7498 410614
rect -7414 410378 -7178 410614
rect -7734 410058 -7498 410294
rect -7414 410058 -7178 410294
rect -7734 374378 -7498 374614
rect -7414 374378 -7178 374614
rect -7734 374058 -7498 374294
rect -7414 374058 -7178 374294
rect -7734 338378 -7498 338614
rect -7414 338378 -7178 338614
rect -7734 338058 -7498 338294
rect -7414 338058 -7178 338294
rect -7734 302378 -7498 302614
rect -7414 302378 -7178 302614
rect -7734 302058 -7498 302294
rect -7414 302058 -7178 302294
rect -7734 266378 -7498 266614
rect -7414 266378 -7178 266614
rect -7734 266058 -7498 266294
rect -7414 266058 -7178 266294
rect -7734 230378 -7498 230614
rect -7414 230378 -7178 230614
rect -7734 230058 -7498 230294
rect -7414 230058 -7178 230294
rect -7734 194378 -7498 194614
rect -7414 194378 -7178 194614
rect -7734 194058 -7498 194294
rect -7414 194058 -7178 194294
rect -7734 158378 -7498 158614
rect -7414 158378 -7178 158614
rect -7734 158058 -7498 158294
rect -7414 158058 -7178 158294
rect -7734 122378 -7498 122614
rect -7414 122378 -7178 122614
rect -7734 122058 -7498 122294
rect -7414 122058 -7178 122294
rect -7734 86378 -7498 86614
rect -7414 86378 -7178 86614
rect -7734 86058 -7498 86294
rect -7414 86058 -7178 86294
rect -7734 50378 -7498 50614
rect -7414 50378 -7178 50614
rect -7734 50058 -7498 50294
rect -7414 50058 -7178 50294
rect -7734 14378 -7498 14614
rect -7414 14378 -7178 14614
rect -7734 14058 -7498 14294
rect -7414 14058 -7178 14294
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 676658 -6538 676894
rect -6454 676658 -6218 676894
rect -6774 676338 -6538 676574
rect -6454 676338 -6218 676574
rect -6774 640658 -6538 640894
rect -6454 640658 -6218 640894
rect -6774 640338 -6538 640574
rect -6454 640338 -6218 640574
rect -6774 604658 -6538 604894
rect -6454 604658 -6218 604894
rect -6774 604338 -6538 604574
rect -6454 604338 -6218 604574
rect -6774 568658 -6538 568894
rect -6454 568658 -6218 568894
rect -6774 568338 -6538 568574
rect -6454 568338 -6218 568574
rect -6774 532658 -6538 532894
rect -6454 532658 -6218 532894
rect -6774 532338 -6538 532574
rect -6454 532338 -6218 532574
rect -6774 496658 -6538 496894
rect -6454 496658 -6218 496894
rect -6774 496338 -6538 496574
rect -6454 496338 -6218 496574
rect -6774 460658 -6538 460894
rect -6454 460658 -6218 460894
rect -6774 460338 -6538 460574
rect -6454 460338 -6218 460574
rect -6774 424658 -6538 424894
rect -6454 424658 -6218 424894
rect -6774 424338 -6538 424574
rect -6454 424338 -6218 424574
rect -6774 388658 -6538 388894
rect -6454 388658 -6218 388894
rect -6774 388338 -6538 388574
rect -6454 388338 -6218 388574
rect -6774 352658 -6538 352894
rect -6454 352658 -6218 352894
rect -6774 352338 -6538 352574
rect -6454 352338 -6218 352574
rect -6774 316658 -6538 316894
rect -6454 316658 -6218 316894
rect -6774 316338 -6538 316574
rect -6454 316338 -6218 316574
rect -6774 280658 -6538 280894
rect -6454 280658 -6218 280894
rect -6774 280338 -6538 280574
rect -6454 280338 -6218 280574
rect -6774 244658 -6538 244894
rect -6454 244658 -6218 244894
rect -6774 244338 -6538 244574
rect -6454 244338 -6218 244574
rect -6774 208658 -6538 208894
rect -6454 208658 -6218 208894
rect -6774 208338 -6538 208574
rect -6454 208338 -6218 208574
rect -6774 172658 -6538 172894
rect -6454 172658 -6218 172894
rect -6774 172338 -6538 172574
rect -6454 172338 -6218 172574
rect -6774 136658 -6538 136894
rect -6454 136658 -6218 136894
rect -6774 136338 -6538 136574
rect -6454 136338 -6218 136574
rect -6774 100658 -6538 100894
rect -6454 100658 -6218 100894
rect -6774 100338 -6538 100574
rect -6454 100338 -6218 100574
rect -6774 64658 -6538 64894
rect -6454 64658 -6218 64894
rect -6774 64338 -6538 64574
rect -6454 64338 -6218 64574
rect -6774 28658 -6538 28894
rect -6454 28658 -6218 28894
rect -6774 28338 -6538 28574
rect -6454 28338 -6218 28574
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect 9266 708442 9502 708678
rect 9586 708442 9822 708678
rect 9266 708122 9502 708358
rect 9586 708122 9822 708358
rect -5814 694658 -5578 694894
rect -5494 694658 -5258 694894
rect -5814 694338 -5578 694574
rect -5494 694338 -5258 694574
rect -5814 658658 -5578 658894
rect -5494 658658 -5258 658894
rect -5814 658338 -5578 658574
rect -5494 658338 -5258 658574
rect -5814 622658 -5578 622894
rect -5494 622658 -5258 622894
rect -5814 622338 -5578 622574
rect -5494 622338 -5258 622574
rect -5814 586658 -5578 586894
rect -5494 586658 -5258 586894
rect -5814 586338 -5578 586574
rect -5494 586338 -5258 586574
rect -5814 550658 -5578 550894
rect -5494 550658 -5258 550894
rect -5814 550338 -5578 550574
rect -5494 550338 -5258 550574
rect -5814 514658 -5578 514894
rect -5494 514658 -5258 514894
rect -5814 514338 -5578 514574
rect -5494 514338 -5258 514574
rect -5814 478658 -5578 478894
rect -5494 478658 -5258 478894
rect -5814 478338 -5578 478574
rect -5494 478338 -5258 478574
rect -5814 442658 -5578 442894
rect -5494 442658 -5258 442894
rect -5814 442338 -5578 442574
rect -5494 442338 -5258 442574
rect -5814 406658 -5578 406894
rect -5494 406658 -5258 406894
rect -5814 406338 -5578 406574
rect -5494 406338 -5258 406574
rect -5814 370658 -5578 370894
rect -5494 370658 -5258 370894
rect -5814 370338 -5578 370574
rect -5494 370338 -5258 370574
rect -5814 334658 -5578 334894
rect -5494 334658 -5258 334894
rect -5814 334338 -5578 334574
rect -5494 334338 -5258 334574
rect -5814 298658 -5578 298894
rect -5494 298658 -5258 298894
rect -5814 298338 -5578 298574
rect -5494 298338 -5258 298574
rect -5814 262658 -5578 262894
rect -5494 262658 -5258 262894
rect -5814 262338 -5578 262574
rect -5494 262338 -5258 262574
rect -5814 226658 -5578 226894
rect -5494 226658 -5258 226894
rect -5814 226338 -5578 226574
rect -5494 226338 -5258 226574
rect -5814 190658 -5578 190894
rect -5494 190658 -5258 190894
rect -5814 190338 -5578 190574
rect -5494 190338 -5258 190574
rect -5814 154658 -5578 154894
rect -5494 154658 -5258 154894
rect -5814 154338 -5578 154574
rect -5494 154338 -5258 154574
rect -5814 118658 -5578 118894
rect -5494 118658 -5258 118894
rect -5814 118338 -5578 118574
rect -5494 118338 -5258 118574
rect -5814 82658 -5578 82894
rect -5494 82658 -5258 82894
rect -5814 82338 -5578 82574
rect -5494 82338 -5258 82574
rect -5814 46658 -5578 46894
rect -5494 46658 -5258 46894
rect -5814 46338 -5578 46574
rect -5494 46338 -5258 46574
rect -5814 10658 -5578 10894
rect -5494 10658 -5258 10894
rect -5814 10338 -5578 10574
rect -5494 10338 -5258 10574
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 672938 -4618 673174
rect -4534 672938 -4298 673174
rect -4854 672618 -4618 672854
rect -4534 672618 -4298 672854
rect -4854 636938 -4618 637174
rect -4534 636938 -4298 637174
rect -4854 636618 -4618 636854
rect -4534 636618 -4298 636854
rect -4854 600938 -4618 601174
rect -4534 600938 -4298 601174
rect -4854 600618 -4618 600854
rect -4534 600618 -4298 600854
rect -4854 564938 -4618 565174
rect -4534 564938 -4298 565174
rect -4854 564618 -4618 564854
rect -4534 564618 -4298 564854
rect -4854 528938 -4618 529174
rect -4534 528938 -4298 529174
rect -4854 528618 -4618 528854
rect -4534 528618 -4298 528854
rect -4854 492938 -4618 493174
rect -4534 492938 -4298 493174
rect -4854 492618 -4618 492854
rect -4534 492618 -4298 492854
rect -4854 456938 -4618 457174
rect -4534 456938 -4298 457174
rect -4854 456618 -4618 456854
rect -4534 456618 -4298 456854
rect -4854 420938 -4618 421174
rect -4534 420938 -4298 421174
rect -4854 420618 -4618 420854
rect -4534 420618 -4298 420854
rect -4854 384938 -4618 385174
rect -4534 384938 -4298 385174
rect -4854 384618 -4618 384854
rect -4534 384618 -4298 384854
rect -4854 348938 -4618 349174
rect -4534 348938 -4298 349174
rect -4854 348618 -4618 348854
rect -4534 348618 -4298 348854
rect -4854 312938 -4618 313174
rect -4534 312938 -4298 313174
rect -4854 312618 -4618 312854
rect -4534 312618 -4298 312854
rect -4854 276938 -4618 277174
rect -4534 276938 -4298 277174
rect -4854 276618 -4618 276854
rect -4534 276618 -4298 276854
rect -4854 240938 -4618 241174
rect -4534 240938 -4298 241174
rect -4854 240618 -4618 240854
rect -4534 240618 -4298 240854
rect -4854 204938 -4618 205174
rect -4534 204938 -4298 205174
rect -4854 204618 -4618 204854
rect -4534 204618 -4298 204854
rect -4854 168938 -4618 169174
rect -4534 168938 -4298 169174
rect -4854 168618 -4618 168854
rect -4534 168618 -4298 168854
rect -4854 132938 -4618 133174
rect -4534 132938 -4298 133174
rect -4854 132618 -4618 132854
rect -4534 132618 -4298 132854
rect -4854 96938 -4618 97174
rect -4534 96938 -4298 97174
rect -4854 96618 -4618 96854
rect -4534 96618 -4298 96854
rect -4854 60938 -4618 61174
rect -4534 60938 -4298 61174
rect -4854 60618 -4618 60854
rect -4534 60618 -4298 60854
rect -4854 24938 -4618 25174
rect -4534 24938 -4298 25174
rect -4854 24618 -4618 24854
rect -4534 24618 -4298 24854
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect 5546 706522 5782 706758
rect 5866 706522 6102 706758
rect 5546 706202 5782 706438
rect 5866 706202 6102 706438
rect -3894 690938 -3658 691174
rect -3574 690938 -3338 691174
rect -3894 690618 -3658 690854
rect -3574 690618 -3338 690854
rect -3894 654938 -3658 655174
rect -3574 654938 -3338 655174
rect -3894 654618 -3658 654854
rect -3574 654618 -3338 654854
rect -3894 618938 -3658 619174
rect -3574 618938 -3338 619174
rect -3894 618618 -3658 618854
rect -3574 618618 -3338 618854
rect -3894 582938 -3658 583174
rect -3574 582938 -3338 583174
rect -3894 582618 -3658 582854
rect -3574 582618 -3338 582854
rect -3894 546938 -3658 547174
rect -3574 546938 -3338 547174
rect -3894 546618 -3658 546854
rect -3574 546618 -3338 546854
rect -3894 510938 -3658 511174
rect -3574 510938 -3338 511174
rect -3894 510618 -3658 510854
rect -3574 510618 -3338 510854
rect -3894 474938 -3658 475174
rect -3574 474938 -3338 475174
rect -3894 474618 -3658 474854
rect -3574 474618 -3338 474854
rect -3894 438938 -3658 439174
rect -3574 438938 -3338 439174
rect -3894 438618 -3658 438854
rect -3574 438618 -3338 438854
rect -3894 402938 -3658 403174
rect -3574 402938 -3338 403174
rect -3894 402618 -3658 402854
rect -3574 402618 -3338 402854
rect -3894 366938 -3658 367174
rect -3574 366938 -3338 367174
rect -3894 366618 -3658 366854
rect -3574 366618 -3338 366854
rect -3894 330938 -3658 331174
rect -3574 330938 -3338 331174
rect -3894 330618 -3658 330854
rect -3574 330618 -3338 330854
rect -3894 294938 -3658 295174
rect -3574 294938 -3338 295174
rect -3894 294618 -3658 294854
rect -3574 294618 -3338 294854
rect -3894 258938 -3658 259174
rect -3574 258938 -3338 259174
rect -3894 258618 -3658 258854
rect -3574 258618 -3338 258854
rect -3894 222938 -3658 223174
rect -3574 222938 -3338 223174
rect -3894 222618 -3658 222854
rect -3574 222618 -3338 222854
rect -3894 186938 -3658 187174
rect -3574 186938 -3338 187174
rect -3894 186618 -3658 186854
rect -3574 186618 -3338 186854
rect -3894 150938 -3658 151174
rect -3574 150938 -3338 151174
rect -3894 150618 -3658 150854
rect -3574 150618 -3338 150854
rect -3894 114938 -3658 115174
rect -3574 114938 -3338 115174
rect -3894 114618 -3658 114854
rect -3574 114618 -3338 114854
rect -3894 78938 -3658 79174
rect -3574 78938 -3338 79174
rect -3894 78618 -3658 78854
rect -3574 78618 -3338 78854
rect -3894 42938 -3658 43174
rect -3574 42938 -3338 43174
rect -3894 42618 -3658 42854
rect -3574 42618 -3338 42854
rect -3894 6938 -3658 7174
rect -3574 6938 -3338 7174
rect -3894 6618 -3658 6854
rect -3574 6618 -3338 6854
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 669218 -2698 669454
rect -2614 669218 -2378 669454
rect -2934 668898 -2698 669134
rect -2614 668898 -2378 669134
rect -2934 633218 -2698 633454
rect -2614 633218 -2378 633454
rect -2934 632898 -2698 633134
rect -2614 632898 -2378 633134
rect -2934 597218 -2698 597454
rect -2614 597218 -2378 597454
rect -2934 596898 -2698 597134
rect -2614 596898 -2378 597134
rect -2934 561218 -2698 561454
rect -2614 561218 -2378 561454
rect -2934 560898 -2698 561134
rect -2614 560898 -2378 561134
rect -2934 525218 -2698 525454
rect -2614 525218 -2378 525454
rect -2934 524898 -2698 525134
rect -2614 524898 -2378 525134
rect -2934 489218 -2698 489454
rect -2614 489218 -2378 489454
rect -2934 488898 -2698 489134
rect -2614 488898 -2378 489134
rect -2934 453218 -2698 453454
rect -2614 453218 -2378 453454
rect -2934 452898 -2698 453134
rect -2614 452898 -2378 453134
rect -2934 417218 -2698 417454
rect -2614 417218 -2378 417454
rect -2934 416898 -2698 417134
rect -2614 416898 -2378 417134
rect -2934 381218 -2698 381454
rect -2614 381218 -2378 381454
rect -2934 380898 -2698 381134
rect -2614 380898 -2378 381134
rect -2934 345218 -2698 345454
rect -2614 345218 -2378 345454
rect -2934 344898 -2698 345134
rect -2614 344898 -2378 345134
rect -2934 309218 -2698 309454
rect -2614 309218 -2378 309454
rect -2934 308898 -2698 309134
rect -2614 308898 -2378 309134
rect -2934 273218 -2698 273454
rect -2614 273218 -2378 273454
rect -2934 272898 -2698 273134
rect -2614 272898 -2378 273134
rect -2934 237218 -2698 237454
rect -2614 237218 -2378 237454
rect -2934 236898 -2698 237134
rect -2614 236898 -2378 237134
rect -2934 201218 -2698 201454
rect -2614 201218 -2378 201454
rect -2934 200898 -2698 201134
rect -2614 200898 -2378 201134
rect -2934 165218 -2698 165454
rect -2614 165218 -2378 165454
rect -2934 164898 -2698 165134
rect -2614 164898 -2378 165134
rect -2934 129218 -2698 129454
rect -2614 129218 -2378 129454
rect -2934 128898 -2698 129134
rect -2614 128898 -2378 129134
rect -2934 93218 -2698 93454
rect -2614 93218 -2378 93454
rect -2934 92898 -2698 93134
rect -2614 92898 -2378 93134
rect -2934 57218 -2698 57454
rect -2614 57218 -2378 57454
rect -2934 56898 -2698 57134
rect -2614 56898 -2378 57134
rect -2934 21218 -2698 21454
rect -2614 21218 -2378 21454
rect -2934 20898 -2698 21134
rect -2614 20898 -2378 21134
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect 5546 690938 5782 691174
rect 5866 690938 6102 691174
rect 5546 690618 5782 690854
rect 5866 690618 6102 690854
rect 5546 654938 5782 655174
rect 5866 654938 6102 655174
rect 5546 654618 5782 654854
rect 5866 654618 6102 654854
rect 5546 618938 5782 619174
rect 5866 618938 6102 619174
rect 5546 618618 5782 618854
rect 5866 618618 6102 618854
rect 5546 582938 5782 583174
rect 5866 582938 6102 583174
rect 5546 582618 5782 582854
rect 5866 582618 6102 582854
rect 5546 546938 5782 547174
rect 5866 546938 6102 547174
rect 5546 546618 5782 546854
rect 5866 546618 6102 546854
rect 5546 510938 5782 511174
rect 5866 510938 6102 511174
rect 5546 510618 5782 510854
rect 5866 510618 6102 510854
rect 5546 474938 5782 475174
rect 5866 474938 6102 475174
rect 5546 474618 5782 474854
rect 5866 474618 6102 474854
rect 5546 438938 5782 439174
rect 5866 438938 6102 439174
rect 5546 438618 5782 438854
rect 5866 438618 6102 438854
rect 5546 402938 5782 403174
rect 5866 402938 6102 403174
rect 5546 402618 5782 402854
rect 5866 402618 6102 402854
rect 5546 366938 5782 367174
rect 5866 366938 6102 367174
rect 5546 366618 5782 366854
rect 5866 366618 6102 366854
rect 5546 330938 5782 331174
rect 5866 330938 6102 331174
rect 5546 330618 5782 330854
rect 5866 330618 6102 330854
rect 5546 294938 5782 295174
rect 5866 294938 6102 295174
rect 5546 294618 5782 294854
rect 5866 294618 6102 294854
rect 5546 258938 5782 259174
rect 5866 258938 6102 259174
rect 5546 258618 5782 258854
rect 5866 258618 6102 258854
rect 5546 222938 5782 223174
rect 5866 222938 6102 223174
rect 5546 222618 5782 222854
rect 5866 222618 6102 222854
rect 5546 186938 5782 187174
rect 5866 186938 6102 187174
rect 5546 186618 5782 186854
rect 5866 186618 6102 186854
rect 5546 150938 5782 151174
rect 5866 150938 6102 151174
rect 5546 150618 5782 150854
rect 5866 150618 6102 150854
rect 5546 114938 5782 115174
rect 5866 114938 6102 115174
rect 5546 114618 5782 114854
rect 5866 114618 6102 114854
rect 5546 78938 5782 79174
rect 5866 78938 6102 79174
rect 5546 78618 5782 78854
rect 5866 78618 6102 78854
rect 5546 42938 5782 43174
rect 5866 42938 6102 43174
rect 5546 42618 5782 42854
rect 5866 42618 6102 42854
rect 5546 6938 5782 7174
rect 5866 6938 6102 7174
rect 5546 6618 5782 6854
rect 5866 6618 6102 6854
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect 5546 -2502 5782 -2266
rect 5866 -2502 6102 -2266
rect 5546 -2822 5782 -2586
rect 5866 -2822 6102 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect 9266 694658 9502 694894
rect 9586 694658 9822 694894
rect 9266 694338 9502 694574
rect 9586 694338 9822 694574
rect 9266 658658 9502 658894
rect 9586 658658 9822 658894
rect 9266 658338 9502 658574
rect 9586 658338 9822 658574
rect 9266 622658 9502 622894
rect 9586 622658 9822 622894
rect 9266 622338 9502 622574
rect 9586 622338 9822 622574
rect 9266 586658 9502 586894
rect 9586 586658 9822 586894
rect 9266 586338 9502 586574
rect 9586 586338 9822 586574
rect 9266 550658 9502 550894
rect 9586 550658 9822 550894
rect 9266 550338 9502 550574
rect 9586 550338 9822 550574
rect 9266 514658 9502 514894
rect 9586 514658 9822 514894
rect 9266 514338 9502 514574
rect 9586 514338 9822 514574
rect 9266 478658 9502 478894
rect 9586 478658 9822 478894
rect 9266 478338 9502 478574
rect 9586 478338 9822 478574
rect 9266 442658 9502 442894
rect 9586 442658 9822 442894
rect 9266 442338 9502 442574
rect 9586 442338 9822 442574
rect 9266 406658 9502 406894
rect 9586 406658 9822 406894
rect 9266 406338 9502 406574
rect 9586 406338 9822 406574
rect 9266 370658 9502 370894
rect 9586 370658 9822 370894
rect 9266 370338 9502 370574
rect 9586 370338 9822 370574
rect 9266 334658 9502 334894
rect 9586 334658 9822 334894
rect 9266 334338 9502 334574
rect 9586 334338 9822 334574
rect 9266 298658 9502 298894
rect 9586 298658 9822 298894
rect 9266 298338 9502 298574
rect 9586 298338 9822 298574
rect 9266 262658 9502 262894
rect 9586 262658 9822 262894
rect 9266 262338 9502 262574
rect 9586 262338 9822 262574
rect 9266 226658 9502 226894
rect 9586 226658 9822 226894
rect 9266 226338 9502 226574
rect 9586 226338 9822 226574
rect 9266 190658 9502 190894
rect 9586 190658 9822 190894
rect 9266 190338 9502 190574
rect 9586 190338 9822 190574
rect 9266 154658 9502 154894
rect 9586 154658 9822 154894
rect 9266 154338 9502 154574
rect 9586 154338 9822 154574
rect 9266 118658 9502 118894
rect 9586 118658 9822 118894
rect 9266 118338 9502 118574
rect 9586 118338 9822 118574
rect 9266 82658 9502 82894
rect 9586 82658 9822 82894
rect 9266 82338 9502 82574
rect 9586 82338 9822 82574
rect 9266 46658 9502 46894
rect 9586 46658 9822 46894
rect 9266 46338 9502 46574
rect 9586 46338 9822 46574
rect 9266 10658 9502 10894
rect 9586 10658 9822 10894
rect 9266 10338 9502 10574
rect 9586 10338 9822 10574
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect 9266 -4422 9502 -4186
rect 9586 -4422 9822 -4186
rect 9266 -4742 9502 -4506
rect 9586 -4742 9822 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect 30986 711322 31222 711558
rect 31306 711322 31542 711558
rect 30986 711002 31222 711238
rect 31306 711002 31542 711238
rect 27266 709402 27502 709638
rect 27586 709402 27822 709638
rect 27266 709082 27502 709318
rect 27586 709082 27822 709318
rect 23546 707482 23782 707718
rect 23866 707482 24102 707718
rect 23546 707162 23782 707398
rect 23866 707162 24102 707398
rect 12986 698378 13222 698614
rect 13306 698378 13542 698614
rect 12986 698058 13222 698294
rect 13306 698058 13542 698294
rect 12986 662378 13222 662614
rect 13306 662378 13542 662614
rect 12986 662058 13222 662294
rect 13306 662058 13542 662294
rect 12986 626378 13222 626614
rect 13306 626378 13542 626614
rect 12986 626058 13222 626294
rect 13306 626058 13542 626294
rect 12986 590378 13222 590614
rect 13306 590378 13542 590614
rect 12986 590058 13222 590294
rect 13306 590058 13542 590294
rect 12986 554378 13222 554614
rect 13306 554378 13542 554614
rect 12986 554058 13222 554294
rect 13306 554058 13542 554294
rect 12986 518378 13222 518614
rect 13306 518378 13542 518614
rect 12986 518058 13222 518294
rect 13306 518058 13542 518294
rect 12986 482378 13222 482614
rect 13306 482378 13542 482614
rect 12986 482058 13222 482294
rect 13306 482058 13542 482294
rect 12986 446378 13222 446614
rect 13306 446378 13542 446614
rect 12986 446058 13222 446294
rect 13306 446058 13542 446294
rect 12986 410378 13222 410614
rect 13306 410378 13542 410614
rect 12986 410058 13222 410294
rect 13306 410058 13542 410294
rect 12986 374378 13222 374614
rect 13306 374378 13542 374614
rect 12986 374058 13222 374294
rect 13306 374058 13542 374294
rect 12986 338378 13222 338614
rect 13306 338378 13542 338614
rect 12986 338058 13222 338294
rect 13306 338058 13542 338294
rect 12986 302378 13222 302614
rect 13306 302378 13542 302614
rect 12986 302058 13222 302294
rect 13306 302058 13542 302294
rect 12986 266378 13222 266614
rect 13306 266378 13542 266614
rect 12986 266058 13222 266294
rect 13306 266058 13542 266294
rect 12986 230378 13222 230614
rect 13306 230378 13542 230614
rect 12986 230058 13222 230294
rect 13306 230058 13542 230294
rect 12986 194378 13222 194614
rect 13306 194378 13542 194614
rect 12986 194058 13222 194294
rect 13306 194058 13542 194294
rect 12986 158378 13222 158614
rect 13306 158378 13542 158614
rect 12986 158058 13222 158294
rect 13306 158058 13542 158294
rect 12986 122378 13222 122614
rect 13306 122378 13542 122614
rect 12986 122058 13222 122294
rect 13306 122058 13542 122294
rect 12986 86378 13222 86614
rect 13306 86378 13542 86614
rect 12986 86058 13222 86294
rect 13306 86058 13542 86294
rect 12986 50378 13222 50614
rect 13306 50378 13542 50614
rect 12986 50058 13222 50294
rect 13306 50058 13542 50294
rect 12986 14378 13222 14614
rect 13306 14378 13542 14614
rect 12986 14058 13222 14294
rect 13306 14058 13542 14294
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect 19826 705562 20062 705798
rect 20146 705562 20382 705798
rect 19826 705242 20062 705478
rect 20146 705242 20382 705478
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -1542 20062 -1306
rect 20146 -1542 20382 -1306
rect 19826 -1862 20062 -1626
rect 20146 -1862 20382 -1626
rect 23546 672938 23782 673174
rect 23866 672938 24102 673174
rect 23546 672618 23782 672854
rect 23866 672618 24102 672854
rect 23546 636938 23782 637174
rect 23866 636938 24102 637174
rect 23546 636618 23782 636854
rect 23866 636618 24102 636854
rect 23546 600938 23782 601174
rect 23866 600938 24102 601174
rect 23546 600618 23782 600854
rect 23866 600618 24102 600854
rect 23546 564938 23782 565174
rect 23866 564938 24102 565174
rect 23546 564618 23782 564854
rect 23866 564618 24102 564854
rect 23546 528938 23782 529174
rect 23866 528938 24102 529174
rect 23546 528618 23782 528854
rect 23866 528618 24102 528854
rect 23546 492938 23782 493174
rect 23866 492938 24102 493174
rect 23546 492618 23782 492854
rect 23866 492618 24102 492854
rect 23546 456938 23782 457174
rect 23866 456938 24102 457174
rect 23546 456618 23782 456854
rect 23866 456618 24102 456854
rect 23546 420938 23782 421174
rect 23866 420938 24102 421174
rect 23546 420618 23782 420854
rect 23866 420618 24102 420854
rect 23546 384938 23782 385174
rect 23866 384938 24102 385174
rect 23546 384618 23782 384854
rect 23866 384618 24102 384854
rect 23546 348938 23782 349174
rect 23866 348938 24102 349174
rect 23546 348618 23782 348854
rect 23866 348618 24102 348854
rect 23546 312938 23782 313174
rect 23866 312938 24102 313174
rect 23546 312618 23782 312854
rect 23866 312618 24102 312854
rect 23546 276938 23782 277174
rect 23866 276938 24102 277174
rect 23546 276618 23782 276854
rect 23866 276618 24102 276854
rect 23546 240938 23782 241174
rect 23866 240938 24102 241174
rect 23546 240618 23782 240854
rect 23866 240618 24102 240854
rect 23546 204938 23782 205174
rect 23866 204938 24102 205174
rect 23546 204618 23782 204854
rect 23866 204618 24102 204854
rect 23546 168938 23782 169174
rect 23866 168938 24102 169174
rect 23546 168618 23782 168854
rect 23866 168618 24102 168854
rect 23546 132938 23782 133174
rect 23866 132938 24102 133174
rect 23546 132618 23782 132854
rect 23866 132618 24102 132854
rect 23546 96938 23782 97174
rect 23866 96938 24102 97174
rect 23546 96618 23782 96854
rect 23866 96618 24102 96854
rect 23546 60938 23782 61174
rect 23866 60938 24102 61174
rect 23546 60618 23782 60854
rect 23866 60618 24102 60854
rect 23546 24938 23782 25174
rect 23866 24938 24102 25174
rect 23546 24618 23782 24854
rect 23866 24618 24102 24854
rect 23546 -3462 23782 -3226
rect 23866 -3462 24102 -3226
rect 23546 -3782 23782 -3546
rect 23866 -3782 24102 -3546
rect 27266 676658 27502 676894
rect 27586 676658 27822 676894
rect 27266 676338 27502 676574
rect 27586 676338 27822 676574
rect 27266 640658 27502 640894
rect 27586 640658 27822 640894
rect 27266 640338 27502 640574
rect 27586 640338 27822 640574
rect 27266 604658 27502 604894
rect 27586 604658 27822 604894
rect 27266 604338 27502 604574
rect 27586 604338 27822 604574
rect 27266 568658 27502 568894
rect 27586 568658 27822 568894
rect 27266 568338 27502 568574
rect 27586 568338 27822 568574
rect 27266 532658 27502 532894
rect 27586 532658 27822 532894
rect 27266 532338 27502 532574
rect 27586 532338 27822 532574
rect 27266 496658 27502 496894
rect 27586 496658 27822 496894
rect 27266 496338 27502 496574
rect 27586 496338 27822 496574
rect 27266 460658 27502 460894
rect 27586 460658 27822 460894
rect 27266 460338 27502 460574
rect 27586 460338 27822 460574
rect 27266 424658 27502 424894
rect 27586 424658 27822 424894
rect 27266 424338 27502 424574
rect 27586 424338 27822 424574
rect 27266 388658 27502 388894
rect 27586 388658 27822 388894
rect 27266 388338 27502 388574
rect 27586 388338 27822 388574
rect 27266 352658 27502 352894
rect 27586 352658 27822 352894
rect 27266 352338 27502 352574
rect 27586 352338 27822 352574
rect 27266 316658 27502 316894
rect 27586 316658 27822 316894
rect 27266 316338 27502 316574
rect 27586 316338 27822 316574
rect 27266 280658 27502 280894
rect 27586 280658 27822 280894
rect 27266 280338 27502 280574
rect 27586 280338 27822 280574
rect 27266 244658 27502 244894
rect 27586 244658 27822 244894
rect 27266 244338 27502 244574
rect 27586 244338 27822 244574
rect 27266 208658 27502 208894
rect 27586 208658 27822 208894
rect 27266 208338 27502 208574
rect 27586 208338 27822 208574
rect 27266 172658 27502 172894
rect 27586 172658 27822 172894
rect 27266 172338 27502 172574
rect 27586 172338 27822 172574
rect 27266 136658 27502 136894
rect 27586 136658 27822 136894
rect 27266 136338 27502 136574
rect 27586 136338 27822 136574
rect 27266 100658 27502 100894
rect 27586 100658 27822 100894
rect 27266 100338 27502 100574
rect 27586 100338 27822 100574
rect 27266 64658 27502 64894
rect 27586 64658 27822 64894
rect 27266 64338 27502 64574
rect 27586 64338 27822 64574
rect 27266 28658 27502 28894
rect 27586 28658 27822 28894
rect 27266 28338 27502 28574
rect 27586 28338 27822 28574
rect 27266 -5382 27502 -5146
rect 27586 -5382 27822 -5146
rect 27266 -5702 27502 -5466
rect 27586 -5702 27822 -5466
rect 48986 710362 49222 710598
rect 49306 710362 49542 710598
rect 48986 710042 49222 710278
rect 49306 710042 49542 710278
rect 45266 708442 45502 708678
rect 45586 708442 45822 708678
rect 45266 708122 45502 708358
rect 45586 708122 45822 708358
rect 41546 706522 41782 706758
rect 41866 706522 42102 706758
rect 41546 706202 41782 706438
rect 41866 706202 42102 706438
rect 30986 680378 31222 680614
rect 31306 680378 31542 680614
rect 30986 680058 31222 680294
rect 31306 680058 31542 680294
rect 30986 644378 31222 644614
rect 31306 644378 31542 644614
rect 30986 644058 31222 644294
rect 31306 644058 31542 644294
rect 30986 608378 31222 608614
rect 31306 608378 31542 608614
rect 30986 608058 31222 608294
rect 31306 608058 31542 608294
rect 30986 572378 31222 572614
rect 31306 572378 31542 572614
rect 30986 572058 31222 572294
rect 31306 572058 31542 572294
rect 30986 536378 31222 536614
rect 31306 536378 31542 536614
rect 30986 536058 31222 536294
rect 31306 536058 31542 536294
rect 30986 500378 31222 500614
rect 31306 500378 31542 500614
rect 30986 500058 31222 500294
rect 31306 500058 31542 500294
rect 30986 464378 31222 464614
rect 31306 464378 31542 464614
rect 30986 464058 31222 464294
rect 31306 464058 31542 464294
rect 30986 428378 31222 428614
rect 31306 428378 31542 428614
rect 30986 428058 31222 428294
rect 31306 428058 31542 428294
rect 30986 392378 31222 392614
rect 31306 392378 31542 392614
rect 30986 392058 31222 392294
rect 31306 392058 31542 392294
rect 30986 356378 31222 356614
rect 31306 356378 31542 356614
rect 30986 356058 31222 356294
rect 31306 356058 31542 356294
rect 30986 320378 31222 320614
rect 31306 320378 31542 320614
rect 30986 320058 31222 320294
rect 31306 320058 31542 320294
rect 30986 284378 31222 284614
rect 31306 284378 31542 284614
rect 30986 284058 31222 284294
rect 31306 284058 31542 284294
rect 30986 248378 31222 248614
rect 31306 248378 31542 248614
rect 30986 248058 31222 248294
rect 31306 248058 31542 248294
rect 30986 212378 31222 212614
rect 31306 212378 31542 212614
rect 30986 212058 31222 212294
rect 31306 212058 31542 212294
rect 30986 176378 31222 176614
rect 31306 176378 31542 176614
rect 30986 176058 31222 176294
rect 31306 176058 31542 176294
rect 30986 140378 31222 140614
rect 31306 140378 31542 140614
rect 30986 140058 31222 140294
rect 31306 140058 31542 140294
rect 30986 104378 31222 104614
rect 31306 104378 31542 104614
rect 30986 104058 31222 104294
rect 31306 104058 31542 104294
rect 30986 68378 31222 68614
rect 31306 68378 31542 68614
rect 30986 68058 31222 68294
rect 31306 68058 31542 68294
rect 30986 32378 31222 32614
rect 31306 32378 31542 32614
rect 30986 32058 31222 32294
rect 31306 32058 31542 32294
rect 12986 -6342 13222 -6106
rect 13306 -6342 13542 -6106
rect 12986 -6662 13222 -6426
rect 13306 -6662 13542 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 41546 690938 41782 691174
rect 41866 690938 42102 691174
rect 41546 690618 41782 690854
rect 41866 690618 42102 690854
rect 41546 654938 41782 655174
rect 41866 654938 42102 655174
rect 41546 654618 41782 654854
rect 41866 654618 42102 654854
rect 41546 618938 41782 619174
rect 41866 618938 42102 619174
rect 41546 618618 41782 618854
rect 41866 618618 42102 618854
rect 41546 582938 41782 583174
rect 41866 582938 42102 583174
rect 41546 582618 41782 582854
rect 41866 582618 42102 582854
rect 41546 546938 41782 547174
rect 41866 546938 42102 547174
rect 41546 546618 41782 546854
rect 41866 546618 42102 546854
rect 41546 510938 41782 511174
rect 41866 510938 42102 511174
rect 41546 510618 41782 510854
rect 41866 510618 42102 510854
rect 41546 474938 41782 475174
rect 41866 474938 42102 475174
rect 41546 474618 41782 474854
rect 41866 474618 42102 474854
rect 41546 438938 41782 439174
rect 41866 438938 42102 439174
rect 41546 438618 41782 438854
rect 41866 438618 42102 438854
rect 41546 402938 41782 403174
rect 41866 402938 42102 403174
rect 41546 402618 41782 402854
rect 41866 402618 42102 402854
rect 41546 366938 41782 367174
rect 41866 366938 42102 367174
rect 41546 366618 41782 366854
rect 41866 366618 42102 366854
rect 41546 330938 41782 331174
rect 41866 330938 42102 331174
rect 41546 330618 41782 330854
rect 41866 330618 42102 330854
rect 41546 294938 41782 295174
rect 41866 294938 42102 295174
rect 41546 294618 41782 294854
rect 41866 294618 42102 294854
rect 41546 258938 41782 259174
rect 41866 258938 42102 259174
rect 41546 258618 41782 258854
rect 41866 258618 42102 258854
rect 41546 222938 41782 223174
rect 41866 222938 42102 223174
rect 41546 222618 41782 222854
rect 41866 222618 42102 222854
rect 41546 186938 41782 187174
rect 41866 186938 42102 187174
rect 41546 186618 41782 186854
rect 41866 186618 42102 186854
rect 41546 150938 41782 151174
rect 41866 150938 42102 151174
rect 41546 150618 41782 150854
rect 41866 150618 42102 150854
rect 41546 114938 41782 115174
rect 41866 114938 42102 115174
rect 41546 114618 41782 114854
rect 41866 114618 42102 114854
rect 41546 78938 41782 79174
rect 41866 78938 42102 79174
rect 41546 78618 41782 78854
rect 41866 78618 42102 78854
rect 41546 42938 41782 43174
rect 41866 42938 42102 43174
rect 41546 42618 41782 42854
rect 41866 42618 42102 42854
rect 41546 6938 41782 7174
rect 41866 6938 42102 7174
rect 41546 6618 41782 6854
rect 41866 6618 42102 6854
rect 41546 -2502 41782 -2266
rect 41866 -2502 42102 -2266
rect 41546 -2822 41782 -2586
rect 41866 -2822 42102 -2586
rect 45266 694658 45502 694894
rect 45586 694658 45822 694894
rect 45266 694338 45502 694574
rect 45586 694338 45822 694574
rect 45266 658658 45502 658894
rect 45586 658658 45822 658894
rect 45266 658338 45502 658574
rect 45586 658338 45822 658574
rect 45266 622658 45502 622894
rect 45586 622658 45822 622894
rect 45266 622338 45502 622574
rect 45586 622338 45822 622574
rect 45266 586658 45502 586894
rect 45586 586658 45822 586894
rect 45266 586338 45502 586574
rect 45586 586338 45822 586574
rect 45266 550658 45502 550894
rect 45586 550658 45822 550894
rect 45266 550338 45502 550574
rect 45586 550338 45822 550574
rect 45266 514658 45502 514894
rect 45586 514658 45822 514894
rect 45266 514338 45502 514574
rect 45586 514338 45822 514574
rect 45266 478658 45502 478894
rect 45586 478658 45822 478894
rect 45266 478338 45502 478574
rect 45586 478338 45822 478574
rect 45266 442658 45502 442894
rect 45586 442658 45822 442894
rect 45266 442338 45502 442574
rect 45586 442338 45822 442574
rect 45266 406658 45502 406894
rect 45586 406658 45822 406894
rect 45266 406338 45502 406574
rect 45586 406338 45822 406574
rect 45266 370658 45502 370894
rect 45586 370658 45822 370894
rect 45266 370338 45502 370574
rect 45586 370338 45822 370574
rect 45266 334658 45502 334894
rect 45586 334658 45822 334894
rect 45266 334338 45502 334574
rect 45586 334338 45822 334574
rect 45266 298658 45502 298894
rect 45586 298658 45822 298894
rect 45266 298338 45502 298574
rect 45586 298338 45822 298574
rect 45266 262658 45502 262894
rect 45586 262658 45822 262894
rect 45266 262338 45502 262574
rect 45586 262338 45822 262574
rect 45266 226658 45502 226894
rect 45586 226658 45822 226894
rect 45266 226338 45502 226574
rect 45586 226338 45822 226574
rect 45266 190658 45502 190894
rect 45586 190658 45822 190894
rect 45266 190338 45502 190574
rect 45586 190338 45822 190574
rect 45266 154658 45502 154894
rect 45586 154658 45822 154894
rect 45266 154338 45502 154574
rect 45586 154338 45822 154574
rect 45266 118658 45502 118894
rect 45586 118658 45822 118894
rect 45266 118338 45502 118574
rect 45586 118338 45822 118574
rect 45266 82658 45502 82894
rect 45586 82658 45822 82894
rect 45266 82338 45502 82574
rect 45586 82338 45822 82574
rect 45266 46658 45502 46894
rect 45586 46658 45822 46894
rect 45266 46338 45502 46574
rect 45586 46338 45822 46574
rect 45266 10658 45502 10894
rect 45586 10658 45822 10894
rect 45266 10338 45502 10574
rect 45586 10338 45822 10574
rect 45266 -4422 45502 -4186
rect 45586 -4422 45822 -4186
rect 45266 -4742 45502 -4506
rect 45586 -4742 45822 -4506
rect 66986 711322 67222 711558
rect 67306 711322 67542 711558
rect 66986 711002 67222 711238
rect 67306 711002 67542 711238
rect 63266 709402 63502 709638
rect 63586 709402 63822 709638
rect 63266 709082 63502 709318
rect 63586 709082 63822 709318
rect 59546 707482 59782 707718
rect 59866 707482 60102 707718
rect 59546 707162 59782 707398
rect 59866 707162 60102 707398
rect 48986 698378 49222 698614
rect 49306 698378 49542 698614
rect 48986 698058 49222 698294
rect 49306 698058 49542 698294
rect 48986 662378 49222 662614
rect 49306 662378 49542 662614
rect 48986 662058 49222 662294
rect 49306 662058 49542 662294
rect 48986 626378 49222 626614
rect 49306 626378 49542 626614
rect 48986 626058 49222 626294
rect 49306 626058 49542 626294
rect 48986 590378 49222 590614
rect 49306 590378 49542 590614
rect 48986 590058 49222 590294
rect 49306 590058 49542 590294
rect 48986 554378 49222 554614
rect 49306 554378 49542 554614
rect 48986 554058 49222 554294
rect 49306 554058 49542 554294
rect 48986 518378 49222 518614
rect 49306 518378 49542 518614
rect 48986 518058 49222 518294
rect 49306 518058 49542 518294
rect 48986 482378 49222 482614
rect 49306 482378 49542 482614
rect 48986 482058 49222 482294
rect 49306 482058 49542 482294
rect 48986 446378 49222 446614
rect 49306 446378 49542 446614
rect 48986 446058 49222 446294
rect 49306 446058 49542 446294
rect 48986 410378 49222 410614
rect 49306 410378 49542 410614
rect 48986 410058 49222 410294
rect 49306 410058 49542 410294
rect 48986 374378 49222 374614
rect 49306 374378 49542 374614
rect 48986 374058 49222 374294
rect 49306 374058 49542 374294
rect 48986 338378 49222 338614
rect 49306 338378 49542 338614
rect 48986 338058 49222 338294
rect 49306 338058 49542 338294
rect 48986 302378 49222 302614
rect 49306 302378 49542 302614
rect 48986 302058 49222 302294
rect 49306 302058 49542 302294
rect 55826 705562 56062 705798
rect 56146 705562 56382 705798
rect 55826 705242 56062 705478
rect 56146 705242 56382 705478
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 55826 381218 56062 381454
rect 56146 381218 56382 381454
rect 55826 380898 56062 381134
rect 56146 380898 56382 381134
rect 55826 345218 56062 345454
rect 56146 345218 56382 345454
rect 55826 344898 56062 345134
rect 56146 344898 56382 345134
rect 55826 309218 56062 309454
rect 56146 309218 56382 309454
rect 55826 308898 56062 309134
rect 56146 308898 56382 309134
rect 48986 266378 49222 266614
rect 49306 266378 49542 266614
rect 48986 266058 49222 266294
rect 49306 266058 49542 266294
rect 48986 230378 49222 230614
rect 49306 230378 49542 230614
rect 48986 230058 49222 230294
rect 49306 230058 49542 230294
rect 48986 194378 49222 194614
rect 49306 194378 49542 194614
rect 48986 194058 49222 194294
rect 49306 194058 49542 194294
rect 48986 158378 49222 158614
rect 49306 158378 49542 158614
rect 48986 158058 49222 158294
rect 49306 158058 49542 158294
rect 48986 122378 49222 122614
rect 49306 122378 49542 122614
rect 48986 122058 49222 122294
rect 49306 122058 49542 122294
rect 48986 86378 49222 86614
rect 49306 86378 49542 86614
rect 48986 86058 49222 86294
rect 49306 86058 49542 86294
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 55826 237218 56062 237454
rect 56146 237218 56382 237454
rect 55826 236898 56062 237134
rect 56146 236898 56382 237134
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 48986 50378 49222 50614
rect 49306 50378 49542 50614
rect 48986 50058 49222 50294
rect 49306 50058 49542 50294
rect 48986 14378 49222 14614
rect 49306 14378 49542 14614
rect 48986 14058 49222 14294
rect 49306 14058 49542 14294
rect 30986 -7302 31222 -7066
rect 31306 -7302 31542 -7066
rect 30986 -7622 31222 -7386
rect 31306 -7622 31542 -7386
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -1542 56062 -1306
rect 56146 -1542 56382 -1306
rect 55826 -1862 56062 -1626
rect 56146 -1862 56382 -1626
rect 59546 672938 59782 673174
rect 59866 672938 60102 673174
rect 59546 672618 59782 672854
rect 59866 672618 60102 672854
rect 59546 636938 59782 637174
rect 59866 636938 60102 637174
rect 59546 636618 59782 636854
rect 59866 636618 60102 636854
rect 59546 600938 59782 601174
rect 59866 600938 60102 601174
rect 59546 600618 59782 600854
rect 59866 600618 60102 600854
rect 59546 564938 59782 565174
rect 59866 564938 60102 565174
rect 59546 564618 59782 564854
rect 59866 564618 60102 564854
rect 59546 528938 59782 529174
rect 59866 528938 60102 529174
rect 59546 528618 59782 528854
rect 59866 528618 60102 528854
rect 59546 492938 59782 493174
rect 59866 492938 60102 493174
rect 59546 492618 59782 492854
rect 59866 492618 60102 492854
rect 59546 456938 59782 457174
rect 59866 456938 60102 457174
rect 59546 456618 59782 456854
rect 59866 456618 60102 456854
rect 59546 420938 59782 421174
rect 59866 420938 60102 421174
rect 59546 420618 59782 420854
rect 59866 420618 60102 420854
rect 59546 384938 59782 385174
rect 59866 384938 60102 385174
rect 59546 384618 59782 384854
rect 59866 384618 60102 384854
rect 59546 348938 59782 349174
rect 59866 348938 60102 349174
rect 59546 348618 59782 348854
rect 59866 348618 60102 348854
rect 63266 676658 63502 676894
rect 63586 676658 63822 676894
rect 63266 676338 63502 676574
rect 63586 676338 63822 676574
rect 63266 640658 63502 640894
rect 63586 640658 63822 640894
rect 63266 640338 63502 640574
rect 63586 640338 63822 640574
rect 63266 604658 63502 604894
rect 63586 604658 63822 604894
rect 63266 604338 63502 604574
rect 63586 604338 63822 604574
rect 84986 710362 85222 710598
rect 85306 710362 85542 710598
rect 84986 710042 85222 710278
rect 85306 710042 85542 710278
rect 81266 708442 81502 708678
rect 81586 708442 81822 708678
rect 81266 708122 81502 708358
rect 81586 708122 81822 708358
rect 77546 706522 77782 706758
rect 77866 706522 78102 706758
rect 77546 706202 77782 706438
rect 77866 706202 78102 706438
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 66986 680378 67222 680614
rect 67306 680378 67542 680614
rect 66986 680058 67222 680294
rect 67306 680058 67542 680294
rect 66986 644378 67222 644614
rect 67306 644378 67542 644614
rect 66986 644058 67222 644294
rect 67306 644058 67542 644294
rect 66986 608378 67222 608614
rect 67306 608378 67542 608614
rect 66986 608058 67222 608294
rect 67306 608058 67542 608294
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 77546 690938 77782 691174
rect 77866 690938 78102 691174
rect 77546 690618 77782 690854
rect 77866 690618 78102 690854
rect 77546 654938 77782 655174
rect 77866 654938 78102 655174
rect 77546 654618 77782 654854
rect 77866 654618 78102 654854
rect 77546 618938 77782 619174
rect 77866 618938 78102 619174
rect 77546 618618 77782 618854
rect 77866 618618 78102 618854
rect 81266 694658 81502 694894
rect 81586 694658 81822 694894
rect 81266 694338 81502 694574
rect 81586 694338 81822 694574
rect 81266 658658 81502 658894
rect 81586 658658 81822 658894
rect 81266 658338 81502 658574
rect 81586 658338 81822 658574
rect 81266 622658 81502 622894
rect 81586 622658 81822 622894
rect 81266 622338 81502 622574
rect 81586 622338 81822 622574
rect 102986 711322 103222 711558
rect 103306 711322 103542 711558
rect 102986 711002 103222 711238
rect 103306 711002 103542 711238
rect 99266 709402 99502 709638
rect 99586 709402 99822 709638
rect 99266 709082 99502 709318
rect 99586 709082 99822 709318
rect 95546 707482 95782 707718
rect 95866 707482 96102 707718
rect 95546 707162 95782 707398
rect 95866 707162 96102 707398
rect 84986 698378 85222 698614
rect 85306 698378 85542 698614
rect 84986 698058 85222 698294
rect 85306 698058 85542 698294
rect 84986 662378 85222 662614
rect 85306 662378 85542 662614
rect 84986 662058 85222 662294
rect 85306 662058 85542 662294
rect 84986 626378 85222 626614
rect 85306 626378 85542 626614
rect 84986 626058 85222 626294
rect 85306 626058 85542 626294
rect 91826 705562 92062 705798
rect 92146 705562 92382 705798
rect 91826 705242 92062 705478
rect 92146 705242 92382 705478
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 91826 633218 92062 633454
rect 92146 633218 92382 633454
rect 91826 632898 92062 633134
rect 92146 632898 92382 633134
rect 91826 597218 92062 597454
rect 92146 597218 92382 597454
rect 91826 596898 92062 597134
rect 92146 596898 92382 597134
rect 72721 579218 72957 579454
rect 72721 578898 72957 579134
rect 78651 579218 78887 579454
rect 78651 578898 78887 579134
rect 84582 579218 84818 579454
rect 84582 578898 84818 579134
rect 63266 568658 63502 568894
rect 63586 568658 63822 568894
rect 63266 568338 63502 568574
rect 63586 568338 63822 568574
rect 75686 561218 75922 561454
rect 75686 560898 75922 561134
rect 81617 561218 81853 561454
rect 81617 560898 81853 561134
rect 63266 532658 63502 532894
rect 63586 532658 63822 532894
rect 63266 532338 63502 532574
rect 63586 532338 63822 532574
rect 66986 536378 67222 536614
rect 67306 536378 67542 536614
rect 66986 536058 67222 536294
rect 67306 536058 67542 536294
rect 63266 496658 63502 496894
rect 63586 496658 63822 496894
rect 63266 496338 63502 496574
rect 63586 496338 63822 496574
rect 63266 460658 63502 460894
rect 63586 460658 63822 460894
rect 63266 460338 63502 460574
rect 63586 460338 63822 460574
rect 63266 424658 63502 424894
rect 63586 424658 63822 424894
rect 63266 424338 63502 424574
rect 63586 424338 63822 424574
rect 72721 543218 72957 543454
rect 72721 542898 72957 543134
rect 78651 543218 78887 543454
rect 78651 542898 78887 543134
rect 84582 543218 84818 543454
rect 84582 542898 84818 543134
rect 66986 500378 67222 500614
rect 67306 500378 67542 500614
rect 66986 500058 67222 500294
rect 67306 500058 67542 500294
rect 66986 464378 67222 464614
rect 67306 464378 67542 464614
rect 66986 464058 67222 464294
rect 67306 464058 67542 464294
rect 63266 388658 63502 388894
rect 63586 388658 63822 388894
rect 63266 388338 63502 388574
rect 63586 388338 63822 388574
rect 63266 352658 63502 352894
rect 63586 352658 63822 352894
rect 63266 352338 63502 352574
rect 63586 352338 63822 352574
rect 59546 312938 59782 313174
rect 59866 312938 60102 313174
rect 59546 312618 59782 312854
rect 59866 312618 60102 312854
rect 59546 276938 59782 277174
rect 59866 276938 60102 277174
rect 59546 276618 59782 276854
rect 59866 276618 60102 276854
rect 59546 240938 59782 241174
rect 59866 240938 60102 241174
rect 59546 240618 59782 240854
rect 59866 240618 60102 240854
rect 59546 204938 59782 205174
rect 59866 204938 60102 205174
rect 59546 204618 59782 204854
rect 59866 204618 60102 204854
rect 59546 168938 59782 169174
rect 59866 168938 60102 169174
rect 59546 168618 59782 168854
rect 59866 168618 60102 168854
rect 59546 132938 59782 133174
rect 59866 132938 60102 133174
rect 59546 132618 59782 132854
rect 59866 132618 60102 132854
rect 59546 96938 59782 97174
rect 59866 96938 60102 97174
rect 59546 96618 59782 96854
rect 59866 96618 60102 96854
rect 63266 316658 63502 316894
rect 63586 316658 63822 316894
rect 63266 316338 63502 316574
rect 63586 316338 63822 316574
rect 63266 280658 63502 280894
rect 63586 280658 63822 280894
rect 63266 280338 63502 280574
rect 63586 280338 63822 280574
rect 63266 244658 63502 244894
rect 63586 244658 63822 244894
rect 63266 244338 63502 244574
rect 63586 244338 63822 244574
rect 66986 356378 67222 356614
rect 67306 356378 67542 356614
rect 66986 356058 67222 356294
rect 67306 356058 67542 356294
rect 73826 507218 74062 507454
rect 74146 507218 74382 507454
rect 73826 506898 74062 507134
rect 74146 506898 74382 507134
rect 73826 471218 74062 471454
rect 74146 471218 74382 471454
rect 73826 470898 74062 471134
rect 74146 470898 74382 471134
rect 77546 510938 77782 511174
rect 77866 510938 78102 511174
rect 77546 510618 77782 510854
rect 77866 510618 78102 510854
rect 77546 474938 77782 475174
rect 77866 474938 78102 475174
rect 77546 474618 77782 474854
rect 77866 474618 78102 474854
rect 81266 514658 81502 514894
rect 81586 514658 81822 514894
rect 81266 514338 81502 514574
rect 81586 514338 81822 514574
rect 81266 478658 81502 478894
rect 81586 478658 81822 478894
rect 81266 478338 81502 478574
rect 81586 478338 81822 478574
rect 84986 518378 85222 518614
rect 85306 518378 85542 518614
rect 84986 518058 85222 518294
rect 85306 518058 85542 518294
rect 84986 482378 85222 482614
rect 85306 482378 85542 482614
rect 84986 482058 85222 482294
rect 85306 482058 85542 482294
rect 63266 208658 63502 208894
rect 63586 208658 63822 208894
rect 63266 208338 63502 208574
rect 63586 208338 63822 208574
rect 63266 172658 63502 172894
rect 63586 172658 63822 172894
rect 63266 172338 63502 172574
rect 63586 172338 63822 172574
rect 63266 136658 63502 136894
rect 63586 136658 63822 136894
rect 63266 136338 63502 136574
rect 63586 136338 63822 136574
rect 63266 100658 63502 100894
rect 63586 100658 63822 100894
rect 63266 100338 63502 100574
rect 63586 100338 63822 100574
rect 59546 60938 59782 61174
rect 59866 60938 60102 61174
rect 59546 60618 59782 60854
rect 59866 60618 60102 60854
rect 59546 24938 59782 25174
rect 59866 24938 60102 25174
rect 59546 24618 59782 24854
rect 59866 24618 60102 24854
rect 59546 -3462 59782 -3226
rect 59866 -3462 60102 -3226
rect 59546 -3782 59782 -3546
rect 59866 -3782 60102 -3546
rect 63266 64658 63502 64894
rect 63586 64658 63822 64894
rect 63266 64338 63502 64574
rect 63586 64338 63822 64574
rect 66986 212378 67222 212614
rect 67306 212378 67542 212614
rect 66986 212058 67222 212294
rect 67306 212058 67542 212294
rect 66986 68378 67222 68614
rect 67306 68378 67542 68614
rect 66986 68058 67222 68294
rect 67306 68058 67542 68294
rect 63266 28658 63502 28894
rect 63586 28658 63822 28894
rect 63266 28338 63502 28574
rect 63586 28338 63822 28574
rect 63266 -5382 63502 -5146
rect 63586 -5382 63822 -5146
rect 63266 -5702 63502 -5466
rect 63586 -5702 63822 -5466
rect 73020 435218 73256 435454
rect 73020 434898 73256 435134
rect 88380 417218 88616 417454
rect 88380 416898 88616 417134
rect 73020 399218 73256 399454
rect 73020 398898 73256 399134
rect 95546 672938 95782 673174
rect 95866 672938 96102 673174
rect 95546 672618 95782 672854
rect 95866 672618 96102 672854
rect 95546 636938 95782 637174
rect 95866 636938 96102 637174
rect 95546 636618 95782 636854
rect 95866 636618 96102 636854
rect 95546 600938 95782 601174
rect 95866 600938 96102 601174
rect 95546 600618 95782 600854
rect 95866 600618 96102 600854
rect 91826 561218 92062 561454
rect 92146 561218 92382 561454
rect 91826 560898 92062 561134
rect 92146 560898 92382 561134
rect 91826 525218 92062 525454
rect 92146 525218 92382 525454
rect 91826 524898 92062 525134
rect 92146 524898 92382 525134
rect 91826 489218 92062 489454
rect 92146 489218 92382 489454
rect 91826 488898 92062 489134
rect 92146 488898 92382 489134
rect 91826 453218 92062 453454
rect 92146 453218 92382 453454
rect 91826 452898 92062 453134
rect 92146 452898 92382 453134
rect 95546 564938 95782 565174
rect 95866 564938 96102 565174
rect 95546 564618 95782 564854
rect 95866 564618 96102 564854
rect 95546 528938 95782 529174
rect 95866 528938 96102 529174
rect 95546 528618 95782 528854
rect 95866 528618 96102 528854
rect 95546 492938 95782 493174
rect 95866 492938 96102 493174
rect 95546 492618 95782 492854
rect 95866 492618 96102 492854
rect 73826 363218 74062 363454
rect 74146 363218 74382 363454
rect 73826 362898 74062 363134
rect 74146 362898 74382 363134
rect 73020 291218 73256 291454
rect 73020 290898 73256 291134
rect 73020 255218 73256 255454
rect 73020 254898 73256 255134
rect 77546 366938 77782 367174
rect 77866 366938 78102 367174
rect 77546 366618 77782 366854
rect 77866 366618 78102 366854
rect 81266 370658 81502 370894
rect 81586 370658 81822 370894
rect 81266 370338 81502 370574
rect 81586 370338 81822 370574
rect 73826 219218 74062 219454
rect 74146 219218 74382 219454
rect 73826 218898 74062 219134
rect 74146 218898 74382 219134
rect 84986 374378 85222 374614
rect 85306 374378 85542 374614
rect 84986 374058 85222 374294
rect 85306 374058 85542 374294
rect 84986 338378 85222 338614
rect 85306 338378 85542 338614
rect 84986 338058 85222 338294
rect 85306 338058 85542 338294
rect 81266 334658 81502 334894
rect 81586 334658 81822 334894
rect 81266 334338 81502 334574
rect 81586 334338 81822 334574
rect 77546 222938 77782 223174
rect 77866 222938 78102 223174
rect 77546 222618 77782 222854
rect 77866 222618 78102 222854
rect 73826 183218 74062 183454
rect 74146 183218 74382 183454
rect 73826 182898 74062 183134
rect 74146 182898 74382 183134
rect 77546 186938 77782 187174
rect 77866 186938 78102 187174
rect 77546 186618 77782 186854
rect 77866 186618 78102 186854
rect 91826 381218 92062 381454
rect 92146 381218 92382 381454
rect 91826 380898 92062 381134
rect 92146 380898 92382 381134
rect 91826 345218 92062 345454
rect 92146 345218 92382 345454
rect 91826 344898 92062 345134
rect 92146 344898 92382 345134
rect 99266 676658 99502 676894
rect 99586 676658 99822 676894
rect 99266 676338 99502 676574
rect 99586 676338 99822 676574
rect 99266 640658 99502 640894
rect 99586 640658 99822 640894
rect 99266 640338 99502 640574
rect 99586 640338 99822 640574
rect 99266 604658 99502 604894
rect 99586 604658 99822 604894
rect 99266 604338 99502 604574
rect 99586 604338 99822 604574
rect 99266 568658 99502 568894
rect 99586 568658 99822 568894
rect 99266 568338 99502 568574
rect 99586 568338 99822 568574
rect 99266 532658 99502 532894
rect 99586 532658 99822 532894
rect 99266 532338 99502 532574
rect 99586 532338 99822 532574
rect 99266 496658 99502 496894
rect 99586 496658 99822 496894
rect 99266 496338 99502 496574
rect 99586 496338 99822 496574
rect 120986 710362 121222 710598
rect 121306 710362 121542 710598
rect 120986 710042 121222 710278
rect 121306 710042 121542 710278
rect 117266 708442 117502 708678
rect 117586 708442 117822 708678
rect 117266 708122 117502 708358
rect 117586 708122 117822 708358
rect 113546 706522 113782 706758
rect 113866 706522 114102 706758
rect 113546 706202 113782 706438
rect 113866 706202 114102 706438
rect 102986 680378 103222 680614
rect 103306 680378 103542 680614
rect 102986 680058 103222 680294
rect 103306 680058 103542 680294
rect 102986 644378 103222 644614
rect 103306 644378 103542 644614
rect 102986 644058 103222 644294
rect 103306 644058 103542 644294
rect 102986 608378 103222 608614
rect 103306 608378 103542 608614
rect 102986 608058 103222 608294
rect 103306 608058 103542 608294
rect 102986 572378 103222 572614
rect 103306 572378 103542 572614
rect 102986 572058 103222 572294
rect 103306 572058 103542 572294
rect 102986 536378 103222 536614
rect 103306 536378 103542 536614
rect 102986 536058 103222 536294
rect 103306 536058 103542 536294
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 109826 615218 110062 615454
rect 110146 615218 110382 615454
rect 109826 614898 110062 615134
rect 110146 614898 110382 615134
rect 109826 579218 110062 579454
rect 110146 579218 110382 579454
rect 109826 578898 110062 579134
rect 110146 578898 110382 579134
rect 109826 543218 110062 543454
rect 110146 543218 110382 543454
rect 109826 542898 110062 543134
rect 110146 542898 110382 543134
rect 102986 500378 103222 500614
rect 103306 500378 103542 500614
rect 102986 500058 103222 500294
rect 103306 500058 103542 500294
rect 102986 464378 103222 464614
rect 103306 464378 103542 464614
rect 99266 460658 99502 460894
rect 99586 460658 99822 460894
rect 99266 460338 99502 460574
rect 99586 460338 99822 460574
rect 95546 456938 95782 457174
rect 95866 456938 96102 457174
rect 95546 456618 95782 456854
rect 95866 456618 96102 456854
rect 95546 384938 95782 385174
rect 95866 384938 96102 385174
rect 95546 384618 95782 384854
rect 95866 384618 96102 384854
rect 95546 348938 95782 349174
rect 95866 348938 96102 349174
rect 95546 348618 95782 348854
rect 95866 348618 96102 348854
rect 102986 464058 103222 464294
rect 103306 464058 103542 464294
rect 103740 435218 103976 435454
rect 103740 434898 103976 435134
rect 103740 399218 103976 399454
rect 103740 398898 103976 399134
rect 109826 507218 110062 507454
rect 110146 507218 110382 507454
rect 109826 506898 110062 507134
rect 110146 506898 110382 507134
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 99266 352658 99502 352894
rect 99586 352658 99822 352894
rect 99266 352338 99502 352574
rect 99586 352338 99822 352574
rect 102986 356378 103222 356614
rect 103306 356378 103542 356614
rect 102986 356058 103222 356294
rect 103306 356058 103542 356294
rect 113546 690938 113782 691174
rect 113866 690938 114102 691174
rect 113546 690618 113782 690854
rect 113866 690618 114102 690854
rect 113546 654938 113782 655174
rect 113866 654938 114102 655174
rect 113546 654618 113782 654854
rect 113866 654618 114102 654854
rect 113546 618938 113782 619174
rect 113866 618938 114102 619174
rect 113546 618618 113782 618854
rect 113866 618618 114102 618854
rect 113546 582938 113782 583174
rect 113866 582938 114102 583174
rect 113546 582618 113782 582854
rect 113866 582618 114102 582854
rect 113546 546938 113782 547174
rect 113866 546938 114102 547174
rect 113546 546618 113782 546854
rect 113866 546618 114102 546854
rect 113546 510938 113782 511174
rect 113866 510938 114102 511174
rect 113546 510618 113782 510854
rect 113866 510618 114102 510854
rect 113546 474938 113782 475174
rect 113866 474938 114102 475174
rect 113546 474618 113782 474854
rect 113866 474618 114102 474854
rect 117266 694658 117502 694894
rect 117586 694658 117822 694894
rect 117266 694338 117502 694574
rect 117586 694338 117822 694574
rect 117266 658658 117502 658894
rect 117586 658658 117822 658894
rect 117266 658338 117502 658574
rect 117586 658338 117822 658574
rect 117266 622658 117502 622894
rect 117586 622658 117822 622894
rect 117266 622338 117502 622574
rect 117586 622338 117822 622574
rect 117266 586658 117502 586894
rect 117586 586658 117822 586894
rect 117266 586338 117502 586574
rect 117586 586338 117822 586574
rect 117266 550658 117502 550894
rect 117586 550658 117822 550894
rect 117266 550338 117502 550574
rect 117586 550338 117822 550574
rect 117266 514658 117502 514894
rect 117586 514658 117822 514894
rect 117266 514338 117502 514574
rect 117586 514338 117822 514574
rect 117266 478658 117502 478894
rect 117586 478658 117822 478894
rect 117266 478338 117502 478574
rect 117586 478338 117822 478574
rect 109826 363218 110062 363454
rect 110146 363218 110382 363454
rect 109826 362898 110062 363134
rect 110146 362898 110382 363134
rect 138986 711322 139222 711558
rect 139306 711322 139542 711558
rect 138986 711002 139222 711238
rect 139306 711002 139542 711238
rect 135266 709402 135502 709638
rect 135586 709402 135822 709638
rect 135266 709082 135502 709318
rect 135586 709082 135822 709318
rect 131546 707482 131782 707718
rect 131866 707482 132102 707718
rect 131546 707162 131782 707398
rect 131866 707162 132102 707398
rect 120986 698378 121222 698614
rect 121306 698378 121542 698614
rect 120986 698058 121222 698294
rect 121306 698058 121542 698294
rect 120986 662378 121222 662614
rect 121306 662378 121542 662614
rect 120986 662058 121222 662294
rect 121306 662058 121542 662294
rect 120986 626378 121222 626614
rect 121306 626378 121542 626614
rect 120986 626058 121222 626294
rect 121306 626058 121542 626294
rect 120986 590378 121222 590614
rect 121306 590378 121542 590614
rect 120986 590058 121222 590294
rect 121306 590058 121542 590294
rect 127826 705562 128062 705798
rect 128146 705562 128382 705798
rect 127826 705242 128062 705478
rect 128146 705242 128382 705478
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 127826 597218 128062 597454
rect 128146 597218 128382 597454
rect 127826 596898 128062 597134
rect 128146 596898 128382 597134
rect 120986 554378 121222 554614
rect 121306 554378 121542 554614
rect 120986 554058 121222 554294
rect 121306 554058 121542 554294
rect 120986 518378 121222 518614
rect 121306 518378 121542 518614
rect 120986 518058 121222 518294
rect 121306 518058 121542 518294
rect 120986 482378 121222 482614
rect 121306 482378 121542 482614
rect 120986 482058 121222 482294
rect 121306 482058 121542 482294
rect 113546 366938 113782 367174
rect 113866 366938 114102 367174
rect 113546 366618 113782 366854
rect 113866 366618 114102 366854
rect 117266 370658 117502 370894
rect 117586 370658 117822 370894
rect 117266 370338 117502 370574
rect 117586 370338 117822 370574
rect 119100 417218 119336 417454
rect 119100 416898 119336 417134
rect 127826 561218 128062 561454
rect 128146 561218 128382 561454
rect 127826 560898 128062 561134
rect 128146 560898 128382 561134
rect 127826 525218 128062 525454
rect 128146 525218 128382 525454
rect 127826 524898 128062 525134
rect 128146 524898 128382 525134
rect 127826 489218 128062 489454
rect 128146 489218 128382 489454
rect 127826 488898 128062 489134
rect 128146 488898 128382 489134
rect 127826 453218 128062 453454
rect 128146 453218 128382 453454
rect 127826 452898 128062 453134
rect 128146 452898 128382 453134
rect 127826 417218 128062 417454
rect 128146 417218 128382 417454
rect 127826 416898 128062 417134
rect 128146 416898 128382 417134
rect 120986 374378 121222 374614
rect 121306 374378 121542 374614
rect 120986 374058 121222 374294
rect 121306 374058 121542 374294
rect 117266 334658 117502 334894
rect 117586 334658 117822 334894
rect 117266 334338 117502 334574
rect 117586 334338 117822 334574
rect 120986 338378 121222 338614
rect 121306 338378 121542 338614
rect 120986 338058 121222 338294
rect 121306 338058 121542 338294
rect 127826 381218 128062 381454
rect 128146 381218 128382 381454
rect 127826 380898 128062 381134
rect 128146 380898 128382 381134
rect 127826 345218 128062 345454
rect 128146 345218 128382 345454
rect 127826 344898 128062 345134
rect 128146 344898 128382 345134
rect 131546 672938 131782 673174
rect 131866 672938 132102 673174
rect 131546 672618 131782 672854
rect 131866 672618 132102 672854
rect 131546 636938 131782 637174
rect 131866 636938 132102 637174
rect 131546 636618 131782 636854
rect 131866 636618 132102 636854
rect 131546 600938 131782 601174
rect 131866 600938 132102 601174
rect 131546 600618 131782 600854
rect 131866 600618 132102 600854
rect 131546 564938 131782 565174
rect 131866 564938 132102 565174
rect 131546 564618 131782 564854
rect 131866 564618 132102 564854
rect 131546 528938 131782 529174
rect 131866 528938 132102 529174
rect 131546 528618 131782 528854
rect 131866 528618 132102 528854
rect 131546 492938 131782 493174
rect 131866 492938 132102 493174
rect 131546 492618 131782 492854
rect 131866 492618 132102 492854
rect 131546 456938 131782 457174
rect 131866 456938 132102 457174
rect 131546 456618 131782 456854
rect 131866 456618 132102 456854
rect 131546 420938 131782 421174
rect 131866 420938 132102 421174
rect 131546 420618 131782 420854
rect 131866 420618 132102 420854
rect 131546 384938 131782 385174
rect 131866 384938 132102 385174
rect 131546 384618 131782 384854
rect 131866 384618 132102 384854
rect 131546 348938 131782 349174
rect 131866 348938 132102 349174
rect 131546 348618 131782 348854
rect 131866 348618 132102 348854
rect 135266 676658 135502 676894
rect 135586 676658 135822 676894
rect 135266 676338 135502 676574
rect 135586 676338 135822 676574
rect 135266 640658 135502 640894
rect 135586 640658 135822 640894
rect 135266 640338 135502 640574
rect 135586 640338 135822 640574
rect 135266 604658 135502 604894
rect 135586 604658 135822 604894
rect 135266 604338 135502 604574
rect 135586 604338 135822 604574
rect 135266 568658 135502 568894
rect 135586 568658 135822 568894
rect 135266 568338 135502 568574
rect 135586 568338 135822 568574
rect 135266 532658 135502 532894
rect 135586 532658 135822 532894
rect 135266 532338 135502 532574
rect 135586 532338 135822 532574
rect 135266 496658 135502 496894
rect 135586 496658 135822 496894
rect 135266 496338 135502 496574
rect 135586 496338 135822 496574
rect 135266 460658 135502 460894
rect 135586 460658 135822 460894
rect 135266 460338 135502 460574
rect 135586 460338 135822 460574
rect 135266 424658 135502 424894
rect 135586 424658 135822 424894
rect 135266 424338 135502 424574
rect 135586 424338 135822 424574
rect 135266 388658 135502 388894
rect 135586 388658 135822 388894
rect 135266 388338 135502 388574
rect 135586 388338 135822 388574
rect 135266 352658 135502 352894
rect 135586 352658 135822 352894
rect 135266 352338 135502 352574
rect 135586 352338 135822 352574
rect 156986 710362 157222 710598
rect 157306 710362 157542 710598
rect 156986 710042 157222 710278
rect 157306 710042 157542 710278
rect 153266 708442 153502 708678
rect 153586 708442 153822 708678
rect 153266 708122 153502 708358
rect 153586 708122 153822 708358
rect 149546 706522 149782 706758
rect 149866 706522 150102 706758
rect 149546 706202 149782 706438
rect 149866 706202 150102 706438
rect 138986 680378 139222 680614
rect 139306 680378 139542 680614
rect 138986 680058 139222 680294
rect 139306 680058 139542 680294
rect 138986 644378 139222 644614
rect 139306 644378 139542 644614
rect 138986 644058 139222 644294
rect 139306 644058 139542 644294
rect 138986 608378 139222 608614
rect 139306 608378 139542 608614
rect 138986 608058 139222 608294
rect 139306 608058 139542 608294
rect 138986 572378 139222 572614
rect 139306 572378 139542 572614
rect 138986 572058 139222 572294
rect 139306 572058 139542 572294
rect 138986 536378 139222 536614
rect 139306 536378 139542 536614
rect 138986 536058 139222 536294
rect 139306 536058 139542 536294
rect 138986 500378 139222 500614
rect 139306 500378 139542 500614
rect 138986 500058 139222 500294
rect 139306 500058 139542 500294
rect 138986 464378 139222 464614
rect 139306 464378 139542 464614
rect 138986 464058 139222 464294
rect 139306 464058 139542 464294
rect 138986 428378 139222 428614
rect 139306 428378 139542 428614
rect 138986 428058 139222 428294
rect 139306 428058 139542 428294
rect 138986 392378 139222 392614
rect 139306 392378 139542 392614
rect 138986 392058 139222 392294
rect 139306 392058 139542 392294
rect 138986 356378 139222 356614
rect 139306 356378 139542 356614
rect 138986 356058 139222 356294
rect 139306 356058 139542 356294
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 145826 543218 146062 543454
rect 146146 543218 146382 543454
rect 145826 542898 146062 543134
rect 146146 542898 146382 543134
rect 145826 507218 146062 507454
rect 146146 507218 146382 507454
rect 145826 506898 146062 507134
rect 146146 506898 146382 507134
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 145826 435218 146062 435454
rect 146146 435218 146382 435454
rect 145826 434898 146062 435134
rect 146146 434898 146382 435134
rect 145826 399218 146062 399454
rect 146146 399218 146382 399454
rect 145826 398898 146062 399134
rect 146146 398898 146382 399134
rect 145826 363218 146062 363454
rect 146146 363218 146382 363454
rect 145826 362898 146062 363134
rect 146146 362898 146382 363134
rect 149546 690938 149782 691174
rect 149866 690938 150102 691174
rect 149546 690618 149782 690854
rect 149866 690618 150102 690854
rect 149546 654938 149782 655174
rect 149866 654938 150102 655174
rect 149546 654618 149782 654854
rect 149866 654618 150102 654854
rect 149546 618938 149782 619174
rect 149866 618938 150102 619174
rect 149546 618618 149782 618854
rect 149866 618618 150102 618854
rect 149546 582938 149782 583174
rect 149866 582938 150102 583174
rect 149546 582618 149782 582854
rect 149866 582618 150102 582854
rect 149546 546938 149782 547174
rect 149866 546938 150102 547174
rect 149546 546618 149782 546854
rect 149866 546618 150102 546854
rect 149546 510938 149782 511174
rect 149866 510938 150102 511174
rect 149546 510618 149782 510854
rect 149866 510618 150102 510854
rect 149546 474938 149782 475174
rect 149866 474938 150102 475174
rect 149546 474618 149782 474854
rect 149866 474618 150102 474854
rect 149546 438938 149782 439174
rect 149866 438938 150102 439174
rect 149546 438618 149782 438854
rect 149866 438618 150102 438854
rect 149546 402938 149782 403174
rect 149866 402938 150102 403174
rect 149546 402618 149782 402854
rect 149866 402618 150102 402854
rect 149546 366938 149782 367174
rect 149866 366938 150102 367174
rect 149546 366618 149782 366854
rect 149866 366618 150102 366854
rect 153266 694658 153502 694894
rect 153586 694658 153822 694894
rect 153266 694338 153502 694574
rect 153586 694338 153822 694574
rect 153266 658658 153502 658894
rect 153586 658658 153822 658894
rect 153266 658338 153502 658574
rect 153586 658338 153822 658574
rect 153266 622658 153502 622894
rect 153586 622658 153822 622894
rect 153266 622338 153502 622574
rect 153586 622338 153822 622574
rect 153266 586658 153502 586894
rect 153586 586658 153822 586894
rect 153266 586338 153502 586574
rect 153586 586338 153822 586574
rect 153266 550658 153502 550894
rect 153586 550658 153822 550894
rect 153266 550338 153502 550574
rect 153586 550338 153822 550574
rect 153266 514658 153502 514894
rect 153586 514658 153822 514894
rect 153266 514338 153502 514574
rect 153586 514338 153822 514574
rect 174986 711322 175222 711558
rect 175306 711322 175542 711558
rect 174986 711002 175222 711238
rect 175306 711002 175542 711238
rect 171266 709402 171502 709638
rect 171586 709402 171822 709638
rect 171266 709082 171502 709318
rect 171586 709082 171822 709318
rect 167546 707482 167782 707718
rect 167866 707482 168102 707718
rect 167546 707162 167782 707398
rect 167866 707162 168102 707398
rect 156986 698378 157222 698614
rect 157306 698378 157542 698614
rect 156986 698058 157222 698294
rect 157306 698058 157542 698294
rect 156986 662378 157222 662614
rect 157306 662378 157542 662614
rect 156986 662058 157222 662294
rect 157306 662058 157542 662294
rect 156986 626378 157222 626614
rect 157306 626378 157542 626614
rect 156986 626058 157222 626294
rect 157306 626058 157542 626294
rect 156986 590378 157222 590614
rect 157306 590378 157542 590614
rect 156986 590058 157222 590294
rect 157306 590058 157542 590294
rect 156986 554378 157222 554614
rect 157306 554378 157542 554614
rect 156986 554058 157222 554294
rect 157306 554058 157542 554294
rect 163826 705562 164062 705798
rect 164146 705562 164382 705798
rect 163826 705242 164062 705478
rect 164146 705242 164382 705478
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 163826 633218 164062 633454
rect 164146 633218 164382 633454
rect 163826 632898 164062 633134
rect 164146 632898 164382 633134
rect 163826 597218 164062 597454
rect 164146 597218 164382 597454
rect 163826 596898 164062 597134
rect 164146 596898 164382 597134
rect 163826 561218 164062 561454
rect 164146 561218 164382 561454
rect 163826 560898 164062 561134
rect 164146 560898 164382 561134
rect 156986 518378 157222 518614
rect 157306 518378 157542 518614
rect 156986 518058 157222 518294
rect 157306 518058 157542 518294
rect 153266 478658 153502 478894
rect 153586 478658 153822 478894
rect 153266 478338 153502 478574
rect 153586 478338 153822 478574
rect 153266 442658 153502 442894
rect 153586 442658 153822 442894
rect 153266 442338 153502 442574
rect 153586 442338 153822 442574
rect 153266 406658 153502 406894
rect 153586 406658 153822 406894
rect 153266 406338 153502 406574
rect 153586 406338 153822 406574
rect 153266 370658 153502 370894
rect 153586 370658 153822 370894
rect 153266 370338 153502 370574
rect 153586 370338 153822 370574
rect 153266 334658 153502 334894
rect 153586 334658 153822 334894
rect 153266 334338 153502 334574
rect 153586 334338 153822 334574
rect 88380 309218 88616 309454
rect 88380 308898 88616 309134
rect 119100 309218 119336 309454
rect 119100 308898 119336 309134
rect 149820 309218 150056 309454
rect 149820 308898 150056 309134
rect 103740 291218 103976 291454
rect 103740 290898 103976 291134
rect 134460 291218 134696 291454
rect 134460 290898 134696 291134
rect 88380 273218 88616 273454
rect 88380 272898 88616 273134
rect 119100 273218 119336 273454
rect 119100 272898 119336 273134
rect 149820 273218 150056 273454
rect 149820 272898 150056 273134
rect 103740 255218 103976 255454
rect 103740 254898 103976 255134
rect 134460 255218 134696 255454
rect 134460 254898 134696 255134
rect 84986 230378 85222 230614
rect 85306 230378 85542 230614
rect 84986 230058 85222 230294
rect 85306 230058 85542 230294
rect 81266 226658 81502 226894
rect 81586 226658 81822 226894
rect 81266 226338 81502 226574
rect 81586 226338 81822 226574
rect 81266 190658 81502 190894
rect 81586 190658 81822 190894
rect 81266 190338 81502 190574
rect 81586 190338 81822 190574
rect 84986 194378 85222 194614
rect 85306 194378 85542 194614
rect 84986 194058 85222 194294
rect 85306 194058 85542 194294
rect 91826 237218 92062 237454
rect 92146 237218 92382 237454
rect 91826 236898 92062 237134
rect 92146 236898 92382 237134
rect 91826 201218 92062 201454
rect 92146 201218 92382 201454
rect 91826 200898 92062 201134
rect 92146 200898 92382 201134
rect 95546 204938 95782 205174
rect 95866 204938 96102 205174
rect 95546 204618 95782 204854
rect 95866 204618 96102 204854
rect 99266 208658 99502 208894
rect 99586 208658 99822 208894
rect 99266 208338 99502 208574
rect 99586 208338 99822 208574
rect 102986 212378 103222 212614
rect 103306 212378 103542 212614
rect 102986 212058 103222 212294
rect 103306 212058 103542 212294
rect 109826 219218 110062 219454
rect 110146 219218 110382 219454
rect 109826 218898 110062 219134
rect 110146 218898 110382 219134
rect 109826 183218 110062 183454
rect 110146 183218 110382 183454
rect 109826 182898 110062 183134
rect 110146 182898 110382 183134
rect 113546 222938 113782 223174
rect 113866 222938 114102 223174
rect 113546 222618 113782 222854
rect 113866 222618 114102 222854
rect 113546 186938 113782 187174
rect 113866 186938 114102 187174
rect 113546 186618 113782 186854
rect 113866 186618 114102 186854
rect 117266 226658 117502 226894
rect 117586 226658 117822 226894
rect 117266 226338 117502 226574
rect 117586 226338 117822 226574
rect 117266 190658 117502 190894
rect 117586 190658 117822 190894
rect 117266 190338 117502 190574
rect 117586 190338 117822 190574
rect 120986 230378 121222 230614
rect 121306 230378 121542 230614
rect 120986 230058 121222 230294
rect 121306 230058 121542 230294
rect 120986 194378 121222 194614
rect 121306 194378 121542 194614
rect 120986 194058 121222 194294
rect 121306 194058 121542 194294
rect 127826 237218 128062 237454
rect 128146 237218 128382 237454
rect 127826 236898 128062 237134
rect 128146 236898 128382 237134
rect 127826 201218 128062 201454
rect 128146 201218 128382 201454
rect 127826 200898 128062 201134
rect 128146 200898 128382 201134
rect 131546 204938 131782 205174
rect 131866 204938 132102 205174
rect 131546 204618 131782 204854
rect 131866 204618 132102 204854
rect 135266 208658 135502 208894
rect 135586 208658 135822 208894
rect 135266 208338 135502 208574
rect 135586 208338 135822 208574
rect 138986 212378 139222 212614
rect 139306 212378 139542 212614
rect 138986 212058 139222 212294
rect 139306 212058 139542 212294
rect 145826 219218 146062 219454
rect 146146 219218 146382 219454
rect 145826 218898 146062 219134
rect 146146 218898 146382 219134
rect 145826 183218 146062 183454
rect 146146 183218 146382 183454
rect 145826 182898 146062 183134
rect 146146 182898 146382 183134
rect 149546 222938 149782 223174
rect 149866 222938 150102 223174
rect 149546 222618 149782 222854
rect 149866 222618 150102 222854
rect 149546 186938 149782 187174
rect 149866 186938 150102 187174
rect 149546 186618 149782 186854
rect 149866 186618 150102 186854
rect 156986 482378 157222 482614
rect 157306 482378 157542 482614
rect 156986 482058 157222 482294
rect 157306 482058 157542 482294
rect 156986 446378 157222 446614
rect 157306 446378 157542 446614
rect 156986 446058 157222 446294
rect 157306 446058 157542 446294
rect 156986 410378 157222 410614
rect 157306 410378 157542 410614
rect 156986 410058 157222 410294
rect 157306 410058 157542 410294
rect 156986 374378 157222 374614
rect 157306 374378 157542 374614
rect 156986 374058 157222 374294
rect 157306 374058 157542 374294
rect 156986 338378 157222 338614
rect 157306 338378 157542 338614
rect 156986 338058 157222 338294
rect 157306 338058 157542 338294
rect 153266 226658 153502 226894
rect 153586 226658 153822 226894
rect 153266 226338 153502 226574
rect 153586 226338 153822 226574
rect 153266 190658 153502 190894
rect 153586 190658 153822 190894
rect 153266 190338 153502 190574
rect 153586 190338 153822 190574
rect 163826 525218 164062 525454
rect 164146 525218 164382 525454
rect 163826 524898 164062 525134
rect 164146 524898 164382 525134
rect 163826 489218 164062 489454
rect 164146 489218 164382 489454
rect 163826 488898 164062 489134
rect 164146 488898 164382 489134
rect 163826 453218 164062 453454
rect 164146 453218 164382 453454
rect 163826 452898 164062 453134
rect 164146 452898 164382 453134
rect 163826 417218 164062 417454
rect 164146 417218 164382 417454
rect 163826 416898 164062 417134
rect 164146 416898 164382 417134
rect 167546 672938 167782 673174
rect 167866 672938 168102 673174
rect 167546 672618 167782 672854
rect 167866 672618 168102 672854
rect 167546 636938 167782 637174
rect 167866 636938 168102 637174
rect 167546 636618 167782 636854
rect 167866 636618 168102 636854
rect 167546 600938 167782 601174
rect 167866 600938 168102 601174
rect 167546 600618 167782 600854
rect 167866 600618 168102 600854
rect 167546 564938 167782 565174
rect 167866 564938 168102 565174
rect 167546 564618 167782 564854
rect 167866 564618 168102 564854
rect 171266 676658 171502 676894
rect 171586 676658 171822 676894
rect 171266 676338 171502 676574
rect 171586 676338 171822 676574
rect 171266 640658 171502 640894
rect 171586 640658 171822 640894
rect 171266 640338 171502 640574
rect 171586 640338 171822 640574
rect 171266 604658 171502 604894
rect 171586 604658 171822 604894
rect 171266 604338 171502 604574
rect 171586 604338 171822 604574
rect 171266 568658 171502 568894
rect 171586 568658 171822 568894
rect 171266 568338 171502 568574
rect 171586 568338 171822 568574
rect 167546 528938 167782 529174
rect 167866 528938 168102 529174
rect 167546 528618 167782 528854
rect 167866 528618 168102 528854
rect 167546 492938 167782 493174
rect 167866 492938 168102 493174
rect 167546 492618 167782 492854
rect 167866 492618 168102 492854
rect 167546 456938 167782 457174
rect 167866 456938 168102 457174
rect 167546 456618 167782 456854
rect 167866 456618 168102 456854
rect 167546 420938 167782 421174
rect 167866 420938 168102 421174
rect 167546 420618 167782 420854
rect 167866 420618 168102 420854
rect 163826 381218 164062 381454
rect 164146 381218 164382 381454
rect 163826 380898 164062 381134
rect 164146 380898 164382 381134
rect 163826 345218 164062 345454
rect 164146 345218 164382 345454
rect 163826 344898 164062 345134
rect 164146 344898 164382 345134
rect 163826 309218 164062 309454
rect 164146 309218 164382 309454
rect 163826 308898 164062 309134
rect 164146 308898 164382 309134
rect 156986 230378 157222 230614
rect 157306 230378 157542 230614
rect 156986 230058 157222 230294
rect 157306 230058 157542 230294
rect 163826 273218 164062 273454
rect 164146 273218 164382 273454
rect 163826 272898 164062 273134
rect 164146 272898 164382 273134
rect 163826 237218 164062 237454
rect 164146 237218 164382 237454
rect 163826 236898 164062 237134
rect 164146 236898 164382 237134
rect 156986 194378 157222 194614
rect 157306 194378 157542 194614
rect 156986 194058 157222 194294
rect 157306 194058 157542 194294
rect 163826 201218 164062 201454
rect 164146 201218 164382 201454
rect 163826 200898 164062 201134
rect 164146 200898 164382 201134
rect 69128 165218 69364 165454
rect 69128 164898 69364 165134
rect 164192 165218 164428 165454
rect 164192 164898 164428 165134
rect 69808 147218 70044 147454
rect 69808 146898 70044 147134
rect 163512 147218 163748 147454
rect 163512 146898 163748 147134
rect 69128 129218 69364 129454
rect 69128 128898 69364 129134
rect 164192 129218 164428 129454
rect 164192 128898 164428 129134
rect 69808 111218 70044 111454
rect 69808 110898 70044 111134
rect 163512 111218 163748 111454
rect 163512 110898 163748 111134
rect 73826 75218 74062 75454
rect 74146 75218 74382 75454
rect 73826 74898 74062 75134
rect 74146 74898 74382 75134
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 66986 32378 67222 32614
rect 67306 32378 67542 32614
rect 66986 32058 67222 32294
rect 67306 32058 67542 32294
rect 48986 -6342 49222 -6106
rect 49306 -6342 49542 -6106
rect 48986 -6662 49222 -6426
rect 49306 -6662 49542 -6426
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 77546 78938 77782 79174
rect 77866 78938 78102 79174
rect 77546 78618 77782 78854
rect 77866 78618 78102 78854
rect 77546 42938 77782 43174
rect 77866 42938 78102 43174
rect 77546 42618 77782 42854
rect 77866 42618 78102 42854
rect 77546 6938 77782 7174
rect 77866 6938 78102 7174
rect 77546 6618 77782 6854
rect 77866 6618 78102 6854
rect 77546 -2502 77782 -2266
rect 77866 -2502 78102 -2266
rect 77546 -2822 77782 -2586
rect 77866 -2822 78102 -2586
rect 81266 82658 81502 82894
rect 81586 82658 81822 82894
rect 81266 82338 81502 82574
rect 81586 82338 81822 82574
rect 81266 46658 81502 46894
rect 81586 46658 81822 46894
rect 81266 46338 81502 46574
rect 81586 46338 81822 46574
rect 81266 10658 81502 10894
rect 81586 10658 81822 10894
rect 81266 10338 81502 10574
rect 81586 10338 81822 10574
rect 81266 -4422 81502 -4186
rect 81586 -4422 81822 -4186
rect 81266 -4742 81502 -4506
rect 81586 -4742 81822 -4506
rect 84986 86378 85222 86614
rect 85306 86378 85542 86614
rect 84986 86058 85222 86294
rect 85306 86058 85542 86294
rect 84986 50378 85222 50614
rect 85306 50378 85542 50614
rect 84986 50058 85222 50294
rect 85306 50058 85542 50294
rect 84986 14378 85222 14614
rect 85306 14378 85542 14614
rect 84986 14058 85222 14294
rect 85306 14058 85542 14294
rect 66986 -7302 67222 -7066
rect 67306 -7302 67542 -7066
rect 66986 -7622 67222 -7386
rect 67306 -7622 67542 -7386
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -1542 92062 -1306
rect 92146 -1542 92382 -1306
rect 91826 -1862 92062 -1626
rect 92146 -1862 92382 -1626
rect 95546 60938 95782 61174
rect 95866 60938 96102 61174
rect 95546 60618 95782 60854
rect 95866 60618 96102 60854
rect 95546 24938 95782 25174
rect 95866 24938 96102 25174
rect 95546 24618 95782 24854
rect 95866 24618 96102 24854
rect 95546 -3462 95782 -3226
rect 95866 -3462 96102 -3226
rect 95546 -3782 95782 -3546
rect 95866 -3782 96102 -3546
rect 99266 64658 99502 64894
rect 99586 64658 99822 64894
rect 99266 64338 99502 64574
rect 99586 64338 99822 64574
rect 99266 28658 99502 28894
rect 99586 28658 99822 28894
rect 99266 28338 99502 28574
rect 99586 28338 99822 28574
rect 99266 -5382 99502 -5146
rect 99586 -5382 99822 -5146
rect 99266 -5702 99502 -5466
rect 99586 -5702 99822 -5466
rect 102986 68378 103222 68614
rect 103306 68378 103542 68614
rect 102986 68058 103222 68294
rect 103306 68058 103542 68294
rect 102986 32378 103222 32614
rect 103306 32378 103542 32614
rect 102986 32058 103222 32294
rect 103306 32058 103542 32294
rect 84986 -6342 85222 -6106
rect 85306 -6342 85542 -6106
rect 84986 -6662 85222 -6426
rect 85306 -6662 85542 -6426
rect 109826 75218 110062 75454
rect 110146 75218 110382 75454
rect 109826 74898 110062 75134
rect 110146 74898 110382 75134
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 113546 78938 113782 79174
rect 113866 78938 114102 79174
rect 113546 78618 113782 78854
rect 113866 78618 114102 78854
rect 113546 42938 113782 43174
rect 113866 42938 114102 43174
rect 113546 42618 113782 42854
rect 113866 42618 114102 42854
rect 113546 6938 113782 7174
rect 113866 6938 114102 7174
rect 113546 6618 113782 6854
rect 113866 6618 114102 6854
rect 113546 -2502 113782 -2266
rect 113866 -2502 114102 -2266
rect 113546 -2822 113782 -2586
rect 113866 -2822 114102 -2586
rect 117266 82658 117502 82894
rect 117586 82658 117822 82894
rect 117266 82338 117502 82574
rect 117586 82338 117822 82574
rect 117266 46658 117502 46894
rect 117586 46658 117822 46894
rect 117266 46338 117502 46574
rect 117586 46338 117822 46574
rect 117266 10658 117502 10894
rect 117586 10658 117822 10894
rect 117266 10338 117502 10574
rect 117586 10338 117822 10574
rect 117266 -4422 117502 -4186
rect 117586 -4422 117822 -4186
rect 117266 -4742 117502 -4506
rect 117586 -4742 117822 -4506
rect 120986 86378 121222 86614
rect 121306 86378 121542 86614
rect 120986 86058 121222 86294
rect 121306 86058 121542 86294
rect 120986 50378 121222 50614
rect 121306 50378 121542 50614
rect 120986 50058 121222 50294
rect 121306 50058 121542 50294
rect 120986 14378 121222 14614
rect 121306 14378 121542 14614
rect 120986 14058 121222 14294
rect 121306 14058 121542 14294
rect 102986 -7302 103222 -7066
rect 103306 -7302 103542 -7066
rect 102986 -7622 103222 -7386
rect 103306 -7622 103542 -7386
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -1542 128062 -1306
rect 128146 -1542 128382 -1306
rect 127826 -1862 128062 -1626
rect 128146 -1862 128382 -1626
rect 131546 60938 131782 61174
rect 131866 60938 132102 61174
rect 131546 60618 131782 60854
rect 131866 60618 132102 60854
rect 131546 24938 131782 25174
rect 131866 24938 132102 25174
rect 131546 24618 131782 24854
rect 131866 24618 132102 24854
rect 131546 -3462 131782 -3226
rect 131866 -3462 132102 -3226
rect 131546 -3782 131782 -3546
rect 131866 -3782 132102 -3546
rect 135266 64658 135502 64894
rect 135586 64658 135822 64894
rect 135266 64338 135502 64574
rect 135586 64338 135822 64574
rect 135266 28658 135502 28894
rect 135586 28658 135822 28894
rect 135266 28338 135502 28574
rect 135586 28338 135822 28574
rect 135266 -5382 135502 -5146
rect 135586 -5382 135822 -5146
rect 135266 -5702 135502 -5466
rect 135586 -5702 135822 -5466
rect 138986 68378 139222 68614
rect 139306 68378 139542 68614
rect 138986 68058 139222 68294
rect 139306 68058 139542 68294
rect 138986 32378 139222 32614
rect 139306 32378 139542 32614
rect 138986 32058 139222 32294
rect 139306 32058 139542 32294
rect 120986 -6342 121222 -6106
rect 121306 -6342 121542 -6106
rect 120986 -6662 121222 -6426
rect 121306 -6662 121542 -6426
rect 145826 75218 146062 75454
rect 146146 75218 146382 75454
rect 145826 74898 146062 75134
rect 146146 74898 146382 75134
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 149546 78938 149782 79174
rect 149866 78938 150102 79174
rect 149546 78618 149782 78854
rect 149866 78618 150102 78854
rect 149546 42938 149782 43174
rect 149866 42938 150102 43174
rect 149546 42618 149782 42854
rect 149866 42618 150102 42854
rect 149546 6938 149782 7174
rect 149866 6938 150102 7174
rect 149546 6618 149782 6854
rect 149866 6618 150102 6854
rect 149546 -2502 149782 -2266
rect 149866 -2502 150102 -2266
rect 149546 -2822 149782 -2586
rect 149866 -2822 150102 -2586
rect 153266 82658 153502 82894
rect 153586 82658 153822 82894
rect 153266 82338 153502 82574
rect 153586 82338 153822 82574
rect 153266 46658 153502 46894
rect 153586 46658 153822 46894
rect 153266 46338 153502 46574
rect 153586 46338 153822 46574
rect 153266 10658 153502 10894
rect 153586 10658 153822 10894
rect 153266 10338 153502 10574
rect 153586 10338 153822 10574
rect 153266 -4422 153502 -4186
rect 153586 -4422 153822 -4186
rect 153266 -4742 153502 -4506
rect 153586 -4742 153822 -4506
rect 156986 86378 157222 86614
rect 157306 86378 157542 86614
rect 156986 86058 157222 86294
rect 157306 86058 157542 86294
rect 156986 50378 157222 50614
rect 157306 50378 157542 50614
rect 156986 50058 157222 50294
rect 157306 50058 157542 50294
rect 156986 14378 157222 14614
rect 157306 14378 157542 14614
rect 156986 14058 157222 14294
rect 157306 14058 157542 14294
rect 138986 -7302 139222 -7066
rect 139306 -7302 139542 -7066
rect 138986 -7622 139222 -7386
rect 139306 -7622 139542 -7386
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 167546 384938 167782 385174
rect 167866 384938 168102 385174
rect 167546 384618 167782 384854
rect 167866 384618 168102 384854
rect 167546 348938 167782 349174
rect 167866 348938 168102 349174
rect 167546 348618 167782 348854
rect 167866 348618 168102 348854
rect 167546 312938 167782 313174
rect 167866 312938 168102 313174
rect 167546 312618 167782 312854
rect 167866 312618 168102 312854
rect 167546 276938 167782 277174
rect 167866 276938 168102 277174
rect 167546 276618 167782 276854
rect 167866 276618 168102 276854
rect 167546 240938 167782 241174
rect 167866 240938 168102 241174
rect 167546 240618 167782 240854
rect 167866 240618 168102 240854
rect 167546 204938 167782 205174
rect 167866 204938 168102 205174
rect 167546 204618 167782 204854
rect 167866 204618 168102 204854
rect 167546 168938 167782 169174
rect 167866 168938 168102 169174
rect 167546 168618 167782 168854
rect 167866 168618 168102 168854
rect 167546 132938 167782 133174
rect 167866 132938 168102 133174
rect 167546 132618 167782 132854
rect 167866 132618 168102 132854
rect 167546 96938 167782 97174
rect 167866 96938 168102 97174
rect 167546 96618 167782 96854
rect 167866 96618 168102 96854
rect 192986 710362 193222 710598
rect 193306 710362 193542 710598
rect 192986 710042 193222 710278
rect 193306 710042 193542 710278
rect 189266 708442 189502 708678
rect 189586 708442 189822 708678
rect 189266 708122 189502 708358
rect 189586 708122 189822 708358
rect 185546 706522 185782 706758
rect 185866 706522 186102 706758
rect 185546 706202 185782 706438
rect 185866 706202 186102 706438
rect 174986 680378 175222 680614
rect 175306 680378 175542 680614
rect 174986 680058 175222 680294
rect 175306 680058 175542 680294
rect 174986 644378 175222 644614
rect 175306 644378 175542 644614
rect 174986 644058 175222 644294
rect 175306 644058 175542 644294
rect 174986 608378 175222 608614
rect 175306 608378 175542 608614
rect 174986 608058 175222 608294
rect 175306 608058 175542 608294
rect 174986 572378 175222 572614
rect 175306 572378 175542 572614
rect 174986 572058 175222 572294
rect 175306 572058 175542 572294
rect 171266 532658 171502 532894
rect 171586 532658 171822 532894
rect 171266 532338 171502 532574
rect 171586 532338 171822 532574
rect 171266 496658 171502 496894
rect 171586 496658 171822 496894
rect 171266 496338 171502 496574
rect 171586 496338 171822 496574
rect 171266 460658 171502 460894
rect 171586 460658 171822 460894
rect 171266 460338 171502 460574
rect 171586 460338 171822 460574
rect 171266 424658 171502 424894
rect 171586 424658 171822 424894
rect 171266 424338 171502 424574
rect 171586 424338 171822 424574
rect 171266 388658 171502 388894
rect 171586 388658 171822 388894
rect 171266 388338 171502 388574
rect 171586 388338 171822 388574
rect 171266 352658 171502 352894
rect 171586 352658 171822 352894
rect 171266 352338 171502 352574
rect 171586 352338 171822 352574
rect 171266 316658 171502 316894
rect 171586 316658 171822 316894
rect 171266 316338 171502 316574
rect 171586 316338 171822 316574
rect 171266 280658 171502 280894
rect 171586 280658 171822 280894
rect 171266 280338 171502 280574
rect 171586 280338 171822 280574
rect 167546 60938 167782 61174
rect 167866 60938 168102 61174
rect 167546 60618 167782 60854
rect 167866 60618 168102 60854
rect 167546 24938 167782 25174
rect 167866 24938 168102 25174
rect 167546 24618 167782 24854
rect 167866 24618 168102 24854
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -1542 164062 -1306
rect 164146 -1542 164382 -1306
rect 163826 -1862 164062 -1626
rect 164146 -1862 164382 -1626
rect 171266 244658 171502 244894
rect 171586 244658 171822 244894
rect 171266 244338 171502 244574
rect 171586 244338 171822 244574
rect 174986 536378 175222 536614
rect 175306 536378 175542 536614
rect 174986 536058 175222 536294
rect 175306 536058 175542 536294
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 181826 543218 182062 543454
rect 182146 543218 182382 543454
rect 181826 542898 182062 543134
rect 182146 542898 182382 543134
rect 174986 500378 175222 500614
rect 175306 500378 175542 500614
rect 174986 500058 175222 500294
rect 175306 500058 175542 500294
rect 174986 464378 175222 464614
rect 175306 464378 175542 464614
rect 174986 464058 175222 464294
rect 175306 464058 175542 464294
rect 174986 428378 175222 428614
rect 175306 428378 175542 428614
rect 174986 428058 175222 428294
rect 175306 428058 175542 428294
rect 174986 392378 175222 392614
rect 175306 392378 175542 392614
rect 174986 392058 175222 392294
rect 175306 392058 175542 392294
rect 174986 356378 175222 356614
rect 175306 356378 175542 356614
rect 174986 356058 175222 356294
rect 175306 356058 175542 356294
rect 174986 320378 175222 320614
rect 175306 320378 175542 320614
rect 174986 320058 175222 320294
rect 175306 320058 175542 320294
rect 171266 208658 171502 208894
rect 171586 208658 171822 208894
rect 171266 208338 171502 208574
rect 171586 208338 171822 208574
rect 171266 172658 171502 172894
rect 171586 172658 171822 172894
rect 171266 172338 171502 172574
rect 171586 172338 171822 172574
rect 171266 136658 171502 136894
rect 171586 136658 171822 136894
rect 171266 136338 171502 136574
rect 171586 136338 171822 136574
rect 171266 100658 171502 100894
rect 171586 100658 171822 100894
rect 171266 100338 171502 100574
rect 171586 100338 171822 100574
rect 171266 64658 171502 64894
rect 171586 64658 171822 64894
rect 171266 64338 171502 64574
rect 171586 64338 171822 64574
rect 171266 28658 171502 28894
rect 171586 28658 171822 28894
rect 171266 28338 171502 28574
rect 171586 28338 171822 28574
rect 167546 -3462 167782 -3226
rect 167866 -3462 168102 -3226
rect 167546 -3782 167782 -3546
rect 167866 -3782 168102 -3546
rect 174986 284378 175222 284614
rect 175306 284378 175542 284614
rect 174986 284058 175222 284294
rect 175306 284058 175542 284294
rect 174986 248378 175222 248614
rect 175306 248378 175542 248614
rect 174986 248058 175222 248294
rect 175306 248058 175542 248294
rect 174986 212378 175222 212614
rect 175306 212378 175542 212614
rect 174986 212058 175222 212294
rect 175306 212058 175542 212294
rect 174986 176378 175222 176614
rect 175306 176378 175542 176614
rect 174986 176058 175222 176294
rect 175306 176058 175542 176294
rect 174986 140378 175222 140614
rect 175306 140378 175542 140614
rect 174986 140058 175222 140294
rect 175306 140058 175542 140294
rect 174986 104378 175222 104614
rect 175306 104378 175542 104614
rect 174986 104058 175222 104294
rect 175306 104058 175542 104294
rect 185546 690938 185782 691174
rect 185866 690938 186102 691174
rect 185546 690618 185782 690854
rect 185866 690618 186102 690854
rect 185546 654938 185782 655174
rect 185866 654938 186102 655174
rect 185546 654618 185782 654854
rect 185866 654618 186102 654854
rect 185546 618938 185782 619174
rect 185866 618938 186102 619174
rect 185546 618618 185782 618854
rect 185866 618618 186102 618854
rect 185546 582938 185782 583174
rect 185866 582938 186102 583174
rect 185546 582618 185782 582854
rect 185866 582618 186102 582854
rect 185546 546938 185782 547174
rect 185866 546938 186102 547174
rect 185546 546618 185782 546854
rect 185866 546618 186102 546854
rect 181826 507218 182062 507454
rect 182146 507218 182382 507454
rect 181826 506898 182062 507134
rect 182146 506898 182382 507134
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 181826 435218 182062 435454
rect 182146 435218 182382 435454
rect 181826 434898 182062 435134
rect 182146 434898 182382 435134
rect 181826 399218 182062 399454
rect 182146 399218 182382 399454
rect 181826 398898 182062 399134
rect 182146 398898 182382 399134
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 174986 68378 175222 68614
rect 175306 68378 175542 68614
rect 174986 68058 175222 68294
rect 175306 68058 175542 68294
rect 174986 32378 175222 32614
rect 175306 32378 175542 32614
rect 174986 32058 175222 32294
rect 175306 32058 175542 32294
rect 171266 -5382 171502 -5146
rect 171586 -5382 171822 -5146
rect 171266 -5702 171502 -5466
rect 171586 -5702 171822 -5466
rect 156986 -6342 157222 -6106
rect 157306 -6342 157542 -6106
rect 156986 -6662 157222 -6426
rect 157306 -6662 157542 -6426
rect 181826 327218 182062 327454
rect 182146 327218 182382 327454
rect 181826 326898 182062 327134
rect 182146 326898 182382 327134
rect 181826 291218 182062 291454
rect 182146 291218 182382 291454
rect 181826 290898 182062 291134
rect 182146 290898 182382 291134
rect 181826 255218 182062 255454
rect 182146 255218 182382 255454
rect 181826 254898 182062 255134
rect 182146 254898 182382 255134
rect 181826 219218 182062 219454
rect 182146 219218 182382 219454
rect 181826 218898 182062 219134
rect 182146 218898 182382 219134
rect 189266 694658 189502 694894
rect 189586 694658 189822 694894
rect 189266 694338 189502 694574
rect 189586 694338 189822 694574
rect 189266 658658 189502 658894
rect 189586 658658 189822 658894
rect 189266 658338 189502 658574
rect 189586 658338 189822 658574
rect 189266 622658 189502 622894
rect 189586 622658 189822 622894
rect 189266 622338 189502 622574
rect 189586 622338 189822 622574
rect 189266 586658 189502 586894
rect 189586 586658 189822 586894
rect 189266 586338 189502 586574
rect 189586 586338 189822 586574
rect 189266 550658 189502 550894
rect 189586 550658 189822 550894
rect 189266 550338 189502 550574
rect 189586 550338 189822 550574
rect 185546 510938 185782 511174
rect 185866 510938 186102 511174
rect 185546 510618 185782 510854
rect 185866 510618 186102 510854
rect 185546 474938 185782 475174
rect 185866 474938 186102 475174
rect 185546 474618 185782 474854
rect 185866 474618 186102 474854
rect 185546 438938 185782 439174
rect 185866 438938 186102 439174
rect 185546 438618 185782 438854
rect 185866 438618 186102 438854
rect 185546 402938 185782 403174
rect 185866 402938 186102 403174
rect 185546 402618 185782 402854
rect 185866 402618 186102 402854
rect 185546 366938 185782 367174
rect 185866 366938 186102 367174
rect 185546 366618 185782 366854
rect 185866 366618 186102 366854
rect 185546 330938 185782 331174
rect 185866 330938 186102 331174
rect 185546 330618 185782 330854
rect 185866 330618 186102 330854
rect 181826 183218 182062 183454
rect 182146 183218 182382 183454
rect 181826 182898 182062 183134
rect 182146 182898 182382 183134
rect 181826 147218 182062 147454
rect 182146 147218 182382 147454
rect 181826 146898 182062 147134
rect 182146 146898 182382 147134
rect 181826 111218 182062 111454
rect 182146 111218 182382 111454
rect 181826 110898 182062 111134
rect 182146 110898 182382 111134
rect 181826 75218 182062 75454
rect 182146 75218 182382 75454
rect 181826 74898 182062 75134
rect 182146 74898 182382 75134
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 185546 294938 185782 295174
rect 185866 294938 186102 295174
rect 185546 294618 185782 294854
rect 185866 294618 186102 294854
rect 185546 258938 185782 259174
rect 185866 258938 186102 259174
rect 185546 258618 185782 258854
rect 185866 258618 186102 258854
rect 185546 222938 185782 223174
rect 185866 222938 186102 223174
rect 185546 222618 185782 222854
rect 185866 222618 186102 222854
rect 185546 186938 185782 187174
rect 185866 186938 186102 187174
rect 185546 186618 185782 186854
rect 185866 186618 186102 186854
rect 210986 711322 211222 711558
rect 211306 711322 211542 711558
rect 210986 711002 211222 711238
rect 211306 711002 211542 711238
rect 207266 709402 207502 709638
rect 207586 709402 207822 709638
rect 207266 709082 207502 709318
rect 207586 709082 207822 709318
rect 203546 707482 203782 707718
rect 203866 707482 204102 707718
rect 203546 707162 203782 707398
rect 203866 707162 204102 707398
rect 192986 698378 193222 698614
rect 193306 698378 193542 698614
rect 192986 698058 193222 698294
rect 193306 698058 193542 698294
rect 192986 662378 193222 662614
rect 193306 662378 193542 662614
rect 192986 662058 193222 662294
rect 193306 662058 193542 662294
rect 192986 626378 193222 626614
rect 193306 626378 193542 626614
rect 192986 626058 193222 626294
rect 193306 626058 193542 626294
rect 192986 590378 193222 590614
rect 193306 590378 193542 590614
rect 192986 590058 193222 590294
rect 193306 590058 193542 590294
rect 192986 554378 193222 554614
rect 193306 554378 193542 554614
rect 192986 554058 193222 554294
rect 193306 554058 193542 554294
rect 189266 514658 189502 514894
rect 189586 514658 189822 514894
rect 189266 514338 189502 514574
rect 189586 514338 189822 514574
rect 189266 478658 189502 478894
rect 189586 478658 189822 478894
rect 189266 478338 189502 478574
rect 189586 478338 189822 478574
rect 189266 442658 189502 442894
rect 189586 442658 189822 442894
rect 189266 442338 189502 442574
rect 189586 442338 189822 442574
rect 189266 406658 189502 406894
rect 189586 406658 189822 406894
rect 189266 406338 189502 406574
rect 189586 406338 189822 406574
rect 189266 370658 189502 370894
rect 189586 370658 189822 370894
rect 189266 370338 189502 370574
rect 189586 370338 189822 370574
rect 189266 334658 189502 334894
rect 189586 334658 189822 334894
rect 189266 334338 189502 334574
rect 189586 334338 189822 334574
rect 189266 298658 189502 298894
rect 189586 298658 189822 298894
rect 189266 298338 189502 298574
rect 189586 298338 189822 298574
rect 189266 262658 189502 262894
rect 189586 262658 189822 262894
rect 189266 262338 189502 262574
rect 189586 262338 189822 262574
rect 189266 226658 189502 226894
rect 189586 226658 189822 226894
rect 189266 226338 189502 226574
rect 189586 226338 189822 226574
rect 189266 190658 189502 190894
rect 189586 190658 189822 190894
rect 189266 190338 189502 190574
rect 189586 190338 189822 190574
rect 185546 150938 185782 151174
rect 185866 150938 186102 151174
rect 185546 150618 185782 150854
rect 185866 150618 186102 150854
rect 185546 114938 185782 115174
rect 185866 114938 186102 115174
rect 185546 114618 185782 114854
rect 185866 114618 186102 114854
rect 185546 78938 185782 79174
rect 185866 78938 186102 79174
rect 185546 78618 185782 78854
rect 185866 78618 186102 78854
rect 185546 42938 185782 43174
rect 185866 42938 186102 43174
rect 185546 42618 185782 42854
rect 185866 42618 186102 42854
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 185546 6938 185782 7174
rect 185866 6938 186102 7174
rect 185546 6618 185782 6854
rect 185866 6618 186102 6854
rect 185546 -2502 185782 -2266
rect 185866 -2502 186102 -2266
rect 185546 -2822 185782 -2586
rect 185866 -2822 186102 -2586
rect 189266 154658 189502 154894
rect 189586 154658 189822 154894
rect 189266 154338 189502 154574
rect 189586 154338 189822 154574
rect 189266 118658 189502 118894
rect 189586 118658 189822 118894
rect 189266 118338 189502 118574
rect 189586 118338 189822 118574
rect 189266 82658 189502 82894
rect 189586 82658 189822 82894
rect 189266 82338 189502 82574
rect 189586 82338 189822 82574
rect 189266 46658 189502 46894
rect 189586 46658 189822 46894
rect 189266 46338 189502 46574
rect 189586 46338 189822 46574
rect 199826 705562 200062 705798
rect 200146 705562 200382 705798
rect 199826 705242 200062 705478
rect 200146 705242 200382 705478
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 199826 633218 200062 633454
rect 200146 633218 200382 633454
rect 199826 632898 200062 633134
rect 200146 632898 200382 633134
rect 199826 597218 200062 597454
rect 200146 597218 200382 597454
rect 199826 596898 200062 597134
rect 200146 596898 200382 597134
rect 199826 561218 200062 561454
rect 200146 561218 200382 561454
rect 199826 560898 200062 561134
rect 200146 560898 200382 561134
rect 192986 518378 193222 518614
rect 193306 518378 193542 518614
rect 192986 518058 193222 518294
rect 193306 518058 193542 518294
rect 192986 482378 193222 482614
rect 193306 482378 193542 482614
rect 192986 482058 193222 482294
rect 193306 482058 193542 482294
rect 192986 446378 193222 446614
rect 193306 446378 193542 446614
rect 192986 446058 193222 446294
rect 193306 446058 193542 446294
rect 192986 410378 193222 410614
rect 193306 410378 193542 410614
rect 192986 410058 193222 410294
rect 193306 410058 193542 410294
rect 192986 374378 193222 374614
rect 193306 374378 193542 374614
rect 192986 374058 193222 374294
rect 193306 374058 193542 374294
rect 192986 338378 193222 338614
rect 193306 338378 193542 338614
rect 192986 338058 193222 338294
rect 193306 338058 193542 338294
rect 192986 302378 193222 302614
rect 193306 302378 193542 302614
rect 192986 302058 193222 302294
rect 193306 302058 193542 302294
rect 192986 266378 193222 266614
rect 193306 266378 193542 266614
rect 192986 266058 193222 266294
rect 193306 266058 193542 266294
rect 192986 230378 193222 230614
rect 193306 230378 193542 230614
rect 192986 230058 193222 230294
rect 193306 230058 193542 230294
rect 203546 672938 203782 673174
rect 203866 672938 204102 673174
rect 203546 672618 203782 672854
rect 203866 672618 204102 672854
rect 203546 636938 203782 637174
rect 203866 636938 204102 637174
rect 203546 636618 203782 636854
rect 203866 636618 204102 636854
rect 203546 600938 203782 601174
rect 203866 600938 204102 601174
rect 203546 600618 203782 600854
rect 203866 600618 204102 600854
rect 203546 564938 203782 565174
rect 203866 564938 204102 565174
rect 203546 564618 203782 564854
rect 203866 564618 204102 564854
rect 207266 676658 207502 676894
rect 207586 676658 207822 676894
rect 207266 676338 207502 676574
rect 207586 676338 207822 676574
rect 207266 640658 207502 640894
rect 207586 640658 207822 640894
rect 207266 640338 207502 640574
rect 207586 640338 207822 640574
rect 207266 604658 207502 604894
rect 207586 604658 207822 604894
rect 207266 604338 207502 604574
rect 207586 604338 207822 604574
rect 207266 568658 207502 568894
rect 207586 568658 207822 568894
rect 207266 568338 207502 568574
rect 207586 568338 207822 568574
rect 228986 710362 229222 710598
rect 229306 710362 229542 710598
rect 228986 710042 229222 710278
rect 229306 710042 229542 710278
rect 225266 708442 225502 708678
rect 225586 708442 225822 708678
rect 225266 708122 225502 708358
rect 225586 708122 225822 708358
rect 221546 706522 221782 706758
rect 221866 706522 222102 706758
rect 221546 706202 221782 706438
rect 221866 706202 222102 706438
rect 210986 680378 211222 680614
rect 211306 680378 211542 680614
rect 210986 680058 211222 680294
rect 211306 680058 211542 680294
rect 210986 644378 211222 644614
rect 211306 644378 211542 644614
rect 210986 644058 211222 644294
rect 211306 644058 211542 644294
rect 210986 608378 211222 608614
rect 211306 608378 211542 608614
rect 210986 608058 211222 608294
rect 211306 608058 211542 608294
rect 210986 572378 211222 572614
rect 211306 572378 211542 572614
rect 210986 572058 211222 572294
rect 211306 572058 211542 572294
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 217826 543218 218062 543454
rect 218146 543218 218382 543454
rect 217826 542898 218062 543134
rect 218146 542898 218382 543134
rect 221546 690938 221782 691174
rect 221866 690938 222102 691174
rect 221546 690618 221782 690854
rect 221866 690618 222102 690854
rect 221546 654938 221782 655174
rect 221866 654938 222102 655174
rect 221546 654618 221782 654854
rect 221866 654618 222102 654854
rect 221546 618938 221782 619174
rect 221866 618938 222102 619174
rect 221546 618618 221782 618854
rect 221866 618618 222102 618854
rect 221546 582938 221782 583174
rect 221866 582938 222102 583174
rect 221546 582618 221782 582854
rect 221866 582618 222102 582854
rect 221546 546938 221782 547174
rect 221866 546938 222102 547174
rect 221546 546618 221782 546854
rect 221866 546618 222102 546854
rect 225266 694658 225502 694894
rect 225586 694658 225822 694894
rect 225266 694338 225502 694574
rect 225586 694338 225822 694574
rect 225266 658658 225502 658894
rect 225586 658658 225822 658894
rect 225266 658338 225502 658574
rect 225586 658338 225822 658574
rect 225266 622658 225502 622894
rect 225586 622658 225822 622894
rect 225266 622338 225502 622574
rect 225586 622338 225822 622574
rect 225266 586658 225502 586894
rect 225586 586658 225822 586894
rect 225266 586338 225502 586574
rect 225586 586338 225822 586574
rect 225266 550658 225502 550894
rect 225586 550658 225822 550894
rect 225266 550338 225502 550574
rect 225586 550338 225822 550574
rect 246986 711322 247222 711558
rect 247306 711322 247542 711558
rect 246986 711002 247222 711238
rect 247306 711002 247542 711238
rect 243266 709402 243502 709638
rect 243586 709402 243822 709638
rect 243266 709082 243502 709318
rect 243586 709082 243822 709318
rect 239546 707482 239782 707718
rect 239866 707482 240102 707718
rect 239546 707162 239782 707398
rect 239866 707162 240102 707398
rect 228986 698378 229222 698614
rect 229306 698378 229542 698614
rect 228986 698058 229222 698294
rect 229306 698058 229542 698294
rect 228986 662378 229222 662614
rect 229306 662378 229542 662614
rect 228986 662058 229222 662294
rect 229306 662058 229542 662294
rect 228986 626378 229222 626614
rect 229306 626378 229542 626614
rect 228986 626058 229222 626294
rect 229306 626058 229542 626294
rect 228986 590378 229222 590614
rect 229306 590378 229542 590614
rect 228986 590058 229222 590294
rect 229306 590058 229542 590294
rect 228986 554378 229222 554614
rect 229306 554378 229542 554614
rect 228986 554058 229222 554294
rect 229306 554058 229542 554294
rect 235826 705562 236062 705798
rect 236146 705562 236382 705798
rect 235826 705242 236062 705478
rect 236146 705242 236382 705478
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 235826 633218 236062 633454
rect 236146 633218 236382 633454
rect 235826 632898 236062 633134
rect 236146 632898 236382 633134
rect 235826 597218 236062 597454
rect 236146 597218 236382 597454
rect 235826 596898 236062 597134
rect 236146 596898 236382 597134
rect 235826 561218 236062 561454
rect 236146 561218 236382 561454
rect 235826 560898 236062 561134
rect 236146 560898 236382 561134
rect 239546 672938 239782 673174
rect 239866 672938 240102 673174
rect 239546 672618 239782 672854
rect 239866 672618 240102 672854
rect 239546 636938 239782 637174
rect 239866 636938 240102 637174
rect 239546 636618 239782 636854
rect 239866 636618 240102 636854
rect 239546 600938 239782 601174
rect 239866 600938 240102 601174
rect 239546 600618 239782 600854
rect 239866 600618 240102 600854
rect 239546 564938 239782 565174
rect 239866 564938 240102 565174
rect 239546 564618 239782 564854
rect 239866 564618 240102 564854
rect 243266 676658 243502 676894
rect 243586 676658 243822 676894
rect 243266 676338 243502 676574
rect 243586 676338 243822 676574
rect 243266 640658 243502 640894
rect 243586 640658 243822 640894
rect 243266 640338 243502 640574
rect 243586 640338 243822 640574
rect 243266 604658 243502 604894
rect 243586 604658 243822 604894
rect 243266 604338 243502 604574
rect 243586 604338 243822 604574
rect 243266 568658 243502 568894
rect 243586 568658 243822 568894
rect 243266 568338 243502 568574
rect 243586 568338 243822 568574
rect 264986 710362 265222 710598
rect 265306 710362 265542 710598
rect 264986 710042 265222 710278
rect 265306 710042 265542 710278
rect 261266 708442 261502 708678
rect 261586 708442 261822 708678
rect 261266 708122 261502 708358
rect 261586 708122 261822 708358
rect 257546 706522 257782 706758
rect 257866 706522 258102 706758
rect 257546 706202 257782 706438
rect 257866 706202 258102 706438
rect 246986 680378 247222 680614
rect 247306 680378 247542 680614
rect 246986 680058 247222 680294
rect 247306 680058 247542 680294
rect 246986 644378 247222 644614
rect 247306 644378 247542 644614
rect 246986 644058 247222 644294
rect 247306 644058 247542 644294
rect 246986 608378 247222 608614
rect 247306 608378 247542 608614
rect 246986 608058 247222 608294
rect 247306 608058 247542 608294
rect 246986 572378 247222 572614
rect 247306 572378 247542 572614
rect 246986 572058 247222 572294
rect 247306 572058 247542 572294
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 253826 615218 254062 615454
rect 254146 615218 254382 615454
rect 253826 614898 254062 615134
rect 254146 614898 254382 615134
rect 253826 579218 254062 579454
rect 254146 579218 254382 579454
rect 253826 578898 254062 579134
rect 254146 578898 254382 579134
rect 253826 543218 254062 543454
rect 254146 543218 254382 543454
rect 253826 542898 254062 543134
rect 254146 542898 254382 543134
rect 257546 690938 257782 691174
rect 257866 690938 258102 691174
rect 257546 690618 257782 690854
rect 257866 690618 258102 690854
rect 257546 654938 257782 655174
rect 257866 654938 258102 655174
rect 257546 654618 257782 654854
rect 257866 654618 258102 654854
rect 257546 618938 257782 619174
rect 257866 618938 258102 619174
rect 257546 618618 257782 618854
rect 257866 618618 258102 618854
rect 257546 582938 257782 583174
rect 257866 582938 258102 583174
rect 257546 582618 257782 582854
rect 257866 582618 258102 582854
rect 257546 546938 257782 547174
rect 257866 546938 258102 547174
rect 257546 546618 257782 546854
rect 257866 546618 258102 546854
rect 261266 694658 261502 694894
rect 261586 694658 261822 694894
rect 261266 694338 261502 694574
rect 261586 694338 261822 694574
rect 261266 658658 261502 658894
rect 261586 658658 261822 658894
rect 261266 658338 261502 658574
rect 261586 658338 261822 658574
rect 261266 622658 261502 622894
rect 261586 622658 261822 622894
rect 261266 622338 261502 622574
rect 261586 622338 261822 622574
rect 261266 586658 261502 586894
rect 261586 586658 261822 586894
rect 261266 586338 261502 586574
rect 261586 586338 261822 586574
rect 261266 550658 261502 550894
rect 261586 550658 261822 550894
rect 261266 550338 261502 550574
rect 261586 550338 261822 550574
rect 282986 711322 283222 711558
rect 283306 711322 283542 711558
rect 282986 711002 283222 711238
rect 283306 711002 283542 711238
rect 279266 709402 279502 709638
rect 279586 709402 279822 709638
rect 279266 709082 279502 709318
rect 279586 709082 279822 709318
rect 275546 707482 275782 707718
rect 275866 707482 276102 707718
rect 275546 707162 275782 707398
rect 275866 707162 276102 707398
rect 264986 698378 265222 698614
rect 265306 698378 265542 698614
rect 264986 698058 265222 698294
rect 265306 698058 265542 698294
rect 264986 662378 265222 662614
rect 265306 662378 265542 662614
rect 264986 662058 265222 662294
rect 265306 662058 265542 662294
rect 264986 626378 265222 626614
rect 265306 626378 265542 626614
rect 264986 626058 265222 626294
rect 265306 626058 265542 626294
rect 264986 590378 265222 590614
rect 265306 590378 265542 590614
rect 264986 590058 265222 590294
rect 265306 590058 265542 590294
rect 264986 554378 265222 554614
rect 265306 554378 265542 554614
rect 264986 554058 265222 554294
rect 265306 554058 265542 554294
rect 271826 705562 272062 705798
rect 272146 705562 272382 705798
rect 271826 705242 272062 705478
rect 272146 705242 272382 705478
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 271826 633218 272062 633454
rect 272146 633218 272382 633454
rect 271826 632898 272062 633134
rect 272146 632898 272382 633134
rect 271826 597218 272062 597454
rect 272146 597218 272382 597454
rect 271826 596898 272062 597134
rect 272146 596898 272382 597134
rect 271826 561218 272062 561454
rect 272146 561218 272382 561454
rect 271826 560898 272062 561134
rect 272146 560898 272382 561134
rect 275546 672938 275782 673174
rect 275866 672938 276102 673174
rect 275546 672618 275782 672854
rect 275866 672618 276102 672854
rect 275546 636938 275782 637174
rect 275866 636938 276102 637174
rect 275546 636618 275782 636854
rect 275866 636618 276102 636854
rect 275546 600938 275782 601174
rect 275866 600938 276102 601174
rect 275546 600618 275782 600854
rect 275866 600618 276102 600854
rect 275546 564938 275782 565174
rect 275866 564938 276102 565174
rect 275546 564618 275782 564854
rect 275866 564618 276102 564854
rect 279266 676658 279502 676894
rect 279586 676658 279822 676894
rect 279266 676338 279502 676574
rect 279586 676338 279822 676574
rect 279266 640658 279502 640894
rect 279586 640658 279822 640894
rect 279266 640338 279502 640574
rect 279586 640338 279822 640574
rect 279266 604658 279502 604894
rect 279586 604658 279822 604894
rect 279266 604338 279502 604574
rect 279586 604338 279822 604574
rect 279266 568658 279502 568894
rect 279586 568658 279822 568894
rect 279266 568338 279502 568574
rect 279586 568338 279822 568574
rect 300986 710362 301222 710598
rect 301306 710362 301542 710598
rect 300986 710042 301222 710278
rect 301306 710042 301542 710278
rect 297266 708442 297502 708678
rect 297586 708442 297822 708678
rect 297266 708122 297502 708358
rect 297586 708122 297822 708358
rect 293546 706522 293782 706758
rect 293866 706522 294102 706758
rect 293546 706202 293782 706438
rect 293866 706202 294102 706438
rect 282986 680378 283222 680614
rect 283306 680378 283542 680614
rect 282986 680058 283222 680294
rect 283306 680058 283542 680294
rect 282986 644378 283222 644614
rect 283306 644378 283542 644614
rect 282986 644058 283222 644294
rect 283306 644058 283542 644294
rect 282986 608378 283222 608614
rect 283306 608378 283542 608614
rect 282986 608058 283222 608294
rect 283306 608058 283542 608294
rect 282986 572378 283222 572614
rect 283306 572378 283542 572614
rect 282986 572058 283222 572294
rect 283306 572058 283542 572294
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 289826 543218 290062 543454
rect 290146 543218 290382 543454
rect 289826 542898 290062 543134
rect 290146 542898 290382 543134
rect 293546 690938 293782 691174
rect 293866 690938 294102 691174
rect 293546 690618 293782 690854
rect 293866 690618 294102 690854
rect 293546 654938 293782 655174
rect 293866 654938 294102 655174
rect 293546 654618 293782 654854
rect 293866 654618 294102 654854
rect 293546 618938 293782 619174
rect 293866 618938 294102 619174
rect 293546 618618 293782 618854
rect 293866 618618 294102 618854
rect 293546 582938 293782 583174
rect 293866 582938 294102 583174
rect 293546 582618 293782 582854
rect 293866 582618 294102 582854
rect 293546 546938 293782 547174
rect 293866 546938 294102 547174
rect 293546 546618 293782 546854
rect 293866 546618 294102 546854
rect 297266 694658 297502 694894
rect 297586 694658 297822 694894
rect 297266 694338 297502 694574
rect 297586 694338 297822 694574
rect 297266 658658 297502 658894
rect 297586 658658 297822 658894
rect 297266 658338 297502 658574
rect 297586 658338 297822 658574
rect 297266 622658 297502 622894
rect 297586 622658 297822 622894
rect 297266 622338 297502 622574
rect 297586 622338 297822 622574
rect 297266 586658 297502 586894
rect 297586 586658 297822 586894
rect 297266 586338 297502 586574
rect 297586 586338 297822 586574
rect 297266 550658 297502 550894
rect 297586 550658 297822 550894
rect 297266 550338 297502 550574
rect 297586 550338 297822 550574
rect 318986 711322 319222 711558
rect 319306 711322 319542 711558
rect 318986 711002 319222 711238
rect 319306 711002 319542 711238
rect 315266 709402 315502 709638
rect 315586 709402 315822 709638
rect 315266 709082 315502 709318
rect 315586 709082 315822 709318
rect 311546 707482 311782 707718
rect 311866 707482 312102 707718
rect 311546 707162 311782 707398
rect 311866 707162 312102 707398
rect 300986 698378 301222 698614
rect 301306 698378 301542 698614
rect 300986 698058 301222 698294
rect 301306 698058 301542 698294
rect 300986 662378 301222 662614
rect 301306 662378 301542 662614
rect 300986 662058 301222 662294
rect 301306 662058 301542 662294
rect 300986 626378 301222 626614
rect 301306 626378 301542 626614
rect 300986 626058 301222 626294
rect 301306 626058 301542 626294
rect 300986 590378 301222 590614
rect 301306 590378 301542 590614
rect 300986 590058 301222 590294
rect 301306 590058 301542 590294
rect 300986 554378 301222 554614
rect 301306 554378 301542 554614
rect 300986 554058 301222 554294
rect 301306 554058 301542 554294
rect 307826 705562 308062 705798
rect 308146 705562 308382 705798
rect 307826 705242 308062 705478
rect 308146 705242 308382 705478
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 307826 561218 308062 561454
rect 308146 561218 308382 561454
rect 307826 560898 308062 561134
rect 308146 560898 308382 561134
rect 311546 672938 311782 673174
rect 311866 672938 312102 673174
rect 311546 672618 311782 672854
rect 311866 672618 312102 672854
rect 311546 636938 311782 637174
rect 311866 636938 312102 637174
rect 311546 636618 311782 636854
rect 311866 636618 312102 636854
rect 311546 600938 311782 601174
rect 311866 600938 312102 601174
rect 311546 600618 311782 600854
rect 311866 600618 312102 600854
rect 311546 564938 311782 565174
rect 311866 564938 312102 565174
rect 311546 564618 311782 564854
rect 311866 564618 312102 564854
rect 315266 676658 315502 676894
rect 315586 676658 315822 676894
rect 315266 676338 315502 676574
rect 315586 676338 315822 676574
rect 315266 640658 315502 640894
rect 315586 640658 315822 640894
rect 315266 640338 315502 640574
rect 315586 640338 315822 640574
rect 315266 604658 315502 604894
rect 315586 604658 315822 604894
rect 315266 604338 315502 604574
rect 315586 604338 315822 604574
rect 315266 568658 315502 568894
rect 315586 568658 315822 568894
rect 315266 568338 315502 568574
rect 315586 568338 315822 568574
rect 336986 710362 337222 710598
rect 337306 710362 337542 710598
rect 336986 710042 337222 710278
rect 337306 710042 337542 710278
rect 333266 708442 333502 708678
rect 333586 708442 333822 708678
rect 333266 708122 333502 708358
rect 333586 708122 333822 708358
rect 329546 706522 329782 706758
rect 329866 706522 330102 706758
rect 329546 706202 329782 706438
rect 329866 706202 330102 706438
rect 318986 680378 319222 680614
rect 319306 680378 319542 680614
rect 318986 680058 319222 680294
rect 319306 680058 319542 680294
rect 318986 644378 319222 644614
rect 319306 644378 319542 644614
rect 318986 644058 319222 644294
rect 319306 644058 319542 644294
rect 318986 608378 319222 608614
rect 319306 608378 319542 608614
rect 318986 608058 319222 608294
rect 319306 608058 319542 608294
rect 318986 572378 319222 572614
rect 319306 572378 319542 572614
rect 318986 572058 319222 572294
rect 319306 572058 319542 572294
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 325826 543218 326062 543454
rect 326146 543218 326382 543454
rect 325826 542898 326062 543134
rect 326146 542898 326382 543134
rect 329546 690938 329782 691174
rect 329866 690938 330102 691174
rect 329546 690618 329782 690854
rect 329866 690618 330102 690854
rect 329546 654938 329782 655174
rect 329866 654938 330102 655174
rect 329546 654618 329782 654854
rect 329866 654618 330102 654854
rect 329546 618938 329782 619174
rect 329866 618938 330102 619174
rect 329546 618618 329782 618854
rect 329866 618618 330102 618854
rect 329546 582938 329782 583174
rect 329866 582938 330102 583174
rect 329546 582618 329782 582854
rect 329866 582618 330102 582854
rect 329546 546938 329782 547174
rect 329866 546938 330102 547174
rect 329546 546618 329782 546854
rect 329866 546618 330102 546854
rect 333266 694658 333502 694894
rect 333586 694658 333822 694894
rect 333266 694338 333502 694574
rect 333586 694338 333822 694574
rect 333266 658658 333502 658894
rect 333586 658658 333822 658894
rect 333266 658338 333502 658574
rect 333586 658338 333822 658574
rect 333266 622658 333502 622894
rect 333586 622658 333822 622894
rect 333266 622338 333502 622574
rect 333586 622338 333822 622574
rect 333266 586658 333502 586894
rect 333586 586658 333822 586894
rect 333266 586338 333502 586574
rect 333586 586338 333822 586574
rect 333266 550658 333502 550894
rect 333586 550658 333822 550894
rect 333266 550338 333502 550574
rect 333586 550338 333822 550574
rect 354986 711322 355222 711558
rect 355306 711322 355542 711558
rect 354986 711002 355222 711238
rect 355306 711002 355542 711238
rect 351266 709402 351502 709638
rect 351586 709402 351822 709638
rect 351266 709082 351502 709318
rect 351586 709082 351822 709318
rect 347546 707482 347782 707718
rect 347866 707482 348102 707718
rect 347546 707162 347782 707398
rect 347866 707162 348102 707398
rect 336986 698378 337222 698614
rect 337306 698378 337542 698614
rect 336986 698058 337222 698294
rect 337306 698058 337542 698294
rect 336986 662378 337222 662614
rect 337306 662378 337542 662614
rect 336986 662058 337222 662294
rect 337306 662058 337542 662294
rect 336986 626378 337222 626614
rect 337306 626378 337542 626614
rect 336986 626058 337222 626294
rect 337306 626058 337542 626294
rect 336986 590378 337222 590614
rect 337306 590378 337542 590614
rect 336986 590058 337222 590294
rect 337306 590058 337542 590294
rect 336986 554378 337222 554614
rect 337306 554378 337542 554614
rect 336986 554058 337222 554294
rect 337306 554058 337542 554294
rect 343826 705562 344062 705798
rect 344146 705562 344382 705798
rect 343826 705242 344062 705478
rect 344146 705242 344382 705478
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 343826 633218 344062 633454
rect 344146 633218 344382 633454
rect 343826 632898 344062 633134
rect 344146 632898 344382 633134
rect 343826 597218 344062 597454
rect 344146 597218 344382 597454
rect 343826 596898 344062 597134
rect 344146 596898 344382 597134
rect 343826 561218 344062 561454
rect 344146 561218 344382 561454
rect 343826 560898 344062 561134
rect 344146 560898 344382 561134
rect 347546 672938 347782 673174
rect 347866 672938 348102 673174
rect 347546 672618 347782 672854
rect 347866 672618 348102 672854
rect 347546 636938 347782 637174
rect 347866 636938 348102 637174
rect 347546 636618 347782 636854
rect 347866 636618 348102 636854
rect 347546 600938 347782 601174
rect 347866 600938 348102 601174
rect 347546 600618 347782 600854
rect 347866 600618 348102 600854
rect 347546 564938 347782 565174
rect 347866 564938 348102 565174
rect 347546 564618 347782 564854
rect 347866 564618 348102 564854
rect 351266 676658 351502 676894
rect 351586 676658 351822 676894
rect 351266 676338 351502 676574
rect 351586 676338 351822 676574
rect 351266 640658 351502 640894
rect 351586 640658 351822 640894
rect 351266 640338 351502 640574
rect 351586 640338 351822 640574
rect 351266 604658 351502 604894
rect 351586 604658 351822 604894
rect 351266 604338 351502 604574
rect 351586 604338 351822 604574
rect 351266 568658 351502 568894
rect 351586 568658 351822 568894
rect 351266 568338 351502 568574
rect 351586 568338 351822 568574
rect 372986 710362 373222 710598
rect 373306 710362 373542 710598
rect 372986 710042 373222 710278
rect 373306 710042 373542 710278
rect 369266 708442 369502 708678
rect 369586 708442 369822 708678
rect 369266 708122 369502 708358
rect 369586 708122 369822 708358
rect 365546 706522 365782 706758
rect 365866 706522 366102 706758
rect 365546 706202 365782 706438
rect 365866 706202 366102 706438
rect 354986 680378 355222 680614
rect 355306 680378 355542 680614
rect 354986 680058 355222 680294
rect 355306 680058 355542 680294
rect 354986 644378 355222 644614
rect 355306 644378 355542 644614
rect 354986 644058 355222 644294
rect 355306 644058 355542 644294
rect 354986 608378 355222 608614
rect 355306 608378 355542 608614
rect 354986 608058 355222 608294
rect 355306 608058 355542 608294
rect 354986 572378 355222 572614
rect 355306 572378 355542 572614
rect 354986 572058 355222 572294
rect 355306 572058 355542 572294
rect 219610 525218 219846 525454
rect 219610 524898 219846 525134
rect 250330 525218 250566 525454
rect 250330 524898 250566 525134
rect 281050 525218 281286 525454
rect 281050 524898 281286 525134
rect 311770 525218 312006 525454
rect 311770 524898 312006 525134
rect 342490 525218 342726 525454
rect 342490 524898 342726 525134
rect 204250 507218 204486 507454
rect 204250 506898 204486 507134
rect 234970 507218 235206 507454
rect 234970 506898 235206 507134
rect 265690 507218 265926 507454
rect 265690 506898 265926 507134
rect 296410 507218 296646 507454
rect 296410 506898 296646 507134
rect 327130 507218 327366 507454
rect 327130 506898 327366 507134
rect 219610 489218 219846 489454
rect 219610 488898 219846 489134
rect 250330 489218 250566 489454
rect 250330 488898 250566 489134
rect 281050 489218 281286 489454
rect 281050 488898 281286 489134
rect 311770 489218 312006 489454
rect 311770 488898 312006 489134
rect 342490 489218 342726 489454
rect 342490 488898 342726 489134
rect 204250 471218 204486 471454
rect 204250 470898 204486 471134
rect 234970 471218 235206 471454
rect 234970 470898 235206 471134
rect 265690 471218 265926 471454
rect 265690 470898 265926 471134
rect 296410 471218 296646 471454
rect 296410 470898 296646 471134
rect 327130 471218 327366 471454
rect 327130 470898 327366 471134
rect 219610 453218 219846 453454
rect 219610 452898 219846 453134
rect 250330 453218 250566 453454
rect 250330 452898 250566 453134
rect 281050 453218 281286 453454
rect 281050 452898 281286 453134
rect 311770 453218 312006 453454
rect 311770 452898 312006 453134
rect 342490 453218 342726 453454
rect 342490 452898 342726 453134
rect 204250 435218 204486 435454
rect 204250 434898 204486 435134
rect 234970 435218 235206 435454
rect 234970 434898 235206 435134
rect 265690 435218 265926 435454
rect 265690 434898 265926 435134
rect 296410 435218 296646 435454
rect 296410 434898 296646 435134
rect 327130 435218 327366 435454
rect 327130 434898 327366 435134
rect 219610 417218 219846 417454
rect 219610 416898 219846 417134
rect 250330 417218 250566 417454
rect 250330 416898 250566 417134
rect 281050 417218 281286 417454
rect 281050 416898 281286 417134
rect 311770 417218 312006 417454
rect 311770 416898 312006 417134
rect 342490 417218 342726 417454
rect 342490 416898 342726 417134
rect 204250 399218 204486 399454
rect 204250 398898 204486 399134
rect 234970 399218 235206 399454
rect 234970 398898 235206 399134
rect 265690 399218 265926 399454
rect 265690 398898 265926 399134
rect 296410 399218 296646 399454
rect 296410 398898 296646 399134
rect 327130 399218 327366 399454
rect 327130 398898 327366 399134
rect 219610 381218 219846 381454
rect 219610 380898 219846 381134
rect 250330 381218 250566 381454
rect 250330 380898 250566 381134
rect 281050 381218 281286 381454
rect 281050 380898 281286 381134
rect 311770 381218 312006 381454
rect 311770 380898 312006 381134
rect 342490 381218 342726 381454
rect 342490 380898 342726 381134
rect 199826 345218 200062 345454
rect 200146 345218 200382 345454
rect 199826 344898 200062 345134
rect 200146 344898 200382 345134
rect 203546 348938 203782 349174
rect 203866 348938 204102 349174
rect 203546 348618 203782 348854
rect 203866 348618 204102 348854
rect 199826 309218 200062 309454
rect 200146 309218 200382 309454
rect 199826 308898 200062 309134
rect 200146 308898 200382 309134
rect 199826 237218 200062 237454
rect 200146 237218 200382 237454
rect 199826 236898 200062 237134
rect 200146 236898 200382 237134
rect 192986 194378 193222 194614
rect 193306 194378 193542 194614
rect 192986 194058 193222 194294
rect 193306 194058 193542 194294
rect 192986 158378 193222 158614
rect 193306 158378 193542 158614
rect 192986 158058 193222 158294
rect 193306 158058 193542 158294
rect 192986 122378 193222 122614
rect 193306 122378 193542 122614
rect 192986 122058 193222 122294
rect 193306 122058 193542 122294
rect 192986 86378 193222 86614
rect 193306 86378 193542 86614
rect 192986 86058 193222 86294
rect 193306 86058 193542 86294
rect 192986 50378 193222 50614
rect 193306 50378 193542 50614
rect 192986 50058 193222 50294
rect 193306 50058 193542 50294
rect 189266 10658 189502 10894
rect 189586 10658 189822 10894
rect 189266 10338 189502 10574
rect 189586 10338 189822 10574
rect 189266 -4422 189502 -4186
rect 189586 -4422 189822 -4186
rect 189266 -4742 189502 -4506
rect 189586 -4742 189822 -4506
rect 192986 14378 193222 14614
rect 193306 14378 193542 14614
rect 192986 14058 193222 14294
rect 193306 14058 193542 14294
rect 174986 -7302 175222 -7066
rect 175306 -7302 175542 -7066
rect 174986 -7622 175222 -7386
rect 175306 -7622 175542 -7386
rect 199826 201218 200062 201454
rect 200146 201218 200382 201454
rect 199826 200898 200062 201134
rect 200146 200898 200382 201134
rect 199826 165218 200062 165454
rect 200146 165218 200382 165454
rect 199826 164898 200062 165134
rect 200146 164898 200382 165134
rect 199826 129218 200062 129454
rect 200146 129218 200382 129454
rect 199826 128898 200062 129134
rect 200146 128898 200382 129134
rect 203546 312938 203782 313174
rect 203866 312938 204102 313174
rect 203546 312618 203782 312854
rect 203866 312618 204102 312854
rect 207266 352658 207502 352894
rect 207586 352658 207822 352894
rect 207266 352338 207502 352574
rect 207586 352338 207822 352574
rect 210986 356378 211222 356614
rect 211306 356378 211542 356614
rect 210986 356058 211222 356294
rect 211306 356058 211542 356294
rect 207266 316658 207502 316894
rect 207586 316658 207822 316894
rect 207266 316338 207502 316574
rect 207586 316338 207822 316574
rect 204450 255218 204686 255454
rect 204450 254898 204686 255134
rect 203546 204938 203782 205174
rect 203866 204938 204102 205174
rect 203546 204618 203782 204854
rect 203866 204618 204102 204854
rect 203546 168938 203782 169174
rect 203866 168938 204102 169174
rect 203546 168618 203782 168854
rect 203866 168618 204102 168854
rect 203546 132938 203782 133174
rect 203866 132938 204102 133174
rect 203546 132618 203782 132854
rect 203866 132618 204102 132854
rect 203546 96938 203782 97174
rect 203866 96938 204102 97174
rect 203546 96618 203782 96854
rect 203866 96618 204102 96854
rect 199826 93218 200062 93454
rect 200146 93218 200382 93454
rect 199826 92898 200062 93134
rect 200146 92898 200382 93134
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -1542 200062 -1306
rect 200146 -1542 200382 -1306
rect 199826 -1862 200062 -1626
rect 200146 -1862 200382 -1626
rect 203546 60938 203782 61174
rect 203866 60938 204102 61174
rect 203546 60618 203782 60854
rect 203866 60618 204102 60854
rect 203546 24938 203782 25174
rect 203866 24938 204102 25174
rect 203546 24618 203782 24854
rect 203866 24618 204102 24854
rect 203546 -3462 203782 -3226
rect 203866 -3462 204102 -3226
rect 203546 -3782 203782 -3546
rect 203866 -3782 204102 -3546
rect 217826 363218 218062 363454
rect 218146 363218 218382 363454
rect 217826 362898 218062 363134
rect 218146 362898 218382 363134
rect 210986 320378 211222 320614
rect 211306 320378 211542 320614
rect 210986 320058 211222 320294
rect 211306 320058 211542 320294
rect 210986 212378 211222 212614
rect 211306 212378 211542 212614
rect 210986 212058 211222 212294
rect 211306 212058 211542 212294
rect 207266 208658 207502 208894
rect 207586 208658 207822 208894
rect 207266 208338 207502 208574
rect 207586 208338 207822 208574
rect 207266 172658 207502 172894
rect 207586 172658 207822 172894
rect 207266 172338 207502 172574
rect 207586 172338 207822 172574
rect 207266 136658 207502 136894
rect 207586 136658 207822 136894
rect 207266 136338 207502 136574
rect 207586 136338 207822 136574
rect 207266 100658 207502 100894
rect 207586 100658 207822 100894
rect 207266 100338 207502 100574
rect 207586 100338 207822 100574
rect 207266 64658 207502 64894
rect 207586 64658 207822 64894
rect 207266 64338 207502 64574
rect 207586 64338 207822 64574
rect 207266 28658 207502 28894
rect 207586 28658 207822 28894
rect 207266 28338 207502 28574
rect 207586 28338 207822 28574
rect 207266 -5382 207502 -5146
rect 207586 -5382 207822 -5146
rect 207266 -5702 207502 -5466
rect 207586 -5702 207822 -5466
rect 217826 327218 218062 327454
rect 218146 327218 218382 327454
rect 217826 326898 218062 327134
rect 218146 326898 218382 327134
rect 210986 176378 211222 176614
rect 211306 176378 211542 176614
rect 210986 176058 211222 176294
rect 211306 176058 211542 176294
rect 210986 140378 211222 140614
rect 211306 140378 211542 140614
rect 210986 140058 211222 140294
rect 211306 140058 211542 140294
rect 210986 104378 211222 104614
rect 211306 104378 211542 104614
rect 210986 104058 211222 104294
rect 211306 104058 211542 104294
rect 225266 370658 225502 370894
rect 225586 370658 225822 370894
rect 225266 370338 225502 370574
rect 225586 370338 225822 370574
rect 221546 366938 221782 367174
rect 221866 366938 222102 367174
rect 221546 366618 221782 366854
rect 221866 366618 222102 366854
rect 221546 330938 221782 331174
rect 221866 330938 222102 331174
rect 221546 330618 221782 330854
rect 221866 330618 222102 330854
rect 217826 291218 218062 291454
rect 218146 291218 218382 291454
rect 217826 290898 218062 291134
rect 218146 290898 218382 291134
rect 221546 294938 221782 295174
rect 221866 294938 222102 295174
rect 221546 294618 221782 294854
rect 221866 294618 222102 294854
rect 219810 273218 220046 273454
rect 219810 272898 220046 273134
rect 217826 219218 218062 219454
rect 218146 219218 218382 219454
rect 217826 218898 218062 219134
rect 218146 218898 218382 219134
rect 221546 222938 221782 223174
rect 221866 222938 222102 223174
rect 221546 222618 221782 222854
rect 221866 222618 222102 222854
rect 217826 183218 218062 183454
rect 218146 183218 218382 183454
rect 217826 182898 218062 183134
rect 218146 182898 218382 183134
rect 221546 186938 221782 187174
rect 221866 186938 222102 187174
rect 221546 186618 221782 186854
rect 221866 186618 222102 186854
rect 225266 334658 225502 334894
rect 225586 334658 225822 334894
rect 225266 334338 225502 334574
rect 225586 334338 225822 334574
rect 228986 374378 229222 374614
rect 229306 374378 229542 374614
rect 228986 374058 229222 374294
rect 229306 374058 229542 374294
rect 228986 338378 229222 338614
rect 229306 338378 229542 338614
rect 228986 338058 229222 338294
rect 229306 338058 229542 338294
rect 225266 298658 225502 298894
rect 225586 298658 225822 298894
rect 225266 298338 225502 298574
rect 225586 298338 225822 298574
rect 225266 226658 225502 226894
rect 225586 226658 225822 226894
rect 225266 226338 225502 226574
rect 225586 226338 225822 226574
rect 225266 190658 225502 190894
rect 225586 190658 225822 190894
rect 225266 190338 225502 190574
rect 225586 190338 225822 190574
rect 228986 302378 229222 302614
rect 229306 302378 229542 302614
rect 228986 302058 229222 302294
rect 229306 302058 229542 302294
rect 228986 230378 229222 230614
rect 229306 230378 229542 230614
rect 228986 230058 229222 230294
rect 229306 230058 229542 230294
rect 228986 194378 229222 194614
rect 229306 194378 229542 194614
rect 228986 194058 229222 194294
rect 229306 194058 229542 194294
rect 221249 165218 221485 165454
rect 221249 164898 221485 165134
rect 224513 165218 224749 165454
rect 224513 164898 224749 165134
rect 219617 147218 219853 147454
rect 219617 146898 219853 147134
rect 222881 147218 223117 147454
rect 222881 146898 223117 147134
rect 226145 147218 226381 147454
rect 226145 146898 226381 147134
rect 235826 345218 236062 345454
rect 236146 345218 236382 345454
rect 235826 344898 236062 345134
rect 236146 344898 236382 345134
rect 235826 309218 236062 309454
rect 236146 309218 236382 309454
rect 235826 308898 236062 309134
rect 236146 308898 236382 309134
rect 239546 348938 239782 349174
rect 239866 348938 240102 349174
rect 239546 348618 239782 348854
rect 239866 348618 240102 348854
rect 239546 312938 239782 313174
rect 239866 312938 240102 313174
rect 239546 312618 239782 312854
rect 239866 312618 240102 312854
rect 235170 255218 235406 255454
rect 235170 254898 235406 255134
rect 235826 237218 236062 237454
rect 236146 237218 236382 237454
rect 235826 236898 236062 237134
rect 236146 236898 236382 237134
rect 235826 201218 236062 201454
rect 236146 201218 236382 201454
rect 235826 200898 236062 201134
rect 236146 200898 236382 201134
rect 235826 165218 236062 165454
rect 236146 165218 236382 165454
rect 235826 164898 236062 165134
rect 236146 164898 236382 165134
rect 221249 129218 221485 129454
rect 221249 128898 221485 129134
rect 224513 129218 224749 129454
rect 224513 128898 224749 129134
rect 219617 111218 219853 111454
rect 219617 110898 219853 111134
rect 222881 111218 223117 111454
rect 222881 110898 223117 111134
rect 226145 111218 226381 111454
rect 226145 110898 226381 111134
rect 210986 68378 211222 68614
rect 211306 68378 211542 68614
rect 210986 68058 211222 68294
rect 211306 68058 211542 68294
rect 210986 32378 211222 32614
rect 211306 32378 211542 32614
rect 210986 32058 211222 32294
rect 211306 32058 211542 32294
rect 192986 -6342 193222 -6106
rect 193306 -6342 193542 -6106
rect 192986 -6662 193222 -6426
rect 193306 -6662 193542 -6426
rect 217826 75218 218062 75454
rect 218146 75218 218382 75454
rect 217826 74898 218062 75134
rect 218146 74898 218382 75134
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 221546 78938 221782 79174
rect 221866 78938 222102 79174
rect 221546 78618 221782 78854
rect 221866 78618 222102 78854
rect 221546 42938 221782 43174
rect 221866 42938 222102 43174
rect 221546 42618 221782 42854
rect 221866 42618 222102 42854
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 225266 82658 225502 82894
rect 225586 82658 225822 82894
rect 225266 82338 225502 82574
rect 225586 82338 225822 82574
rect 225266 46658 225502 46894
rect 225586 46658 225822 46894
rect 225266 46338 225502 46574
rect 225586 46338 225822 46574
rect 221546 6938 221782 7174
rect 221866 6938 222102 7174
rect 221546 6618 221782 6854
rect 221866 6618 222102 6854
rect 221546 -2502 221782 -2266
rect 221866 -2502 222102 -2266
rect 221546 -2822 221782 -2586
rect 221866 -2822 222102 -2586
rect 225266 10658 225502 10894
rect 225586 10658 225822 10894
rect 225266 10338 225502 10574
rect 225586 10338 225822 10574
rect 228986 86378 229222 86614
rect 229306 86378 229542 86614
rect 228986 86058 229222 86294
rect 229306 86058 229542 86294
rect 228986 50378 229222 50614
rect 229306 50378 229542 50614
rect 228986 50058 229222 50294
rect 229306 50058 229542 50294
rect 239546 204938 239782 205174
rect 239866 204938 240102 205174
rect 239546 204618 239782 204854
rect 239866 204618 240102 204854
rect 243266 352658 243502 352894
rect 243586 352658 243822 352894
rect 243266 352338 243502 352574
rect 243586 352338 243822 352574
rect 243266 316658 243502 316894
rect 243586 316658 243822 316894
rect 243266 316338 243502 316574
rect 243586 316338 243822 316574
rect 246986 356378 247222 356614
rect 247306 356378 247542 356614
rect 246986 356058 247222 356294
rect 247306 356058 247542 356294
rect 253826 363218 254062 363454
rect 254146 363218 254382 363454
rect 253826 362898 254062 363134
rect 254146 362898 254382 363134
rect 246986 320378 247222 320614
rect 247306 320378 247542 320614
rect 246986 320058 247222 320294
rect 247306 320058 247542 320294
rect 246986 284378 247222 284614
rect 247306 284378 247542 284614
rect 246986 284058 247222 284294
rect 247306 284058 247542 284294
rect 246986 248378 247222 248614
rect 247306 248378 247542 248614
rect 246986 248058 247222 248294
rect 247306 248058 247542 248294
rect 243266 208658 243502 208894
rect 243586 208658 243822 208894
rect 243266 208338 243502 208574
rect 243586 208338 243822 208574
rect 239546 168938 239782 169174
rect 239866 168938 240102 169174
rect 239546 168618 239782 168854
rect 239866 168618 240102 168854
rect 235826 129218 236062 129454
rect 236146 129218 236382 129454
rect 235826 128898 236062 129134
rect 236146 128898 236382 129134
rect 239546 132938 239782 133174
rect 239866 132938 240102 133174
rect 239546 132618 239782 132854
rect 239866 132618 240102 132854
rect 235826 93218 236062 93454
rect 236146 93218 236382 93454
rect 235826 92898 236062 93134
rect 236146 92898 236382 93134
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 228986 14378 229222 14614
rect 229306 14378 229542 14614
rect 228986 14058 229222 14294
rect 229306 14058 229542 14294
rect 225266 -4422 225502 -4186
rect 225586 -4422 225822 -4186
rect 225266 -4742 225502 -4506
rect 225586 -4742 225822 -4506
rect 210986 -7302 211222 -7066
rect 211306 -7302 211542 -7066
rect 210986 -7622 211222 -7386
rect 211306 -7622 211542 -7386
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -1542 236062 -1306
rect 236146 -1542 236382 -1306
rect 235826 -1862 236062 -1626
rect 236146 -1862 236382 -1626
rect 239546 96938 239782 97174
rect 239866 96938 240102 97174
rect 239546 96618 239782 96854
rect 239866 96618 240102 96854
rect 239546 60938 239782 61174
rect 239866 60938 240102 61174
rect 239546 60618 239782 60854
rect 239866 60618 240102 60854
rect 239546 24938 239782 25174
rect 239866 24938 240102 25174
rect 239546 24618 239782 24854
rect 239866 24618 240102 24854
rect 243266 172658 243502 172894
rect 243586 172658 243822 172894
rect 246986 212378 247222 212614
rect 247306 212378 247542 212614
rect 246986 212058 247222 212294
rect 247306 212058 247542 212294
rect 243266 172338 243502 172574
rect 243586 172338 243822 172574
rect 243266 136658 243502 136894
rect 243586 136658 243822 136894
rect 243266 136338 243502 136574
rect 243586 136338 243822 136574
rect 243266 100658 243502 100894
rect 243586 100658 243822 100894
rect 243266 100338 243502 100574
rect 243586 100338 243822 100574
rect 243266 64658 243502 64894
rect 243586 64658 243822 64894
rect 243266 64338 243502 64574
rect 243586 64338 243822 64574
rect 243266 28658 243502 28894
rect 243586 28658 243822 28894
rect 243266 28338 243502 28574
rect 243586 28338 243822 28574
rect 239546 -3462 239782 -3226
rect 239866 -3462 240102 -3226
rect 239546 -3782 239782 -3546
rect 239866 -3782 240102 -3546
rect 246986 176378 247222 176614
rect 247306 176378 247542 176614
rect 246986 176058 247222 176294
rect 247306 176058 247542 176294
rect 246986 140378 247222 140614
rect 247306 140378 247542 140614
rect 246986 140058 247222 140294
rect 247306 140058 247542 140294
rect 246986 104378 247222 104614
rect 247306 104378 247542 104614
rect 246986 104058 247222 104294
rect 247306 104058 247542 104294
rect 246986 68378 247222 68614
rect 247306 68378 247542 68614
rect 246986 68058 247222 68294
rect 247306 68058 247542 68294
rect 246986 32378 247222 32614
rect 247306 32378 247542 32614
rect 246986 32058 247222 32294
rect 247306 32058 247542 32294
rect 243266 -5382 243502 -5146
rect 243586 -5382 243822 -5146
rect 243266 -5702 243502 -5466
rect 243586 -5702 243822 -5466
rect 228986 -6342 229222 -6106
rect 229306 -6342 229542 -6106
rect 228986 -6662 229222 -6426
rect 229306 -6662 229542 -6426
rect 257546 366938 257782 367174
rect 257866 366938 258102 367174
rect 257546 366618 257782 366854
rect 257866 366618 258102 366854
rect 257546 330938 257782 331174
rect 257866 330938 258102 331174
rect 257546 330618 257782 330854
rect 257866 330618 258102 330854
rect 253826 327218 254062 327454
rect 254146 327218 254382 327454
rect 253826 326898 254062 327134
rect 254146 326898 254382 327134
rect 253826 291218 254062 291454
rect 254146 291218 254382 291454
rect 253826 290898 254062 291134
rect 254146 290898 254382 291134
rect 257546 294938 257782 295174
rect 257866 294938 258102 295174
rect 257546 294618 257782 294854
rect 257866 294618 258102 294854
rect 253826 255218 254062 255454
rect 254146 255218 254382 255454
rect 253826 254898 254062 255134
rect 254146 254898 254382 255134
rect 253826 219218 254062 219454
rect 254146 219218 254382 219454
rect 253826 218898 254062 219134
rect 254146 218898 254382 219134
rect 253826 183218 254062 183454
rect 254146 183218 254382 183454
rect 253826 182898 254062 183134
rect 254146 182898 254382 183134
rect 257546 258938 257782 259174
rect 257866 258938 258102 259174
rect 257546 258618 257782 258854
rect 257866 258618 258102 258854
rect 257546 222938 257782 223174
rect 257866 222938 258102 223174
rect 257546 222618 257782 222854
rect 257866 222618 258102 222854
rect 261266 370658 261502 370894
rect 261586 370658 261822 370894
rect 261266 370338 261502 370574
rect 261586 370338 261822 370574
rect 261266 334658 261502 334894
rect 261586 334658 261822 334894
rect 261266 334338 261502 334574
rect 261586 334338 261822 334574
rect 264986 374378 265222 374614
rect 265306 374378 265542 374614
rect 264986 374058 265222 374294
rect 265306 374058 265542 374294
rect 264986 338378 265222 338614
rect 265306 338378 265542 338614
rect 264986 338058 265222 338294
rect 265306 338058 265542 338294
rect 261266 298658 261502 298894
rect 261586 298658 261822 298894
rect 261266 298338 261502 298574
rect 261586 298338 261822 298574
rect 261266 262658 261502 262894
rect 261586 262658 261822 262894
rect 261266 262338 261502 262574
rect 261586 262338 261822 262574
rect 261266 226658 261502 226894
rect 261586 226658 261822 226894
rect 261266 226338 261502 226574
rect 261586 226338 261822 226574
rect 257546 186938 257782 187174
rect 257866 186938 258102 187174
rect 257546 186618 257782 186854
rect 257866 186618 258102 186854
rect 253826 147218 254062 147454
rect 254146 147218 254382 147454
rect 253826 146898 254062 147134
rect 254146 146898 254382 147134
rect 253826 111218 254062 111454
rect 254146 111218 254382 111454
rect 253826 110898 254062 111134
rect 254146 110898 254382 111134
rect 257546 150938 257782 151174
rect 257866 150938 258102 151174
rect 257546 150618 257782 150854
rect 257866 150618 258102 150854
rect 257546 114938 257782 115174
rect 257866 114938 258102 115174
rect 257546 114618 257782 114854
rect 257866 114618 258102 114854
rect 253826 75218 254062 75454
rect 254146 75218 254382 75454
rect 253826 74898 254062 75134
rect 254146 74898 254382 75134
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 257546 78938 257782 79174
rect 257866 78938 258102 79174
rect 257546 78618 257782 78854
rect 257866 78618 258102 78854
rect 257546 42938 257782 43174
rect 257866 42938 258102 43174
rect 257546 42618 257782 42854
rect 257866 42618 258102 42854
rect 261266 190658 261502 190894
rect 261586 190658 261822 190894
rect 261266 190338 261502 190574
rect 261586 190338 261822 190574
rect 261266 154658 261502 154894
rect 261586 154658 261822 154894
rect 261266 154338 261502 154574
rect 261586 154338 261822 154574
rect 261266 118658 261502 118894
rect 261586 118658 261822 118894
rect 261266 118338 261502 118574
rect 261586 118338 261822 118574
rect 261266 82658 261502 82894
rect 261586 82658 261822 82894
rect 261266 82338 261502 82574
rect 261586 82338 261822 82574
rect 264986 302378 265222 302614
rect 265306 302378 265542 302614
rect 264986 302058 265222 302294
rect 265306 302058 265542 302294
rect 264986 266378 265222 266614
rect 265306 266378 265542 266614
rect 264986 266058 265222 266294
rect 265306 266058 265542 266294
rect 264986 230378 265222 230614
rect 265306 230378 265542 230614
rect 264986 230058 265222 230294
rect 265306 230058 265542 230294
rect 264986 194378 265222 194614
rect 265306 194378 265542 194614
rect 264986 194058 265222 194294
rect 265306 194058 265542 194294
rect 271826 345218 272062 345454
rect 272146 345218 272382 345454
rect 271826 344898 272062 345134
rect 272146 344898 272382 345134
rect 271826 309218 272062 309454
rect 272146 309218 272382 309454
rect 271826 308898 272062 309134
rect 272146 308898 272382 309134
rect 271826 273218 272062 273454
rect 272146 273218 272382 273454
rect 271826 272898 272062 273134
rect 272146 272898 272382 273134
rect 271826 237218 272062 237454
rect 272146 237218 272382 237454
rect 271826 236898 272062 237134
rect 272146 236898 272382 237134
rect 271826 201218 272062 201454
rect 272146 201218 272382 201454
rect 271826 200898 272062 201134
rect 272146 200898 272382 201134
rect 275546 348938 275782 349174
rect 275866 348938 276102 349174
rect 275546 348618 275782 348854
rect 275866 348618 276102 348854
rect 279266 352658 279502 352894
rect 279586 352658 279822 352894
rect 279266 352338 279502 352574
rect 279586 352338 279822 352574
rect 279266 316658 279502 316894
rect 279586 316658 279822 316894
rect 279266 316338 279502 316574
rect 279586 316338 279822 316574
rect 275546 312938 275782 313174
rect 275866 312938 276102 313174
rect 275546 312618 275782 312854
rect 275866 312618 276102 312854
rect 275546 276938 275782 277174
rect 275866 276938 276102 277174
rect 275546 276618 275782 276854
rect 275866 276618 276102 276854
rect 275546 240938 275782 241174
rect 275866 240938 276102 241174
rect 275546 240618 275782 240854
rect 275866 240618 276102 240854
rect 275546 204938 275782 205174
rect 275866 204938 276102 205174
rect 275546 204618 275782 204854
rect 275866 204618 276102 204854
rect 282986 356378 283222 356614
rect 283306 356378 283542 356614
rect 282986 356058 283222 356294
rect 283306 356058 283542 356294
rect 282986 320378 283222 320614
rect 283306 320378 283542 320614
rect 282986 320058 283222 320294
rect 283306 320058 283542 320294
rect 279266 280658 279502 280894
rect 279586 280658 279822 280894
rect 279266 280338 279502 280574
rect 279586 280338 279822 280574
rect 279266 244658 279502 244894
rect 279586 244658 279822 244894
rect 279266 244338 279502 244574
rect 279586 244338 279822 244574
rect 279266 208658 279502 208894
rect 279586 208658 279822 208894
rect 279266 208338 279502 208574
rect 279586 208338 279822 208574
rect 272249 165218 272485 165454
rect 272249 164898 272485 165134
rect 275513 165218 275749 165454
rect 275513 164898 275749 165134
rect 264986 158378 265222 158614
rect 265306 158378 265542 158614
rect 264986 158058 265222 158294
rect 265306 158058 265542 158294
rect 261266 46658 261502 46894
rect 261586 46658 261822 46894
rect 261266 46338 261502 46574
rect 261586 46338 261822 46574
rect 257546 6938 257782 7174
rect 257866 6938 258102 7174
rect 257546 6618 257782 6854
rect 257866 6618 258102 6854
rect 257546 -2502 257782 -2266
rect 257866 -2502 258102 -2266
rect 257546 -2822 257782 -2586
rect 257866 -2822 258102 -2586
rect 270617 147218 270853 147454
rect 270617 146898 270853 147134
rect 273881 147218 274117 147454
rect 273881 146898 274117 147134
rect 277145 147218 277381 147454
rect 277145 146898 277381 147134
rect 264986 122378 265222 122614
rect 265306 122378 265542 122614
rect 264986 122058 265222 122294
rect 265306 122058 265542 122294
rect 264986 86378 265222 86614
rect 265306 86378 265542 86614
rect 264986 86058 265222 86294
rect 265306 86058 265542 86294
rect 264986 50378 265222 50614
rect 265306 50378 265542 50614
rect 264986 50058 265222 50294
rect 265306 50058 265542 50294
rect 261266 10658 261502 10894
rect 261586 10658 261822 10894
rect 261266 10338 261502 10574
rect 261586 10338 261822 10574
rect 261266 -4422 261502 -4186
rect 261586 -4422 261822 -4186
rect 261266 -4742 261502 -4506
rect 261586 -4742 261822 -4506
rect 272249 129218 272485 129454
rect 272249 128898 272485 129134
rect 275513 129218 275749 129454
rect 275513 128898 275749 129134
rect 282986 284378 283222 284614
rect 283306 284378 283542 284614
rect 282986 284058 283222 284294
rect 283306 284058 283542 284294
rect 282986 248378 283222 248614
rect 283306 248378 283542 248614
rect 282986 248058 283222 248294
rect 283306 248058 283542 248294
rect 282986 212378 283222 212614
rect 283306 212378 283542 212614
rect 282986 212058 283222 212294
rect 283306 212058 283542 212294
rect 282986 176378 283222 176614
rect 283306 176378 283542 176614
rect 282986 176058 283222 176294
rect 283306 176058 283542 176294
rect 282986 140378 283222 140614
rect 283306 140378 283542 140614
rect 282986 140058 283222 140294
rect 283306 140058 283542 140294
rect 270617 111218 270853 111454
rect 270617 110898 270853 111134
rect 273881 111218 274117 111454
rect 273881 110898 274117 111134
rect 277145 111218 277381 111454
rect 277145 110898 277381 111134
rect 282986 104378 283222 104614
rect 283306 104378 283542 104614
rect 282986 104058 283222 104294
rect 283306 104058 283542 104294
rect 271826 93218 272062 93454
rect 272146 93218 272382 93454
rect 271826 92898 272062 93134
rect 272146 92898 272382 93134
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 264986 14378 265222 14614
rect 265306 14378 265542 14614
rect 264986 14058 265222 14294
rect 265306 14058 265542 14294
rect 246986 -7302 247222 -7066
rect 247306 -7302 247542 -7066
rect 246986 -7622 247222 -7386
rect 247306 -7622 247542 -7386
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -1542 272062 -1306
rect 272146 -1542 272382 -1306
rect 271826 -1862 272062 -1626
rect 272146 -1862 272382 -1626
rect 275546 60938 275782 61174
rect 275866 60938 276102 61174
rect 275546 60618 275782 60854
rect 275866 60618 276102 60854
rect 275546 24938 275782 25174
rect 275866 24938 276102 25174
rect 275546 24618 275782 24854
rect 275866 24618 276102 24854
rect 275546 -3462 275782 -3226
rect 275866 -3462 276102 -3226
rect 275546 -3782 275782 -3546
rect 275866 -3782 276102 -3546
rect 279266 64658 279502 64894
rect 279586 64658 279822 64894
rect 279266 64338 279502 64574
rect 279586 64338 279822 64574
rect 279266 28658 279502 28894
rect 279586 28658 279822 28894
rect 279266 28338 279502 28574
rect 279586 28338 279822 28574
rect 279266 -5382 279502 -5146
rect 279586 -5382 279822 -5146
rect 279266 -5702 279502 -5466
rect 279586 -5702 279822 -5466
rect 282986 68378 283222 68614
rect 283306 68378 283542 68614
rect 282986 68058 283222 68294
rect 283306 68058 283542 68294
rect 282986 32378 283222 32614
rect 283306 32378 283542 32614
rect 282986 32058 283222 32294
rect 283306 32058 283542 32294
rect 264986 -6342 265222 -6106
rect 265306 -6342 265542 -6106
rect 264986 -6662 265222 -6426
rect 265306 -6662 265542 -6426
rect 289826 363218 290062 363454
rect 290146 363218 290382 363454
rect 289826 362898 290062 363134
rect 290146 362898 290382 363134
rect 289826 327218 290062 327454
rect 290146 327218 290382 327454
rect 289826 326898 290062 327134
rect 290146 326898 290382 327134
rect 293546 366938 293782 367174
rect 293866 366938 294102 367174
rect 293546 366618 293782 366854
rect 293866 366618 294102 366854
rect 297266 370658 297502 370894
rect 297586 370658 297822 370894
rect 297266 370338 297502 370574
rect 297586 370338 297822 370574
rect 293546 330938 293782 331174
rect 293866 330938 294102 331174
rect 293546 330618 293782 330854
rect 293866 330618 294102 330854
rect 289826 291218 290062 291454
rect 290146 291218 290382 291454
rect 289826 290898 290062 291134
rect 290146 290898 290382 291134
rect 289826 255218 290062 255454
rect 290146 255218 290382 255454
rect 289826 254898 290062 255134
rect 290146 254898 290382 255134
rect 289826 219218 290062 219454
rect 290146 219218 290382 219454
rect 289826 218898 290062 219134
rect 290146 218898 290382 219134
rect 289826 183218 290062 183454
rect 290146 183218 290382 183454
rect 289826 182898 290062 183134
rect 290146 182898 290382 183134
rect 289826 147218 290062 147454
rect 290146 147218 290382 147454
rect 289826 146898 290062 147134
rect 290146 146898 290382 147134
rect 289826 111218 290062 111454
rect 290146 111218 290382 111454
rect 289826 110898 290062 111134
rect 290146 110898 290382 111134
rect 289826 75218 290062 75454
rect 290146 75218 290382 75454
rect 289826 74898 290062 75134
rect 290146 74898 290382 75134
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 293546 294938 293782 295174
rect 293866 294938 294102 295174
rect 293546 294618 293782 294854
rect 293866 294618 294102 294854
rect 293546 258938 293782 259174
rect 293866 258938 294102 259174
rect 293546 258618 293782 258854
rect 293866 258618 294102 258854
rect 293546 222938 293782 223174
rect 293866 222938 294102 223174
rect 293546 222618 293782 222854
rect 293866 222618 294102 222854
rect 293546 186938 293782 187174
rect 293866 186938 294102 187174
rect 293546 186618 293782 186854
rect 293866 186618 294102 186854
rect 293546 150938 293782 151174
rect 293866 150938 294102 151174
rect 293546 150618 293782 150854
rect 293866 150618 294102 150854
rect 293546 114938 293782 115174
rect 293866 114938 294102 115174
rect 293546 114618 293782 114854
rect 293866 114618 294102 114854
rect 293546 78938 293782 79174
rect 293866 78938 294102 79174
rect 293546 78618 293782 78854
rect 293866 78618 294102 78854
rect 293546 42938 293782 43174
rect 293866 42938 294102 43174
rect 293546 42618 293782 42854
rect 293866 42618 294102 42854
rect 297266 334658 297502 334894
rect 297586 334658 297822 334894
rect 297266 334338 297502 334574
rect 297586 334338 297822 334574
rect 297266 298658 297502 298894
rect 297586 298658 297822 298894
rect 297266 298338 297502 298574
rect 297586 298338 297822 298574
rect 297266 262658 297502 262894
rect 297586 262658 297822 262894
rect 297266 262338 297502 262574
rect 297586 262338 297822 262574
rect 297266 226658 297502 226894
rect 297586 226658 297822 226894
rect 297266 226338 297502 226574
rect 297586 226338 297822 226574
rect 300986 374378 301222 374614
rect 301306 374378 301542 374614
rect 300986 374058 301222 374294
rect 301306 374058 301542 374294
rect 300986 338378 301222 338614
rect 301306 338378 301542 338614
rect 300986 338058 301222 338294
rect 301306 338058 301542 338294
rect 300986 302378 301222 302614
rect 301306 302378 301542 302614
rect 300986 302058 301222 302294
rect 301306 302058 301542 302294
rect 300986 266378 301222 266614
rect 301306 266378 301542 266614
rect 300986 266058 301222 266294
rect 301306 266058 301542 266294
rect 300986 230378 301222 230614
rect 301306 230378 301542 230614
rect 300986 230058 301222 230294
rect 301306 230058 301542 230294
rect 297266 190658 297502 190894
rect 297586 190658 297822 190894
rect 297266 190338 297502 190574
rect 297586 190338 297822 190574
rect 297266 154658 297502 154894
rect 297586 154658 297822 154894
rect 297266 154338 297502 154574
rect 297586 154338 297822 154574
rect 297266 118658 297502 118894
rect 297586 118658 297822 118894
rect 297266 118338 297502 118574
rect 297586 118338 297822 118574
rect 297266 82658 297502 82894
rect 297586 82658 297822 82894
rect 297266 82338 297502 82574
rect 297586 82338 297822 82574
rect 297266 46658 297502 46894
rect 297586 46658 297822 46894
rect 297266 46338 297502 46574
rect 297586 46338 297822 46574
rect 293546 6938 293782 7174
rect 293866 6938 294102 7174
rect 293546 6618 293782 6854
rect 293866 6618 294102 6854
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 293546 -2502 293782 -2266
rect 293866 -2502 294102 -2266
rect 293546 -2822 293782 -2586
rect 293866 -2822 294102 -2586
rect 297266 10658 297502 10894
rect 297586 10658 297822 10894
rect 297266 10338 297502 10574
rect 297586 10338 297822 10574
rect 300986 194378 301222 194614
rect 301306 194378 301542 194614
rect 300986 194058 301222 194294
rect 301306 194058 301542 194294
rect 300986 158378 301222 158614
rect 301306 158378 301542 158614
rect 300986 158058 301222 158294
rect 301306 158058 301542 158294
rect 300986 122378 301222 122614
rect 301306 122378 301542 122614
rect 300986 122058 301222 122294
rect 301306 122058 301542 122294
rect 300986 86378 301222 86614
rect 301306 86378 301542 86614
rect 300986 86058 301222 86294
rect 301306 86058 301542 86294
rect 300986 50378 301222 50614
rect 301306 50378 301542 50614
rect 300986 50058 301222 50294
rect 301306 50058 301542 50294
rect 300986 14378 301222 14614
rect 301306 14378 301542 14614
rect 300986 14058 301222 14294
rect 301306 14058 301542 14294
rect 297266 -4422 297502 -4186
rect 297586 -4422 297822 -4186
rect 297266 -4742 297502 -4506
rect 297586 -4742 297822 -4506
rect 282986 -7302 283222 -7066
rect 283306 -7302 283542 -7066
rect 282986 -7622 283222 -7386
rect 283306 -7622 283542 -7386
rect 307826 345218 308062 345454
rect 308146 345218 308382 345454
rect 307826 344898 308062 345134
rect 308146 344898 308382 345134
rect 307826 309218 308062 309454
rect 308146 309218 308382 309454
rect 307826 308898 308062 309134
rect 308146 308898 308382 309134
rect 307826 273218 308062 273454
rect 308146 273218 308382 273454
rect 307826 272898 308062 273134
rect 308146 272898 308382 273134
rect 307826 237218 308062 237454
rect 308146 237218 308382 237454
rect 307826 236898 308062 237134
rect 308146 236898 308382 237134
rect 307826 201218 308062 201454
rect 308146 201218 308382 201454
rect 307826 200898 308062 201134
rect 308146 200898 308382 201134
rect 307826 165218 308062 165454
rect 308146 165218 308382 165454
rect 307826 164898 308062 165134
rect 308146 164898 308382 165134
rect 307826 129218 308062 129454
rect 308146 129218 308382 129454
rect 307826 128898 308062 129134
rect 308146 128898 308382 129134
rect 307826 93218 308062 93454
rect 308146 93218 308382 93454
rect 307826 92898 308062 93134
rect 308146 92898 308382 93134
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -1542 308062 -1306
rect 308146 -1542 308382 -1306
rect 307826 -1862 308062 -1626
rect 308146 -1862 308382 -1626
rect 311546 348938 311782 349174
rect 311866 348938 312102 349174
rect 311546 348618 311782 348854
rect 311866 348618 312102 348854
rect 311546 312938 311782 313174
rect 311866 312938 312102 313174
rect 311546 312618 311782 312854
rect 311866 312618 312102 312854
rect 311546 276938 311782 277174
rect 311866 276938 312102 277174
rect 311546 276618 311782 276854
rect 311866 276618 312102 276854
rect 311546 240938 311782 241174
rect 311866 240938 312102 241174
rect 311546 240618 311782 240854
rect 311866 240618 312102 240854
rect 311546 204938 311782 205174
rect 311866 204938 312102 205174
rect 311546 204618 311782 204854
rect 311866 204618 312102 204854
rect 311546 168938 311782 169174
rect 311866 168938 312102 169174
rect 311546 168618 311782 168854
rect 311866 168618 312102 168854
rect 311546 132938 311782 133174
rect 311866 132938 312102 133174
rect 311546 132618 311782 132854
rect 311866 132618 312102 132854
rect 311546 96938 311782 97174
rect 311866 96938 312102 97174
rect 311546 96618 311782 96854
rect 311866 96618 312102 96854
rect 311546 60938 311782 61174
rect 311866 60938 312102 61174
rect 311546 60618 311782 60854
rect 311866 60618 312102 60854
rect 311546 24938 311782 25174
rect 311866 24938 312102 25174
rect 311546 24618 311782 24854
rect 311866 24618 312102 24854
rect 311546 -3462 311782 -3226
rect 311866 -3462 312102 -3226
rect 311546 -3782 311782 -3546
rect 311866 -3782 312102 -3546
rect 315266 352658 315502 352894
rect 315586 352658 315822 352894
rect 315266 352338 315502 352574
rect 315586 352338 315822 352574
rect 315266 316658 315502 316894
rect 315586 316658 315822 316894
rect 315266 316338 315502 316574
rect 315586 316338 315822 316574
rect 315266 280658 315502 280894
rect 315586 280658 315822 280894
rect 315266 280338 315502 280574
rect 315586 280338 315822 280574
rect 315266 244658 315502 244894
rect 315586 244658 315822 244894
rect 315266 244338 315502 244574
rect 315586 244338 315822 244574
rect 315266 208658 315502 208894
rect 315586 208658 315822 208894
rect 315266 208338 315502 208574
rect 315586 208338 315822 208574
rect 315266 172658 315502 172894
rect 315586 172658 315822 172894
rect 315266 172338 315502 172574
rect 315586 172338 315822 172574
rect 315266 136658 315502 136894
rect 315586 136658 315822 136894
rect 315266 136338 315502 136574
rect 315586 136338 315822 136574
rect 315266 100658 315502 100894
rect 315586 100658 315822 100894
rect 315266 100338 315502 100574
rect 315586 100338 315822 100574
rect 315266 64658 315502 64894
rect 315586 64658 315822 64894
rect 315266 64338 315502 64574
rect 315586 64338 315822 64574
rect 315266 28658 315502 28894
rect 315586 28658 315822 28894
rect 315266 28338 315502 28574
rect 315586 28338 315822 28574
rect 315266 -5382 315502 -5146
rect 315586 -5382 315822 -5146
rect 315266 -5702 315502 -5466
rect 315586 -5702 315822 -5466
rect 318986 356378 319222 356614
rect 319306 356378 319542 356614
rect 318986 356058 319222 356294
rect 319306 356058 319542 356294
rect 318986 320378 319222 320614
rect 319306 320378 319542 320614
rect 318986 320058 319222 320294
rect 319306 320058 319542 320294
rect 318986 284378 319222 284614
rect 319306 284378 319542 284614
rect 318986 284058 319222 284294
rect 319306 284058 319542 284294
rect 318986 248378 319222 248614
rect 319306 248378 319542 248614
rect 318986 248058 319222 248294
rect 319306 248058 319542 248294
rect 318986 212378 319222 212614
rect 319306 212378 319542 212614
rect 318986 212058 319222 212294
rect 319306 212058 319542 212294
rect 318986 176378 319222 176614
rect 319306 176378 319542 176614
rect 318986 176058 319222 176294
rect 319306 176058 319542 176294
rect 318986 140378 319222 140614
rect 319306 140378 319542 140614
rect 318986 140058 319222 140294
rect 319306 140058 319542 140294
rect 318986 104378 319222 104614
rect 319306 104378 319542 104614
rect 318986 104058 319222 104294
rect 319306 104058 319542 104294
rect 318986 68378 319222 68614
rect 319306 68378 319542 68614
rect 318986 68058 319222 68294
rect 319306 68058 319542 68294
rect 318986 32378 319222 32614
rect 319306 32378 319542 32614
rect 318986 32058 319222 32294
rect 319306 32058 319542 32294
rect 300986 -6342 301222 -6106
rect 301306 -6342 301542 -6106
rect 300986 -6662 301222 -6426
rect 301306 -6662 301542 -6426
rect 325826 363218 326062 363454
rect 326146 363218 326382 363454
rect 325826 362898 326062 363134
rect 326146 362898 326382 363134
rect 325826 327218 326062 327454
rect 326146 327218 326382 327454
rect 325826 326898 326062 327134
rect 326146 326898 326382 327134
rect 325826 291218 326062 291454
rect 326146 291218 326382 291454
rect 325826 290898 326062 291134
rect 326146 290898 326382 291134
rect 325826 255218 326062 255454
rect 326146 255218 326382 255454
rect 325826 254898 326062 255134
rect 326146 254898 326382 255134
rect 325826 219218 326062 219454
rect 326146 219218 326382 219454
rect 325826 218898 326062 219134
rect 326146 218898 326382 219134
rect 325826 183218 326062 183454
rect 326146 183218 326382 183454
rect 325826 182898 326062 183134
rect 326146 182898 326382 183134
rect 325826 147218 326062 147454
rect 326146 147218 326382 147454
rect 325826 146898 326062 147134
rect 326146 146898 326382 147134
rect 325826 111218 326062 111454
rect 326146 111218 326382 111454
rect 325826 110898 326062 111134
rect 326146 110898 326382 111134
rect 325826 75218 326062 75454
rect 326146 75218 326382 75454
rect 325826 74898 326062 75134
rect 326146 74898 326382 75134
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 329546 366938 329782 367174
rect 329866 366938 330102 367174
rect 329546 366618 329782 366854
rect 329866 366618 330102 366854
rect 329546 330938 329782 331174
rect 329866 330938 330102 331174
rect 329546 330618 329782 330854
rect 329866 330618 330102 330854
rect 329546 294938 329782 295174
rect 329866 294938 330102 295174
rect 329546 294618 329782 294854
rect 329866 294618 330102 294854
rect 329546 258938 329782 259174
rect 329866 258938 330102 259174
rect 329546 258618 329782 258854
rect 329866 258618 330102 258854
rect 329546 222938 329782 223174
rect 329866 222938 330102 223174
rect 329546 222618 329782 222854
rect 329866 222618 330102 222854
rect 329546 186938 329782 187174
rect 329866 186938 330102 187174
rect 329546 186618 329782 186854
rect 329866 186618 330102 186854
rect 329546 150938 329782 151174
rect 329866 150938 330102 151174
rect 329546 150618 329782 150854
rect 329866 150618 330102 150854
rect 329546 114938 329782 115174
rect 329866 114938 330102 115174
rect 329546 114618 329782 114854
rect 329866 114618 330102 114854
rect 329546 78938 329782 79174
rect 329866 78938 330102 79174
rect 329546 78618 329782 78854
rect 329866 78618 330102 78854
rect 329546 42938 329782 43174
rect 329866 42938 330102 43174
rect 329546 42618 329782 42854
rect 329866 42618 330102 42854
rect 329546 6938 329782 7174
rect 329866 6938 330102 7174
rect 329546 6618 329782 6854
rect 329866 6618 330102 6854
rect 329546 -2502 329782 -2266
rect 329866 -2502 330102 -2266
rect 329546 -2822 329782 -2586
rect 329866 -2822 330102 -2586
rect 333266 370658 333502 370894
rect 333586 370658 333822 370894
rect 333266 370338 333502 370574
rect 333586 370338 333822 370574
rect 333266 334658 333502 334894
rect 333586 334658 333822 334894
rect 333266 334338 333502 334574
rect 333586 334338 333822 334574
rect 333266 298658 333502 298894
rect 333586 298658 333822 298894
rect 333266 298338 333502 298574
rect 333586 298338 333822 298574
rect 333266 262658 333502 262894
rect 333586 262658 333822 262894
rect 333266 262338 333502 262574
rect 333586 262338 333822 262574
rect 333266 226658 333502 226894
rect 333586 226658 333822 226894
rect 333266 226338 333502 226574
rect 333586 226338 333822 226574
rect 333266 190658 333502 190894
rect 333586 190658 333822 190894
rect 333266 190338 333502 190574
rect 333586 190338 333822 190574
rect 333266 154658 333502 154894
rect 333586 154658 333822 154894
rect 333266 154338 333502 154574
rect 333586 154338 333822 154574
rect 333266 118658 333502 118894
rect 333586 118658 333822 118894
rect 333266 118338 333502 118574
rect 333586 118338 333822 118574
rect 333266 82658 333502 82894
rect 333586 82658 333822 82894
rect 333266 82338 333502 82574
rect 333586 82338 333822 82574
rect 333266 46658 333502 46894
rect 333586 46658 333822 46894
rect 333266 46338 333502 46574
rect 333586 46338 333822 46574
rect 333266 10658 333502 10894
rect 333586 10658 333822 10894
rect 333266 10338 333502 10574
rect 333586 10338 333822 10574
rect 333266 -4422 333502 -4186
rect 333586 -4422 333822 -4186
rect 333266 -4742 333502 -4506
rect 333586 -4742 333822 -4506
rect 336986 374378 337222 374614
rect 337306 374378 337542 374614
rect 336986 374058 337222 374294
rect 337306 374058 337542 374294
rect 336986 338378 337222 338614
rect 337306 338378 337542 338614
rect 336986 338058 337222 338294
rect 337306 338058 337542 338294
rect 336986 302378 337222 302614
rect 337306 302378 337542 302614
rect 336986 302058 337222 302294
rect 337306 302058 337542 302294
rect 336986 266378 337222 266614
rect 337306 266378 337542 266614
rect 336986 266058 337222 266294
rect 337306 266058 337542 266294
rect 336986 230378 337222 230614
rect 337306 230378 337542 230614
rect 336986 230058 337222 230294
rect 337306 230058 337542 230294
rect 336986 194378 337222 194614
rect 337306 194378 337542 194614
rect 336986 194058 337222 194294
rect 337306 194058 337542 194294
rect 336986 158378 337222 158614
rect 337306 158378 337542 158614
rect 336986 158058 337222 158294
rect 337306 158058 337542 158294
rect 336986 122378 337222 122614
rect 337306 122378 337542 122614
rect 336986 122058 337222 122294
rect 337306 122058 337542 122294
rect 336986 86378 337222 86614
rect 337306 86378 337542 86614
rect 336986 86058 337222 86294
rect 337306 86058 337542 86294
rect 336986 50378 337222 50614
rect 337306 50378 337542 50614
rect 336986 50058 337222 50294
rect 337306 50058 337542 50294
rect 336986 14378 337222 14614
rect 337306 14378 337542 14614
rect 336986 14058 337222 14294
rect 337306 14058 337542 14294
rect 318986 -7302 319222 -7066
rect 319306 -7302 319542 -7066
rect 318986 -7622 319222 -7386
rect 319306 -7622 319542 -7386
rect 343826 345218 344062 345454
rect 344146 345218 344382 345454
rect 343826 344898 344062 345134
rect 344146 344898 344382 345134
rect 343826 309218 344062 309454
rect 344146 309218 344382 309454
rect 343826 308898 344062 309134
rect 344146 308898 344382 309134
rect 343826 273218 344062 273454
rect 344146 273218 344382 273454
rect 343826 272898 344062 273134
rect 344146 272898 344382 273134
rect 343826 237218 344062 237454
rect 344146 237218 344382 237454
rect 343826 236898 344062 237134
rect 344146 236898 344382 237134
rect 343826 201218 344062 201454
rect 344146 201218 344382 201454
rect 343826 200898 344062 201134
rect 344146 200898 344382 201134
rect 343826 165218 344062 165454
rect 344146 165218 344382 165454
rect 343826 164898 344062 165134
rect 344146 164898 344382 165134
rect 343826 129218 344062 129454
rect 344146 129218 344382 129454
rect 343826 128898 344062 129134
rect 344146 128898 344382 129134
rect 343826 93218 344062 93454
rect 344146 93218 344382 93454
rect 343826 92898 344062 93134
rect 344146 92898 344382 93134
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -1542 344062 -1306
rect 344146 -1542 344382 -1306
rect 343826 -1862 344062 -1626
rect 344146 -1862 344382 -1626
rect 347546 348938 347782 349174
rect 347866 348938 348102 349174
rect 347546 348618 347782 348854
rect 347866 348618 348102 348854
rect 347546 312938 347782 313174
rect 347866 312938 348102 313174
rect 347546 312618 347782 312854
rect 347866 312618 348102 312854
rect 347546 276938 347782 277174
rect 347866 276938 348102 277174
rect 347546 276618 347782 276854
rect 347866 276618 348102 276854
rect 347546 240938 347782 241174
rect 347866 240938 348102 241174
rect 347546 240618 347782 240854
rect 347866 240618 348102 240854
rect 347546 204938 347782 205174
rect 347866 204938 348102 205174
rect 347546 204618 347782 204854
rect 347866 204618 348102 204854
rect 347546 168938 347782 169174
rect 347866 168938 348102 169174
rect 347546 168618 347782 168854
rect 347866 168618 348102 168854
rect 347546 132938 347782 133174
rect 347866 132938 348102 133174
rect 347546 132618 347782 132854
rect 347866 132618 348102 132854
rect 347546 96938 347782 97174
rect 347866 96938 348102 97174
rect 347546 96618 347782 96854
rect 347866 96618 348102 96854
rect 347546 60938 347782 61174
rect 347866 60938 348102 61174
rect 347546 60618 347782 60854
rect 347866 60618 348102 60854
rect 347546 24938 347782 25174
rect 347866 24938 348102 25174
rect 347546 24618 347782 24854
rect 347866 24618 348102 24854
rect 347546 -3462 347782 -3226
rect 347866 -3462 348102 -3226
rect 347546 -3782 347782 -3546
rect 347866 -3782 348102 -3546
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 361826 543218 362062 543454
rect 362146 543218 362382 543454
rect 361826 542898 362062 543134
rect 362146 542898 362382 543134
rect 354986 356378 355222 356614
rect 355306 356378 355542 356614
rect 354986 356058 355222 356294
rect 355306 356058 355542 356294
rect 351266 352658 351502 352894
rect 351586 352658 351822 352894
rect 351266 352338 351502 352574
rect 351586 352338 351822 352574
rect 351266 316658 351502 316894
rect 351586 316658 351822 316894
rect 351266 316338 351502 316574
rect 351586 316338 351822 316574
rect 351266 280658 351502 280894
rect 351586 280658 351822 280894
rect 351266 280338 351502 280574
rect 351586 280338 351822 280574
rect 351266 244658 351502 244894
rect 351586 244658 351822 244894
rect 351266 244338 351502 244574
rect 351586 244338 351822 244574
rect 351266 208658 351502 208894
rect 351586 208658 351822 208894
rect 351266 208338 351502 208574
rect 351586 208338 351822 208574
rect 351266 172658 351502 172894
rect 351586 172658 351822 172894
rect 351266 172338 351502 172574
rect 351586 172338 351822 172574
rect 351266 136658 351502 136894
rect 351586 136658 351822 136894
rect 351266 136338 351502 136574
rect 351586 136338 351822 136574
rect 351266 100658 351502 100894
rect 351586 100658 351822 100894
rect 351266 100338 351502 100574
rect 351586 100338 351822 100574
rect 351266 64658 351502 64894
rect 351586 64658 351822 64894
rect 351266 64338 351502 64574
rect 351586 64338 351822 64574
rect 351266 28658 351502 28894
rect 351586 28658 351822 28894
rect 351266 28338 351502 28574
rect 351586 28338 351822 28574
rect 351266 -5382 351502 -5146
rect 351586 -5382 351822 -5146
rect 351266 -5702 351502 -5466
rect 351586 -5702 351822 -5466
rect 354986 320378 355222 320614
rect 355306 320378 355542 320614
rect 354986 320058 355222 320294
rect 355306 320058 355542 320294
rect 354986 284378 355222 284614
rect 355306 284378 355542 284614
rect 354986 284058 355222 284294
rect 355306 284058 355542 284294
rect 354986 248378 355222 248614
rect 355306 248378 355542 248614
rect 354986 248058 355222 248294
rect 355306 248058 355542 248294
rect 354986 212378 355222 212614
rect 355306 212378 355542 212614
rect 354986 212058 355222 212294
rect 355306 212058 355542 212294
rect 354986 176378 355222 176614
rect 355306 176378 355542 176614
rect 354986 176058 355222 176294
rect 355306 176058 355542 176294
rect 354986 140378 355222 140614
rect 355306 140378 355542 140614
rect 354986 140058 355222 140294
rect 355306 140058 355542 140294
rect 354986 104378 355222 104614
rect 355306 104378 355542 104614
rect 354986 104058 355222 104294
rect 355306 104058 355542 104294
rect 354986 68378 355222 68614
rect 355306 68378 355542 68614
rect 354986 68058 355222 68294
rect 355306 68058 355542 68294
rect 354986 32378 355222 32614
rect 355306 32378 355542 32614
rect 354986 32058 355222 32294
rect 355306 32058 355542 32294
rect 336986 -6342 337222 -6106
rect 337306 -6342 337542 -6106
rect 336986 -6662 337222 -6426
rect 337306 -6662 337542 -6426
rect 365546 690938 365782 691174
rect 365866 690938 366102 691174
rect 365546 690618 365782 690854
rect 365866 690618 366102 690854
rect 365546 654938 365782 655174
rect 365866 654938 366102 655174
rect 365546 654618 365782 654854
rect 365866 654618 366102 654854
rect 365546 618938 365782 619174
rect 365866 618938 366102 619174
rect 365546 618618 365782 618854
rect 365866 618618 366102 618854
rect 365546 582938 365782 583174
rect 365866 582938 366102 583174
rect 365546 582618 365782 582854
rect 365866 582618 366102 582854
rect 365546 546938 365782 547174
rect 365866 546938 366102 547174
rect 365546 546618 365782 546854
rect 365866 546618 366102 546854
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 361826 435218 362062 435454
rect 362146 435218 362382 435454
rect 361826 434898 362062 435134
rect 362146 434898 362382 435134
rect 361826 399218 362062 399454
rect 362146 399218 362382 399454
rect 361826 398898 362062 399134
rect 362146 398898 362382 399134
rect 361826 363218 362062 363454
rect 362146 363218 362382 363454
rect 361826 362898 362062 363134
rect 362146 362898 362382 363134
rect 361826 327218 362062 327454
rect 362146 327218 362382 327454
rect 361826 326898 362062 327134
rect 362146 326898 362382 327134
rect 361826 291218 362062 291454
rect 362146 291218 362382 291454
rect 361826 290898 362062 291134
rect 362146 290898 362382 291134
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 361826 219218 362062 219454
rect 362146 219218 362382 219454
rect 361826 218898 362062 219134
rect 362146 218898 362382 219134
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 365546 510938 365782 511174
rect 365866 510938 366102 511174
rect 365546 510618 365782 510854
rect 365866 510618 366102 510854
rect 365546 474938 365782 475174
rect 365866 474938 366102 475174
rect 365546 474618 365782 474854
rect 365866 474618 366102 474854
rect 365546 438938 365782 439174
rect 365866 438938 366102 439174
rect 365546 438618 365782 438854
rect 365866 438618 366102 438854
rect 365546 402938 365782 403174
rect 365866 402938 366102 403174
rect 365546 402618 365782 402854
rect 365866 402618 366102 402854
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 365546 366938 365782 367174
rect 365866 366938 366102 367174
rect 365546 366618 365782 366854
rect 365866 366618 366102 366854
rect 365546 330938 365782 331174
rect 365866 330938 366102 331174
rect 365546 330618 365782 330854
rect 365866 330618 366102 330854
rect 365546 294938 365782 295174
rect 365866 294938 366102 295174
rect 365546 294618 365782 294854
rect 365866 294618 366102 294854
rect 365546 258938 365782 259174
rect 365866 258938 366102 259174
rect 365546 258618 365782 258854
rect 365866 258618 366102 258854
rect 365546 222938 365782 223174
rect 365866 222938 366102 223174
rect 365546 222618 365782 222854
rect 365866 222618 366102 222854
rect 365546 186938 365782 187174
rect 365866 186938 366102 187174
rect 365546 186618 365782 186854
rect 365866 186618 366102 186854
rect 365546 150938 365782 151174
rect 365866 150938 366102 151174
rect 365546 150618 365782 150854
rect 365866 150618 366102 150854
rect 365546 114938 365782 115174
rect 365866 114938 366102 115174
rect 365546 114618 365782 114854
rect 365866 114618 366102 114854
rect 365546 78938 365782 79174
rect 365866 78938 366102 79174
rect 365546 78618 365782 78854
rect 365866 78618 366102 78854
rect 365546 42938 365782 43174
rect 365866 42938 366102 43174
rect 365546 42618 365782 42854
rect 365866 42618 366102 42854
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 365546 6938 365782 7174
rect 365866 6938 366102 7174
rect 365546 6618 365782 6854
rect 365866 6618 366102 6854
rect 365546 -2502 365782 -2266
rect 365866 -2502 366102 -2266
rect 365546 -2822 365782 -2586
rect 365866 -2822 366102 -2586
rect 369266 694658 369502 694894
rect 369586 694658 369822 694894
rect 369266 694338 369502 694574
rect 369586 694338 369822 694574
rect 369266 658658 369502 658894
rect 369586 658658 369822 658894
rect 369266 658338 369502 658574
rect 369586 658338 369822 658574
rect 369266 622658 369502 622894
rect 369586 622658 369822 622894
rect 369266 622338 369502 622574
rect 369586 622338 369822 622574
rect 369266 586658 369502 586894
rect 369586 586658 369822 586894
rect 369266 586338 369502 586574
rect 369586 586338 369822 586574
rect 369266 550658 369502 550894
rect 369586 550658 369822 550894
rect 369266 550338 369502 550574
rect 369586 550338 369822 550574
rect 369266 514658 369502 514894
rect 369586 514658 369822 514894
rect 369266 514338 369502 514574
rect 369586 514338 369822 514574
rect 369266 478658 369502 478894
rect 369586 478658 369822 478894
rect 369266 478338 369502 478574
rect 369586 478338 369822 478574
rect 369266 442658 369502 442894
rect 369586 442658 369822 442894
rect 369266 442338 369502 442574
rect 369586 442338 369822 442574
rect 369266 406658 369502 406894
rect 369586 406658 369822 406894
rect 369266 406338 369502 406574
rect 369586 406338 369822 406574
rect 369266 370658 369502 370894
rect 369586 370658 369822 370894
rect 369266 370338 369502 370574
rect 369586 370338 369822 370574
rect 369266 334658 369502 334894
rect 369586 334658 369822 334894
rect 369266 334338 369502 334574
rect 369586 334338 369822 334574
rect 369266 298658 369502 298894
rect 369586 298658 369822 298894
rect 369266 298338 369502 298574
rect 369586 298338 369822 298574
rect 369266 262658 369502 262894
rect 369586 262658 369822 262894
rect 369266 262338 369502 262574
rect 369586 262338 369822 262574
rect 369266 226658 369502 226894
rect 369586 226658 369822 226894
rect 369266 226338 369502 226574
rect 369586 226338 369822 226574
rect 369266 190658 369502 190894
rect 369586 190658 369822 190894
rect 369266 190338 369502 190574
rect 369586 190338 369822 190574
rect 369266 154658 369502 154894
rect 369586 154658 369822 154894
rect 369266 154338 369502 154574
rect 369586 154338 369822 154574
rect 369266 118658 369502 118894
rect 369586 118658 369822 118894
rect 369266 118338 369502 118574
rect 369586 118338 369822 118574
rect 369266 82658 369502 82894
rect 369586 82658 369822 82894
rect 369266 82338 369502 82574
rect 369586 82338 369822 82574
rect 369266 46658 369502 46894
rect 369586 46658 369822 46894
rect 369266 46338 369502 46574
rect 369586 46338 369822 46574
rect 369266 10658 369502 10894
rect 369586 10658 369822 10894
rect 369266 10338 369502 10574
rect 369586 10338 369822 10574
rect 369266 -4422 369502 -4186
rect 369586 -4422 369822 -4186
rect 369266 -4742 369502 -4506
rect 369586 -4742 369822 -4506
rect 390986 711322 391222 711558
rect 391306 711322 391542 711558
rect 390986 711002 391222 711238
rect 391306 711002 391542 711238
rect 387266 709402 387502 709638
rect 387586 709402 387822 709638
rect 387266 709082 387502 709318
rect 387586 709082 387822 709318
rect 383546 707482 383782 707718
rect 383866 707482 384102 707718
rect 383546 707162 383782 707398
rect 383866 707162 384102 707398
rect 372986 698378 373222 698614
rect 373306 698378 373542 698614
rect 372986 698058 373222 698294
rect 373306 698058 373542 698294
rect 372986 662378 373222 662614
rect 373306 662378 373542 662614
rect 372986 662058 373222 662294
rect 373306 662058 373542 662294
rect 372986 626378 373222 626614
rect 373306 626378 373542 626614
rect 372986 626058 373222 626294
rect 373306 626058 373542 626294
rect 372986 590378 373222 590614
rect 373306 590378 373542 590614
rect 372986 590058 373222 590294
rect 373306 590058 373542 590294
rect 372986 554378 373222 554614
rect 373306 554378 373542 554614
rect 372986 554058 373222 554294
rect 373306 554058 373542 554294
rect 372986 518378 373222 518614
rect 373306 518378 373542 518614
rect 372986 518058 373222 518294
rect 373306 518058 373542 518294
rect 372986 482378 373222 482614
rect 373306 482378 373542 482614
rect 372986 482058 373222 482294
rect 373306 482058 373542 482294
rect 372986 446378 373222 446614
rect 373306 446378 373542 446614
rect 372986 446058 373222 446294
rect 373306 446058 373542 446294
rect 372986 410378 373222 410614
rect 373306 410378 373542 410614
rect 372986 410058 373222 410294
rect 373306 410058 373542 410294
rect 372986 374378 373222 374614
rect 373306 374378 373542 374614
rect 372986 374058 373222 374294
rect 373306 374058 373542 374294
rect 372986 338378 373222 338614
rect 373306 338378 373542 338614
rect 372986 338058 373222 338294
rect 373306 338058 373542 338294
rect 372986 302378 373222 302614
rect 373306 302378 373542 302614
rect 372986 302058 373222 302294
rect 373306 302058 373542 302294
rect 372986 266378 373222 266614
rect 373306 266378 373542 266614
rect 372986 266058 373222 266294
rect 373306 266058 373542 266294
rect 372986 230378 373222 230614
rect 373306 230378 373542 230614
rect 372986 230058 373222 230294
rect 373306 230058 373542 230294
rect 372986 194378 373222 194614
rect 373306 194378 373542 194614
rect 372986 194058 373222 194294
rect 373306 194058 373542 194294
rect 372986 158378 373222 158614
rect 373306 158378 373542 158614
rect 372986 158058 373222 158294
rect 373306 158058 373542 158294
rect 372986 122378 373222 122614
rect 373306 122378 373542 122614
rect 372986 122058 373222 122294
rect 373306 122058 373542 122294
rect 372986 86378 373222 86614
rect 373306 86378 373542 86614
rect 372986 86058 373222 86294
rect 373306 86058 373542 86294
rect 372986 50378 373222 50614
rect 373306 50378 373542 50614
rect 372986 50058 373222 50294
rect 373306 50058 373542 50294
rect 372986 14378 373222 14614
rect 373306 14378 373542 14614
rect 372986 14058 373222 14294
rect 373306 14058 373542 14294
rect 354986 -7302 355222 -7066
rect 355306 -7302 355542 -7066
rect 354986 -7622 355222 -7386
rect 355306 -7622 355542 -7386
rect 379826 705562 380062 705798
rect 380146 705562 380382 705798
rect 379826 705242 380062 705478
rect 380146 705242 380382 705478
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 379826 633218 380062 633454
rect 380146 633218 380382 633454
rect 379826 632898 380062 633134
rect 380146 632898 380382 633134
rect 379826 597218 380062 597454
rect 380146 597218 380382 597454
rect 379826 596898 380062 597134
rect 380146 596898 380382 597134
rect 379826 561218 380062 561454
rect 380146 561218 380382 561454
rect 379826 560898 380062 561134
rect 380146 560898 380382 561134
rect 379826 525218 380062 525454
rect 380146 525218 380382 525454
rect 379826 524898 380062 525134
rect 380146 524898 380382 525134
rect 379826 489218 380062 489454
rect 380146 489218 380382 489454
rect 379826 488898 380062 489134
rect 380146 488898 380382 489134
rect 379826 453218 380062 453454
rect 380146 453218 380382 453454
rect 379826 452898 380062 453134
rect 380146 452898 380382 453134
rect 379826 417218 380062 417454
rect 380146 417218 380382 417454
rect 379826 416898 380062 417134
rect 380146 416898 380382 417134
rect 379826 381218 380062 381454
rect 380146 381218 380382 381454
rect 379826 380898 380062 381134
rect 380146 380898 380382 381134
rect 379826 345218 380062 345454
rect 380146 345218 380382 345454
rect 379826 344898 380062 345134
rect 380146 344898 380382 345134
rect 379826 309218 380062 309454
rect 380146 309218 380382 309454
rect 379826 308898 380062 309134
rect 380146 308898 380382 309134
rect 379826 273218 380062 273454
rect 380146 273218 380382 273454
rect 379826 272898 380062 273134
rect 380146 272898 380382 273134
rect 379826 237218 380062 237454
rect 380146 237218 380382 237454
rect 379826 236898 380062 237134
rect 380146 236898 380382 237134
rect 379826 201218 380062 201454
rect 380146 201218 380382 201454
rect 379826 200898 380062 201134
rect 380146 200898 380382 201134
rect 379826 165218 380062 165454
rect 380146 165218 380382 165454
rect 379826 164898 380062 165134
rect 380146 164898 380382 165134
rect 379826 129218 380062 129454
rect 380146 129218 380382 129454
rect 379826 128898 380062 129134
rect 380146 128898 380382 129134
rect 379826 93218 380062 93454
rect 380146 93218 380382 93454
rect 379826 92898 380062 93134
rect 380146 92898 380382 93134
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -1542 380062 -1306
rect 380146 -1542 380382 -1306
rect 379826 -1862 380062 -1626
rect 380146 -1862 380382 -1626
rect 383546 672938 383782 673174
rect 383866 672938 384102 673174
rect 383546 672618 383782 672854
rect 383866 672618 384102 672854
rect 383546 636938 383782 637174
rect 383866 636938 384102 637174
rect 383546 636618 383782 636854
rect 383866 636618 384102 636854
rect 383546 600938 383782 601174
rect 383866 600938 384102 601174
rect 383546 600618 383782 600854
rect 383866 600618 384102 600854
rect 383546 564938 383782 565174
rect 383866 564938 384102 565174
rect 383546 564618 383782 564854
rect 383866 564618 384102 564854
rect 383546 528938 383782 529174
rect 383866 528938 384102 529174
rect 383546 528618 383782 528854
rect 383866 528618 384102 528854
rect 383546 492938 383782 493174
rect 383866 492938 384102 493174
rect 383546 492618 383782 492854
rect 383866 492618 384102 492854
rect 383546 456938 383782 457174
rect 383866 456938 384102 457174
rect 383546 456618 383782 456854
rect 383866 456618 384102 456854
rect 383546 420938 383782 421174
rect 383866 420938 384102 421174
rect 383546 420618 383782 420854
rect 383866 420618 384102 420854
rect 383546 384938 383782 385174
rect 383866 384938 384102 385174
rect 383546 384618 383782 384854
rect 383866 384618 384102 384854
rect 383546 348938 383782 349174
rect 383866 348938 384102 349174
rect 383546 348618 383782 348854
rect 383866 348618 384102 348854
rect 383546 312938 383782 313174
rect 383866 312938 384102 313174
rect 383546 312618 383782 312854
rect 383866 312618 384102 312854
rect 383546 276938 383782 277174
rect 383866 276938 384102 277174
rect 383546 276618 383782 276854
rect 383866 276618 384102 276854
rect 383546 240938 383782 241174
rect 383866 240938 384102 241174
rect 383546 240618 383782 240854
rect 383866 240618 384102 240854
rect 383546 204938 383782 205174
rect 383866 204938 384102 205174
rect 383546 204618 383782 204854
rect 383866 204618 384102 204854
rect 383546 168938 383782 169174
rect 383866 168938 384102 169174
rect 383546 168618 383782 168854
rect 383866 168618 384102 168854
rect 383546 132938 383782 133174
rect 383866 132938 384102 133174
rect 383546 132618 383782 132854
rect 383866 132618 384102 132854
rect 383546 96938 383782 97174
rect 383866 96938 384102 97174
rect 383546 96618 383782 96854
rect 383866 96618 384102 96854
rect 383546 60938 383782 61174
rect 383866 60938 384102 61174
rect 383546 60618 383782 60854
rect 383866 60618 384102 60854
rect 383546 24938 383782 25174
rect 383866 24938 384102 25174
rect 383546 24618 383782 24854
rect 383866 24618 384102 24854
rect 383546 -3462 383782 -3226
rect 383866 -3462 384102 -3226
rect 383546 -3782 383782 -3546
rect 383866 -3782 384102 -3546
rect 387266 676658 387502 676894
rect 387586 676658 387822 676894
rect 387266 676338 387502 676574
rect 387586 676338 387822 676574
rect 387266 640658 387502 640894
rect 387586 640658 387822 640894
rect 387266 640338 387502 640574
rect 387586 640338 387822 640574
rect 387266 604658 387502 604894
rect 387586 604658 387822 604894
rect 387266 604338 387502 604574
rect 387586 604338 387822 604574
rect 387266 568658 387502 568894
rect 387586 568658 387822 568894
rect 387266 568338 387502 568574
rect 387586 568338 387822 568574
rect 387266 532658 387502 532894
rect 387586 532658 387822 532894
rect 387266 532338 387502 532574
rect 387586 532338 387822 532574
rect 387266 496658 387502 496894
rect 387586 496658 387822 496894
rect 387266 496338 387502 496574
rect 387586 496338 387822 496574
rect 387266 460658 387502 460894
rect 387586 460658 387822 460894
rect 387266 460338 387502 460574
rect 387586 460338 387822 460574
rect 387266 424658 387502 424894
rect 387586 424658 387822 424894
rect 387266 424338 387502 424574
rect 387586 424338 387822 424574
rect 387266 388658 387502 388894
rect 387586 388658 387822 388894
rect 387266 388338 387502 388574
rect 387586 388338 387822 388574
rect 387266 352658 387502 352894
rect 387586 352658 387822 352894
rect 387266 352338 387502 352574
rect 387586 352338 387822 352574
rect 387266 316658 387502 316894
rect 387586 316658 387822 316894
rect 387266 316338 387502 316574
rect 387586 316338 387822 316574
rect 387266 280658 387502 280894
rect 387586 280658 387822 280894
rect 387266 280338 387502 280574
rect 387586 280338 387822 280574
rect 387266 244658 387502 244894
rect 387586 244658 387822 244894
rect 387266 244338 387502 244574
rect 387586 244338 387822 244574
rect 387266 208658 387502 208894
rect 387586 208658 387822 208894
rect 387266 208338 387502 208574
rect 387586 208338 387822 208574
rect 387266 172658 387502 172894
rect 387586 172658 387822 172894
rect 387266 172338 387502 172574
rect 387586 172338 387822 172574
rect 387266 136658 387502 136894
rect 387586 136658 387822 136894
rect 387266 136338 387502 136574
rect 387586 136338 387822 136574
rect 387266 100658 387502 100894
rect 387586 100658 387822 100894
rect 387266 100338 387502 100574
rect 387586 100338 387822 100574
rect 387266 64658 387502 64894
rect 387586 64658 387822 64894
rect 387266 64338 387502 64574
rect 387586 64338 387822 64574
rect 387266 28658 387502 28894
rect 387586 28658 387822 28894
rect 387266 28338 387502 28574
rect 387586 28338 387822 28574
rect 387266 -5382 387502 -5146
rect 387586 -5382 387822 -5146
rect 387266 -5702 387502 -5466
rect 387586 -5702 387822 -5466
rect 408986 710362 409222 710598
rect 409306 710362 409542 710598
rect 408986 710042 409222 710278
rect 409306 710042 409542 710278
rect 405266 708442 405502 708678
rect 405586 708442 405822 708678
rect 405266 708122 405502 708358
rect 405586 708122 405822 708358
rect 401546 706522 401782 706758
rect 401866 706522 402102 706758
rect 401546 706202 401782 706438
rect 401866 706202 402102 706438
rect 390986 680378 391222 680614
rect 391306 680378 391542 680614
rect 390986 680058 391222 680294
rect 391306 680058 391542 680294
rect 390986 644378 391222 644614
rect 391306 644378 391542 644614
rect 390986 644058 391222 644294
rect 391306 644058 391542 644294
rect 390986 608378 391222 608614
rect 391306 608378 391542 608614
rect 390986 608058 391222 608294
rect 391306 608058 391542 608294
rect 390986 572378 391222 572614
rect 391306 572378 391542 572614
rect 390986 572058 391222 572294
rect 391306 572058 391542 572294
rect 390986 536378 391222 536614
rect 391306 536378 391542 536614
rect 390986 536058 391222 536294
rect 391306 536058 391542 536294
rect 390986 500378 391222 500614
rect 391306 500378 391542 500614
rect 390986 500058 391222 500294
rect 391306 500058 391542 500294
rect 390986 464378 391222 464614
rect 391306 464378 391542 464614
rect 390986 464058 391222 464294
rect 391306 464058 391542 464294
rect 390986 428378 391222 428614
rect 391306 428378 391542 428614
rect 390986 428058 391222 428294
rect 391306 428058 391542 428294
rect 390986 392378 391222 392614
rect 391306 392378 391542 392614
rect 390986 392058 391222 392294
rect 391306 392058 391542 392294
rect 390986 356378 391222 356614
rect 391306 356378 391542 356614
rect 390986 356058 391222 356294
rect 391306 356058 391542 356294
rect 390986 320378 391222 320614
rect 391306 320378 391542 320614
rect 390986 320058 391222 320294
rect 391306 320058 391542 320294
rect 390986 284378 391222 284614
rect 391306 284378 391542 284614
rect 390986 284058 391222 284294
rect 391306 284058 391542 284294
rect 390986 248378 391222 248614
rect 391306 248378 391542 248614
rect 390986 248058 391222 248294
rect 391306 248058 391542 248294
rect 390986 212378 391222 212614
rect 391306 212378 391542 212614
rect 390986 212058 391222 212294
rect 391306 212058 391542 212294
rect 390986 176378 391222 176614
rect 391306 176378 391542 176614
rect 390986 176058 391222 176294
rect 391306 176058 391542 176294
rect 390986 140378 391222 140614
rect 391306 140378 391542 140614
rect 390986 140058 391222 140294
rect 391306 140058 391542 140294
rect 390986 104378 391222 104614
rect 391306 104378 391542 104614
rect 390986 104058 391222 104294
rect 391306 104058 391542 104294
rect 390986 68378 391222 68614
rect 391306 68378 391542 68614
rect 390986 68058 391222 68294
rect 391306 68058 391542 68294
rect 390986 32378 391222 32614
rect 391306 32378 391542 32614
rect 390986 32058 391222 32294
rect 391306 32058 391542 32294
rect 372986 -6342 373222 -6106
rect 373306 -6342 373542 -6106
rect 372986 -6662 373222 -6426
rect 373306 -6662 373542 -6426
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 397826 543218 398062 543454
rect 398146 543218 398382 543454
rect 397826 542898 398062 543134
rect 398146 542898 398382 543134
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 397826 435218 398062 435454
rect 398146 435218 398382 435454
rect 397826 434898 398062 435134
rect 398146 434898 398382 435134
rect 397826 399218 398062 399454
rect 398146 399218 398382 399454
rect 397826 398898 398062 399134
rect 398146 398898 398382 399134
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 397826 327218 398062 327454
rect 398146 327218 398382 327454
rect 397826 326898 398062 327134
rect 398146 326898 398382 327134
rect 397826 291218 398062 291454
rect 398146 291218 398382 291454
rect 397826 290898 398062 291134
rect 398146 290898 398382 291134
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 397826 219218 398062 219454
rect 398146 219218 398382 219454
rect 397826 218898 398062 219134
rect 398146 218898 398382 219134
rect 397826 183218 398062 183454
rect 398146 183218 398382 183454
rect 397826 182898 398062 183134
rect 398146 182898 398382 183134
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 397826 111218 398062 111454
rect 398146 111218 398382 111454
rect 397826 110898 398062 111134
rect 398146 110898 398382 111134
rect 397826 75218 398062 75454
rect 398146 75218 398382 75454
rect 397826 74898 398062 75134
rect 398146 74898 398382 75134
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 401546 690938 401782 691174
rect 401866 690938 402102 691174
rect 401546 690618 401782 690854
rect 401866 690618 402102 690854
rect 401546 654938 401782 655174
rect 401866 654938 402102 655174
rect 401546 654618 401782 654854
rect 401866 654618 402102 654854
rect 401546 618938 401782 619174
rect 401866 618938 402102 619174
rect 401546 618618 401782 618854
rect 401866 618618 402102 618854
rect 401546 582938 401782 583174
rect 401866 582938 402102 583174
rect 401546 582618 401782 582854
rect 401866 582618 402102 582854
rect 401546 546938 401782 547174
rect 401866 546938 402102 547174
rect 401546 546618 401782 546854
rect 401866 546618 402102 546854
rect 401546 510938 401782 511174
rect 401866 510938 402102 511174
rect 401546 510618 401782 510854
rect 401866 510618 402102 510854
rect 401546 474938 401782 475174
rect 401866 474938 402102 475174
rect 401546 474618 401782 474854
rect 401866 474618 402102 474854
rect 401546 438938 401782 439174
rect 401866 438938 402102 439174
rect 401546 438618 401782 438854
rect 401866 438618 402102 438854
rect 401546 402938 401782 403174
rect 401866 402938 402102 403174
rect 401546 402618 401782 402854
rect 401866 402618 402102 402854
rect 401546 366938 401782 367174
rect 401866 366938 402102 367174
rect 401546 366618 401782 366854
rect 401866 366618 402102 366854
rect 401546 330938 401782 331174
rect 401866 330938 402102 331174
rect 401546 330618 401782 330854
rect 401866 330618 402102 330854
rect 401546 294938 401782 295174
rect 401866 294938 402102 295174
rect 401546 294618 401782 294854
rect 401866 294618 402102 294854
rect 401546 258938 401782 259174
rect 401866 258938 402102 259174
rect 401546 258618 401782 258854
rect 401866 258618 402102 258854
rect 401546 222938 401782 223174
rect 401866 222938 402102 223174
rect 401546 222618 401782 222854
rect 401866 222618 402102 222854
rect 401546 186938 401782 187174
rect 401866 186938 402102 187174
rect 401546 186618 401782 186854
rect 401866 186618 402102 186854
rect 401546 150938 401782 151174
rect 401866 150938 402102 151174
rect 401546 150618 401782 150854
rect 401866 150618 402102 150854
rect 401546 114938 401782 115174
rect 401866 114938 402102 115174
rect 401546 114618 401782 114854
rect 401866 114618 402102 114854
rect 401546 78938 401782 79174
rect 401866 78938 402102 79174
rect 401546 78618 401782 78854
rect 401866 78618 402102 78854
rect 401546 42938 401782 43174
rect 401866 42938 402102 43174
rect 401546 42618 401782 42854
rect 401866 42618 402102 42854
rect 401546 6938 401782 7174
rect 401866 6938 402102 7174
rect 401546 6618 401782 6854
rect 401866 6618 402102 6854
rect 401546 -2502 401782 -2266
rect 401866 -2502 402102 -2266
rect 401546 -2822 401782 -2586
rect 401866 -2822 402102 -2586
rect 405266 694658 405502 694894
rect 405586 694658 405822 694894
rect 405266 694338 405502 694574
rect 405586 694338 405822 694574
rect 405266 658658 405502 658894
rect 405586 658658 405822 658894
rect 405266 658338 405502 658574
rect 405586 658338 405822 658574
rect 405266 622658 405502 622894
rect 405586 622658 405822 622894
rect 405266 622338 405502 622574
rect 405586 622338 405822 622574
rect 405266 586658 405502 586894
rect 405586 586658 405822 586894
rect 405266 586338 405502 586574
rect 405586 586338 405822 586574
rect 405266 550658 405502 550894
rect 405586 550658 405822 550894
rect 405266 550338 405502 550574
rect 405586 550338 405822 550574
rect 405266 514658 405502 514894
rect 405586 514658 405822 514894
rect 405266 514338 405502 514574
rect 405586 514338 405822 514574
rect 405266 478658 405502 478894
rect 405586 478658 405822 478894
rect 405266 478338 405502 478574
rect 405586 478338 405822 478574
rect 405266 442658 405502 442894
rect 405586 442658 405822 442894
rect 405266 442338 405502 442574
rect 405586 442338 405822 442574
rect 405266 406658 405502 406894
rect 405586 406658 405822 406894
rect 405266 406338 405502 406574
rect 405586 406338 405822 406574
rect 405266 370658 405502 370894
rect 405586 370658 405822 370894
rect 405266 370338 405502 370574
rect 405586 370338 405822 370574
rect 405266 334658 405502 334894
rect 405586 334658 405822 334894
rect 405266 334338 405502 334574
rect 405586 334338 405822 334574
rect 405266 298658 405502 298894
rect 405586 298658 405822 298894
rect 405266 298338 405502 298574
rect 405586 298338 405822 298574
rect 405266 262658 405502 262894
rect 405586 262658 405822 262894
rect 405266 262338 405502 262574
rect 405586 262338 405822 262574
rect 405266 226658 405502 226894
rect 405586 226658 405822 226894
rect 405266 226338 405502 226574
rect 405586 226338 405822 226574
rect 405266 190658 405502 190894
rect 405586 190658 405822 190894
rect 405266 190338 405502 190574
rect 405586 190338 405822 190574
rect 405266 154658 405502 154894
rect 405586 154658 405822 154894
rect 405266 154338 405502 154574
rect 405586 154338 405822 154574
rect 405266 118658 405502 118894
rect 405586 118658 405822 118894
rect 405266 118338 405502 118574
rect 405586 118338 405822 118574
rect 405266 82658 405502 82894
rect 405586 82658 405822 82894
rect 405266 82338 405502 82574
rect 405586 82338 405822 82574
rect 405266 46658 405502 46894
rect 405586 46658 405822 46894
rect 405266 46338 405502 46574
rect 405586 46338 405822 46574
rect 405266 10658 405502 10894
rect 405586 10658 405822 10894
rect 405266 10338 405502 10574
rect 405586 10338 405822 10574
rect 405266 -4422 405502 -4186
rect 405586 -4422 405822 -4186
rect 405266 -4742 405502 -4506
rect 405586 -4742 405822 -4506
rect 426986 711322 427222 711558
rect 427306 711322 427542 711558
rect 426986 711002 427222 711238
rect 427306 711002 427542 711238
rect 423266 709402 423502 709638
rect 423586 709402 423822 709638
rect 423266 709082 423502 709318
rect 423586 709082 423822 709318
rect 419546 707482 419782 707718
rect 419866 707482 420102 707718
rect 419546 707162 419782 707398
rect 419866 707162 420102 707398
rect 408986 698378 409222 698614
rect 409306 698378 409542 698614
rect 408986 698058 409222 698294
rect 409306 698058 409542 698294
rect 408986 662378 409222 662614
rect 409306 662378 409542 662614
rect 408986 662058 409222 662294
rect 409306 662058 409542 662294
rect 408986 626378 409222 626614
rect 409306 626378 409542 626614
rect 408986 626058 409222 626294
rect 409306 626058 409542 626294
rect 408986 590378 409222 590614
rect 409306 590378 409542 590614
rect 408986 590058 409222 590294
rect 409306 590058 409542 590294
rect 408986 554378 409222 554614
rect 409306 554378 409542 554614
rect 408986 554058 409222 554294
rect 409306 554058 409542 554294
rect 408986 518378 409222 518614
rect 409306 518378 409542 518614
rect 408986 518058 409222 518294
rect 409306 518058 409542 518294
rect 408986 482378 409222 482614
rect 409306 482378 409542 482614
rect 408986 482058 409222 482294
rect 409306 482058 409542 482294
rect 408986 446378 409222 446614
rect 409306 446378 409542 446614
rect 408986 446058 409222 446294
rect 409306 446058 409542 446294
rect 408986 410378 409222 410614
rect 409306 410378 409542 410614
rect 408986 410058 409222 410294
rect 409306 410058 409542 410294
rect 408986 374378 409222 374614
rect 409306 374378 409542 374614
rect 408986 374058 409222 374294
rect 409306 374058 409542 374294
rect 408986 338378 409222 338614
rect 409306 338378 409542 338614
rect 408986 338058 409222 338294
rect 409306 338058 409542 338294
rect 408986 302378 409222 302614
rect 409306 302378 409542 302614
rect 408986 302058 409222 302294
rect 409306 302058 409542 302294
rect 408986 266378 409222 266614
rect 409306 266378 409542 266614
rect 408986 266058 409222 266294
rect 409306 266058 409542 266294
rect 408986 230378 409222 230614
rect 409306 230378 409542 230614
rect 408986 230058 409222 230294
rect 409306 230058 409542 230294
rect 408986 194378 409222 194614
rect 409306 194378 409542 194614
rect 408986 194058 409222 194294
rect 409306 194058 409542 194294
rect 408986 158378 409222 158614
rect 409306 158378 409542 158614
rect 408986 158058 409222 158294
rect 409306 158058 409542 158294
rect 408986 122378 409222 122614
rect 409306 122378 409542 122614
rect 408986 122058 409222 122294
rect 409306 122058 409542 122294
rect 408986 86378 409222 86614
rect 409306 86378 409542 86614
rect 408986 86058 409222 86294
rect 409306 86058 409542 86294
rect 408986 50378 409222 50614
rect 409306 50378 409542 50614
rect 408986 50058 409222 50294
rect 409306 50058 409542 50294
rect 408986 14378 409222 14614
rect 409306 14378 409542 14614
rect 408986 14058 409222 14294
rect 409306 14058 409542 14294
rect 390986 -7302 391222 -7066
rect 391306 -7302 391542 -7066
rect 390986 -7622 391222 -7386
rect 391306 -7622 391542 -7386
rect 415826 705562 416062 705798
rect 416146 705562 416382 705798
rect 415826 705242 416062 705478
rect 416146 705242 416382 705478
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 415826 633218 416062 633454
rect 416146 633218 416382 633454
rect 415826 632898 416062 633134
rect 416146 632898 416382 633134
rect 415826 597218 416062 597454
rect 416146 597218 416382 597454
rect 415826 596898 416062 597134
rect 416146 596898 416382 597134
rect 415826 561218 416062 561454
rect 416146 561218 416382 561454
rect 415826 560898 416062 561134
rect 416146 560898 416382 561134
rect 415826 525218 416062 525454
rect 416146 525218 416382 525454
rect 415826 524898 416062 525134
rect 416146 524898 416382 525134
rect 415826 489218 416062 489454
rect 416146 489218 416382 489454
rect 415826 488898 416062 489134
rect 416146 488898 416382 489134
rect 415826 453218 416062 453454
rect 416146 453218 416382 453454
rect 415826 452898 416062 453134
rect 416146 452898 416382 453134
rect 415826 417218 416062 417454
rect 416146 417218 416382 417454
rect 415826 416898 416062 417134
rect 416146 416898 416382 417134
rect 415826 381218 416062 381454
rect 416146 381218 416382 381454
rect 415826 380898 416062 381134
rect 416146 380898 416382 381134
rect 415826 345218 416062 345454
rect 416146 345218 416382 345454
rect 415826 344898 416062 345134
rect 416146 344898 416382 345134
rect 415826 309218 416062 309454
rect 416146 309218 416382 309454
rect 415826 308898 416062 309134
rect 416146 308898 416382 309134
rect 415826 273218 416062 273454
rect 416146 273218 416382 273454
rect 415826 272898 416062 273134
rect 416146 272898 416382 273134
rect 415826 237218 416062 237454
rect 416146 237218 416382 237454
rect 415826 236898 416062 237134
rect 416146 236898 416382 237134
rect 415826 201218 416062 201454
rect 416146 201218 416382 201454
rect 415826 200898 416062 201134
rect 416146 200898 416382 201134
rect 415826 165218 416062 165454
rect 416146 165218 416382 165454
rect 415826 164898 416062 165134
rect 416146 164898 416382 165134
rect 415826 129218 416062 129454
rect 416146 129218 416382 129454
rect 415826 128898 416062 129134
rect 416146 128898 416382 129134
rect 415826 93218 416062 93454
rect 416146 93218 416382 93454
rect 415826 92898 416062 93134
rect 416146 92898 416382 93134
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -1542 416062 -1306
rect 416146 -1542 416382 -1306
rect 415826 -1862 416062 -1626
rect 416146 -1862 416382 -1626
rect 419546 672938 419782 673174
rect 419866 672938 420102 673174
rect 419546 672618 419782 672854
rect 419866 672618 420102 672854
rect 419546 636938 419782 637174
rect 419866 636938 420102 637174
rect 419546 636618 419782 636854
rect 419866 636618 420102 636854
rect 419546 600938 419782 601174
rect 419866 600938 420102 601174
rect 419546 600618 419782 600854
rect 419866 600618 420102 600854
rect 419546 564938 419782 565174
rect 419866 564938 420102 565174
rect 419546 564618 419782 564854
rect 419866 564618 420102 564854
rect 419546 528938 419782 529174
rect 419866 528938 420102 529174
rect 419546 528618 419782 528854
rect 419866 528618 420102 528854
rect 419546 492938 419782 493174
rect 419866 492938 420102 493174
rect 419546 492618 419782 492854
rect 419866 492618 420102 492854
rect 419546 456938 419782 457174
rect 419866 456938 420102 457174
rect 419546 456618 419782 456854
rect 419866 456618 420102 456854
rect 419546 420938 419782 421174
rect 419866 420938 420102 421174
rect 419546 420618 419782 420854
rect 419866 420618 420102 420854
rect 419546 384938 419782 385174
rect 419866 384938 420102 385174
rect 419546 384618 419782 384854
rect 419866 384618 420102 384854
rect 419546 348938 419782 349174
rect 419866 348938 420102 349174
rect 419546 348618 419782 348854
rect 419866 348618 420102 348854
rect 419546 312938 419782 313174
rect 419866 312938 420102 313174
rect 419546 312618 419782 312854
rect 419866 312618 420102 312854
rect 419546 276938 419782 277174
rect 419866 276938 420102 277174
rect 419546 276618 419782 276854
rect 419866 276618 420102 276854
rect 419546 240938 419782 241174
rect 419866 240938 420102 241174
rect 419546 240618 419782 240854
rect 419866 240618 420102 240854
rect 419546 204938 419782 205174
rect 419866 204938 420102 205174
rect 419546 204618 419782 204854
rect 419866 204618 420102 204854
rect 419546 168938 419782 169174
rect 419866 168938 420102 169174
rect 419546 168618 419782 168854
rect 419866 168618 420102 168854
rect 419546 132938 419782 133174
rect 419866 132938 420102 133174
rect 419546 132618 419782 132854
rect 419866 132618 420102 132854
rect 419546 96938 419782 97174
rect 419866 96938 420102 97174
rect 419546 96618 419782 96854
rect 419866 96618 420102 96854
rect 419546 60938 419782 61174
rect 419866 60938 420102 61174
rect 419546 60618 419782 60854
rect 419866 60618 420102 60854
rect 419546 24938 419782 25174
rect 419866 24938 420102 25174
rect 419546 24618 419782 24854
rect 419866 24618 420102 24854
rect 419546 -3462 419782 -3226
rect 419866 -3462 420102 -3226
rect 419546 -3782 419782 -3546
rect 419866 -3782 420102 -3546
rect 423266 676658 423502 676894
rect 423586 676658 423822 676894
rect 423266 676338 423502 676574
rect 423586 676338 423822 676574
rect 423266 640658 423502 640894
rect 423586 640658 423822 640894
rect 423266 640338 423502 640574
rect 423586 640338 423822 640574
rect 423266 604658 423502 604894
rect 423586 604658 423822 604894
rect 423266 604338 423502 604574
rect 423586 604338 423822 604574
rect 423266 568658 423502 568894
rect 423586 568658 423822 568894
rect 423266 568338 423502 568574
rect 423586 568338 423822 568574
rect 423266 532658 423502 532894
rect 423586 532658 423822 532894
rect 423266 532338 423502 532574
rect 423586 532338 423822 532574
rect 423266 496658 423502 496894
rect 423586 496658 423822 496894
rect 423266 496338 423502 496574
rect 423586 496338 423822 496574
rect 423266 460658 423502 460894
rect 423586 460658 423822 460894
rect 423266 460338 423502 460574
rect 423586 460338 423822 460574
rect 423266 424658 423502 424894
rect 423586 424658 423822 424894
rect 423266 424338 423502 424574
rect 423586 424338 423822 424574
rect 423266 388658 423502 388894
rect 423586 388658 423822 388894
rect 423266 388338 423502 388574
rect 423586 388338 423822 388574
rect 423266 352658 423502 352894
rect 423586 352658 423822 352894
rect 423266 352338 423502 352574
rect 423586 352338 423822 352574
rect 423266 316658 423502 316894
rect 423586 316658 423822 316894
rect 423266 316338 423502 316574
rect 423586 316338 423822 316574
rect 423266 280658 423502 280894
rect 423586 280658 423822 280894
rect 423266 280338 423502 280574
rect 423586 280338 423822 280574
rect 423266 244658 423502 244894
rect 423586 244658 423822 244894
rect 423266 244338 423502 244574
rect 423586 244338 423822 244574
rect 423266 208658 423502 208894
rect 423586 208658 423822 208894
rect 423266 208338 423502 208574
rect 423586 208338 423822 208574
rect 423266 172658 423502 172894
rect 423586 172658 423822 172894
rect 423266 172338 423502 172574
rect 423586 172338 423822 172574
rect 423266 136658 423502 136894
rect 423586 136658 423822 136894
rect 423266 136338 423502 136574
rect 423586 136338 423822 136574
rect 423266 100658 423502 100894
rect 423586 100658 423822 100894
rect 423266 100338 423502 100574
rect 423586 100338 423822 100574
rect 423266 64658 423502 64894
rect 423586 64658 423822 64894
rect 423266 64338 423502 64574
rect 423586 64338 423822 64574
rect 423266 28658 423502 28894
rect 423586 28658 423822 28894
rect 423266 28338 423502 28574
rect 423586 28338 423822 28574
rect 423266 -5382 423502 -5146
rect 423586 -5382 423822 -5146
rect 423266 -5702 423502 -5466
rect 423586 -5702 423822 -5466
rect 444986 710362 445222 710598
rect 445306 710362 445542 710598
rect 444986 710042 445222 710278
rect 445306 710042 445542 710278
rect 441266 708442 441502 708678
rect 441586 708442 441822 708678
rect 441266 708122 441502 708358
rect 441586 708122 441822 708358
rect 437546 706522 437782 706758
rect 437866 706522 438102 706758
rect 437546 706202 437782 706438
rect 437866 706202 438102 706438
rect 426986 680378 427222 680614
rect 427306 680378 427542 680614
rect 426986 680058 427222 680294
rect 427306 680058 427542 680294
rect 426986 644378 427222 644614
rect 427306 644378 427542 644614
rect 426986 644058 427222 644294
rect 427306 644058 427542 644294
rect 426986 608378 427222 608614
rect 427306 608378 427542 608614
rect 426986 608058 427222 608294
rect 427306 608058 427542 608294
rect 426986 572378 427222 572614
rect 427306 572378 427542 572614
rect 426986 572058 427222 572294
rect 427306 572058 427542 572294
rect 426986 536378 427222 536614
rect 427306 536378 427542 536614
rect 426986 536058 427222 536294
rect 427306 536058 427542 536294
rect 426986 500378 427222 500614
rect 427306 500378 427542 500614
rect 426986 500058 427222 500294
rect 427306 500058 427542 500294
rect 426986 464378 427222 464614
rect 427306 464378 427542 464614
rect 426986 464058 427222 464294
rect 427306 464058 427542 464294
rect 426986 428378 427222 428614
rect 427306 428378 427542 428614
rect 426986 428058 427222 428294
rect 427306 428058 427542 428294
rect 426986 392378 427222 392614
rect 427306 392378 427542 392614
rect 426986 392058 427222 392294
rect 427306 392058 427542 392294
rect 426986 356378 427222 356614
rect 427306 356378 427542 356614
rect 426986 356058 427222 356294
rect 427306 356058 427542 356294
rect 426986 320378 427222 320614
rect 427306 320378 427542 320614
rect 426986 320058 427222 320294
rect 427306 320058 427542 320294
rect 426986 284378 427222 284614
rect 427306 284378 427542 284614
rect 426986 284058 427222 284294
rect 427306 284058 427542 284294
rect 426986 248378 427222 248614
rect 427306 248378 427542 248614
rect 426986 248058 427222 248294
rect 427306 248058 427542 248294
rect 426986 212378 427222 212614
rect 427306 212378 427542 212614
rect 426986 212058 427222 212294
rect 427306 212058 427542 212294
rect 426986 176378 427222 176614
rect 427306 176378 427542 176614
rect 426986 176058 427222 176294
rect 427306 176058 427542 176294
rect 426986 140378 427222 140614
rect 427306 140378 427542 140614
rect 426986 140058 427222 140294
rect 427306 140058 427542 140294
rect 426986 104378 427222 104614
rect 427306 104378 427542 104614
rect 426986 104058 427222 104294
rect 427306 104058 427542 104294
rect 426986 68378 427222 68614
rect 427306 68378 427542 68614
rect 426986 68058 427222 68294
rect 427306 68058 427542 68294
rect 426986 32378 427222 32614
rect 427306 32378 427542 32614
rect 426986 32058 427222 32294
rect 427306 32058 427542 32294
rect 408986 -6342 409222 -6106
rect 409306 -6342 409542 -6106
rect 408986 -6662 409222 -6426
rect 409306 -6662 409542 -6426
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 433826 435218 434062 435454
rect 434146 435218 434382 435454
rect 433826 434898 434062 435134
rect 434146 434898 434382 435134
rect 433826 399218 434062 399454
rect 434146 399218 434382 399454
rect 433826 398898 434062 399134
rect 434146 398898 434382 399134
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 433826 291218 434062 291454
rect 434146 291218 434382 291454
rect 433826 290898 434062 291134
rect 434146 290898 434382 291134
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 433826 219218 434062 219454
rect 434146 219218 434382 219454
rect 433826 218898 434062 219134
rect 434146 218898 434382 219134
rect 433826 183218 434062 183454
rect 434146 183218 434382 183454
rect 433826 182898 434062 183134
rect 434146 182898 434382 183134
rect 433826 147218 434062 147454
rect 434146 147218 434382 147454
rect 433826 146898 434062 147134
rect 434146 146898 434382 147134
rect 433826 111218 434062 111454
rect 434146 111218 434382 111454
rect 433826 110898 434062 111134
rect 434146 110898 434382 111134
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 437546 690938 437782 691174
rect 437866 690938 438102 691174
rect 437546 690618 437782 690854
rect 437866 690618 438102 690854
rect 437546 654938 437782 655174
rect 437866 654938 438102 655174
rect 437546 654618 437782 654854
rect 437866 654618 438102 654854
rect 437546 618938 437782 619174
rect 437866 618938 438102 619174
rect 437546 618618 437782 618854
rect 437866 618618 438102 618854
rect 437546 582938 437782 583174
rect 437866 582938 438102 583174
rect 437546 582618 437782 582854
rect 437866 582618 438102 582854
rect 437546 546938 437782 547174
rect 437866 546938 438102 547174
rect 437546 546618 437782 546854
rect 437866 546618 438102 546854
rect 437546 510938 437782 511174
rect 437866 510938 438102 511174
rect 437546 510618 437782 510854
rect 437866 510618 438102 510854
rect 437546 474938 437782 475174
rect 437866 474938 438102 475174
rect 437546 474618 437782 474854
rect 437866 474618 438102 474854
rect 437546 438938 437782 439174
rect 437866 438938 438102 439174
rect 437546 438618 437782 438854
rect 437866 438618 438102 438854
rect 437546 402938 437782 403174
rect 437866 402938 438102 403174
rect 437546 402618 437782 402854
rect 437866 402618 438102 402854
rect 437546 366938 437782 367174
rect 437866 366938 438102 367174
rect 437546 366618 437782 366854
rect 437866 366618 438102 366854
rect 437546 330938 437782 331174
rect 437866 330938 438102 331174
rect 437546 330618 437782 330854
rect 437866 330618 438102 330854
rect 437546 294938 437782 295174
rect 437866 294938 438102 295174
rect 437546 294618 437782 294854
rect 437866 294618 438102 294854
rect 437546 258938 437782 259174
rect 437866 258938 438102 259174
rect 437546 258618 437782 258854
rect 437866 258618 438102 258854
rect 437546 222938 437782 223174
rect 437866 222938 438102 223174
rect 437546 222618 437782 222854
rect 437866 222618 438102 222854
rect 437546 186938 437782 187174
rect 437866 186938 438102 187174
rect 437546 186618 437782 186854
rect 437866 186618 438102 186854
rect 437546 150938 437782 151174
rect 437866 150938 438102 151174
rect 437546 150618 437782 150854
rect 437866 150618 438102 150854
rect 437546 114938 437782 115174
rect 437866 114938 438102 115174
rect 437546 114618 437782 114854
rect 437866 114618 438102 114854
rect 437546 78938 437782 79174
rect 437866 78938 438102 79174
rect 437546 78618 437782 78854
rect 437866 78618 438102 78854
rect 437546 42938 437782 43174
rect 437866 42938 438102 43174
rect 437546 42618 437782 42854
rect 437866 42618 438102 42854
rect 437546 6938 437782 7174
rect 437866 6938 438102 7174
rect 437546 6618 437782 6854
rect 437866 6618 438102 6854
rect 437546 -2502 437782 -2266
rect 437866 -2502 438102 -2266
rect 437546 -2822 437782 -2586
rect 437866 -2822 438102 -2586
rect 441266 694658 441502 694894
rect 441586 694658 441822 694894
rect 441266 694338 441502 694574
rect 441586 694338 441822 694574
rect 441266 658658 441502 658894
rect 441586 658658 441822 658894
rect 441266 658338 441502 658574
rect 441586 658338 441822 658574
rect 441266 622658 441502 622894
rect 441586 622658 441822 622894
rect 441266 622338 441502 622574
rect 441586 622338 441822 622574
rect 441266 586658 441502 586894
rect 441586 586658 441822 586894
rect 441266 586338 441502 586574
rect 441586 586338 441822 586574
rect 441266 550658 441502 550894
rect 441586 550658 441822 550894
rect 441266 550338 441502 550574
rect 441586 550338 441822 550574
rect 441266 514658 441502 514894
rect 441586 514658 441822 514894
rect 441266 514338 441502 514574
rect 441586 514338 441822 514574
rect 441266 478658 441502 478894
rect 441586 478658 441822 478894
rect 441266 478338 441502 478574
rect 441586 478338 441822 478574
rect 441266 442658 441502 442894
rect 441586 442658 441822 442894
rect 441266 442338 441502 442574
rect 441586 442338 441822 442574
rect 441266 406658 441502 406894
rect 441586 406658 441822 406894
rect 441266 406338 441502 406574
rect 441586 406338 441822 406574
rect 441266 370658 441502 370894
rect 441586 370658 441822 370894
rect 441266 370338 441502 370574
rect 441586 370338 441822 370574
rect 441266 334658 441502 334894
rect 441586 334658 441822 334894
rect 441266 334338 441502 334574
rect 441586 334338 441822 334574
rect 441266 298658 441502 298894
rect 441586 298658 441822 298894
rect 441266 298338 441502 298574
rect 441586 298338 441822 298574
rect 441266 262658 441502 262894
rect 441586 262658 441822 262894
rect 441266 262338 441502 262574
rect 441586 262338 441822 262574
rect 441266 226658 441502 226894
rect 441586 226658 441822 226894
rect 441266 226338 441502 226574
rect 441586 226338 441822 226574
rect 441266 190658 441502 190894
rect 441586 190658 441822 190894
rect 441266 190338 441502 190574
rect 441586 190338 441822 190574
rect 441266 154658 441502 154894
rect 441586 154658 441822 154894
rect 441266 154338 441502 154574
rect 441586 154338 441822 154574
rect 441266 118658 441502 118894
rect 441586 118658 441822 118894
rect 441266 118338 441502 118574
rect 441586 118338 441822 118574
rect 441266 82658 441502 82894
rect 441586 82658 441822 82894
rect 441266 82338 441502 82574
rect 441586 82338 441822 82574
rect 441266 46658 441502 46894
rect 441586 46658 441822 46894
rect 441266 46338 441502 46574
rect 441586 46338 441822 46574
rect 441266 10658 441502 10894
rect 441586 10658 441822 10894
rect 441266 10338 441502 10574
rect 441586 10338 441822 10574
rect 441266 -4422 441502 -4186
rect 441586 -4422 441822 -4186
rect 441266 -4742 441502 -4506
rect 441586 -4742 441822 -4506
rect 462986 711322 463222 711558
rect 463306 711322 463542 711558
rect 462986 711002 463222 711238
rect 463306 711002 463542 711238
rect 459266 709402 459502 709638
rect 459586 709402 459822 709638
rect 459266 709082 459502 709318
rect 459586 709082 459822 709318
rect 455546 707482 455782 707718
rect 455866 707482 456102 707718
rect 455546 707162 455782 707398
rect 455866 707162 456102 707398
rect 444986 698378 445222 698614
rect 445306 698378 445542 698614
rect 444986 698058 445222 698294
rect 445306 698058 445542 698294
rect 444986 662378 445222 662614
rect 445306 662378 445542 662614
rect 444986 662058 445222 662294
rect 445306 662058 445542 662294
rect 444986 626378 445222 626614
rect 445306 626378 445542 626614
rect 444986 626058 445222 626294
rect 445306 626058 445542 626294
rect 444986 590378 445222 590614
rect 445306 590378 445542 590614
rect 444986 590058 445222 590294
rect 445306 590058 445542 590294
rect 444986 554378 445222 554614
rect 445306 554378 445542 554614
rect 444986 554058 445222 554294
rect 445306 554058 445542 554294
rect 444986 518378 445222 518614
rect 445306 518378 445542 518614
rect 444986 518058 445222 518294
rect 445306 518058 445542 518294
rect 444986 482378 445222 482614
rect 445306 482378 445542 482614
rect 444986 482058 445222 482294
rect 445306 482058 445542 482294
rect 444986 446378 445222 446614
rect 445306 446378 445542 446614
rect 444986 446058 445222 446294
rect 445306 446058 445542 446294
rect 444986 410378 445222 410614
rect 445306 410378 445542 410614
rect 444986 410058 445222 410294
rect 445306 410058 445542 410294
rect 444986 374378 445222 374614
rect 445306 374378 445542 374614
rect 444986 374058 445222 374294
rect 445306 374058 445542 374294
rect 444986 338378 445222 338614
rect 445306 338378 445542 338614
rect 444986 338058 445222 338294
rect 445306 338058 445542 338294
rect 444986 302378 445222 302614
rect 445306 302378 445542 302614
rect 444986 302058 445222 302294
rect 445306 302058 445542 302294
rect 444986 266378 445222 266614
rect 445306 266378 445542 266614
rect 444986 266058 445222 266294
rect 445306 266058 445542 266294
rect 444986 230378 445222 230614
rect 445306 230378 445542 230614
rect 444986 230058 445222 230294
rect 445306 230058 445542 230294
rect 444986 194378 445222 194614
rect 445306 194378 445542 194614
rect 444986 194058 445222 194294
rect 445306 194058 445542 194294
rect 444986 158378 445222 158614
rect 445306 158378 445542 158614
rect 444986 158058 445222 158294
rect 445306 158058 445542 158294
rect 444986 122378 445222 122614
rect 445306 122378 445542 122614
rect 444986 122058 445222 122294
rect 445306 122058 445542 122294
rect 444986 86378 445222 86614
rect 445306 86378 445542 86614
rect 444986 86058 445222 86294
rect 445306 86058 445542 86294
rect 444986 50378 445222 50614
rect 445306 50378 445542 50614
rect 444986 50058 445222 50294
rect 445306 50058 445542 50294
rect 444986 14378 445222 14614
rect 445306 14378 445542 14614
rect 444986 14058 445222 14294
rect 445306 14058 445542 14294
rect 426986 -7302 427222 -7066
rect 427306 -7302 427542 -7066
rect 426986 -7622 427222 -7386
rect 427306 -7622 427542 -7386
rect 451826 705562 452062 705798
rect 452146 705562 452382 705798
rect 451826 705242 452062 705478
rect 452146 705242 452382 705478
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 451826 561218 452062 561454
rect 452146 561218 452382 561454
rect 451826 560898 452062 561134
rect 452146 560898 452382 561134
rect 451826 525218 452062 525454
rect 452146 525218 452382 525454
rect 451826 524898 452062 525134
rect 452146 524898 452382 525134
rect 451826 489218 452062 489454
rect 452146 489218 452382 489454
rect 451826 488898 452062 489134
rect 452146 488898 452382 489134
rect 451826 453218 452062 453454
rect 452146 453218 452382 453454
rect 451826 452898 452062 453134
rect 452146 452898 452382 453134
rect 451826 417218 452062 417454
rect 452146 417218 452382 417454
rect 451826 416898 452062 417134
rect 452146 416898 452382 417134
rect 451826 381218 452062 381454
rect 452146 381218 452382 381454
rect 451826 380898 452062 381134
rect 452146 380898 452382 381134
rect 451826 345218 452062 345454
rect 452146 345218 452382 345454
rect 451826 344898 452062 345134
rect 452146 344898 452382 345134
rect 451826 309218 452062 309454
rect 452146 309218 452382 309454
rect 451826 308898 452062 309134
rect 452146 308898 452382 309134
rect 451826 273218 452062 273454
rect 452146 273218 452382 273454
rect 451826 272898 452062 273134
rect 452146 272898 452382 273134
rect 451826 237218 452062 237454
rect 452146 237218 452382 237454
rect 451826 236898 452062 237134
rect 452146 236898 452382 237134
rect 451826 201218 452062 201454
rect 452146 201218 452382 201454
rect 451826 200898 452062 201134
rect 452146 200898 452382 201134
rect 451826 165218 452062 165454
rect 452146 165218 452382 165454
rect 451826 164898 452062 165134
rect 452146 164898 452382 165134
rect 451826 129218 452062 129454
rect 452146 129218 452382 129454
rect 451826 128898 452062 129134
rect 452146 128898 452382 129134
rect 451826 93218 452062 93454
rect 452146 93218 452382 93454
rect 451826 92898 452062 93134
rect 452146 92898 452382 93134
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -1542 452062 -1306
rect 452146 -1542 452382 -1306
rect 451826 -1862 452062 -1626
rect 452146 -1862 452382 -1626
rect 455546 672938 455782 673174
rect 455866 672938 456102 673174
rect 455546 672618 455782 672854
rect 455866 672618 456102 672854
rect 455546 636938 455782 637174
rect 455866 636938 456102 637174
rect 455546 636618 455782 636854
rect 455866 636618 456102 636854
rect 455546 600938 455782 601174
rect 455866 600938 456102 601174
rect 455546 600618 455782 600854
rect 455866 600618 456102 600854
rect 455546 564938 455782 565174
rect 455866 564938 456102 565174
rect 455546 564618 455782 564854
rect 455866 564618 456102 564854
rect 455546 528938 455782 529174
rect 455866 528938 456102 529174
rect 455546 528618 455782 528854
rect 455866 528618 456102 528854
rect 455546 492938 455782 493174
rect 455866 492938 456102 493174
rect 455546 492618 455782 492854
rect 455866 492618 456102 492854
rect 455546 456938 455782 457174
rect 455866 456938 456102 457174
rect 455546 456618 455782 456854
rect 455866 456618 456102 456854
rect 455546 420938 455782 421174
rect 455866 420938 456102 421174
rect 455546 420618 455782 420854
rect 455866 420618 456102 420854
rect 455546 384938 455782 385174
rect 455866 384938 456102 385174
rect 455546 384618 455782 384854
rect 455866 384618 456102 384854
rect 455546 348938 455782 349174
rect 455866 348938 456102 349174
rect 455546 348618 455782 348854
rect 455866 348618 456102 348854
rect 455546 312938 455782 313174
rect 455866 312938 456102 313174
rect 455546 312618 455782 312854
rect 455866 312618 456102 312854
rect 455546 276938 455782 277174
rect 455866 276938 456102 277174
rect 455546 276618 455782 276854
rect 455866 276618 456102 276854
rect 455546 240938 455782 241174
rect 455866 240938 456102 241174
rect 455546 240618 455782 240854
rect 455866 240618 456102 240854
rect 455546 204938 455782 205174
rect 455866 204938 456102 205174
rect 455546 204618 455782 204854
rect 455866 204618 456102 204854
rect 455546 168938 455782 169174
rect 455866 168938 456102 169174
rect 455546 168618 455782 168854
rect 455866 168618 456102 168854
rect 455546 132938 455782 133174
rect 455866 132938 456102 133174
rect 455546 132618 455782 132854
rect 455866 132618 456102 132854
rect 455546 96938 455782 97174
rect 455866 96938 456102 97174
rect 455546 96618 455782 96854
rect 455866 96618 456102 96854
rect 455546 60938 455782 61174
rect 455866 60938 456102 61174
rect 455546 60618 455782 60854
rect 455866 60618 456102 60854
rect 455546 24938 455782 25174
rect 455866 24938 456102 25174
rect 455546 24618 455782 24854
rect 455866 24618 456102 24854
rect 455546 -3462 455782 -3226
rect 455866 -3462 456102 -3226
rect 455546 -3782 455782 -3546
rect 455866 -3782 456102 -3546
rect 459266 676658 459502 676894
rect 459586 676658 459822 676894
rect 459266 676338 459502 676574
rect 459586 676338 459822 676574
rect 459266 640658 459502 640894
rect 459586 640658 459822 640894
rect 459266 640338 459502 640574
rect 459586 640338 459822 640574
rect 459266 604658 459502 604894
rect 459586 604658 459822 604894
rect 459266 604338 459502 604574
rect 459586 604338 459822 604574
rect 459266 568658 459502 568894
rect 459586 568658 459822 568894
rect 459266 568338 459502 568574
rect 459586 568338 459822 568574
rect 459266 532658 459502 532894
rect 459586 532658 459822 532894
rect 459266 532338 459502 532574
rect 459586 532338 459822 532574
rect 459266 496658 459502 496894
rect 459586 496658 459822 496894
rect 459266 496338 459502 496574
rect 459586 496338 459822 496574
rect 459266 460658 459502 460894
rect 459586 460658 459822 460894
rect 459266 460338 459502 460574
rect 459586 460338 459822 460574
rect 459266 424658 459502 424894
rect 459586 424658 459822 424894
rect 459266 424338 459502 424574
rect 459586 424338 459822 424574
rect 459266 388658 459502 388894
rect 459586 388658 459822 388894
rect 459266 388338 459502 388574
rect 459586 388338 459822 388574
rect 459266 352658 459502 352894
rect 459586 352658 459822 352894
rect 459266 352338 459502 352574
rect 459586 352338 459822 352574
rect 459266 316658 459502 316894
rect 459586 316658 459822 316894
rect 459266 316338 459502 316574
rect 459586 316338 459822 316574
rect 459266 280658 459502 280894
rect 459586 280658 459822 280894
rect 459266 280338 459502 280574
rect 459586 280338 459822 280574
rect 459266 244658 459502 244894
rect 459586 244658 459822 244894
rect 459266 244338 459502 244574
rect 459586 244338 459822 244574
rect 459266 208658 459502 208894
rect 459586 208658 459822 208894
rect 459266 208338 459502 208574
rect 459586 208338 459822 208574
rect 459266 172658 459502 172894
rect 459586 172658 459822 172894
rect 459266 172338 459502 172574
rect 459586 172338 459822 172574
rect 459266 136658 459502 136894
rect 459586 136658 459822 136894
rect 459266 136338 459502 136574
rect 459586 136338 459822 136574
rect 459266 100658 459502 100894
rect 459586 100658 459822 100894
rect 459266 100338 459502 100574
rect 459586 100338 459822 100574
rect 459266 64658 459502 64894
rect 459586 64658 459822 64894
rect 459266 64338 459502 64574
rect 459586 64338 459822 64574
rect 459266 28658 459502 28894
rect 459586 28658 459822 28894
rect 459266 28338 459502 28574
rect 459586 28338 459822 28574
rect 459266 -5382 459502 -5146
rect 459586 -5382 459822 -5146
rect 459266 -5702 459502 -5466
rect 459586 -5702 459822 -5466
rect 480986 710362 481222 710598
rect 481306 710362 481542 710598
rect 480986 710042 481222 710278
rect 481306 710042 481542 710278
rect 477266 708442 477502 708678
rect 477586 708442 477822 708678
rect 477266 708122 477502 708358
rect 477586 708122 477822 708358
rect 473546 706522 473782 706758
rect 473866 706522 474102 706758
rect 473546 706202 473782 706438
rect 473866 706202 474102 706438
rect 462986 680378 463222 680614
rect 463306 680378 463542 680614
rect 462986 680058 463222 680294
rect 463306 680058 463542 680294
rect 462986 644378 463222 644614
rect 463306 644378 463542 644614
rect 462986 644058 463222 644294
rect 463306 644058 463542 644294
rect 462986 608378 463222 608614
rect 463306 608378 463542 608614
rect 462986 608058 463222 608294
rect 463306 608058 463542 608294
rect 462986 572378 463222 572614
rect 463306 572378 463542 572614
rect 462986 572058 463222 572294
rect 463306 572058 463542 572294
rect 462986 536378 463222 536614
rect 463306 536378 463542 536614
rect 462986 536058 463222 536294
rect 463306 536058 463542 536294
rect 462986 500378 463222 500614
rect 463306 500378 463542 500614
rect 462986 500058 463222 500294
rect 463306 500058 463542 500294
rect 462986 464378 463222 464614
rect 463306 464378 463542 464614
rect 462986 464058 463222 464294
rect 463306 464058 463542 464294
rect 462986 428378 463222 428614
rect 463306 428378 463542 428614
rect 462986 428058 463222 428294
rect 463306 428058 463542 428294
rect 462986 392378 463222 392614
rect 463306 392378 463542 392614
rect 462986 392058 463222 392294
rect 463306 392058 463542 392294
rect 462986 356378 463222 356614
rect 463306 356378 463542 356614
rect 462986 356058 463222 356294
rect 463306 356058 463542 356294
rect 462986 320378 463222 320614
rect 463306 320378 463542 320614
rect 462986 320058 463222 320294
rect 463306 320058 463542 320294
rect 462986 284378 463222 284614
rect 463306 284378 463542 284614
rect 462986 284058 463222 284294
rect 463306 284058 463542 284294
rect 462986 248378 463222 248614
rect 463306 248378 463542 248614
rect 462986 248058 463222 248294
rect 463306 248058 463542 248294
rect 462986 212378 463222 212614
rect 463306 212378 463542 212614
rect 462986 212058 463222 212294
rect 463306 212058 463542 212294
rect 462986 176378 463222 176614
rect 463306 176378 463542 176614
rect 462986 176058 463222 176294
rect 463306 176058 463542 176294
rect 462986 140378 463222 140614
rect 463306 140378 463542 140614
rect 462986 140058 463222 140294
rect 463306 140058 463542 140294
rect 462986 104378 463222 104614
rect 463306 104378 463542 104614
rect 462986 104058 463222 104294
rect 463306 104058 463542 104294
rect 462986 68378 463222 68614
rect 463306 68378 463542 68614
rect 462986 68058 463222 68294
rect 463306 68058 463542 68294
rect 462986 32378 463222 32614
rect 463306 32378 463542 32614
rect 462986 32058 463222 32294
rect 463306 32058 463542 32294
rect 444986 -6342 445222 -6106
rect 445306 -6342 445542 -6106
rect 444986 -6662 445222 -6426
rect 445306 -6662 445542 -6426
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 469826 327218 470062 327454
rect 470146 327218 470382 327454
rect 469826 326898 470062 327134
rect 470146 326898 470382 327134
rect 469826 291218 470062 291454
rect 470146 291218 470382 291454
rect 469826 290898 470062 291134
rect 470146 290898 470382 291134
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 469826 219218 470062 219454
rect 470146 219218 470382 219454
rect 469826 218898 470062 219134
rect 470146 218898 470382 219134
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 473546 690938 473782 691174
rect 473866 690938 474102 691174
rect 473546 690618 473782 690854
rect 473866 690618 474102 690854
rect 473546 654938 473782 655174
rect 473866 654938 474102 655174
rect 473546 654618 473782 654854
rect 473866 654618 474102 654854
rect 473546 618938 473782 619174
rect 473866 618938 474102 619174
rect 473546 618618 473782 618854
rect 473866 618618 474102 618854
rect 473546 582938 473782 583174
rect 473866 582938 474102 583174
rect 473546 582618 473782 582854
rect 473866 582618 474102 582854
rect 473546 546938 473782 547174
rect 473866 546938 474102 547174
rect 473546 546618 473782 546854
rect 473866 546618 474102 546854
rect 473546 510938 473782 511174
rect 473866 510938 474102 511174
rect 473546 510618 473782 510854
rect 473866 510618 474102 510854
rect 473546 474938 473782 475174
rect 473866 474938 474102 475174
rect 473546 474618 473782 474854
rect 473866 474618 474102 474854
rect 473546 438938 473782 439174
rect 473866 438938 474102 439174
rect 473546 438618 473782 438854
rect 473866 438618 474102 438854
rect 473546 402938 473782 403174
rect 473866 402938 474102 403174
rect 473546 402618 473782 402854
rect 473866 402618 474102 402854
rect 473546 366938 473782 367174
rect 473866 366938 474102 367174
rect 473546 366618 473782 366854
rect 473866 366618 474102 366854
rect 473546 330938 473782 331174
rect 473866 330938 474102 331174
rect 473546 330618 473782 330854
rect 473866 330618 474102 330854
rect 473546 294938 473782 295174
rect 473866 294938 474102 295174
rect 473546 294618 473782 294854
rect 473866 294618 474102 294854
rect 473546 258938 473782 259174
rect 473866 258938 474102 259174
rect 473546 258618 473782 258854
rect 473866 258618 474102 258854
rect 473546 222938 473782 223174
rect 473866 222938 474102 223174
rect 473546 222618 473782 222854
rect 473866 222618 474102 222854
rect 473546 186938 473782 187174
rect 473866 186938 474102 187174
rect 473546 186618 473782 186854
rect 473866 186618 474102 186854
rect 473546 150938 473782 151174
rect 473866 150938 474102 151174
rect 473546 150618 473782 150854
rect 473866 150618 474102 150854
rect 473546 114938 473782 115174
rect 473866 114938 474102 115174
rect 473546 114618 473782 114854
rect 473866 114618 474102 114854
rect 473546 78938 473782 79174
rect 473866 78938 474102 79174
rect 473546 78618 473782 78854
rect 473866 78618 474102 78854
rect 473546 42938 473782 43174
rect 473866 42938 474102 43174
rect 473546 42618 473782 42854
rect 473866 42618 474102 42854
rect 473546 6938 473782 7174
rect 473866 6938 474102 7174
rect 473546 6618 473782 6854
rect 473866 6618 474102 6854
rect 473546 -2502 473782 -2266
rect 473866 -2502 474102 -2266
rect 473546 -2822 473782 -2586
rect 473866 -2822 474102 -2586
rect 477266 694658 477502 694894
rect 477586 694658 477822 694894
rect 477266 694338 477502 694574
rect 477586 694338 477822 694574
rect 477266 658658 477502 658894
rect 477586 658658 477822 658894
rect 477266 658338 477502 658574
rect 477586 658338 477822 658574
rect 477266 622658 477502 622894
rect 477586 622658 477822 622894
rect 477266 622338 477502 622574
rect 477586 622338 477822 622574
rect 477266 586658 477502 586894
rect 477586 586658 477822 586894
rect 477266 586338 477502 586574
rect 477586 586338 477822 586574
rect 477266 550658 477502 550894
rect 477586 550658 477822 550894
rect 477266 550338 477502 550574
rect 477586 550338 477822 550574
rect 477266 514658 477502 514894
rect 477586 514658 477822 514894
rect 477266 514338 477502 514574
rect 477586 514338 477822 514574
rect 477266 478658 477502 478894
rect 477586 478658 477822 478894
rect 477266 478338 477502 478574
rect 477586 478338 477822 478574
rect 477266 442658 477502 442894
rect 477586 442658 477822 442894
rect 477266 442338 477502 442574
rect 477586 442338 477822 442574
rect 477266 406658 477502 406894
rect 477586 406658 477822 406894
rect 477266 406338 477502 406574
rect 477586 406338 477822 406574
rect 477266 370658 477502 370894
rect 477586 370658 477822 370894
rect 477266 370338 477502 370574
rect 477586 370338 477822 370574
rect 477266 334658 477502 334894
rect 477586 334658 477822 334894
rect 477266 334338 477502 334574
rect 477586 334338 477822 334574
rect 477266 298658 477502 298894
rect 477586 298658 477822 298894
rect 477266 298338 477502 298574
rect 477586 298338 477822 298574
rect 477266 262658 477502 262894
rect 477586 262658 477822 262894
rect 477266 262338 477502 262574
rect 477586 262338 477822 262574
rect 477266 226658 477502 226894
rect 477586 226658 477822 226894
rect 477266 226338 477502 226574
rect 477586 226338 477822 226574
rect 477266 190658 477502 190894
rect 477586 190658 477822 190894
rect 477266 190338 477502 190574
rect 477586 190338 477822 190574
rect 477266 154658 477502 154894
rect 477586 154658 477822 154894
rect 477266 154338 477502 154574
rect 477586 154338 477822 154574
rect 477266 118658 477502 118894
rect 477586 118658 477822 118894
rect 477266 118338 477502 118574
rect 477586 118338 477822 118574
rect 477266 82658 477502 82894
rect 477586 82658 477822 82894
rect 477266 82338 477502 82574
rect 477586 82338 477822 82574
rect 477266 46658 477502 46894
rect 477586 46658 477822 46894
rect 477266 46338 477502 46574
rect 477586 46338 477822 46574
rect 477266 10658 477502 10894
rect 477586 10658 477822 10894
rect 477266 10338 477502 10574
rect 477586 10338 477822 10574
rect 477266 -4422 477502 -4186
rect 477586 -4422 477822 -4186
rect 477266 -4742 477502 -4506
rect 477586 -4742 477822 -4506
rect 498986 711322 499222 711558
rect 499306 711322 499542 711558
rect 498986 711002 499222 711238
rect 499306 711002 499542 711238
rect 495266 709402 495502 709638
rect 495586 709402 495822 709638
rect 495266 709082 495502 709318
rect 495586 709082 495822 709318
rect 491546 707482 491782 707718
rect 491866 707482 492102 707718
rect 491546 707162 491782 707398
rect 491866 707162 492102 707398
rect 480986 698378 481222 698614
rect 481306 698378 481542 698614
rect 480986 698058 481222 698294
rect 481306 698058 481542 698294
rect 480986 662378 481222 662614
rect 481306 662378 481542 662614
rect 480986 662058 481222 662294
rect 481306 662058 481542 662294
rect 480986 626378 481222 626614
rect 481306 626378 481542 626614
rect 480986 626058 481222 626294
rect 481306 626058 481542 626294
rect 480986 590378 481222 590614
rect 481306 590378 481542 590614
rect 480986 590058 481222 590294
rect 481306 590058 481542 590294
rect 480986 554378 481222 554614
rect 481306 554378 481542 554614
rect 480986 554058 481222 554294
rect 481306 554058 481542 554294
rect 480986 518378 481222 518614
rect 481306 518378 481542 518614
rect 480986 518058 481222 518294
rect 481306 518058 481542 518294
rect 480986 482378 481222 482614
rect 481306 482378 481542 482614
rect 480986 482058 481222 482294
rect 481306 482058 481542 482294
rect 480986 446378 481222 446614
rect 481306 446378 481542 446614
rect 480986 446058 481222 446294
rect 481306 446058 481542 446294
rect 480986 410378 481222 410614
rect 481306 410378 481542 410614
rect 480986 410058 481222 410294
rect 481306 410058 481542 410294
rect 480986 374378 481222 374614
rect 481306 374378 481542 374614
rect 480986 374058 481222 374294
rect 481306 374058 481542 374294
rect 480986 338378 481222 338614
rect 481306 338378 481542 338614
rect 480986 338058 481222 338294
rect 481306 338058 481542 338294
rect 480986 302378 481222 302614
rect 481306 302378 481542 302614
rect 480986 302058 481222 302294
rect 481306 302058 481542 302294
rect 480986 266378 481222 266614
rect 481306 266378 481542 266614
rect 480986 266058 481222 266294
rect 481306 266058 481542 266294
rect 480986 230378 481222 230614
rect 481306 230378 481542 230614
rect 480986 230058 481222 230294
rect 481306 230058 481542 230294
rect 480986 194378 481222 194614
rect 481306 194378 481542 194614
rect 480986 194058 481222 194294
rect 481306 194058 481542 194294
rect 480986 158378 481222 158614
rect 481306 158378 481542 158614
rect 480986 158058 481222 158294
rect 481306 158058 481542 158294
rect 480986 122378 481222 122614
rect 481306 122378 481542 122614
rect 480986 122058 481222 122294
rect 481306 122058 481542 122294
rect 480986 86378 481222 86614
rect 481306 86378 481542 86614
rect 480986 86058 481222 86294
rect 481306 86058 481542 86294
rect 480986 50378 481222 50614
rect 481306 50378 481542 50614
rect 480986 50058 481222 50294
rect 481306 50058 481542 50294
rect 480986 14378 481222 14614
rect 481306 14378 481542 14614
rect 480986 14058 481222 14294
rect 481306 14058 481542 14294
rect 462986 -7302 463222 -7066
rect 463306 -7302 463542 -7066
rect 462986 -7622 463222 -7386
rect 463306 -7622 463542 -7386
rect 487826 705562 488062 705798
rect 488146 705562 488382 705798
rect 487826 705242 488062 705478
rect 488146 705242 488382 705478
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 487826 633218 488062 633454
rect 488146 633218 488382 633454
rect 487826 632898 488062 633134
rect 488146 632898 488382 633134
rect 487826 597218 488062 597454
rect 488146 597218 488382 597454
rect 487826 596898 488062 597134
rect 488146 596898 488382 597134
rect 487826 561218 488062 561454
rect 488146 561218 488382 561454
rect 487826 560898 488062 561134
rect 488146 560898 488382 561134
rect 487826 525218 488062 525454
rect 488146 525218 488382 525454
rect 487826 524898 488062 525134
rect 488146 524898 488382 525134
rect 487826 489218 488062 489454
rect 488146 489218 488382 489454
rect 487826 488898 488062 489134
rect 488146 488898 488382 489134
rect 487826 453218 488062 453454
rect 488146 453218 488382 453454
rect 487826 452898 488062 453134
rect 488146 452898 488382 453134
rect 487826 417218 488062 417454
rect 488146 417218 488382 417454
rect 487826 416898 488062 417134
rect 488146 416898 488382 417134
rect 487826 381218 488062 381454
rect 488146 381218 488382 381454
rect 487826 380898 488062 381134
rect 488146 380898 488382 381134
rect 487826 345218 488062 345454
rect 488146 345218 488382 345454
rect 487826 344898 488062 345134
rect 488146 344898 488382 345134
rect 487826 309218 488062 309454
rect 488146 309218 488382 309454
rect 487826 308898 488062 309134
rect 488146 308898 488382 309134
rect 487826 273218 488062 273454
rect 488146 273218 488382 273454
rect 487826 272898 488062 273134
rect 488146 272898 488382 273134
rect 487826 237218 488062 237454
rect 488146 237218 488382 237454
rect 487826 236898 488062 237134
rect 488146 236898 488382 237134
rect 487826 201218 488062 201454
rect 488146 201218 488382 201454
rect 487826 200898 488062 201134
rect 488146 200898 488382 201134
rect 487826 165218 488062 165454
rect 488146 165218 488382 165454
rect 487826 164898 488062 165134
rect 488146 164898 488382 165134
rect 487826 129218 488062 129454
rect 488146 129218 488382 129454
rect 487826 128898 488062 129134
rect 488146 128898 488382 129134
rect 487826 93218 488062 93454
rect 488146 93218 488382 93454
rect 487826 92898 488062 93134
rect 488146 92898 488382 93134
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -1542 488062 -1306
rect 488146 -1542 488382 -1306
rect 487826 -1862 488062 -1626
rect 488146 -1862 488382 -1626
rect 491546 672938 491782 673174
rect 491866 672938 492102 673174
rect 491546 672618 491782 672854
rect 491866 672618 492102 672854
rect 491546 636938 491782 637174
rect 491866 636938 492102 637174
rect 491546 636618 491782 636854
rect 491866 636618 492102 636854
rect 491546 600938 491782 601174
rect 491866 600938 492102 601174
rect 491546 600618 491782 600854
rect 491866 600618 492102 600854
rect 491546 564938 491782 565174
rect 491866 564938 492102 565174
rect 491546 564618 491782 564854
rect 491866 564618 492102 564854
rect 491546 528938 491782 529174
rect 491866 528938 492102 529174
rect 491546 528618 491782 528854
rect 491866 528618 492102 528854
rect 491546 492938 491782 493174
rect 491866 492938 492102 493174
rect 491546 492618 491782 492854
rect 491866 492618 492102 492854
rect 491546 456938 491782 457174
rect 491866 456938 492102 457174
rect 491546 456618 491782 456854
rect 491866 456618 492102 456854
rect 491546 420938 491782 421174
rect 491866 420938 492102 421174
rect 491546 420618 491782 420854
rect 491866 420618 492102 420854
rect 491546 384938 491782 385174
rect 491866 384938 492102 385174
rect 491546 384618 491782 384854
rect 491866 384618 492102 384854
rect 491546 348938 491782 349174
rect 491866 348938 492102 349174
rect 491546 348618 491782 348854
rect 491866 348618 492102 348854
rect 491546 312938 491782 313174
rect 491866 312938 492102 313174
rect 491546 312618 491782 312854
rect 491866 312618 492102 312854
rect 491546 276938 491782 277174
rect 491866 276938 492102 277174
rect 491546 276618 491782 276854
rect 491866 276618 492102 276854
rect 491546 240938 491782 241174
rect 491866 240938 492102 241174
rect 491546 240618 491782 240854
rect 491866 240618 492102 240854
rect 491546 204938 491782 205174
rect 491866 204938 492102 205174
rect 491546 204618 491782 204854
rect 491866 204618 492102 204854
rect 491546 168938 491782 169174
rect 491866 168938 492102 169174
rect 491546 168618 491782 168854
rect 491866 168618 492102 168854
rect 491546 132938 491782 133174
rect 491866 132938 492102 133174
rect 491546 132618 491782 132854
rect 491866 132618 492102 132854
rect 491546 96938 491782 97174
rect 491866 96938 492102 97174
rect 491546 96618 491782 96854
rect 491866 96618 492102 96854
rect 491546 60938 491782 61174
rect 491866 60938 492102 61174
rect 491546 60618 491782 60854
rect 491866 60618 492102 60854
rect 491546 24938 491782 25174
rect 491866 24938 492102 25174
rect 491546 24618 491782 24854
rect 491866 24618 492102 24854
rect 491546 -3462 491782 -3226
rect 491866 -3462 492102 -3226
rect 491546 -3782 491782 -3546
rect 491866 -3782 492102 -3546
rect 495266 676658 495502 676894
rect 495586 676658 495822 676894
rect 495266 676338 495502 676574
rect 495586 676338 495822 676574
rect 495266 640658 495502 640894
rect 495586 640658 495822 640894
rect 495266 640338 495502 640574
rect 495586 640338 495822 640574
rect 495266 604658 495502 604894
rect 495586 604658 495822 604894
rect 495266 604338 495502 604574
rect 495586 604338 495822 604574
rect 495266 568658 495502 568894
rect 495586 568658 495822 568894
rect 495266 568338 495502 568574
rect 495586 568338 495822 568574
rect 495266 532658 495502 532894
rect 495586 532658 495822 532894
rect 495266 532338 495502 532574
rect 495586 532338 495822 532574
rect 495266 496658 495502 496894
rect 495586 496658 495822 496894
rect 495266 496338 495502 496574
rect 495586 496338 495822 496574
rect 495266 460658 495502 460894
rect 495586 460658 495822 460894
rect 495266 460338 495502 460574
rect 495586 460338 495822 460574
rect 495266 424658 495502 424894
rect 495586 424658 495822 424894
rect 495266 424338 495502 424574
rect 495586 424338 495822 424574
rect 495266 388658 495502 388894
rect 495586 388658 495822 388894
rect 495266 388338 495502 388574
rect 495586 388338 495822 388574
rect 495266 352658 495502 352894
rect 495586 352658 495822 352894
rect 495266 352338 495502 352574
rect 495586 352338 495822 352574
rect 495266 316658 495502 316894
rect 495586 316658 495822 316894
rect 495266 316338 495502 316574
rect 495586 316338 495822 316574
rect 495266 280658 495502 280894
rect 495586 280658 495822 280894
rect 495266 280338 495502 280574
rect 495586 280338 495822 280574
rect 495266 244658 495502 244894
rect 495586 244658 495822 244894
rect 495266 244338 495502 244574
rect 495586 244338 495822 244574
rect 495266 208658 495502 208894
rect 495586 208658 495822 208894
rect 495266 208338 495502 208574
rect 495586 208338 495822 208574
rect 495266 172658 495502 172894
rect 495586 172658 495822 172894
rect 495266 172338 495502 172574
rect 495586 172338 495822 172574
rect 495266 136658 495502 136894
rect 495586 136658 495822 136894
rect 495266 136338 495502 136574
rect 495586 136338 495822 136574
rect 495266 100658 495502 100894
rect 495586 100658 495822 100894
rect 495266 100338 495502 100574
rect 495586 100338 495822 100574
rect 495266 64658 495502 64894
rect 495586 64658 495822 64894
rect 495266 64338 495502 64574
rect 495586 64338 495822 64574
rect 495266 28658 495502 28894
rect 495586 28658 495822 28894
rect 495266 28338 495502 28574
rect 495586 28338 495822 28574
rect 495266 -5382 495502 -5146
rect 495586 -5382 495822 -5146
rect 495266 -5702 495502 -5466
rect 495586 -5702 495822 -5466
rect 516986 710362 517222 710598
rect 517306 710362 517542 710598
rect 516986 710042 517222 710278
rect 517306 710042 517542 710278
rect 513266 708442 513502 708678
rect 513586 708442 513822 708678
rect 513266 708122 513502 708358
rect 513586 708122 513822 708358
rect 509546 706522 509782 706758
rect 509866 706522 510102 706758
rect 509546 706202 509782 706438
rect 509866 706202 510102 706438
rect 498986 680378 499222 680614
rect 499306 680378 499542 680614
rect 498986 680058 499222 680294
rect 499306 680058 499542 680294
rect 498986 644378 499222 644614
rect 499306 644378 499542 644614
rect 498986 644058 499222 644294
rect 499306 644058 499542 644294
rect 498986 608378 499222 608614
rect 499306 608378 499542 608614
rect 498986 608058 499222 608294
rect 499306 608058 499542 608294
rect 498986 572378 499222 572614
rect 499306 572378 499542 572614
rect 498986 572058 499222 572294
rect 499306 572058 499542 572294
rect 498986 536378 499222 536614
rect 499306 536378 499542 536614
rect 498986 536058 499222 536294
rect 499306 536058 499542 536294
rect 498986 500378 499222 500614
rect 499306 500378 499542 500614
rect 498986 500058 499222 500294
rect 499306 500058 499542 500294
rect 498986 464378 499222 464614
rect 499306 464378 499542 464614
rect 498986 464058 499222 464294
rect 499306 464058 499542 464294
rect 498986 428378 499222 428614
rect 499306 428378 499542 428614
rect 498986 428058 499222 428294
rect 499306 428058 499542 428294
rect 498986 392378 499222 392614
rect 499306 392378 499542 392614
rect 498986 392058 499222 392294
rect 499306 392058 499542 392294
rect 498986 356378 499222 356614
rect 499306 356378 499542 356614
rect 498986 356058 499222 356294
rect 499306 356058 499542 356294
rect 498986 320378 499222 320614
rect 499306 320378 499542 320614
rect 498986 320058 499222 320294
rect 499306 320058 499542 320294
rect 498986 284378 499222 284614
rect 499306 284378 499542 284614
rect 498986 284058 499222 284294
rect 499306 284058 499542 284294
rect 498986 248378 499222 248614
rect 499306 248378 499542 248614
rect 498986 248058 499222 248294
rect 499306 248058 499542 248294
rect 498986 212378 499222 212614
rect 499306 212378 499542 212614
rect 498986 212058 499222 212294
rect 499306 212058 499542 212294
rect 498986 176378 499222 176614
rect 499306 176378 499542 176614
rect 498986 176058 499222 176294
rect 499306 176058 499542 176294
rect 498986 140378 499222 140614
rect 499306 140378 499542 140614
rect 498986 140058 499222 140294
rect 499306 140058 499542 140294
rect 498986 104378 499222 104614
rect 499306 104378 499542 104614
rect 498986 104058 499222 104294
rect 499306 104058 499542 104294
rect 498986 68378 499222 68614
rect 499306 68378 499542 68614
rect 498986 68058 499222 68294
rect 499306 68058 499542 68294
rect 498986 32378 499222 32614
rect 499306 32378 499542 32614
rect 498986 32058 499222 32294
rect 499306 32058 499542 32294
rect 480986 -6342 481222 -6106
rect 481306 -6342 481542 -6106
rect 480986 -6662 481222 -6426
rect 481306 -6662 481542 -6426
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 509546 690938 509782 691174
rect 509866 690938 510102 691174
rect 509546 690618 509782 690854
rect 509866 690618 510102 690854
rect 509546 654938 509782 655174
rect 509866 654938 510102 655174
rect 509546 654618 509782 654854
rect 509866 654618 510102 654854
rect 509546 618938 509782 619174
rect 509866 618938 510102 619174
rect 509546 618618 509782 618854
rect 509866 618618 510102 618854
rect 509546 582938 509782 583174
rect 509866 582938 510102 583174
rect 509546 582618 509782 582854
rect 509866 582618 510102 582854
rect 509546 546938 509782 547174
rect 509866 546938 510102 547174
rect 509546 546618 509782 546854
rect 509866 546618 510102 546854
rect 509546 510938 509782 511174
rect 509866 510938 510102 511174
rect 509546 510618 509782 510854
rect 509866 510618 510102 510854
rect 509546 474938 509782 475174
rect 509866 474938 510102 475174
rect 509546 474618 509782 474854
rect 509866 474618 510102 474854
rect 509546 438938 509782 439174
rect 509866 438938 510102 439174
rect 509546 438618 509782 438854
rect 509866 438618 510102 438854
rect 509546 402938 509782 403174
rect 509866 402938 510102 403174
rect 509546 402618 509782 402854
rect 509866 402618 510102 402854
rect 509546 366938 509782 367174
rect 509866 366938 510102 367174
rect 509546 366618 509782 366854
rect 509866 366618 510102 366854
rect 509546 330938 509782 331174
rect 509866 330938 510102 331174
rect 509546 330618 509782 330854
rect 509866 330618 510102 330854
rect 509546 294938 509782 295174
rect 509866 294938 510102 295174
rect 509546 294618 509782 294854
rect 509866 294618 510102 294854
rect 509546 258938 509782 259174
rect 509866 258938 510102 259174
rect 509546 258618 509782 258854
rect 509866 258618 510102 258854
rect 509546 222938 509782 223174
rect 509866 222938 510102 223174
rect 509546 222618 509782 222854
rect 509866 222618 510102 222854
rect 509546 186938 509782 187174
rect 509866 186938 510102 187174
rect 509546 186618 509782 186854
rect 509866 186618 510102 186854
rect 509546 150938 509782 151174
rect 509866 150938 510102 151174
rect 509546 150618 509782 150854
rect 509866 150618 510102 150854
rect 509546 114938 509782 115174
rect 509866 114938 510102 115174
rect 509546 114618 509782 114854
rect 509866 114618 510102 114854
rect 509546 78938 509782 79174
rect 509866 78938 510102 79174
rect 509546 78618 509782 78854
rect 509866 78618 510102 78854
rect 509546 42938 509782 43174
rect 509866 42938 510102 43174
rect 509546 42618 509782 42854
rect 509866 42618 510102 42854
rect 509546 6938 509782 7174
rect 509866 6938 510102 7174
rect 509546 6618 509782 6854
rect 509866 6618 510102 6854
rect 509546 -2502 509782 -2266
rect 509866 -2502 510102 -2266
rect 509546 -2822 509782 -2586
rect 509866 -2822 510102 -2586
rect 513266 694658 513502 694894
rect 513586 694658 513822 694894
rect 513266 694338 513502 694574
rect 513586 694338 513822 694574
rect 513266 658658 513502 658894
rect 513586 658658 513822 658894
rect 513266 658338 513502 658574
rect 513586 658338 513822 658574
rect 513266 622658 513502 622894
rect 513586 622658 513822 622894
rect 513266 622338 513502 622574
rect 513586 622338 513822 622574
rect 513266 586658 513502 586894
rect 513586 586658 513822 586894
rect 513266 586338 513502 586574
rect 513586 586338 513822 586574
rect 513266 550658 513502 550894
rect 513586 550658 513822 550894
rect 513266 550338 513502 550574
rect 513586 550338 513822 550574
rect 513266 514658 513502 514894
rect 513586 514658 513822 514894
rect 513266 514338 513502 514574
rect 513586 514338 513822 514574
rect 513266 478658 513502 478894
rect 513586 478658 513822 478894
rect 513266 478338 513502 478574
rect 513586 478338 513822 478574
rect 513266 442658 513502 442894
rect 513586 442658 513822 442894
rect 513266 442338 513502 442574
rect 513586 442338 513822 442574
rect 513266 406658 513502 406894
rect 513586 406658 513822 406894
rect 513266 406338 513502 406574
rect 513586 406338 513822 406574
rect 513266 370658 513502 370894
rect 513586 370658 513822 370894
rect 513266 370338 513502 370574
rect 513586 370338 513822 370574
rect 513266 334658 513502 334894
rect 513586 334658 513822 334894
rect 513266 334338 513502 334574
rect 513586 334338 513822 334574
rect 513266 298658 513502 298894
rect 513586 298658 513822 298894
rect 513266 298338 513502 298574
rect 513586 298338 513822 298574
rect 513266 262658 513502 262894
rect 513586 262658 513822 262894
rect 513266 262338 513502 262574
rect 513586 262338 513822 262574
rect 513266 226658 513502 226894
rect 513586 226658 513822 226894
rect 513266 226338 513502 226574
rect 513586 226338 513822 226574
rect 513266 190658 513502 190894
rect 513586 190658 513822 190894
rect 513266 190338 513502 190574
rect 513586 190338 513822 190574
rect 513266 154658 513502 154894
rect 513586 154658 513822 154894
rect 513266 154338 513502 154574
rect 513586 154338 513822 154574
rect 513266 118658 513502 118894
rect 513586 118658 513822 118894
rect 513266 118338 513502 118574
rect 513586 118338 513822 118574
rect 513266 82658 513502 82894
rect 513586 82658 513822 82894
rect 513266 82338 513502 82574
rect 513586 82338 513822 82574
rect 513266 46658 513502 46894
rect 513586 46658 513822 46894
rect 513266 46338 513502 46574
rect 513586 46338 513822 46574
rect 513266 10658 513502 10894
rect 513586 10658 513822 10894
rect 513266 10338 513502 10574
rect 513586 10338 513822 10574
rect 513266 -4422 513502 -4186
rect 513586 -4422 513822 -4186
rect 513266 -4742 513502 -4506
rect 513586 -4742 513822 -4506
rect 534986 711322 535222 711558
rect 535306 711322 535542 711558
rect 534986 711002 535222 711238
rect 535306 711002 535542 711238
rect 531266 709402 531502 709638
rect 531586 709402 531822 709638
rect 531266 709082 531502 709318
rect 531586 709082 531822 709318
rect 527546 707482 527782 707718
rect 527866 707482 528102 707718
rect 527546 707162 527782 707398
rect 527866 707162 528102 707398
rect 516986 698378 517222 698614
rect 517306 698378 517542 698614
rect 516986 698058 517222 698294
rect 517306 698058 517542 698294
rect 516986 662378 517222 662614
rect 517306 662378 517542 662614
rect 516986 662058 517222 662294
rect 517306 662058 517542 662294
rect 516986 626378 517222 626614
rect 517306 626378 517542 626614
rect 516986 626058 517222 626294
rect 517306 626058 517542 626294
rect 516986 590378 517222 590614
rect 517306 590378 517542 590614
rect 516986 590058 517222 590294
rect 517306 590058 517542 590294
rect 516986 554378 517222 554614
rect 517306 554378 517542 554614
rect 516986 554058 517222 554294
rect 517306 554058 517542 554294
rect 516986 518378 517222 518614
rect 517306 518378 517542 518614
rect 516986 518058 517222 518294
rect 517306 518058 517542 518294
rect 516986 482378 517222 482614
rect 517306 482378 517542 482614
rect 516986 482058 517222 482294
rect 517306 482058 517542 482294
rect 516986 446378 517222 446614
rect 517306 446378 517542 446614
rect 516986 446058 517222 446294
rect 517306 446058 517542 446294
rect 516986 410378 517222 410614
rect 517306 410378 517542 410614
rect 516986 410058 517222 410294
rect 517306 410058 517542 410294
rect 516986 374378 517222 374614
rect 517306 374378 517542 374614
rect 516986 374058 517222 374294
rect 517306 374058 517542 374294
rect 516986 338378 517222 338614
rect 517306 338378 517542 338614
rect 516986 338058 517222 338294
rect 517306 338058 517542 338294
rect 516986 302378 517222 302614
rect 517306 302378 517542 302614
rect 516986 302058 517222 302294
rect 517306 302058 517542 302294
rect 516986 266378 517222 266614
rect 517306 266378 517542 266614
rect 516986 266058 517222 266294
rect 517306 266058 517542 266294
rect 516986 230378 517222 230614
rect 517306 230378 517542 230614
rect 516986 230058 517222 230294
rect 517306 230058 517542 230294
rect 516986 194378 517222 194614
rect 517306 194378 517542 194614
rect 516986 194058 517222 194294
rect 517306 194058 517542 194294
rect 516986 158378 517222 158614
rect 517306 158378 517542 158614
rect 516986 158058 517222 158294
rect 517306 158058 517542 158294
rect 516986 122378 517222 122614
rect 517306 122378 517542 122614
rect 516986 122058 517222 122294
rect 517306 122058 517542 122294
rect 516986 86378 517222 86614
rect 517306 86378 517542 86614
rect 516986 86058 517222 86294
rect 517306 86058 517542 86294
rect 516986 50378 517222 50614
rect 517306 50378 517542 50614
rect 516986 50058 517222 50294
rect 517306 50058 517542 50294
rect 516986 14378 517222 14614
rect 517306 14378 517542 14614
rect 516986 14058 517222 14294
rect 517306 14058 517542 14294
rect 498986 -7302 499222 -7066
rect 499306 -7302 499542 -7066
rect 498986 -7622 499222 -7386
rect 499306 -7622 499542 -7386
rect 523826 705562 524062 705798
rect 524146 705562 524382 705798
rect 523826 705242 524062 705478
rect 524146 705242 524382 705478
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -1542 524062 -1306
rect 524146 -1542 524382 -1306
rect 523826 -1862 524062 -1626
rect 524146 -1862 524382 -1626
rect 527546 672938 527782 673174
rect 527866 672938 528102 673174
rect 527546 672618 527782 672854
rect 527866 672618 528102 672854
rect 527546 636938 527782 637174
rect 527866 636938 528102 637174
rect 527546 636618 527782 636854
rect 527866 636618 528102 636854
rect 527546 600938 527782 601174
rect 527866 600938 528102 601174
rect 527546 600618 527782 600854
rect 527866 600618 528102 600854
rect 527546 564938 527782 565174
rect 527866 564938 528102 565174
rect 527546 564618 527782 564854
rect 527866 564618 528102 564854
rect 527546 528938 527782 529174
rect 527866 528938 528102 529174
rect 527546 528618 527782 528854
rect 527866 528618 528102 528854
rect 527546 492938 527782 493174
rect 527866 492938 528102 493174
rect 527546 492618 527782 492854
rect 527866 492618 528102 492854
rect 527546 456938 527782 457174
rect 527866 456938 528102 457174
rect 527546 456618 527782 456854
rect 527866 456618 528102 456854
rect 527546 420938 527782 421174
rect 527866 420938 528102 421174
rect 527546 420618 527782 420854
rect 527866 420618 528102 420854
rect 527546 384938 527782 385174
rect 527866 384938 528102 385174
rect 527546 384618 527782 384854
rect 527866 384618 528102 384854
rect 527546 348938 527782 349174
rect 527866 348938 528102 349174
rect 527546 348618 527782 348854
rect 527866 348618 528102 348854
rect 527546 312938 527782 313174
rect 527866 312938 528102 313174
rect 527546 312618 527782 312854
rect 527866 312618 528102 312854
rect 527546 276938 527782 277174
rect 527866 276938 528102 277174
rect 527546 276618 527782 276854
rect 527866 276618 528102 276854
rect 527546 240938 527782 241174
rect 527866 240938 528102 241174
rect 527546 240618 527782 240854
rect 527866 240618 528102 240854
rect 527546 204938 527782 205174
rect 527866 204938 528102 205174
rect 527546 204618 527782 204854
rect 527866 204618 528102 204854
rect 527546 168938 527782 169174
rect 527866 168938 528102 169174
rect 527546 168618 527782 168854
rect 527866 168618 528102 168854
rect 527546 132938 527782 133174
rect 527866 132938 528102 133174
rect 527546 132618 527782 132854
rect 527866 132618 528102 132854
rect 527546 96938 527782 97174
rect 527866 96938 528102 97174
rect 527546 96618 527782 96854
rect 527866 96618 528102 96854
rect 527546 60938 527782 61174
rect 527866 60938 528102 61174
rect 527546 60618 527782 60854
rect 527866 60618 528102 60854
rect 527546 24938 527782 25174
rect 527866 24938 528102 25174
rect 527546 24618 527782 24854
rect 527866 24618 528102 24854
rect 527546 -3462 527782 -3226
rect 527866 -3462 528102 -3226
rect 527546 -3782 527782 -3546
rect 527866 -3782 528102 -3546
rect 531266 676658 531502 676894
rect 531586 676658 531822 676894
rect 531266 676338 531502 676574
rect 531586 676338 531822 676574
rect 531266 640658 531502 640894
rect 531586 640658 531822 640894
rect 531266 640338 531502 640574
rect 531586 640338 531822 640574
rect 531266 604658 531502 604894
rect 531586 604658 531822 604894
rect 531266 604338 531502 604574
rect 531586 604338 531822 604574
rect 531266 568658 531502 568894
rect 531586 568658 531822 568894
rect 531266 568338 531502 568574
rect 531586 568338 531822 568574
rect 531266 532658 531502 532894
rect 531586 532658 531822 532894
rect 531266 532338 531502 532574
rect 531586 532338 531822 532574
rect 531266 496658 531502 496894
rect 531586 496658 531822 496894
rect 531266 496338 531502 496574
rect 531586 496338 531822 496574
rect 531266 460658 531502 460894
rect 531586 460658 531822 460894
rect 531266 460338 531502 460574
rect 531586 460338 531822 460574
rect 531266 424658 531502 424894
rect 531586 424658 531822 424894
rect 531266 424338 531502 424574
rect 531586 424338 531822 424574
rect 531266 388658 531502 388894
rect 531586 388658 531822 388894
rect 531266 388338 531502 388574
rect 531586 388338 531822 388574
rect 531266 352658 531502 352894
rect 531586 352658 531822 352894
rect 531266 352338 531502 352574
rect 531586 352338 531822 352574
rect 531266 316658 531502 316894
rect 531586 316658 531822 316894
rect 531266 316338 531502 316574
rect 531586 316338 531822 316574
rect 531266 280658 531502 280894
rect 531586 280658 531822 280894
rect 531266 280338 531502 280574
rect 531586 280338 531822 280574
rect 531266 244658 531502 244894
rect 531586 244658 531822 244894
rect 531266 244338 531502 244574
rect 531586 244338 531822 244574
rect 531266 208658 531502 208894
rect 531586 208658 531822 208894
rect 531266 208338 531502 208574
rect 531586 208338 531822 208574
rect 531266 172658 531502 172894
rect 531586 172658 531822 172894
rect 531266 172338 531502 172574
rect 531586 172338 531822 172574
rect 531266 136658 531502 136894
rect 531586 136658 531822 136894
rect 531266 136338 531502 136574
rect 531586 136338 531822 136574
rect 531266 100658 531502 100894
rect 531586 100658 531822 100894
rect 531266 100338 531502 100574
rect 531586 100338 531822 100574
rect 531266 64658 531502 64894
rect 531586 64658 531822 64894
rect 531266 64338 531502 64574
rect 531586 64338 531822 64574
rect 531266 28658 531502 28894
rect 531586 28658 531822 28894
rect 531266 28338 531502 28574
rect 531586 28338 531822 28574
rect 531266 -5382 531502 -5146
rect 531586 -5382 531822 -5146
rect 531266 -5702 531502 -5466
rect 531586 -5702 531822 -5466
rect 552986 710362 553222 710598
rect 553306 710362 553542 710598
rect 552986 710042 553222 710278
rect 553306 710042 553542 710278
rect 549266 708442 549502 708678
rect 549586 708442 549822 708678
rect 549266 708122 549502 708358
rect 549586 708122 549822 708358
rect 545546 706522 545782 706758
rect 545866 706522 546102 706758
rect 545546 706202 545782 706438
rect 545866 706202 546102 706438
rect 534986 680378 535222 680614
rect 535306 680378 535542 680614
rect 534986 680058 535222 680294
rect 535306 680058 535542 680294
rect 534986 644378 535222 644614
rect 535306 644378 535542 644614
rect 534986 644058 535222 644294
rect 535306 644058 535542 644294
rect 534986 608378 535222 608614
rect 535306 608378 535542 608614
rect 534986 608058 535222 608294
rect 535306 608058 535542 608294
rect 534986 572378 535222 572614
rect 535306 572378 535542 572614
rect 534986 572058 535222 572294
rect 535306 572058 535542 572294
rect 534986 536378 535222 536614
rect 535306 536378 535542 536614
rect 534986 536058 535222 536294
rect 535306 536058 535542 536294
rect 534986 500378 535222 500614
rect 535306 500378 535542 500614
rect 534986 500058 535222 500294
rect 535306 500058 535542 500294
rect 534986 464378 535222 464614
rect 535306 464378 535542 464614
rect 534986 464058 535222 464294
rect 535306 464058 535542 464294
rect 534986 428378 535222 428614
rect 535306 428378 535542 428614
rect 534986 428058 535222 428294
rect 535306 428058 535542 428294
rect 534986 392378 535222 392614
rect 535306 392378 535542 392614
rect 534986 392058 535222 392294
rect 535306 392058 535542 392294
rect 534986 356378 535222 356614
rect 535306 356378 535542 356614
rect 534986 356058 535222 356294
rect 535306 356058 535542 356294
rect 534986 320378 535222 320614
rect 535306 320378 535542 320614
rect 534986 320058 535222 320294
rect 535306 320058 535542 320294
rect 534986 284378 535222 284614
rect 535306 284378 535542 284614
rect 534986 284058 535222 284294
rect 535306 284058 535542 284294
rect 534986 248378 535222 248614
rect 535306 248378 535542 248614
rect 534986 248058 535222 248294
rect 535306 248058 535542 248294
rect 534986 212378 535222 212614
rect 535306 212378 535542 212614
rect 534986 212058 535222 212294
rect 535306 212058 535542 212294
rect 534986 176378 535222 176614
rect 535306 176378 535542 176614
rect 534986 176058 535222 176294
rect 535306 176058 535542 176294
rect 534986 140378 535222 140614
rect 535306 140378 535542 140614
rect 534986 140058 535222 140294
rect 535306 140058 535542 140294
rect 534986 104378 535222 104614
rect 535306 104378 535542 104614
rect 534986 104058 535222 104294
rect 535306 104058 535542 104294
rect 534986 68378 535222 68614
rect 535306 68378 535542 68614
rect 534986 68058 535222 68294
rect 535306 68058 535542 68294
rect 534986 32378 535222 32614
rect 535306 32378 535542 32614
rect 534986 32058 535222 32294
rect 535306 32058 535542 32294
rect 516986 -6342 517222 -6106
rect 517306 -6342 517542 -6106
rect 516986 -6662 517222 -6426
rect 517306 -6662 517542 -6426
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 545546 690938 545782 691174
rect 545866 690938 546102 691174
rect 545546 690618 545782 690854
rect 545866 690618 546102 690854
rect 545546 654938 545782 655174
rect 545866 654938 546102 655174
rect 545546 654618 545782 654854
rect 545866 654618 546102 654854
rect 545546 618938 545782 619174
rect 545866 618938 546102 619174
rect 545546 618618 545782 618854
rect 545866 618618 546102 618854
rect 545546 582938 545782 583174
rect 545866 582938 546102 583174
rect 545546 582618 545782 582854
rect 545866 582618 546102 582854
rect 545546 546938 545782 547174
rect 545866 546938 546102 547174
rect 545546 546618 545782 546854
rect 545866 546618 546102 546854
rect 545546 510938 545782 511174
rect 545866 510938 546102 511174
rect 545546 510618 545782 510854
rect 545866 510618 546102 510854
rect 545546 474938 545782 475174
rect 545866 474938 546102 475174
rect 545546 474618 545782 474854
rect 545866 474618 546102 474854
rect 545546 438938 545782 439174
rect 545866 438938 546102 439174
rect 545546 438618 545782 438854
rect 545866 438618 546102 438854
rect 545546 402938 545782 403174
rect 545866 402938 546102 403174
rect 545546 402618 545782 402854
rect 545866 402618 546102 402854
rect 545546 366938 545782 367174
rect 545866 366938 546102 367174
rect 545546 366618 545782 366854
rect 545866 366618 546102 366854
rect 545546 330938 545782 331174
rect 545866 330938 546102 331174
rect 545546 330618 545782 330854
rect 545866 330618 546102 330854
rect 545546 294938 545782 295174
rect 545866 294938 546102 295174
rect 545546 294618 545782 294854
rect 545866 294618 546102 294854
rect 545546 258938 545782 259174
rect 545866 258938 546102 259174
rect 545546 258618 545782 258854
rect 545866 258618 546102 258854
rect 545546 222938 545782 223174
rect 545866 222938 546102 223174
rect 545546 222618 545782 222854
rect 545866 222618 546102 222854
rect 545546 186938 545782 187174
rect 545866 186938 546102 187174
rect 545546 186618 545782 186854
rect 545866 186618 546102 186854
rect 545546 150938 545782 151174
rect 545866 150938 546102 151174
rect 545546 150618 545782 150854
rect 545866 150618 546102 150854
rect 545546 114938 545782 115174
rect 545866 114938 546102 115174
rect 545546 114618 545782 114854
rect 545866 114618 546102 114854
rect 545546 78938 545782 79174
rect 545866 78938 546102 79174
rect 545546 78618 545782 78854
rect 545866 78618 546102 78854
rect 545546 42938 545782 43174
rect 545866 42938 546102 43174
rect 545546 42618 545782 42854
rect 545866 42618 546102 42854
rect 545546 6938 545782 7174
rect 545866 6938 546102 7174
rect 545546 6618 545782 6854
rect 545866 6618 546102 6854
rect 545546 -2502 545782 -2266
rect 545866 -2502 546102 -2266
rect 545546 -2822 545782 -2586
rect 545866 -2822 546102 -2586
rect 549266 694658 549502 694894
rect 549586 694658 549822 694894
rect 549266 694338 549502 694574
rect 549586 694338 549822 694574
rect 549266 658658 549502 658894
rect 549586 658658 549822 658894
rect 549266 658338 549502 658574
rect 549586 658338 549822 658574
rect 549266 622658 549502 622894
rect 549586 622658 549822 622894
rect 549266 622338 549502 622574
rect 549586 622338 549822 622574
rect 549266 586658 549502 586894
rect 549586 586658 549822 586894
rect 549266 586338 549502 586574
rect 549586 586338 549822 586574
rect 549266 550658 549502 550894
rect 549586 550658 549822 550894
rect 549266 550338 549502 550574
rect 549586 550338 549822 550574
rect 549266 514658 549502 514894
rect 549586 514658 549822 514894
rect 549266 514338 549502 514574
rect 549586 514338 549822 514574
rect 549266 478658 549502 478894
rect 549586 478658 549822 478894
rect 549266 478338 549502 478574
rect 549586 478338 549822 478574
rect 549266 442658 549502 442894
rect 549586 442658 549822 442894
rect 549266 442338 549502 442574
rect 549586 442338 549822 442574
rect 549266 406658 549502 406894
rect 549586 406658 549822 406894
rect 549266 406338 549502 406574
rect 549586 406338 549822 406574
rect 549266 370658 549502 370894
rect 549586 370658 549822 370894
rect 549266 370338 549502 370574
rect 549586 370338 549822 370574
rect 549266 334658 549502 334894
rect 549586 334658 549822 334894
rect 549266 334338 549502 334574
rect 549586 334338 549822 334574
rect 549266 298658 549502 298894
rect 549586 298658 549822 298894
rect 549266 298338 549502 298574
rect 549586 298338 549822 298574
rect 549266 262658 549502 262894
rect 549586 262658 549822 262894
rect 549266 262338 549502 262574
rect 549586 262338 549822 262574
rect 549266 226658 549502 226894
rect 549586 226658 549822 226894
rect 549266 226338 549502 226574
rect 549586 226338 549822 226574
rect 549266 190658 549502 190894
rect 549586 190658 549822 190894
rect 549266 190338 549502 190574
rect 549586 190338 549822 190574
rect 549266 154658 549502 154894
rect 549586 154658 549822 154894
rect 549266 154338 549502 154574
rect 549586 154338 549822 154574
rect 549266 118658 549502 118894
rect 549586 118658 549822 118894
rect 549266 118338 549502 118574
rect 549586 118338 549822 118574
rect 549266 82658 549502 82894
rect 549586 82658 549822 82894
rect 549266 82338 549502 82574
rect 549586 82338 549822 82574
rect 549266 46658 549502 46894
rect 549586 46658 549822 46894
rect 549266 46338 549502 46574
rect 549586 46338 549822 46574
rect 549266 10658 549502 10894
rect 549586 10658 549822 10894
rect 549266 10338 549502 10574
rect 549586 10338 549822 10574
rect 549266 -4422 549502 -4186
rect 549586 -4422 549822 -4186
rect 549266 -4742 549502 -4506
rect 549586 -4742 549822 -4506
rect 570986 711322 571222 711558
rect 571306 711322 571542 711558
rect 570986 711002 571222 711238
rect 571306 711002 571542 711238
rect 567266 709402 567502 709638
rect 567586 709402 567822 709638
rect 567266 709082 567502 709318
rect 567586 709082 567822 709318
rect 563546 707482 563782 707718
rect 563866 707482 564102 707718
rect 563546 707162 563782 707398
rect 563866 707162 564102 707398
rect 552986 698378 553222 698614
rect 553306 698378 553542 698614
rect 552986 698058 553222 698294
rect 553306 698058 553542 698294
rect 552986 662378 553222 662614
rect 553306 662378 553542 662614
rect 552986 662058 553222 662294
rect 553306 662058 553542 662294
rect 552986 626378 553222 626614
rect 553306 626378 553542 626614
rect 552986 626058 553222 626294
rect 553306 626058 553542 626294
rect 552986 590378 553222 590614
rect 553306 590378 553542 590614
rect 552986 590058 553222 590294
rect 553306 590058 553542 590294
rect 552986 554378 553222 554614
rect 553306 554378 553542 554614
rect 552986 554058 553222 554294
rect 553306 554058 553542 554294
rect 552986 518378 553222 518614
rect 553306 518378 553542 518614
rect 552986 518058 553222 518294
rect 553306 518058 553542 518294
rect 552986 482378 553222 482614
rect 553306 482378 553542 482614
rect 552986 482058 553222 482294
rect 553306 482058 553542 482294
rect 552986 446378 553222 446614
rect 553306 446378 553542 446614
rect 552986 446058 553222 446294
rect 553306 446058 553542 446294
rect 552986 410378 553222 410614
rect 553306 410378 553542 410614
rect 552986 410058 553222 410294
rect 553306 410058 553542 410294
rect 552986 374378 553222 374614
rect 553306 374378 553542 374614
rect 552986 374058 553222 374294
rect 553306 374058 553542 374294
rect 552986 338378 553222 338614
rect 553306 338378 553542 338614
rect 552986 338058 553222 338294
rect 553306 338058 553542 338294
rect 552986 302378 553222 302614
rect 553306 302378 553542 302614
rect 552986 302058 553222 302294
rect 553306 302058 553542 302294
rect 552986 266378 553222 266614
rect 553306 266378 553542 266614
rect 552986 266058 553222 266294
rect 553306 266058 553542 266294
rect 552986 230378 553222 230614
rect 553306 230378 553542 230614
rect 552986 230058 553222 230294
rect 553306 230058 553542 230294
rect 552986 194378 553222 194614
rect 553306 194378 553542 194614
rect 552986 194058 553222 194294
rect 553306 194058 553542 194294
rect 552986 158378 553222 158614
rect 553306 158378 553542 158614
rect 552986 158058 553222 158294
rect 553306 158058 553542 158294
rect 552986 122378 553222 122614
rect 553306 122378 553542 122614
rect 552986 122058 553222 122294
rect 553306 122058 553542 122294
rect 552986 86378 553222 86614
rect 553306 86378 553542 86614
rect 552986 86058 553222 86294
rect 553306 86058 553542 86294
rect 552986 50378 553222 50614
rect 553306 50378 553542 50614
rect 552986 50058 553222 50294
rect 553306 50058 553542 50294
rect 552986 14378 553222 14614
rect 553306 14378 553542 14614
rect 552986 14058 553222 14294
rect 553306 14058 553542 14294
rect 534986 -7302 535222 -7066
rect 535306 -7302 535542 -7066
rect 534986 -7622 535222 -7386
rect 535306 -7622 535542 -7386
rect 559826 705562 560062 705798
rect 560146 705562 560382 705798
rect 559826 705242 560062 705478
rect 560146 705242 560382 705478
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -1542 560062 -1306
rect 560146 -1542 560382 -1306
rect 559826 -1862 560062 -1626
rect 560146 -1862 560382 -1626
rect 563546 672938 563782 673174
rect 563866 672938 564102 673174
rect 563546 672618 563782 672854
rect 563866 672618 564102 672854
rect 563546 636938 563782 637174
rect 563866 636938 564102 637174
rect 563546 636618 563782 636854
rect 563866 636618 564102 636854
rect 563546 600938 563782 601174
rect 563866 600938 564102 601174
rect 563546 600618 563782 600854
rect 563866 600618 564102 600854
rect 563546 564938 563782 565174
rect 563866 564938 564102 565174
rect 563546 564618 563782 564854
rect 563866 564618 564102 564854
rect 563546 528938 563782 529174
rect 563866 528938 564102 529174
rect 563546 528618 563782 528854
rect 563866 528618 564102 528854
rect 563546 492938 563782 493174
rect 563866 492938 564102 493174
rect 563546 492618 563782 492854
rect 563866 492618 564102 492854
rect 563546 456938 563782 457174
rect 563866 456938 564102 457174
rect 563546 456618 563782 456854
rect 563866 456618 564102 456854
rect 563546 420938 563782 421174
rect 563866 420938 564102 421174
rect 563546 420618 563782 420854
rect 563866 420618 564102 420854
rect 563546 384938 563782 385174
rect 563866 384938 564102 385174
rect 563546 384618 563782 384854
rect 563866 384618 564102 384854
rect 563546 348938 563782 349174
rect 563866 348938 564102 349174
rect 563546 348618 563782 348854
rect 563866 348618 564102 348854
rect 563546 312938 563782 313174
rect 563866 312938 564102 313174
rect 563546 312618 563782 312854
rect 563866 312618 564102 312854
rect 563546 276938 563782 277174
rect 563866 276938 564102 277174
rect 563546 276618 563782 276854
rect 563866 276618 564102 276854
rect 563546 240938 563782 241174
rect 563866 240938 564102 241174
rect 563546 240618 563782 240854
rect 563866 240618 564102 240854
rect 563546 204938 563782 205174
rect 563866 204938 564102 205174
rect 563546 204618 563782 204854
rect 563866 204618 564102 204854
rect 563546 168938 563782 169174
rect 563866 168938 564102 169174
rect 563546 168618 563782 168854
rect 563866 168618 564102 168854
rect 563546 132938 563782 133174
rect 563866 132938 564102 133174
rect 563546 132618 563782 132854
rect 563866 132618 564102 132854
rect 563546 96938 563782 97174
rect 563866 96938 564102 97174
rect 563546 96618 563782 96854
rect 563866 96618 564102 96854
rect 563546 60938 563782 61174
rect 563866 60938 564102 61174
rect 563546 60618 563782 60854
rect 563866 60618 564102 60854
rect 563546 24938 563782 25174
rect 563866 24938 564102 25174
rect 563546 24618 563782 24854
rect 563866 24618 564102 24854
rect 563546 -3462 563782 -3226
rect 563866 -3462 564102 -3226
rect 563546 -3782 563782 -3546
rect 563866 -3782 564102 -3546
rect 567266 676658 567502 676894
rect 567586 676658 567822 676894
rect 567266 676338 567502 676574
rect 567586 676338 567822 676574
rect 567266 640658 567502 640894
rect 567586 640658 567822 640894
rect 567266 640338 567502 640574
rect 567586 640338 567822 640574
rect 567266 604658 567502 604894
rect 567586 604658 567822 604894
rect 567266 604338 567502 604574
rect 567586 604338 567822 604574
rect 567266 568658 567502 568894
rect 567586 568658 567822 568894
rect 567266 568338 567502 568574
rect 567586 568338 567822 568574
rect 567266 532658 567502 532894
rect 567586 532658 567822 532894
rect 567266 532338 567502 532574
rect 567586 532338 567822 532574
rect 567266 496658 567502 496894
rect 567586 496658 567822 496894
rect 567266 496338 567502 496574
rect 567586 496338 567822 496574
rect 567266 460658 567502 460894
rect 567586 460658 567822 460894
rect 567266 460338 567502 460574
rect 567586 460338 567822 460574
rect 567266 424658 567502 424894
rect 567586 424658 567822 424894
rect 567266 424338 567502 424574
rect 567586 424338 567822 424574
rect 567266 388658 567502 388894
rect 567586 388658 567822 388894
rect 567266 388338 567502 388574
rect 567586 388338 567822 388574
rect 567266 352658 567502 352894
rect 567586 352658 567822 352894
rect 567266 352338 567502 352574
rect 567586 352338 567822 352574
rect 567266 316658 567502 316894
rect 567586 316658 567822 316894
rect 567266 316338 567502 316574
rect 567586 316338 567822 316574
rect 567266 280658 567502 280894
rect 567586 280658 567822 280894
rect 567266 280338 567502 280574
rect 567586 280338 567822 280574
rect 567266 244658 567502 244894
rect 567586 244658 567822 244894
rect 567266 244338 567502 244574
rect 567586 244338 567822 244574
rect 567266 208658 567502 208894
rect 567586 208658 567822 208894
rect 567266 208338 567502 208574
rect 567586 208338 567822 208574
rect 567266 172658 567502 172894
rect 567586 172658 567822 172894
rect 567266 172338 567502 172574
rect 567586 172338 567822 172574
rect 567266 136658 567502 136894
rect 567586 136658 567822 136894
rect 567266 136338 567502 136574
rect 567586 136338 567822 136574
rect 567266 100658 567502 100894
rect 567586 100658 567822 100894
rect 567266 100338 567502 100574
rect 567586 100338 567822 100574
rect 567266 64658 567502 64894
rect 567586 64658 567822 64894
rect 567266 64338 567502 64574
rect 567586 64338 567822 64574
rect 567266 28658 567502 28894
rect 567586 28658 567822 28894
rect 567266 28338 567502 28574
rect 567586 28338 567822 28574
rect 567266 -5382 567502 -5146
rect 567586 -5382 567822 -5146
rect 567266 -5702 567502 -5466
rect 567586 -5702 567822 -5466
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 581546 706522 581782 706758
rect 581866 706522 582102 706758
rect 581546 706202 581782 706438
rect 581866 706202 582102 706438
rect 570986 680378 571222 680614
rect 571306 680378 571542 680614
rect 570986 680058 571222 680294
rect 571306 680058 571542 680294
rect 570986 644378 571222 644614
rect 571306 644378 571542 644614
rect 570986 644058 571222 644294
rect 571306 644058 571542 644294
rect 570986 608378 571222 608614
rect 571306 608378 571542 608614
rect 570986 608058 571222 608294
rect 571306 608058 571542 608294
rect 570986 572378 571222 572614
rect 571306 572378 571542 572614
rect 570986 572058 571222 572294
rect 571306 572058 571542 572294
rect 570986 536378 571222 536614
rect 571306 536378 571542 536614
rect 570986 536058 571222 536294
rect 571306 536058 571542 536294
rect 570986 500378 571222 500614
rect 571306 500378 571542 500614
rect 570986 500058 571222 500294
rect 571306 500058 571542 500294
rect 570986 464378 571222 464614
rect 571306 464378 571542 464614
rect 570986 464058 571222 464294
rect 571306 464058 571542 464294
rect 570986 428378 571222 428614
rect 571306 428378 571542 428614
rect 570986 428058 571222 428294
rect 571306 428058 571542 428294
rect 570986 392378 571222 392614
rect 571306 392378 571542 392614
rect 570986 392058 571222 392294
rect 571306 392058 571542 392294
rect 570986 356378 571222 356614
rect 571306 356378 571542 356614
rect 570986 356058 571222 356294
rect 571306 356058 571542 356294
rect 570986 320378 571222 320614
rect 571306 320378 571542 320614
rect 570986 320058 571222 320294
rect 571306 320058 571542 320294
rect 570986 284378 571222 284614
rect 571306 284378 571542 284614
rect 570986 284058 571222 284294
rect 571306 284058 571542 284294
rect 570986 248378 571222 248614
rect 571306 248378 571542 248614
rect 570986 248058 571222 248294
rect 571306 248058 571542 248294
rect 570986 212378 571222 212614
rect 571306 212378 571542 212614
rect 570986 212058 571222 212294
rect 571306 212058 571542 212294
rect 570986 176378 571222 176614
rect 571306 176378 571542 176614
rect 570986 176058 571222 176294
rect 571306 176058 571542 176294
rect 570986 140378 571222 140614
rect 571306 140378 571542 140614
rect 570986 140058 571222 140294
rect 571306 140058 571542 140294
rect 570986 104378 571222 104614
rect 571306 104378 571542 104614
rect 570986 104058 571222 104294
rect 571306 104058 571542 104294
rect 570986 68378 571222 68614
rect 571306 68378 571542 68614
rect 570986 68058 571222 68294
rect 571306 68058 571542 68294
rect 570986 32378 571222 32614
rect 571306 32378 571542 32614
rect 570986 32058 571222 32294
rect 571306 32058 571542 32294
rect 552986 -6342 553222 -6106
rect 553306 -6342 553542 -6106
rect 552986 -6662 553222 -6426
rect 553306 -6662 553542 -6426
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581546 690938 581782 691174
rect 581866 690938 582102 691174
rect 581546 690618 581782 690854
rect 581866 690618 582102 690854
rect 581546 654938 581782 655174
rect 581866 654938 582102 655174
rect 581546 654618 581782 654854
rect 581866 654618 582102 654854
rect 581546 618938 581782 619174
rect 581866 618938 582102 619174
rect 581546 618618 581782 618854
rect 581866 618618 582102 618854
rect 581546 582938 581782 583174
rect 581866 582938 582102 583174
rect 581546 582618 581782 582854
rect 581866 582618 582102 582854
rect 581546 546938 581782 547174
rect 581866 546938 582102 547174
rect 581546 546618 581782 546854
rect 581866 546618 582102 546854
rect 581546 510938 581782 511174
rect 581866 510938 582102 511174
rect 581546 510618 581782 510854
rect 581866 510618 582102 510854
rect 581546 474938 581782 475174
rect 581866 474938 582102 475174
rect 581546 474618 581782 474854
rect 581866 474618 582102 474854
rect 581546 438938 581782 439174
rect 581866 438938 582102 439174
rect 581546 438618 581782 438854
rect 581866 438618 582102 438854
rect 581546 402938 581782 403174
rect 581866 402938 582102 403174
rect 581546 402618 581782 402854
rect 581866 402618 582102 402854
rect 581546 366938 581782 367174
rect 581866 366938 582102 367174
rect 581546 366618 581782 366854
rect 581866 366618 582102 366854
rect 581546 330938 581782 331174
rect 581866 330938 582102 331174
rect 581546 330618 581782 330854
rect 581866 330618 582102 330854
rect 581546 294938 581782 295174
rect 581866 294938 582102 295174
rect 581546 294618 581782 294854
rect 581866 294618 582102 294854
rect 581546 258938 581782 259174
rect 581866 258938 582102 259174
rect 581546 258618 581782 258854
rect 581866 258618 582102 258854
rect 581546 222938 581782 223174
rect 581866 222938 582102 223174
rect 581546 222618 581782 222854
rect 581866 222618 582102 222854
rect 581546 186938 581782 187174
rect 581866 186938 582102 187174
rect 581546 186618 581782 186854
rect 581866 186618 582102 186854
rect 581546 150938 581782 151174
rect 581866 150938 582102 151174
rect 581546 150618 581782 150854
rect 581866 150618 582102 150854
rect 581546 114938 581782 115174
rect 581866 114938 582102 115174
rect 581546 114618 581782 114854
rect 581866 114618 582102 114854
rect 581546 78938 581782 79174
rect 581866 78938 582102 79174
rect 581546 78618 581782 78854
rect 581866 78618 582102 78854
rect 581546 42938 581782 43174
rect 581866 42938 582102 43174
rect 581546 42618 581782 42854
rect 581866 42618 582102 42854
rect 581546 6938 581782 7174
rect 581866 6938 582102 7174
rect 581546 6618 581782 6854
rect 581866 6618 582102 6854
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 669218 586538 669454
rect 586622 669218 586858 669454
rect 586302 668898 586538 669134
rect 586622 668898 586858 669134
rect 586302 633218 586538 633454
rect 586622 633218 586858 633454
rect 586302 632898 586538 633134
rect 586622 632898 586858 633134
rect 586302 597218 586538 597454
rect 586622 597218 586858 597454
rect 586302 596898 586538 597134
rect 586622 596898 586858 597134
rect 586302 561218 586538 561454
rect 586622 561218 586858 561454
rect 586302 560898 586538 561134
rect 586622 560898 586858 561134
rect 586302 525218 586538 525454
rect 586622 525218 586858 525454
rect 586302 524898 586538 525134
rect 586622 524898 586858 525134
rect 586302 489218 586538 489454
rect 586622 489218 586858 489454
rect 586302 488898 586538 489134
rect 586622 488898 586858 489134
rect 586302 453218 586538 453454
rect 586622 453218 586858 453454
rect 586302 452898 586538 453134
rect 586622 452898 586858 453134
rect 586302 417218 586538 417454
rect 586622 417218 586858 417454
rect 586302 416898 586538 417134
rect 586622 416898 586858 417134
rect 586302 381218 586538 381454
rect 586622 381218 586858 381454
rect 586302 380898 586538 381134
rect 586622 380898 586858 381134
rect 586302 345218 586538 345454
rect 586622 345218 586858 345454
rect 586302 344898 586538 345134
rect 586622 344898 586858 345134
rect 586302 309218 586538 309454
rect 586622 309218 586858 309454
rect 586302 308898 586538 309134
rect 586622 308898 586858 309134
rect 586302 273218 586538 273454
rect 586622 273218 586858 273454
rect 586302 272898 586538 273134
rect 586622 272898 586858 273134
rect 586302 237218 586538 237454
rect 586622 237218 586858 237454
rect 586302 236898 586538 237134
rect 586622 236898 586858 237134
rect 586302 201218 586538 201454
rect 586622 201218 586858 201454
rect 586302 200898 586538 201134
rect 586622 200898 586858 201134
rect 586302 165218 586538 165454
rect 586622 165218 586858 165454
rect 586302 164898 586538 165134
rect 586622 164898 586858 165134
rect 586302 129218 586538 129454
rect 586622 129218 586858 129454
rect 586302 128898 586538 129134
rect 586622 128898 586858 129134
rect 586302 93218 586538 93454
rect 586622 93218 586858 93454
rect 586302 92898 586538 93134
rect 586622 92898 586858 93134
rect 586302 57218 586538 57454
rect 586622 57218 586858 57454
rect 586302 56898 586538 57134
rect 586622 56898 586858 57134
rect 586302 21218 586538 21454
rect 586622 21218 586858 21454
rect 586302 20898 586538 21134
rect 586622 20898 586858 21134
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 690938 587498 691174
rect 587582 690938 587818 691174
rect 587262 690618 587498 690854
rect 587582 690618 587818 690854
rect 587262 654938 587498 655174
rect 587582 654938 587818 655174
rect 587262 654618 587498 654854
rect 587582 654618 587818 654854
rect 587262 618938 587498 619174
rect 587582 618938 587818 619174
rect 587262 618618 587498 618854
rect 587582 618618 587818 618854
rect 587262 582938 587498 583174
rect 587582 582938 587818 583174
rect 587262 582618 587498 582854
rect 587582 582618 587818 582854
rect 587262 546938 587498 547174
rect 587582 546938 587818 547174
rect 587262 546618 587498 546854
rect 587582 546618 587818 546854
rect 587262 510938 587498 511174
rect 587582 510938 587818 511174
rect 587262 510618 587498 510854
rect 587582 510618 587818 510854
rect 587262 474938 587498 475174
rect 587582 474938 587818 475174
rect 587262 474618 587498 474854
rect 587582 474618 587818 474854
rect 587262 438938 587498 439174
rect 587582 438938 587818 439174
rect 587262 438618 587498 438854
rect 587582 438618 587818 438854
rect 587262 402938 587498 403174
rect 587582 402938 587818 403174
rect 587262 402618 587498 402854
rect 587582 402618 587818 402854
rect 587262 366938 587498 367174
rect 587582 366938 587818 367174
rect 587262 366618 587498 366854
rect 587582 366618 587818 366854
rect 587262 330938 587498 331174
rect 587582 330938 587818 331174
rect 587262 330618 587498 330854
rect 587582 330618 587818 330854
rect 587262 294938 587498 295174
rect 587582 294938 587818 295174
rect 587262 294618 587498 294854
rect 587582 294618 587818 294854
rect 587262 258938 587498 259174
rect 587582 258938 587818 259174
rect 587262 258618 587498 258854
rect 587582 258618 587818 258854
rect 587262 222938 587498 223174
rect 587582 222938 587818 223174
rect 587262 222618 587498 222854
rect 587582 222618 587818 222854
rect 587262 186938 587498 187174
rect 587582 186938 587818 187174
rect 587262 186618 587498 186854
rect 587582 186618 587818 186854
rect 587262 150938 587498 151174
rect 587582 150938 587818 151174
rect 587262 150618 587498 150854
rect 587582 150618 587818 150854
rect 587262 114938 587498 115174
rect 587582 114938 587818 115174
rect 587262 114618 587498 114854
rect 587582 114618 587818 114854
rect 587262 78938 587498 79174
rect 587582 78938 587818 79174
rect 587262 78618 587498 78854
rect 587582 78618 587818 78854
rect 587262 42938 587498 43174
rect 587582 42938 587818 43174
rect 587262 42618 587498 42854
rect 587582 42618 587818 42854
rect 587262 6938 587498 7174
rect 587582 6938 587818 7174
rect 587262 6618 587498 6854
rect 587582 6618 587818 6854
rect 581546 -2502 581782 -2266
rect 581866 -2502 582102 -2266
rect 581546 -2822 581782 -2586
rect 581866 -2822 582102 -2586
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 672938 588458 673174
rect 588542 672938 588778 673174
rect 588222 672618 588458 672854
rect 588542 672618 588778 672854
rect 588222 636938 588458 637174
rect 588542 636938 588778 637174
rect 588222 636618 588458 636854
rect 588542 636618 588778 636854
rect 588222 600938 588458 601174
rect 588542 600938 588778 601174
rect 588222 600618 588458 600854
rect 588542 600618 588778 600854
rect 588222 564938 588458 565174
rect 588542 564938 588778 565174
rect 588222 564618 588458 564854
rect 588542 564618 588778 564854
rect 588222 528938 588458 529174
rect 588542 528938 588778 529174
rect 588222 528618 588458 528854
rect 588542 528618 588778 528854
rect 588222 492938 588458 493174
rect 588542 492938 588778 493174
rect 588222 492618 588458 492854
rect 588542 492618 588778 492854
rect 588222 456938 588458 457174
rect 588542 456938 588778 457174
rect 588222 456618 588458 456854
rect 588542 456618 588778 456854
rect 588222 420938 588458 421174
rect 588542 420938 588778 421174
rect 588222 420618 588458 420854
rect 588542 420618 588778 420854
rect 588222 384938 588458 385174
rect 588542 384938 588778 385174
rect 588222 384618 588458 384854
rect 588542 384618 588778 384854
rect 588222 348938 588458 349174
rect 588542 348938 588778 349174
rect 588222 348618 588458 348854
rect 588542 348618 588778 348854
rect 588222 312938 588458 313174
rect 588542 312938 588778 313174
rect 588222 312618 588458 312854
rect 588542 312618 588778 312854
rect 588222 276938 588458 277174
rect 588542 276938 588778 277174
rect 588222 276618 588458 276854
rect 588542 276618 588778 276854
rect 588222 240938 588458 241174
rect 588542 240938 588778 241174
rect 588222 240618 588458 240854
rect 588542 240618 588778 240854
rect 588222 204938 588458 205174
rect 588542 204938 588778 205174
rect 588222 204618 588458 204854
rect 588542 204618 588778 204854
rect 588222 168938 588458 169174
rect 588542 168938 588778 169174
rect 588222 168618 588458 168854
rect 588542 168618 588778 168854
rect 588222 132938 588458 133174
rect 588542 132938 588778 133174
rect 588222 132618 588458 132854
rect 588542 132618 588778 132854
rect 588222 96938 588458 97174
rect 588542 96938 588778 97174
rect 588222 96618 588458 96854
rect 588542 96618 588778 96854
rect 588222 60938 588458 61174
rect 588542 60938 588778 61174
rect 588222 60618 588458 60854
rect 588542 60618 588778 60854
rect 588222 24938 588458 25174
rect 588542 24938 588778 25174
rect 588222 24618 588458 24854
rect 588542 24618 588778 24854
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 694658 589418 694894
rect 589502 694658 589738 694894
rect 589182 694338 589418 694574
rect 589502 694338 589738 694574
rect 589182 658658 589418 658894
rect 589502 658658 589738 658894
rect 589182 658338 589418 658574
rect 589502 658338 589738 658574
rect 589182 622658 589418 622894
rect 589502 622658 589738 622894
rect 589182 622338 589418 622574
rect 589502 622338 589738 622574
rect 589182 586658 589418 586894
rect 589502 586658 589738 586894
rect 589182 586338 589418 586574
rect 589502 586338 589738 586574
rect 589182 550658 589418 550894
rect 589502 550658 589738 550894
rect 589182 550338 589418 550574
rect 589502 550338 589738 550574
rect 589182 514658 589418 514894
rect 589502 514658 589738 514894
rect 589182 514338 589418 514574
rect 589502 514338 589738 514574
rect 589182 478658 589418 478894
rect 589502 478658 589738 478894
rect 589182 478338 589418 478574
rect 589502 478338 589738 478574
rect 589182 442658 589418 442894
rect 589502 442658 589738 442894
rect 589182 442338 589418 442574
rect 589502 442338 589738 442574
rect 589182 406658 589418 406894
rect 589502 406658 589738 406894
rect 589182 406338 589418 406574
rect 589502 406338 589738 406574
rect 589182 370658 589418 370894
rect 589502 370658 589738 370894
rect 589182 370338 589418 370574
rect 589502 370338 589738 370574
rect 589182 334658 589418 334894
rect 589502 334658 589738 334894
rect 589182 334338 589418 334574
rect 589502 334338 589738 334574
rect 589182 298658 589418 298894
rect 589502 298658 589738 298894
rect 589182 298338 589418 298574
rect 589502 298338 589738 298574
rect 589182 262658 589418 262894
rect 589502 262658 589738 262894
rect 589182 262338 589418 262574
rect 589502 262338 589738 262574
rect 589182 226658 589418 226894
rect 589502 226658 589738 226894
rect 589182 226338 589418 226574
rect 589502 226338 589738 226574
rect 589182 190658 589418 190894
rect 589502 190658 589738 190894
rect 589182 190338 589418 190574
rect 589502 190338 589738 190574
rect 589182 154658 589418 154894
rect 589502 154658 589738 154894
rect 589182 154338 589418 154574
rect 589502 154338 589738 154574
rect 589182 118658 589418 118894
rect 589502 118658 589738 118894
rect 589182 118338 589418 118574
rect 589502 118338 589738 118574
rect 589182 82658 589418 82894
rect 589502 82658 589738 82894
rect 589182 82338 589418 82574
rect 589502 82338 589738 82574
rect 589182 46658 589418 46894
rect 589502 46658 589738 46894
rect 589182 46338 589418 46574
rect 589502 46338 589738 46574
rect 589182 10658 589418 10894
rect 589502 10658 589738 10894
rect 589182 10338 589418 10574
rect 589502 10338 589738 10574
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 676658 590378 676894
rect 590462 676658 590698 676894
rect 590142 676338 590378 676574
rect 590462 676338 590698 676574
rect 590142 640658 590378 640894
rect 590462 640658 590698 640894
rect 590142 640338 590378 640574
rect 590462 640338 590698 640574
rect 590142 604658 590378 604894
rect 590462 604658 590698 604894
rect 590142 604338 590378 604574
rect 590462 604338 590698 604574
rect 590142 568658 590378 568894
rect 590462 568658 590698 568894
rect 590142 568338 590378 568574
rect 590462 568338 590698 568574
rect 590142 532658 590378 532894
rect 590462 532658 590698 532894
rect 590142 532338 590378 532574
rect 590462 532338 590698 532574
rect 590142 496658 590378 496894
rect 590462 496658 590698 496894
rect 590142 496338 590378 496574
rect 590462 496338 590698 496574
rect 590142 460658 590378 460894
rect 590462 460658 590698 460894
rect 590142 460338 590378 460574
rect 590462 460338 590698 460574
rect 590142 424658 590378 424894
rect 590462 424658 590698 424894
rect 590142 424338 590378 424574
rect 590462 424338 590698 424574
rect 590142 388658 590378 388894
rect 590462 388658 590698 388894
rect 590142 388338 590378 388574
rect 590462 388338 590698 388574
rect 590142 352658 590378 352894
rect 590462 352658 590698 352894
rect 590142 352338 590378 352574
rect 590462 352338 590698 352574
rect 590142 316658 590378 316894
rect 590462 316658 590698 316894
rect 590142 316338 590378 316574
rect 590462 316338 590698 316574
rect 590142 280658 590378 280894
rect 590462 280658 590698 280894
rect 590142 280338 590378 280574
rect 590462 280338 590698 280574
rect 590142 244658 590378 244894
rect 590462 244658 590698 244894
rect 590142 244338 590378 244574
rect 590462 244338 590698 244574
rect 590142 208658 590378 208894
rect 590462 208658 590698 208894
rect 590142 208338 590378 208574
rect 590462 208338 590698 208574
rect 590142 172658 590378 172894
rect 590462 172658 590698 172894
rect 590142 172338 590378 172574
rect 590462 172338 590698 172574
rect 590142 136658 590378 136894
rect 590462 136658 590698 136894
rect 590142 136338 590378 136574
rect 590462 136338 590698 136574
rect 590142 100658 590378 100894
rect 590462 100658 590698 100894
rect 590142 100338 590378 100574
rect 590462 100338 590698 100574
rect 590142 64658 590378 64894
rect 590462 64658 590698 64894
rect 590142 64338 590378 64574
rect 590462 64338 590698 64574
rect 590142 28658 590378 28894
rect 590462 28658 590698 28894
rect 590142 28338 590378 28574
rect 590462 28338 590698 28574
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 698378 591338 698614
rect 591422 698378 591658 698614
rect 591102 698058 591338 698294
rect 591422 698058 591658 698294
rect 591102 662378 591338 662614
rect 591422 662378 591658 662614
rect 591102 662058 591338 662294
rect 591422 662058 591658 662294
rect 591102 626378 591338 626614
rect 591422 626378 591658 626614
rect 591102 626058 591338 626294
rect 591422 626058 591658 626294
rect 591102 590378 591338 590614
rect 591422 590378 591658 590614
rect 591102 590058 591338 590294
rect 591422 590058 591658 590294
rect 591102 554378 591338 554614
rect 591422 554378 591658 554614
rect 591102 554058 591338 554294
rect 591422 554058 591658 554294
rect 591102 518378 591338 518614
rect 591422 518378 591658 518614
rect 591102 518058 591338 518294
rect 591422 518058 591658 518294
rect 591102 482378 591338 482614
rect 591422 482378 591658 482614
rect 591102 482058 591338 482294
rect 591422 482058 591658 482294
rect 591102 446378 591338 446614
rect 591422 446378 591658 446614
rect 591102 446058 591338 446294
rect 591422 446058 591658 446294
rect 591102 410378 591338 410614
rect 591422 410378 591658 410614
rect 591102 410058 591338 410294
rect 591422 410058 591658 410294
rect 591102 374378 591338 374614
rect 591422 374378 591658 374614
rect 591102 374058 591338 374294
rect 591422 374058 591658 374294
rect 591102 338378 591338 338614
rect 591422 338378 591658 338614
rect 591102 338058 591338 338294
rect 591422 338058 591658 338294
rect 591102 302378 591338 302614
rect 591422 302378 591658 302614
rect 591102 302058 591338 302294
rect 591422 302058 591658 302294
rect 591102 266378 591338 266614
rect 591422 266378 591658 266614
rect 591102 266058 591338 266294
rect 591422 266058 591658 266294
rect 591102 230378 591338 230614
rect 591422 230378 591658 230614
rect 591102 230058 591338 230294
rect 591422 230058 591658 230294
rect 591102 194378 591338 194614
rect 591422 194378 591658 194614
rect 591102 194058 591338 194294
rect 591422 194058 591658 194294
rect 591102 158378 591338 158614
rect 591422 158378 591658 158614
rect 591102 158058 591338 158294
rect 591422 158058 591658 158294
rect 591102 122378 591338 122614
rect 591422 122378 591658 122614
rect 591102 122058 591338 122294
rect 591422 122058 591658 122294
rect 591102 86378 591338 86614
rect 591422 86378 591658 86614
rect 591102 86058 591338 86294
rect 591422 86058 591658 86294
rect 591102 50378 591338 50614
rect 591422 50378 591658 50614
rect 591102 50058 591338 50294
rect 591422 50058 591658 50294
rect 591102 14378 591338 14614
rect 591422 14378 591658 14614
rect 591102 14058 591338 14294
rect 591422 14058 591658 14294
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 680378 592298 680614
rect 592382 680378 592618 680614
rect 592062 680058 592298 680294
rect 592382 680058 592618 680294
rect 592062 644378 592298 644614
rect 592382 644378 592618 644614
rect 592062 644058 592298 644294
rect 592382 644058 592618 644294
rect 592062 608378 592298 608614
rect 592382 608378 592618 608614
rect 592062 608058 592298 608294
rect 592382 608058 592618 608294
rect 592062 572378 592298 572614
rect 592382 572378 592618 572614
rect 592062 572058 592298 572294
rect 592382 572058 592618 572294
rect 592062 536378 592298 536614
rect 592382 536378 592618 536614
rect 592062 536058 592298 536294
rect 592382 536058 592618 536294
rect 592062 500378 592298 500614
rect 592382 500378 592618 500614
rect 592062 500058 592298 500294
rect 592382 500058 592618 500294
rect 592062 464378 592298 464614
rect 592382 464378 592618 464614
rect 592062 464058 592298 464294
rect 592382 464058 592618 464294
rect 592062 428378 592298 428614
rect 592382 428378 592618 428614
rect 592062 428058 592298 428294
rect 592382 428058 592618 428294
rect 592062 392378 592298 392614
rect 592382 392378 592618 392614
rect 592062 392058 592298 392294
rect 592382 392058 592618 392294
rect 592062 356378 592298 356614
rect 592382 356378 592618 356614
rect 592062 356058 592298 356294
rect 592382 356058 592618 356294
rect 592062 320378 592298 320614
rect 592382 320378 592618 320614
rect 592062 320058 592298 320294
rect 592382 320058 592618 320294
rect 592062 284378 592298 284614
rect 592382 284378 592618 284614
rect 592062 284058 592298 284294
rect 592382 284058 592618 284294
rect 592062 248378 592298 248614
rect 592382 248378 592618 248614
rect 592062 248058 592298 248294
rect 592382 248058 592618 248294
rect 592062 212378 592298 212614
rect 592382 212378 592618 212614
rect 592062 212058 592298 212294
rect 592382 212058 592618 212294
rect 592062 176378 592298 176614
rect 592382 176378 592618 176614
rect 592062 176058 592298 176294
rect 592382 176058 592618 176294
rect 592062 140378 592298 140614
rect 592382 140378 592618 140614
rect 592062 140058 592298 140294
rect 592382 140058 592618 140294
rect 592062 104378 592298 104614
rect 592382 104378 592618 104614
rect 592062 104058 592298 104294
rect 592382 104058 592618 104294
rect 592062 68378 592298 68614
rect 592382 68378 592618 68614
rect 592062 68058 592298 68294
rect 592382 68058 592618 68294
rect 592062 32378 592298 32614
rect 592382 32378 592618 32614
rect 592062 32058 592298 32294
rect 592382 32058 592618 32294
rect 570986 -7302 571222 -7066
rect 571306 -7302 571542 -7066
rect 570986 -7622 571222 -7386
rect 571306 -7622 571542 -7386
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 592650 698614
rect -8726 698294 592650 698378
rect -8726 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 592650 698294
rect -8726 698026 592650 698058
rect -6806 694894 590730 694926
rect -6806 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 590730 694894
rect -6806 694574 590730 694658
rect -6806 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 590730 694574
rect -6806 694306 590730 694338
rect -4886 691174 588810 691206
rect -4886 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 588810 691174
rect -4886 690854 588810 690938
rect -4886 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 588810 690854
rect -4886 690586 588810 690618
rect -2966 687454 586890 687486
rect -2966 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 586890 687454
rect -2966 687134 586890 687218
rect -2966 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 586890 687134
rect -2966 686866 586890 686898
rect -8726 680614 592650 680646
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect -8726 680294 592650 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect -8726 680026 592650 680058
rect -6806 676894 590730 676926
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect -6806 676574 590730 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect -6806 676306 590730 676338
rect -4886 673174 588810 673206
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect -4886 672854 588810 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect -4886 672586 588810 672618
rect -2966 669454 586890 669486
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect -2966 669134 586890 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect -2966 668866 586890 668898
rect -8726 662614 592650 662646
rect -8726 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 592650 662614
rect -8726 662294 592650 662378
rect -8726 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 592650 662294
rect -8726 662026 592650 662058
rect -6806 658894 590730 658926
rect -6806 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 590730 658894
rect -6806 658574 590730 658658
rect -6806 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 590730 658574
rect -6806 658306 590730 658338
rect -4886 655174 588810 655206
rect -4886 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 588810 655174
rect -4886 654854 588810 654938
rect -4886 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 588810 654854
rect -4886 654586 588810 654618
rect -2966 651454 586890 651486
rect -2966 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 586890 651454
rect -2966 651134 586890 651218
rect -2966 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 586890 651134
rect -2966 650866 586890 650898
rect -8726 644614 592650 644646
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect -8726 644294 592650 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect -8726 644026 592650 644058
rect -6806 640894 590730 640926
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect -6806 640574 590730 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect -6806 640306 590730 640338
rect -4886 637174 588810 637206
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect -4886 636854 588810 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect -4886 636586 588810 636618
rect -2966 633454 586890 633486
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect -2966 633134 586890 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect -2966 632866 586890 632898
rect -8726 626614 592650 626646
rect -8726 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 592650 626614
rect -8726 626294 592650 626378
rect -8726 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 592650 626294
rect -8726 626026 592650 626058
rect -6806 622894 590730 622926
rect -6806 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 590730 622894
rect -6806 622574 590730 622658
rect -6806 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 590730 622574
rect -6806 622306 590730 622338
rect -4886 619174 588810 619206
rect -4886 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 588810 619174
rect -4886 618854 588810 618938
rect -4886 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 588810 618854
rect -4886 618586 588810 618618
rect -2966 615454 586890 615486
rect -2966 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 586890 615454
rect -2966 615134 586890 615218
rect -2966 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 586890 615134
rect -2966 614866 586890 614898
rect -8726 608614 592650 608646
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect -8726 608294 592650 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect -8726 608026 592650 608058
rect -6806 604894 590730 604926
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect -6806 604574 590730 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect -6806 604306 590730 604338
rect -4886 601174 588810 601206
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect -4886 600854 588810 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect -4886 600586 588810 600618
rect -2966 597454 586890 597486
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect -2966 597134 586890 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect -2966 596866 586890 596898
rect -8726 590614 592650 590646
rect -8726 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 592650 590614
rect -8726 590294 592650 590378
rect -8726 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 592650 590294
rect -8726 590026 592650 590058
rect -6806 586894 590730 586926
rect -6806 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 590730 586894
rect -6806 586574 590730 586658
rect -6806 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 590730 586574
rect -6806 586306 590730 586338
rect -4886 583174 588810 583206
rect -4886 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 588810 583174
rect -4886 582854 588810 582938
rect -4886 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 588810 582854
rect -4886 582586 588810 582618
rect -2966 579454 586890 579486
rect -2966 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 72721 579454
rect 72957 579218 78651 579454
rect 78887 579218 84582 579454
rect 84818 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 586890 579454
rect -2966 579134 586890 579218
rect -2966 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 72721 579134
rect 72957 578898 78651 579134
rect 78887 578898 84582 579134
rect 84818 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 586890 579134
rect -2966 578866 586890 578898
rect -8726 572614 592650 572646
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect -8726 572294 592650 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect -8726 572026 592650 572058
rect -6806 568894 590730 568926
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect -6806 568574 590730 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect -6806 568306 590730 568338
rect -4886 565174 588810 565206
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 95546 565174
rect 95782 564938 95866 565174
rect 96102 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 419546 565174
rect 419782 564938 419866 565174
rect 420102 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect -4886 564854 588810 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 95546 564854
rect 95782 564618 95866 564854
rect 96102 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 419546 564854
rect 419782 564618 419866 564854
rect 420102 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect -4886 564586 588810 564618
rect -2966 561454 586890 561486
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 75686 561454
rect 75922 561218 81617 561454
rect 81853 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect -2966 561134 586890 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 75686 561134
rect 75922 560898 81617 561134
rect 81853 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect -2966 560866 586890 560898
rect -8726 554614 592650 554646
rect -8726 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 592650 554614
rect -8726 554294 592650 554378
rect -8726 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 592650 554294
rect -8726 554026 592650 554058
rect -6806 550894 590730 550926
rect -6806 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 590730 550894
rect -6806 550574 590730 550658
rect -6806 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 590730 550574
rect -6806 550306 590730 550338
rect -4886 547174 588810 547206
rect -4886 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 588810 547174
rect -4886 546854 588810 546938
rect -4886 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 588810 546854
rect -4886 546586 588810 546618
rect -2966 543454 586890 543486
rect -2966 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 72721 543454
rect 72957 543218 78651 543454
rect 78887 543218 84582 543454
rect 84818 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 586890 543454
rect -2966 543134 586890 543218
rect -2966 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 72721 543134
rect 72957 542898 78651 543134
rect 78887 542898 84582 543134
rect 84818 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 586890 543134
rect -2966 542866 586890 542898
rect -8726 536614 592650 536646
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 102986 536614
rect 103222 536378 103306 536614
rect 103542 536378 138986 536614
rect 139222 536378 139306 536614
rect 139542 536378 174986 536614
rect 175222 536378 175306 536614
rect 175542 536378 390986 536614
rect 391222 536378 391306 536614
rect 391542 536378 426986 536614
rect 427222 536378 427306 536614
rect 427542 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect -8726 536294 592650 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 102986 536294
rect 103222 536058 103306 536294
rect 103542 536058 138986 536294
rect 139222 536058 139306 536294
rect 139542 536058 174986 536294
rect 175222 536058 175306 536294
rect 175542 536058 390986 536294
rect 391222 536058 391306 536294
rect 391542 536058 426986 536294
rect 427222 536058 427306 536294
rect 427542 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect -8726 536026 592650 536058
rect -6806 532894 590730 532926
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 99266 532894
rect 99502 532658 99586 532894
rect 99822 532658 135266 532894
rect 135502 532658 135586 532894
rect 135822 532658 171266 532894
rect 171502 532658 171586 532894
rect 171822 532658 387266 532894
rect 387502 532658 387586 532894
rect 387822 532658 423266 532894
rect 423502 532658 423586 532894
rect 423822 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect -6806 532574 590730 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 99266 532574
rect 99502 532338 99586 532574
rect 99822 532338 135266 532574
rect 135502 532338 135586 532574
rect 135822 532338 171266 532574
rect 171502 532338 171586 532574
rect 171822 532338 387266 532574
rect 387502 532338 387586 532574
rect 387822 532338 423266 532574
rect 423502 532338 423586 532574
rect 423822 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect -6806 532306 590730 532338
rect -4886 529174 588810 529206
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 95546 529174
rect 95782 528938 95866 529174
rect 96102 528938 131546 529174
rect 131782 528938 131866 529174
rect 132102 528938 167546 529174
rect 167782 528938 167866 529174
rect 168102 528938 383546 529174
rect 383782 528938 383866 529174
rect 384102 528938 419546 529174
rect 419782 528938 419866 529174
rect 420102 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect -4886 528854 588810 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 95546 528854
rect 95782 528618 95866 528854
rect 96102 528618 131546 528854
rect 131782 528618 131866 528854
rect 132102 528618 167546 528854
rect 167782 528618 167866 528854
rect 168102 528618 383546 528854
rect 383782 528618 383866 528854
rect 384102 528618 419546 528854
rect 419782 528618 419866 528854
rect 420102 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect -4886 528586 588810 528618
rect -2966 525454 586890 525486
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 219610 525454
rect 219846 525218 250330 525454
rect 250566 525218 281050 525454
rect 281286 525218 311770 525454
rect 312006 525218 342490 525454
rect 342726 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect -2966 525134 586890 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 219610 525134
rect 219846 524898 250330 525134
rect 250566 524898 281050 525134
rect 281286 524898 311770 525134
rect 312006 524898 342490 525134
rect 342726 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect -2966 524866 586890 524898
rect -8726 518614 592650 518646
rect -8726 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 592650 518614
rect -8726 518294 592650 518378
rect -8726 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 592650 518294
rect -8726 518026 592650 518058
rect -6806 514894 590730 514926
rect -6806 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 590730 514894
rect -6806 514574 590730 514658
rect -6806 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 590730 514574
rect -6806 514306 590730 514338
rect -4886 511174 588810 511206
rect -4886 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 588810 511174
rect -4886 510854 588810 510938
rect -4886 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 588810 510854
rect -4886 510586 588810 510618
rect -2966 507454 586890 507486
rect -2966 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 204250 507454
rect 204486 507218 234970 507454
rect 235206 507218 265690 507454
rect 265926 507218 296410 507454
rect 296646 507218 327130 507454
rect 327366 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 586890 507454
rect -2966 507134 586890 507218
rect -2966 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 204250 507134
rect 204486 506898 234970 507134
rect 235206 506898 265690 507134
rect 265926 506898 296410 507134
rect 296646 506898 327130 507134
rect 327366 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 586890 507134
rect -2966 506866 586890 506898
rect -8726 500614 592650 500646
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 102986 500614
rect 103222 500378 103306 500614
rect 103542 500378 138986 500614
rect 139222 500378 139306 500614
rect 139542 500378 174986 500614
rect 175222 500378 175306 500614
rect 175542 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect -8726 500294 592650 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 102986 500294
rect 103222 500058 103306 500294
rect 103542 500058 138986 500294
rect 139222 500058 139306 500294
rect 139542 500058 174986 500294
rect 175222 500058 175306 500294
rect 175542 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect -8726 500026 592650 500058
rect -6806 496894 590730 496926
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 99266 496894
rect 99502 496658 99586 496894
rect 99822 496658 135266 496894
rect 135502 496658 135586 496894
rect 135822 496658 171266 496894
rect 171502 496658 171586 496894
rect 171822 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect -6806 496574 590730 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 99266 496574
rect 99502 496338 99586 496574
rect 99822 496338 135266 496574
rect 135502 496338 135586 496574
rect 135822 496338 171266 496574
rect 171502 496338 171586 496574
rect 171822 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect -6806 496306 590730 496338
rect -4886 493174 588810 493206
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 95546 493174
rect 95782 492938 95866 493174
rect 96102 492938 131546 493174
rect 131782 492938 131866 493174
rect 132102 492938 167546 493174
rect 167782 492938 167866 493174
rect 168102 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect -4886 492854 588810 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 95546 492854
rect 95782 492618 95866 492854
rect 96102 492618 131546 492854
rect 131782 492618 131866 492854
rect 132102 492618 167546 492854
rect 167782 492618 167866 492854
rect 168102 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect -4886 492586 588810 492618
rect -2966 489454 586890 489486
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 219610 489454
rect 219846 489218 250330 489454
rect 250566 489218 281050 489454
rect 281286 489218 311770 489454
rect 312006 489218 342490 489454
rect 342726 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect -2966 489134 586890 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 219610 489134
rect 219846 488898 250330 489134
rect 250566 488898 281050 489134
rect 281286 488898 311770 489134
rect 312006 488898 342490 489134
rect 342726 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect -2966 488866 586890 488898
rect -8726 482614 592650 482646
rect -8726 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 592650 482614
rect -8726 482294 592650 482378
rect -8726 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 592650 482294
rect -8726 482026 592650 482058
rect -6806 478894 590730 478926
rect -6806 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 590730 478894
rect -6806 478574 590730 478658
rect -6806 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 590730 478574
rect -6806 478306 590730 478338
rect -4886 475174 588810 475206
rect -4886 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 588810 475174
rect -4886 474854 588810 474938
rect -4886 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 588810 474854
rect -4886 474586 588810 474618
rect -2966 471454 586890 471486
rect -2966 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 204250 471454
rect 204486 471218 234970 471454
rect 235206 471218 265690 471454
rect 265926 471218 296410 471454
rect 296646 471218 327130 471454
rect 327366 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 586890 471454
rect -2966 471134 586890 471218
rect -2966 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 204250 471134
rect 204486 470898 234970 471134
rect 235206 470898 265690 471134
rect 265926 470898 296410 471134
rect 296646 470898 327130 471134
rect 327366 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 586890 471134
rect -2966 470866 586890 470898
rect -8726 464614 592650 464646
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 66986 464614
rect 67222 464378 67306 464614
rect 67542 464378 102986 464614
rect 103222 464378 103306 464614
rect 103542 464378 138986 464614
rect 139222 464378 139306 464614
rect 139542 464378 174986 464614
rect 175222 464378 175306 464614
rect 175542 464378 390986 464614
rect 391222 464378 391306 464614
rect 391542 464378 426986 464614
rect 427222 464378 427306 464614
rect 427542 464378 462986 464614
rect 463222 464378 463306 464614
rect 463542 464378 498986 464614
rect 499222 464378 499306 464614
rect 499542 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect -8726 464294 592650 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 66986 464294
rect 67222 464058 67306 464294
rect 67542 464058 102986 464294
rect 103222 464058 103306 464294
rect 103542 464058 138986 464294
rect 139222 464058 139306 464294
rect 139542 464058 174986 464294
rect 175222 464058 175306 464294
rect 175542 464058 390986 464294
rect 391222 464058 391306 464294
rect 391542 464058 426986 464294
rect 427222 464058 427306 464294
rect 427542 464058 462986 464294
rect 463222 464058 463306 464294
rect 463542 464058 498986 464294
rect 499222 464058 499306 464294
rect 499542 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect -8726 464026 592650 464058
rect -6806 460894 590730 460926
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 63266 460894
rect 63502 460658 63586 460894
rect 63822 460658 99266 460894
rect 99502 460658 99586 460894
rect 99822 460658 135266 460894
rect 135502 460658 135586 460894
rect 135822 460658 171266 460894
rect 171502 460658 171586 460894
rect 171822 460658 387266 460894
rect 387502 460658 387586 460894
rect 387822 460658 423266 460894
rect 423502 460658 423586 460894
rect 423822 460658 459266 460894
rect 459502 460658 459586 460894
rect 459822 460658 495266 460894
rect 495502 460658 495586 460894
rect 495822 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect -6806 460574 590730 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 63266 460574
rect 63502 460338 63586 460574
rect 63822 460338 99266 460574
rect 99502 460338 99586 460574
rect 99822 460338 135266 460574
rect 135502 460338 135586 460574
rect 135822 460338 171266 460574
rect 171502 460338 171586 460574
rect 171822 460338 387266 460574
rect 387502 460338 387586 460574
rect 387822 460338 423266 460574
rect 423502 460338 423586 460574
rect 423822 460338 459266 460574
rect 459502 460338 459586 460574
rect 459822 460338 495266 460574
rect 495502 460338 495586 460574
rect 495822 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect -6806 460306 590730 460338
rect -4886 457174 588810 457206
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 59546 457174
rect 59782 456938 59866 457174
rect 60102 456938 95546 457174
rect 95782 456938 95866 457174
rect 96102 456938 131546 457174
rect 131782 456938 131866 457174
rect 132102 456938 167546 457174
rect 167782 456938 167866 457174
rect 168102 456938 383546 457174
rect 383782 456938 383866 457174
rect 384102 456938 419546 457174
rect 419782 456938 419866 457174
rect 420102 456938 455546 457174
rect 455782 456938 455866 457174
rect 456102 456938 491546 457174
rect 491782 456938 491866 457174
rect 492102 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect -4886 456854 588810 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 59546 456854
rect 59782 456618 59866 456854
rect 60102 456618 95546 456854
rect 95782 456618 95866 456854
rect 96102 456618 131546 456854
rect 131782 456618 131866 456854
rect 132102 456618 167546 456854
rect 167782 456618 167866 456854
rect 168102 456618 383546 456854
rect 383782 456618 383866 456854
rect 384102 456618 419546 456854
rect 419782 456618 419866 456854
rect 420102 456618 455546 456854
rect 455782 456618 455866 456854
rect 456102 456618 491546 456854
rect 491782 456618 491866 456854
rect 492102 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect -4886 456586 588810 456618
rect -2966 453454 586890 453486
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 219610 453454
rect 219846 453218 250330 453454
rect 250566 453218 281050 453454
rect 281286 453218 311770 453454
rect 312006 453218 342490 453454
rect 342726 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect -2966 453134 586890 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 219610 453134
rect 219846 452898 250330 453134
rect 250566 452898 281050 453134
rect 281286 452898 311770 453134
rect 312006 452898 342490 453134
rect 342726 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect -2966 452866 586890 452898
rect -8726 446614 592650 446646
rect -8726 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 156986 446614
rect 157222 446378 157306 446614
rect 157542 446378 192986 446614
rect 193222 446378 193306 446614
rect 193542 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 592650 446614
rect -8726 446294 592650 446378
rect -8726 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 156986 446294
rect 157222 446058 157306 446294
rect 157542 446058 192986 446294
rect 193222 446058 193306 446294
rect 193542 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 592650 446294
rect -8726 446026 592650 446058
rect -6806 442894 590730 442926
rect -6806 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 153266 442894
rect 153502 442658 153586 442894
rect 153822 442658 189266 442894
rect 189502 442658 189586 442894
rect 189822 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 441266 442894
rect 441502 442658 441586 442894
rect 441822 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 590730 442894
rect -6806 442574 590730 442658
rect -6806 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 153266 442574
rect 153502 442338 153586 442574
rect 153822 442338 189266 442574
rect 189502 442338 189586 442574
rect 189822 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 441266 442574
rect 441502 442338 441586 442574
rect 441822 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 590730 442574
rect -6806 442306 590730 442338
rect -4886 439174 588810 439206
rect -4886 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 149546 439174
rect 149782 438938 149866 439174
rect 150102 438938 185546 439174
rect 185782 438938 185866 439174
rect 186102 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 437546 439174
rect 437782 438938 437866 439174
rect 438102 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 588810 439174
rect -4886 438854 588810 438938
rect -4886 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 149546 438854
rect 149782 438618 149866 438854
rect 150102 438618 185546 438854
rect 185782 438618 185866 438854
rect 186102 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 437546 438854
rect 437782 438618 437866 438854
rect 438102 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 588810 438854
rect -4886 438586 588810 438618
rect -2966 435454 586890 435486
rect -2966 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 73020 435454
rect 73256 435218 103740 435454
rect 103976 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 204250 435454
rect 204486 435218 234970 435454
rect 235206 435218 265690 435454
rect 265926 435218 296410 435454
rect 296646 435218 327130 435454
rect 327366 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 586890 435454
rect -2966 435134 586890 435218
rect -2966 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 73020 435134
rect 73256 434898 103740 435134
rect 103976 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 204250 435134
rect 204486 434898 234970 435134
rect 235206 434898 265690 435134
rect 265926 434898 296410 435134
rect 296646 434898 327130 435134
rect 327366 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 586890 435134
rect -2966 434866 586890 434898
rect -8726 428614 592650 428646
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 138986 428614
rect 139222 428378 139306 428614
rect 139542 428378 174986 428614
rect 175222 428378 175306 428614
rect 175542 428378 390986 428614
rect 391222 428378 391306 428614
rect 391542 428378 426986 428614
rect 427222 428378 427306 428614
rect 427542 428378 462986 428614
rect 463222 428378 463306 428614
rect 463542 428378 498986 428614
rect 499222 428378 499306 428614
rect 499542 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect -8726 428294 592650 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 138986 428294
rect 139222 428058 139306 428294
rect 139542 428058 174986 428294
rect 175222 428058 175306 428294
rect 175542 428058 390986 428294
rect 391222 428058 391306 428294
rect 391542 428058 426986 428294
rect 427222 428058 427306 428294
rect 427542 428058 462986 428294
rect 463222 428058 463306 428294
rect 463542 428058 498986 428294
rect 499222 428058 499306 428294
rect 499542 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect -8726 428026 592650 428058
rect -6806 424894 590730 424926
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 63266 424894
rect 63502 424658 63586 424894
rect 63822 424658 135266 424894
rect 135502 424658 135586 424894
rect 135822 424658 171266 424894
rect 171502 424658 171586 424894
rect 171822 424658 387266 424894
rect 387502 424658 387586 424894
rect 387822 424658 423266 424894
rect 423502 424658 423586 424894
rect 423822 424658 459266 424894
rect 459502 424658 459586 424894
rect 459822 424658 495266 424894
rect 495502 424658 495586 424894
rect 495822 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect -6806 424574 590730 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 63266 424574
rect 63502 424338 63586 424574
rect 63822 424338 135266 424574
rect 135502 424338 135586 424574
rect 135822 424338 171266 424574
rect 171502 424338 171586 424574
rect 171822 424338 387266 424574
rect 387502 424338 387586 424574
rect 387822 424338 423266 424574
rect 423502 424338 423586 424574
rect 423822 424338 459266 424574
rect 459502 424338 459586 424574
rect 459822 424338 495266 424574
rect 495502 424338 495586 424574
rect 495822 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect -6806 424306 590730 424338
rect -4886 421174 588810 421206
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 59546 421174
rect 59782 420938 59866 421174
rect 60102 420938 131546 421174
rect 131782 420938 131866 421174
rect 132102 420938 167546 421174
rect 167782 420938 167866 421174
rect 168102 420938 383546 421174
rect 383782 420938 383866 421174
rect 384102 420938 419546 421174
rect 419782 420938 419866 421174
rect 420102 420938 455546 421174
rect 455782 420938 455866 421174
rect 456102 420938 491546 421174
rect 491782 420938 491866 421174
rect 492102 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect -4886 420854 588810 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 59546 420854
rect 59782 420618 59866 420854
rect 60102 420618 131546 420854
rect 131782 420618 131866 420854
rect 132102 420618 167546 420854
rect 167782 420618 167866 420854
rect 168102 420618 383546 420854
rect 383782 420618 383866 420854
rect 384102 420618 419546 420854
rect 419782 420618 419866 420854
rect 420102 420618 455546 420854
rect 455782 420618 455866 420854
rect 456102 420618 491546 420854
rect 491782 420618 491866 420854
rect 492102 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect -4886 420586 588810 420618
rect -2966 417454 586890 417486
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 88380 417454
rect 88616 417218 119100 417454
rect 119336 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 219610 417454
rect 219846 417218 250330 417454
rect 250566 417218 281050 417454
rect 281286 417218 311770 417454
rect 312006 417218 342490 417454
rect 342726 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect -2966 417134 586890 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 88380 417134
rect 88616 416898 119100 417134
rect 119336 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 219610 417134
rect 219846 416898 250330 417134
rect 250566 416898 281050 417134
rect 281286 416898 311770 417134
rect 312006 416898 342490 417134
rect 342726 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect -2966 416866 586890 416898
rect -8726 410614 592650 410646
rect -8726 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 156986 410614
rect 157222 410378 157306 410614
rect 157542 410378 192986 410614
rect 193222 410378 193306 410614
rect 193542 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 408986 410614
rect 409222 410378 409306 410614
rect 409542 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 592650 410614
rect -8726 410294 592650 410378
rect -8726 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 156986 410294
rect 157222 410058 157306 410294
rect 157542 410058 192986 410294
rect 193222 410058 193306 410294
rect 193542 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 408986 410294
rect 409222 410058 409306 410294
rect 409542 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 592650 410294
rect -8726 410026 592650 410058
rect -6806 406894 590730 406926
rect -6806 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 153266 406894
rect 153502 406658 153586 406894
rect 153822 406658 189266 406894
rect 189502 406658 189586 406894
rect 189822 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 405266 406894
rect 405502 406658 405586 406894
rect 405822 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 590730 406894
rect -6806 406574 590730 406658
rect -6806 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 153266 406574
rect 153502 406338 153586 406574
rect 153822 406338 189266 406574
rect 189502 406338 189586 406574
rect 189822 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 405266 406574
rect 405502 406338 405586 406574
rect 405822 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 590730 406574
rect -6806 406306 590730 406338
rect -4886 403174 588810 403206
rect -4886 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 149546 403174
rect 149782 402938 149866 403174
rect 150102 402938 185546 403174
rect 185782 402938 185866 403174
rect 186102 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 588810 403174
rect -4886 402854 588810 402938
rect -4886 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 149546 402854
rect 149782 402618 149866 402854
rect 150102 402618 185546 402854
rect 185782 402618 185866 402854
rect 186102 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 588810 402854
rect -4886 402586 588810 402618
rect -2966 399454 586890 399486
rect -2966 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 73020 399454
rect 73256 399218 103740 399454
rect 103976 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 204250 399454
rect 204486 399218 234970 399454
rect 235206 399218 265690 399454
rect 265926 399218 296410 399454
rect 296646 399218 327130 399454
rect 327366 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 586890 399454
rect -2966 399134 586890 399218
rect -2966 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 73020 399134
rect 73256 398898 103740 399134
rect 103976 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 204250 399134
rect 204486 398898 234970 399134
rect 235206 398898 265690 399134
rect 265926 398898 296410 399134
rect 296646 398898 327130 399134
rect 327366 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 586890 399134
rect -2966 398866 586890 398898
rect -8726 392614 592650 392646
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 138986 392614
rect 139222 392378 139306 392614
rect 139542 392378 174986 392614
rect 175222 392378 175306 392614
rect 175542 392378 390986 392614
rect 391222 392378 391306 392614
rect 391542 392378 426986 392614
rect 427222 392378 427306 392614
rect 427542 392378 462986 392614
rect 463222 392378 463306 392614
rect 463542 392378 498986 392614
rect 499222 392378 499306 392614
rect 499542 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect -8726 392294 592650 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 138986 392294
rect 139222 392058 139306 392294
rect 139542 392058 174986 392294
rect 175222 392058 175306 392294
rect 175542 392058 390986 392294
rect 391222 392058 391306 392294
rect 391542 392058 426986 392294
rect 427222 392058 427306 392294
rect 427542 392058 462986 392294
rect 463222 392058 463306 392294
rect 463542 392058 498986 392294
rect 499222 392058 499306 392294
rect 499542 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect -8726 392026 592650 392058
rect -6806 388894 590730 388926
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 63266 388894
rect 63502 388658 63586 388894
rect 63822 388658 135266 388894
rect 135502 388658 135586 388894
rect 135822 388658 171266 388894
rect 171502 388658 171586 388894
rect 171822 388658 387266 388894
rect 387502 388658 387586 388894
rect 387822 388658 423266 388894
rect 423502 388658 423586 388894
rect 423822 388658 459266 388894
rect 459502 388658 459586 388894
rect 459822 388658 495266 388894
rect 495502 388658 495586 388894
rect 495822 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect -6806 388574 590730 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 63266 388574
rect 63502 388338 63586 388574
rect 63822 388338 135266 388574
rect 135502 388338 135586 388574
rect 135822 388338 171266 388574
rect 171502 388338 171586 388574
rect 171822 388338 387266 388574
rect 387502 388338 387586 388574
rect 387822 388338 423266 388574
rect 423502 388338 423586 388574
rect 423822 388338 459266 388574
rect 459502 388338 459586 388574
rect 459822 388338 495266 388574
rect 495502 388338 495586 388574
rect 495822 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect -6806 388306 590730 388338
rect -4886 385174 588810 385206
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 59546 385174
rect 59782 384938 59866 385174
rect 60102 384938 95546 385174
rect 95782 384938 95866 385174
rect 96102 384938 131546 385174
rect 131782 384938 131866 385174
rect 132102 384938 167546 385174
rect 167782 384938 167866 385174
rect 168102 384938 383546 385174
rect 383782 384938 383866 385174
rect 384102 384938 419546 385174
rect 419782 384938 419866 385174
rect 420102 384938 455546 385174
rect 455782 384938 455866 385174
rect 456102 384938 491546 385174
rect 491782 384938 491866 385174
rect 492102 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect -4886 384854 588810 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 59546 384854
rect 59782 384618 59866 384854
rect 60102 384618 95546 384854
rect 95782 384618 95866 384854
rect 96102 384618 131546 384854
rect 131782 384618 131866 384854
rect 132102 384618 167546 384854
rect 167782 384618 167866 384854
rect 168102 384618 383546 384854
rect 383782 384618 383866 384854
rect 384102 384618 419546 384854
rect 419782 384618 419866 384854
rect 420102 384618 455546 384854
rect 455782 384618 455866 384854
rect 456102 384618 491546 384854
rect 491782 384618 491866 384854
rect 492102 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect -4886 384586 588810 384618
rect -2966 381454 586890 381486
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 219610 381454
rect 219846 381218 250330 381454
rect 250566 381218 281050 381454
rect 281286 381218 311770 381454
rect 312006 381218 342490 381454
rect 342726 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect -2966 381134 586890 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 219610 381134
rect 219846 380898 250330 381134
rect 250566 380898 281050 381134
rect 281286 380898 311770 381134
rect 312006 380898 342490 381134
rect 342726 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect -2966 380866 586890 380898
rect -8726 374614 592650 374646
rect -8726 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 84986 374614
rect 85222 374378 85306 374614
rect 85542 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 228986 374614
rect 229222 374378 229306 374614
rect 229542 374378 264986 374614
rect 265222 374378 265306 374614
rect 265542 374378 300986 374614
rect 301222 374378 301306 374614
rect 301542 374378 336986 374614
rect 337222 374378 337306 374614
rect 337542 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 592650 374614
rect -8726 374294 592650 374378
rect -8726 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 84986 374294
rect 85222 374058 85306 374294
rect 85542 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 228986 374294
rect 229222 374058 229306 374294
rect 229542 374058 264986 374294
rect 265222 374058 265306 374294
rect 265542 374058 300986 374294
rect 301222 374058 301306 374294
rect 301542 374058 336986 374294
rect 337222 374058 337306 374294
rect 337542 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 592650 374294
rect -8726 374026 592650 374058
rect -6806 370894 590730 370926
rect -6806 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 81266 370894
rect 81502 370658 81586 370894
rect 81822 370658 117266 370894
rect 117502 370658 117586 370894
rect 117822 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 225266 370894
rect 225502 370658 225586 370894
rect 225822 370658 261266 370894
rect 261502 370658 261586 370894
rect 261822 370658 297266 370894
rect 297502 370658 297586 370894
rect 297822 370658 333266 370894
rect 333502 370658 333586 370894
rect 333822 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 590730 370894
rect -6806 370574 590730 370658
rect -6806 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 81266 370574
rect 81502 370338 81586 370574
rect 81822 370338 117266 370574
rect 117502 370338 117586 370574
rect 117822 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 225266 370574
rect 225502 370338 225586 370574
rect 225822 370338 261266 370574
rect 261502 370338 261586 370574
rect 261822 370338 297266 370574
rect 297502 370338 297586 370574
rect 297822 370338 333266 370574
rect 333502 370338 333586 370574
rect 333822 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 590730 370574
rect -6806 370306 590730 370338
rect -4886 367174 588810 367206
rect -4886 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 77546 367174
rect 77782 366938 77866 367174
rect 78102 366938 113546 367174
rect 113782 366938 113866 367174
rect 114102 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 257546 367174
rect 257782 366938 257866 367174
rect 258102 366938 293546 367174
rect 293782 366938 293866 367174
rect 294102 366938 329546 367174
rect 329782 366938 329866 367174
rect 330102 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 588810 367174
rect -4886 366854 588810 366938
rect -4886 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 77546 366854
rect 77782 366618 77866 366854
rect 78102 366618 113546 366854
rect 113782 366618 113866 366854
rect 114102 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 257546 366854
rect 257782 366618 257866 366854
rect 258102 366618 293546 366854
rect 293782 366618 293866 366854
rect 294102 366618 329546 366854
rect 329782 366618 329866 366854
rect 330102 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 588810 366854
rect -4886 366586 588810 366618
rect -2966 363454 586890 363486
rect -2966 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 586890 363454
rect -2966 363134 586890 363218
rect -2966 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 586890 363134
rect -2966 362866 586890 362898
rect -8726 356614 592650 356646
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 66986 356614
rect 67222 356378 67306 356614
rect 67542 356378 102986 356614
rect 103222 356378 103306 356614
rect 103542 356378 138986 356614
rect 139222 356378 139306 356614
rect 139542 356378 174986 356614
rect 175222 356378 175306 356614
rect 175542 356378 210986 356614
rect 211222 356378 211306 356614
rect 211542 356378 246986 356614
rect 247222 356378 247306 356614
rect 247542 356378 282986 356614
rect 283222 356378 283306 356614
rect 283542 356378 318986 356614
rect 319222 356378 319306 356614
rect 319542 356378 354986 356614
rect 355222 356378 355306 356614
rect 355542 356378 390986 356614
rect 391222 356378 391306 356614
rect 391542 356378 426986 356614
rect 427222 356378 427306 356614
rect 427542 356378 462986 356614
rect 463222 356378 463306 356614
rect 463542 356378 498986 356614
rect 499222 356378 499306 356614
rect 499542 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect -8726 356294 592650 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 66986 356294
rect 67222 356058 67306 356294
rect 67542 356058 102986 356294
rect 103222 356058 103306 356294
rect 103542 356058 138986 356294
rect 139222 356058 139306 356294
rect 139542 356058 174986 356294
rect 175222 356058 175306 356294
rect 175542 356058 210986 356294
rect 211222 356058 211306 356294
rect 211542 356058 246986 356294
rect 247222 356058 247306 356294
rect 247542 356058 282986 356294
rect 283222 356058 283306 356294
rect 283542 356058 318986 356294
rect 319222 356058 319306 356294
rect 319542 356058 354986 356294
rect 355222 356058 355306 356294
rect 355542 356058 390986 356294
rect 391222 356058 391306 356294
rect 391542 356058 426986 356294
rect 427222 356058 427306 356294
rect 427542 356058 462986 356294
rect 463222 356058 463306 356294
rect 463542 356058 498986 356294
rect 499222 356058 499306 356294
rect 499542 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect -8726 356026 592650 356058
rect -6806 352894 590730 352926
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 63266 352894
rect 63502 352658 63586 352894
rect 63822 352658 99266 352894
rect 99502 352658 99586 352894
rect 99822 352658 135266 352894
rect 135502 352658 135586 352894
rect 135822 352658 171266 352894
rect 171502 352658 171586 352894
rect 171822 352658 207266 352894
rect 207502 352658 207586 352894
rect 207822 352658 243266 352894
rect 243502 352658 243586 352894
rect 243822 352658 279266 352894
rect 279502 352658 279586 352894
rect 279822 352658 315266 352894
rect 315502 352658 315586 352894
rect 315822 352658 351266 352894
rect 351502 352658 351586 352894
rect 351822 352658 387266 352894
rect 387502 352658 387586 352894
rect 387822 352658 423266 352894
rect 423502 352658 423586 352894
rect 423822 352658 459266 352894
rect 459502 352658 459586 352894
rect 459822 352658 495266 352894
rect 495502 352658 495586 352894
rect 495822 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect -6806 352574 590730 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 63266 352574
rect 63502 352338 63586 352574
rect 63822 352338 99266 352574
rect 99502 352338 99586 352574
rect 99822 352338 135266 352574
rect 135502 352338 135586 352574
rect 135822 352338 171266 352574
rect 171502 352338 171586 352574
rect 171822 352338 207266 352574
rect 207502 352338 207586 352574
rect 207822 352338 243266 352574
rect 243502 352338 243586 352574
rect 243822 352338 279266 352574
rect 279502 352338 279586 352574
rect 279822 352338 315266 352574
rect 315502 352338 315586 352574
rect 315822 352338 351266 352574
rect 351502 352338 351586 352574
rect 351822 352338 387266 352574
rect 387502 352338 387586 352574
rect 387822 352338 423266 352574
rect 423502 352338 423586 352574
rect 423822 352338 459266 352574
rect 459502 352338 459586 352574
rect 459822 352338 495266 352574
rect 495502 352338 495586 352574
rect 495822 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect -6806 352306 590730 352338
rect -4886 349174 588810 349206
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 59546 349174
rect 59782 348938 59866 349174
rect 60102 348938 95546 349174
rect 95782 348938 95866 349174
rect 96102 348938 131546 349174
rect 131782 348938 131866 349174
rect 132102 348938 167546 349174
rect 167782 348938 167866 349174
rect 168102 348938 203546 349174
rect 203782 348938 203866 349174
rect 204102 348938 239546 349174
rect 239782 348938 239866 349174
rect 240102 348938 275546 349174
rect 275782 348938 275866 349174
rect 276102 348938 311546 349174
rect 311782 348938 311866 349174
rect 312102 348938 347546 349174
rect 347782 348938 347866 349174
rect 348102 348938 383546 349174
rect 383782 348938 383866 349174
rect 384102 348938 419546 349174
rect 419782 348938 419866 349174
rect 420102 348938 455546 349174
rect 455782 348938 455866 349174
rect 456102 348938 491546 349174
rect 491782 348938 491866 349174
rect 492102 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect -4886 348854 588810 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 59546 348854
rect 59782 348618 59866 348854
rect 60102 348618 95546 348854
rect 95782 348618 95866 348854
rect 96102 348618 131546 348854
rect 131782 348618 131866 348854
rect 132102 348618 167546 348854
rect 167782 348618 167866 348854
rect 168102 348618 203546 348854
rect 203782 348618 203866 348854
rect 204102 348618 239546 348854
rect 239782 348618 239866 348854
rect 240102 348618 275546 348854
rect 275782 348618 275866 348854
rect 276102 348618 311546 348854
rect 311782 348618 311866 348854
rect 312102 348618 347546 348854
rect 347782 348618 347866 348854
rect 348102 348618 383546 348854
rect 383782 348618 383866 348854
rect 384102 348618 419546 348854
rect 419782 348618 419866 348854
rect 420102 348618 455546 348854
rect 455782 348618 455866 348854
rect 456102 348618 491546 348854
rect 491782 348618 491866 348854
rect 492102 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect -4886 348586 588810 348618
rect -2966 345454 586890 345486
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect -2966 345134 586890 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect -2966 344866 586890 344898
rect -8726 338614 592650 338646
rect -8726 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 84986 338614
rect 85222 338378 85306 338614
rect 85542 338378 120986 338614
rect 121222 338378 121306 338614
rect 121542 338378 156986 338614
rect 157222 338378 157306 338614
rect 157542 338378 192986 338614
rect 193222 338378 193306 338614
rect 193542 338378 228986 338614
rect 229222 338378 229306 338614
rect 229542 338378 264986 338614
rect 265222 338378 265306 338614
rect 265542 338378 300986 338614
rect 301222 338378 301306 338614
rect 301542 338378 336986 338614
rect 337222 338378 337306 338614
rect 337542 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 480986 338614
rect 481222 338378 481306 338614
rect 481542 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 592650 338614
rect -8726 338294 592650 338378
rect -8726 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 84986 338294
rect 85222 338058 85306 338294
rect 85542 338058 120986 338294
rect 121222 338058 121306 338294
rect 121542 338058 156986 338294
rect 157222 338058 157306 338294
rect 157542 338058 192986 338294
rect 193222 338058 193306 338294
rect 193542 338058 228986 338294
rect 229222 338058 229306 338294
rect 229542 338058 264986 338294
rect 265222 338058 265306 338294
rect 265542 338058 300986 338294
rect 301222 338058 301306 338294
rect 301542 338058 336986 338294
rect 337222 338058 337306 338294
rect 337542 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 480986 338294
rect 481222 338058 481306 338294
rect 481542 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 592650 338294
rect -8726 338026 592650 338058
rect -6806 334894 590730 334926
rect -6806 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 81266 334894
rect 81502 334658 81586 334894
rect 81822 334658 117266 334894
rect 117502 334658 117586 334894
rect 117822 334658 153266 334894
rect 153502 334658 153586 334894
rect 153822 334658 189266 334894
rect 189502 334658 189586 334894
rect 189822 334658 225266 334894
rect 225502 334658 225586 334894
rect 225822 334658 261266 334894
rect 261502 334658 261586 334894
rect 261822 334658 297266 334894
rect 297502 334658 297586 334894
rect 297822 334658 333266 334894
rect 333502 334658 333586 334894
rect 333822 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 405266 334894
rect 405502 334658 405586 334894
rect 405822 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 477266 334894
rect 477502 334658 477586 334894
rect 477822 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 590730 334894
rect -6806 334574 590730 334658
rect -6806 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 81266 334574
rect 81502 334338 81586 334574
rect 81822 334338 117266 334574
rect 117502 334338 117586 334574
rect 117822 334338 153266 334574
rect 153502 334338 153586 334574
rect 153822 334338 189266 334574
rect 189502 334338 189586 334574
rect 189822 334338 225266 334574
rect 225502 334338 225586 334574
rect 225822 334338 261266 334574
rect 261502 334338 261586 334574
rect 261822 334338 297266 334574
rect 297502 334338 297586 334574
rect 297822 334338 333266 334574
rect 333502 334338 333586 334574
rect 333822 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 405266 334574
rect 405502 334338 405586 334574
rect 405822 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 477266 334574
rect 477502 334338 477586 334574
rect 477822 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 590730 334574
rect -6806 334306 590730 334338
rect -4886 331174 588810 331206
rect -4886 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 185546 331174
rect 185782 330938 185866 331174
rect 186102 330938 221546 331174
rect 221782 330938 221866 331174
rect 222102 330938 257546 331174
rect 257782 330938 257866 331174
rect 258102 330938 293546 331174
rect 293782 330938 293866 331174
rect 294102 330938 329546 331174
rect 329782 330938 329866 331174
rect 330102 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 588810 331174
rect -4886 330854 588810 330938
rect -4886 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 185546 330854
rect 185782 330618 185866 330854
rect 186102 330618 221546 330854
rect 221782 330618 221866 330854
rect 222102 330618 257546 330854
rect 257782 330618 257866 330854
rect 258102 330618 293546 330854
rect 293782 330618 293866 330854
rect 294102 330618 329546 330854
rect 329782 330618 329866 330854
rect 330102 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 588810 330854
rect -4886 330586 588810 330618
rect -2966 327454 586890 327486
rect -2966 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 586890 327454
rect -2966 327134 586890 327218
rect -2966 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 586890 327134
rect -2966 326866 586890 326898
rect -8726 320614 592650 320646
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 174986 320614
rect 175222 320378 175306 320614
rect 175542 320378 210986 320614
rect 211222 320378 211306 320614
rect 211542 320378 246986 320614
rect 247222 320378 247306 320614
rect 247542 320378 282986 320614
rect 283222 320378 283306 320614
rect 283542 320378 318986 320614
rect 319222 320378 319306 320614
rect 319542 320378 354986 320614
rect 355222 320378 355306 320614
rect 355542 320378 390986 320614
rect 391222 320378 391306 320614
rect 391542 320378 426986 320614
rect 427222 320378 427306 320614
rect 427542 320378 462986 320614
rect 463222 320378 463306 320614
rect 463542 320378 498986 320614
rect 499222 320378 499306 320614
rect 499542 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect -8726 320294 592650 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 174986 320294
rect 175222 320058 175306 320294
rect 175542 320058 210986 320294
rect 211222 320058 211306 320294
rect 211542 320058 246986 320294
rect 247222 320058 247306 320294
rect 247542 320058 282986 320294
rect 283222 320058 283306 320294
rect 283542 320058 318986 320294
rect 319222 320058 319306 320294
rect 319542 320058 354986 320294
rect 355222 320058 355306 320294
rect 355542 320058 390986 320294
rect 391222 320058 391306 320294
rect 391542 320058 426986 320294
rect 427222 320058 427306 320294
rect 427542 320058 462986 320294
rect 463222 320058 463306 320294
rect 463542 320058 498986 320294
rect 499222 320058 499306 320294
rect 499542 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect -8726 320026 592650 320058
rect -6806 316894 590730 316926
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 63266 316894
rect 63502 316658 63586 316894
rect 63822 316658 171266 316894
rect 171502 316658 171586 316894
rect 171822 316658 207266 316894
rect 207502 316658 207586 316894
rect 207822 316658 243266 316894
rect 243502 316658 243586 316894
rect 243822 316658 279266 316894
rect 279502 316658 279586 316894
rect 279822 316658 315266 316894
rect 315502 316658 315586 316894
rect 315822 316658 351266 316894
rect 351502 316658 351586 316894
rect 351822 316658 387266 316894
rect 387502 316658 387586 316894
rect 387822 316658 423266 316894
rect 423502 316658 423586 316894
rect 423822 316658 459266 316894
rect 459502 316658 459586 316894
rect 459822 316658 495266 316894
rect 495502 316658 495586 316894
rect 495822 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect -6806 316574 590730 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 63266 316574
rect 63502 316338 63586 316574
rect 63822 316338 171266 316574
rect 171502 316338 171586 316574
rect 171822 316338 207266 316574
rect 207502 316338 207586 316574
rect 207822 316338 243266 316574
rect 243502 316338 243586 316574
rect 243822 316338 279266 316574
rect 279502 316338 279586 316574
rect 279822 316338 315266 316574
rect 315502 316338 315586 316574
rect 315822 316338 351266 316574
rect 351502 316338 351586 316574
rect 351822 316338 387266 316574
rect 387502 316338 387586 316574
rect 387822 316338 423266 316574
rect 423502 316338 423586 316574
rect 423822 316338 459266 316574
rect 459502 316338 459586 316574
rect 459822 316338 495266 316574
rect 495502 316338 495586 316574
rect 495822 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect -6806 316306 590730 316338
rect -4886 313174 588810 313206
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 59546 313174
rect 59782 312938 59866 313174
rect 60102 312938 167546 313174
rect 167782 312938 167866 313174
rect 168102 312938 203546 313174
rect 203782 312938 203866 313174
rect 204102 312938 239546 313174
rect 239782 312938 239866 313174
rect 240102 312938 275546 313174
rect 275782 312938 275866 313174
rect 276102 312938 311546 313174
rect 311782 312938 311866 313174
rect 312102 312938 347546 313174
rect 347782 312938 347866 313174
rect 348102 312938 383546 313174
rect 383782 312938 383866 313174
rect 384102 312938 419546 313174
rect 419782 312938 419866 313174
rect 420102 312938 455546 313174
rect 455782 312938 455866 313174
rect 456102 312938 491546 313174
rect 491782 312938 491866 313174
rect 492102 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect -4886 312854 588810 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 59546 312854
rect 59782 312618 59866 312854
rect 60102 312618 167546 312854
rect 167782 312618 167866 312854
rect 168102 312618 203546 312854
rect 203782 312618 203866 312854
rect 204102 312618 239546 312854
rect 239782 312618 239866 312854
rect 240102 312618 275546 312854
rect 275782 312618 275866 312854
rect 276102 312618 311546 312854
rect 311782 312618 311866 312854
rect 312102 312618 347546 312854
rect 347782 312618 347866 312854
rect 348102 312618 383546 312854
rect 383782 312618 383866 312854
rect 384102 312618 419546 312854
rect 419782 312618 419866 312854
rect 420102 312618 455546 312854
rect 455782 312618 455866 312854
rect 456102 312618 491546 312854
rect 491782 312618 491866 312854
rect 492102 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect -4886 312586 588810 312618
rect -2966 309454 586890 309486
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 88380 309454
rect 88616 309218 119100 309454
rect 119336 309218 149820 309454
rect 150056 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect -2966 309134 586890 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 88380 309134
rect 88616 308898 119100 309134
rect 119336 308898 149820 309134
rect 150056 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect -2966 308866 586890 308898
rect -8726 302614 592650 302646
rect -8726 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 192986 302614
rect 193222 302378 193306 302614
rect 193542 302378 228986 302614
rect 229222 302378 229306 302614
rect 229542 302378 264986 302614
rect 265222 302378 265306 302614
rect 265542 302378 300986 302614
rect 301222 302378 301306 302614
rect 301542 302378 336986 302614
rect 337222 302378 337306 302614
rect 337542 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 408986 302614
rect 409222 302378 409306 302614
rect 409542 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 592650 302614
rect -8726 302294 592650 302378
rect -8726 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 192986 302294
rect 193222 302058 193306 302294
rect 193542 302058 228986 302294
rect 229222 302058 229306 302294
rect 229542 302058 264986 302294
rect 265222 302058 265306 302294
rect 265542 302058 300986 302294
rect 301222 302058 301306 302294
rect 301542 302058 336986 302294
rect 337222 302058 337306 302294
rect 337542 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 408986 302294
rect 409222 302058 409306 302294
rect 409542 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 592650 302294
rect -8726 302026 592650 302058
rect -6806 298894 590730 298926
rect -6806 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 189266 298894
rect 189502 298658 189586 298894
rect 189822 298658 225266 298894
rect 225502 298658 225586 298894
rect 225822 298658 261266 298894
rect 261502 298658 261586 298894
rect 261822 298658 297266 298894
rect 297502 298658 297586 298894
rect 297822 298658 333266 298894
rect 333502 298658 333586 298894
rect 333822 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 405266 298894
rect 405502 298658 405586 298894
rect 405822 298658 441266 298894
rect 441502 298658 441586 298894
rect 441822 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 590730 298894
rect -6806 298574 590730 298658
rect -6806 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 189266 298574
rect 189502 298338 189586 298574
rect 189822 298338 225266 298574
rect 225502 298338 225586 298574
rect 225822 298338 261266 298574
rect 261502 298338 261586 298574
rect 261822 298338 297266 298574
rect 297502 298338 297586 298574
rect 297822 298338 333266 298574
rect 333502 298338 333586 298574
rect 333822 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 405266 298574
rect 405502 298338 405586 298574
rect 405822 298338 441266 298574
rect 441502 298338 441586 298574
rect 441822 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 590730 298574
rect -6806 298306 590730 298338
rect -4886 295174 588810 295206
rect -4886 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 185546 295174
rect 185782 294938 185866 295174
rect 186102 294938 221546 295174
rect 221782 294938 221866 295174
rect 222102 294938 257546 295174
rect 257782 294938 257866 295174
rect 258102 294938 293546 295174
rect 293782 294938 293866 295174
rect 294102 294938 329546 295174
rect 329782 294938 329866 295174
rect 330102 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 588810 295174
rect -4886 294854 588810 294938
rect -4886 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 185546 294854
rect 185782 294618 185866 294854
rect 186102 294618 221546 294854
rect 221782 294618 221866 294854
rect 222102 294618 257546 294854
rect 257782 294618 257866 294854
rect 258102 294618 293546 294854
rect 293782 294618 293866 294854
rect 294102 294618 329546 294854
rect 329782 294618 329866 294854
rect 330102 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 588810 294854
rect -4886 294586 588810 294618
rect -2966 291454 586890 291486
rect -2966 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 73020 291454
rect 73256 291218 103740 291454
rect 103976 291218 134460 291454
rect 134696 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 586890 291454
rect -2966 291134 586890 291218
rect -2966 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 73020 291134
rect 73256 290898 103740 291134
rect 103976 290898 134460 291134
rect 134696 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 586890 291134
rect -2966 290866 586890 290898
rect -8726 284614 592650 284646
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 174986 284614
rect 175222 284378 175306 284614
rect 175542 284378 246986 284614
rect 247222 284378 247306 284614
rect 247542 284378 282986 284614
rect 283222 284378 283306 284614
rect 283542 284378 318986 284614
rect 319222 284378 319306 284614
rect 319542 284378 354986 284614
rect 355222 284378 355306 284614
rect 355542 284378 390986 284614
rect 391222 284378 391306 284614
rect 391542 284378 426986 284614
rect 427222 284378 427306 284614
rect 427542 284378 462986 284614
rect 463222 284378 463306 284614
rect 463542 284378 498986 284614
rect 499222 284378 499306 284614
rect 499542 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect -8726 284294 592650 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 174986 284294
rect 175222 284058 175306 284294
rect 175542 284058 246986 284294
rect 247222 284058 247306 284294
rect 247542 284058 282986 284294
rect 283222 284058 283306 284294
rect 283542 284058 318986 284294
rect 319222 284058 319306 284294
rect 319542 284058 354986 284294
rect 355222 284058 355306 284294
rect 355542 284058 390986 284294
rect 391222 284058 391306 284294
rect 391542 284058 426986 284294
rect 427222 284058 427306 284294
rect 427542 284058 462986 284294
rect 463222 284058 463306 284294
rect 463542 284058 498986 284294
rect 499222 284058 499306 284294
rect 499542 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect -8726 284026 592650 284058
rect -6806 280894 590730 280926
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 63266 280894
rect 63502 280658 63586 280894
rect 63822 280658 171266 280894
rect 171502 280658 171586 280894
rect 171822 280658 279266 280894
rect 279502 280658 279586 280894
rect 279822 280658 315266 280894
rect 315502 280658 315586 280894
rect 315822 280658 351266 280894
rect 351502 280658 351586 280894
rect 351822 280658 387266 280894
rect 387502 280658 387586 280894
rect 387822 280658 423266 280894
rect 423502 280658 423586 280894
rect 423822 280658 459266 280894
rect 459502 280658 459586 280894
rect 459822 280658 495266 280894
rect 495502 280658 495586 280894
rect 495822 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect -6806 280574 590730 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 63266 280574
rect 63502 280338 63586 280574
rect 63822 280338 171266 280574
rect 171502 280338 171586 280574
rect 171822 280338 279266 280574
rect 279502 280338 279586 280574
rect 279822 280338 315266 280574
rect 315502 280338 315586 280574
rect 315822 280338 351266 280574
rect 351502 280338 351586 280574
rect 351822 280338 387266 280574
rect 387502 280338 387586 280574
rect 387822 280338 423266 280574
rect 423502 280338 423586 280574
rect 423822 280338 459266 280574
rect 459502 280338 459586 280574
rect 459822 280338 495266 280574
rect 495502 280338 495586 280574
rect 495822 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect -6806 280306 590730 280338
rect -4886 277174 588810 277206
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 59546 277174
rect 59782 276938 59866 277174
rect 60102 276938 167546 277174
rect 167782 276938 167866 277174
rect 168102 276938 275546 277174
rect 275782 276938 275866 277174
rect 276102 276938 311546 277174
rect 311782 276938 311866 277174
rect 312102 276938 347546 277174
rect 347782 276938 347866 277174
rect 348102 276938 383546 277174
rect 383782 276938 383866 277174
rect 384102 276938 419546 277174
rect 419782 276938 419866 277174
rect 420102 276938 455546 277174
rect 455782 276938 455866 277174
rect 456102 276938 491546 277174
rect 491782 276938 491866 277174
rect 492102 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect -4886 276854 588810 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 59546 276854
rect 59782 276618 59866 276854
rect 60102 276618 167546 276854
rect 167782 276618 167866 276854
rect 168102 276618 275546 276854
rect 275782 276618 275866 276854
rect 276102 276618 311546 276854
rect 311782 276618 311866 276854
rect 312102 276618 347546 276854
rect 347782 276618 347866 276854
rect 348102 276618 383546 276854
rect 383782 276618 383866 276854
rect 384102 276618 419546 276854
rect 419782 276618 419866 276854
rect 420102 276618 455546 276854
rect 455782 276618 455866 276854
rect 456102 276618 491546 276854
rect 491782 276618 491866 276854
rect 492102 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect -4886 276586 588810 276618
rect -2966 273454 586890 273486
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 88380 273454
rect 88616 273218 119100 273454
rect 119336 273218 149820 273454
rect 150056 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 219810 273454
rect 220046 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect -2966 273134 586890 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 88380 273134
rect 88616 272898 119100 273134
rect 119336 272898 149820 273134
rect 150056 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 219810 273134
rect 220046 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect -2966 272866 586890 272898
rect -8726 266614 592650 266646
rect -8726 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 192986 266614
rect 193222 266378 193306 266614
rect 193542 266378 264986 266614
rect 265222 266378 265306 266614
rect 265542 266378 300986 266614
rect 301222 266378 301306 266614
rect 301542 266378 336986 266614
rect 337222 266378 337306 266614
rect 337542 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 592650 266614
rect -8726 266294 592650 266378
rect -8726 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 192986 266294
rect 193222 266058 193306 266294
rect 193542 266058 264986 266294
rect 265222 266058 265306 266294
rect 265542 266058 300986 266294
rect 301222 266058 301306 266294
rect 301542 266058 336986 266294
rect 337222 266058 337306 266294
rect 337542 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 592650 266294
rect -8726 266026 592650 266058
rect -6806 262894 590730 262926
rect -6806 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 261266 262894
rect 261502 262658 261586 262894
rect 261822 262658 297266 262894
rect 297502 262658 297586 262894
rect 297822 262658 333266 262894
rect 333502 262658 333586 262894
rect 333822 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 590730 262894
rect -6806 262574 590730 262658
rect -6806 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 261266 262574
rect 261502 262338 261586 262574
rect 261822 262338 297266 262574
rect 297502 262338 297586 262574
rect 297822 262338 333266 262574
rect 333502 262338 333586 262574
rect 333822 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 590730 262574
rect -6806 262306 590730 262338
rect -4886 259174 588810 259206
rect -4886 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 257546 259174
rect 257782 258938 257866 259174
rect 258102 258938 293546 259174
rect 293782 258938 293866 259174
rect 294102 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 588810 259174
rect -4886 258854 588810 258938
rect -4886 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 257546 258854
rect 257782 258618 257866 258854
rect 258102 258618 293546 258854
rect 293782 258618 293866 258854
rect 294102 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 588810 258854
rect -4886 258586 588810 258618
rect -2966 255454 586890 255486
rect -2966 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 73020 255454
rect 73256 255218 103740 255454
rect 103976 255218 134460 255454
rect 134696 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 204450 255454
rect 204686 255218 235170 255454
rect 235406 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 586890 255454
rect -2966 255134 586890 255218
rect -2966 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 73020 255134
rect 73256 254898 103740 255134
rect 103976 254898 134460 255134
rect 134696 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 204450 255134
rect 204686 254898 235170 255134
rect 235406 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 586890 255134
rect -2966 254866 586890 254898
rect -8726 248614 592650 248646
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 174986 248614
rect 175222 248378 175306 248614
rect 175542 248378 246986 248614
rect 247222 248378 247306 248614
rect 247542 248378 282986 248614
rect 283222 248378 283306 248614
rect 283542 248378 318986 248614
rect 319222 248378 319306 248614
rect 319542 248378 354986 248614
rect 355222 248378 355306 248614
rect 355542 248378 390986 248614
rect 391222 248378 391306 248614
rect 391542 248378 426986 248614
rect 427222 248378 427306 248614
rect 427542 248378 462986 248614
rect 463222 248378 463306 248614
rect 463542 248378 498986 248614
rect 499222 248378 499306 248614
rect 499542 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect -8726 248294 592650 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 174986 248294
rect 175222 248058 175306 248294
rect 175542 248058 246986 248294
rect 247222 248058 247306 248294
rect 247542 248058 282986 248294
rect 283222 248058 283306 248294
rect 283542 248058 318986 248294
rect 319222 248058 319306 248294
rect 319542 248058 354986 248294
rect 355222 248058 355306 248294
rect 355542 248058 390986 248294
rect 391222 248058 391306 248294
rect 391542 248058 426986 248294
rect 427222 248058 427306 248294
rect 427542 248058 462986 248294
rect 463222 248058 463306 248294
rect 463542 248058 498986 248294
rect 499222 248058 499306 248294
rect 499542 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect -8726 248026 592650 248058
rect -6806 244894 590730 244926
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 63266 244894
rect 63502 244658 63586 244894
rect 63822 244658 171266 244894
rect 171502 244658 171586 244894
rect 171822 244658 279266 244894
rect 279502 244658 279586 244894
rect 279822 244658 315266 244894
rect 315502 244658 315586 244894
rect 315822 244658 351266 244894
rect 351502 244658 351586 244894
rect 351822 244658 387266 244894
rect 387502 244658 387586 244894
rect 387822 244658 423266 244894
rect 423502 244658 423586 244894
rect 423822 244658 459266 244894
rect 459502 244658 459586 244894
rect 459822 244658 495266 244894
rect 495502 244658 495586 244894
rect 495822 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect -6806 244574 590730 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 63266 244574
rect 63502 244338 63586 244574
rect 63822 244338 171266 244574
rect 171502 244338 171586 244574
rect 171822 244338 279266 244574
rect 279502 244338 279586 244574
rect 279822 244338 315266 244574
rect 315502 244338 315586 244574
rect 315822 244338 351266 244574
rect 351502 244338 351586 244574
rect 351822 244338 387266 244574
rect 387502 244338 387586 244574
rect 387822 244338 423266 244574
rect 423502 244338 423586 244574
rect 423822 244338 459266 244574
rect 459502 244338 459586 244574
rect 459822 244338 495266 244574
rect 495502 244338 495586 244574
rect 495822 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect -6806 244306 590730 244338
rect -4886 241174 588810 241206
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 59546 241174
rect 59782 240938 59866 241174
rect 60102 240938 167546 241174
rect 167782 240938 167866 241174
rect 168102 240938 275546 241174
rect 275782 240938 275866 241174
rect 276102 240938 311546 241174
rect 311782 240938 311866 241174
rect 312102 240938 347546 241174
rect 347782 240938 347866 241174
rect 348102 240938 383546 241174
rect 383782 240938 383866 241174
rect 384102 240938 419546 241174
rect 419782 240938 419866 241174
rect 420102 240938 455546 241174
rect 455782 240938 455866 241174
rect 456102 240938 491546 241174
rect 491782 240938 491866 241174
rect 492102 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect -4886 240854 588810 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 59546 240854
rect 59782 240618 59866 240854
rect 60102 240618 167546 240854
rect 167782 240618 167866 240854
rect 168102 240618 275546 240854
rect 275782 240618 275866 240854
rect 276102 240618 311546 240854
rect 311782 240618 311866 240854
rect 312102 240618 347546 240854
rect 347782 240618 347866 240854
rect 348102 240618 383546 240854
rect 383782 240618 383866 240854
rect 384102 240618 419546 240854
rect 419782 240618 419866 240854
rect 420102 240618 455546 240854
rect 455782 240618 455866 240854
rect 456102 240618 491546 240854
rect 491782 240618 491866 240854
rect 492102 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect -4886 240586 588810 240618
rect -2966 237454 586890 237486
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect -2966 237134 586890 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect -2966 236866 586890 236898
rect -8726 230614 592650 230646
rect -8726 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 84986 230614
rect 85222 230378 85306 230614
rect 85542 230378 120986 230614
rect 121222 230378 121306 230614
rect 121542 230378 156986 230614
rect 157222 230378 157306 230614
rect 157542 230378 192986 230614
rect 193222 230378 193306 230614
rect 193542 230378 228986 230614
rect 229222 230378 229306 230614
rect 229542 230378 264986 230614
rect 265222 230378 265306 230614
rect 265542 230378 300986 230614
rect 301222 230378 301306 230614
rect 301542 230378 336986 230614
rect 337222 230378 337306 230614
rect 337542 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 592650 230614
rect -8726 230294 592650 230378
rect -8726 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 84986 230294
rect 85222 230058 85306 230294
rect 85542 230058 120986 230294
rect 121222 230058 121306 230294
rect 121542 230058 156986 230294
rect 157222 230058 157306 230294
rect 157542 230058 192986 230294
rect 193222 230058 193306 230294
rect 193542 230058 228986 230294
rect 229222 230058 229306 230294
rect 229542 230058 264986 230294
rect 265222 230058 265306 230294
rect 265542 230058 300986 230294
rect 301222 230058 301306 230294
rect 301542 230058 336986 230294
rect 337222 230058 337306 230294
rect 337542 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 592650 230294
rect -8726 230026 592650 230058
rect -6806 226894 590730 226926
rect -6806 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 81266 226894
rect 81502 226658 81586 226894
rect 81822 226658 117266 226894
rect 117502 226658 117586 226894
rect 117822 226658 153266 226894
rect 153502 226658 153586 226894
rect 153822 226658 189266 226894
rect 189502 226658 189586 226894
rect 189822 226658 225266 226894
rect 225502 226658 225586 226894
rect 225822 226658 261266 226894
rect 261502 226658 261586 226894
rect 261822 226658 297266 226894
rect 297502 226658 297586 226894
rect 297822 226658 333266 226894
rect 333502 226658 333586 226894
rect 333822 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 405266 226894
rect 405502 226658 405586 226894
rect 405822 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 590730 226894
rect -6806 226574 590730 226658
rect -6806 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 81266 226574
rect 81502 226338 81586 226574
rect 81822 226338 117266 226574
rect 117502 226338 117586 226574
rect 117822 226338 153266 226574
rect 153502 226338 153586 226574
rect 153822 226338 189266 226574
rect 189502 226338 189586 226574
rect 189822 226338 225266 226574
rect 225502 226338 225586 226574
rect 225822 226338 261266 226574
rect 261502 226338 261586 226574
rect 261822 226338 297266 226574
rect 297502 226338 297586 226574
rect 297822 226338 333266 226574
rect 333502 226338 333586 226574
rect 333822 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 405266 226574
rect 405502 226338 405586 226574
rect 405822 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 590730 226574
rect -6806 226306 590730 226338
rect -4886 223174 588810 223206
rect -4886 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 77546 223174
rect 77782 222938 77866 223174
rect 78102 222938 113546 223174
rect 113782 222938 113866 223174
rect 114102 222938 149546 223174
rect 149782 222938 149866 223174
rect 150102 222938 185546 223174
rect 185782 222938 185866 223174
rect 186102 222938 221546 223174
rect 221782 222938 221866 223174
rect 222102 222938 257546 223174
rect 257782 222938 257866 223174
rect 258102 222938 293546 223174
rect 293782 222938 293866 223174
rect 294102 222938 329546 223174
rect 329782 222938 329866 223174
rect 330102 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 588810 223174
rect -4886 222854 588810 222938
rect -4886 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 77546 222854
rect 77782 222618 77866 222854
rect 78102 222618 113546 222854
rect 113782 222618 113866 222854
rect 114102 222618 149546 222854
rect 149782 222618 149866 222854
rect 150102 222618 185546 222854
rect 185782 222618 185866 222854
rect 186102 222618 221546 222854
rect 221782 222618 221866 222854
rect 222102 222618 257546 222854
rect 257782 222618 257866 222854
rect 258102 222618 293546 222854
rect 293782 222618 293866 222854
rect 294102 222618 329546 222854
rect 329782 222618 329866 222854
rect 330102 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 588810 222854
rect -4886 222586 588810 222618
rect -2966 219454 586890 219486
rect -2966 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 586890 219454
rect -2966 219134 586890 219218
rect -2966 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 586890 219134
rect -2966 218866 586890 218898
rect -8726 212614 592650 212646
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 66986 212614
rect 67222 212378 67306 212614
rect 67542 212378 102986 212614
rect 103222 212378 103306 212614
rect 103542 212378 138986 212614
rect 139222 212378 139306 212614
rect 139542 212378 174986 212614
rect 175222 212378 175306 212614
rect 175542 212378 210986 212614
rect 211222 212378 211306 212614
rect 211542 212378 246986 212614
rect 247222 212378 247306 212614
rect 247542 212378 282986 212614
rect 283222 212378 283306 212614
rect 283542 212378 318986 212614
rect 319222 212378 319306 212614
rect 319542 212378 354986 212614
rect 355222 212378 355306 212614
rect 355542 212378 390986 212614
rect 391222 212378 391306 212614
rect 391542 212378 426986 212614
rect 427222 212378 427306 212614
rect 427542 212378 462986 212614
rect 463222 212378 463306 212614
rect 463542 212378 498986 212614
rect 499222 212378 499306 212614
rect 499542 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect -8726 212294 592650 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 66986 212294
rect 67222 212058 67306 212294
rect 67542 212058 102986 212294
rect 103222 212058 103306 212294
rect 103542 212058 138986 212294
rect 139222 212058 139306 212294
rect 139542 212058 174986 212294
rect 175222 212058 175306 212294
rect 175542 212058 210986 212294
rect 211222 212058 211306 212294
rect 211542 212058 246986 212294
rect 247222 212058 247306 212294
rect 247542 212058 282986 212294
rect 283222 212058 283306 212294
rect 283542 212058 318986 212294
rect 319222 212058 319306 212294
rect 319542 212058 354986 212294
rect 355222 212058 355306 212294
rect 355542 212058 390986 212294
rect 391222 212058 391306 212294
rect 391542 212058 426986 212294
rect 427222 212058 427306 212294
rect 427542 212058 462986 212294
rect 463222 212058 463306 212294
rect 463542 212058 498986 212294
rect 499222 212058 499306 212294
rect 499542 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect -8726 212026 592650 212058
rect -6806 208894 590730 208926
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 63266 208894
rect 63502 208658 63586 208894
rect 63822 208658 99266 208894
rect 99502 208658 99586 208894
rect 99822 208658 135266 208894
rect 135502 208658 135586 208894
rect 135822 208658 171266 208894
rect 171502 208658 171586 208894
rect 171822 208658 207266 208894
rect 207502 208658 207586 208894
rect 207822 208658 243266 208894
rect 243502 208658 243586 208894
rect 243822 208658 279266 208894
rect 279502 208658 279586 208894
rect 279822 208658 315266 208894
rect 315502 208658 315586 208894
rect 315822 208658 351266 208894
rect 351502 208658 351586 208894
rect 351822 208658 387266 208894
rect 387502 208658 387586 208894
rect 387822 208658 423266 208894
rect 423502 208658 423586 208894
rect 423822 208658 459266 208894
rect 459502 208658 459586 208894
rect 459822 208658 495266 208894
rect 495502 208658 495586 208894
rect 495822 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect -6806 208574 590730 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 63266 208574
rect 63502 208338 63586 208574
rect 63822 208338 99266 208574
rect 99502 208338 99586 208574
rect 99822 208338 135266 208574
rect 135502 208338 135586 208574
rect 135822 208338 171266 208574
rect 171502 208338 171586 208574
rect 171822 208338 207266 208574
rect 207502 208338 207586 208574
rect 207822 208338 243266 208574
rect 243502 208338 243586 208574
rect 243822 208338 279266 208574
rect 279502 208338 279586 208574
rect 279822 208338 315266 208574
rect 315502 208338 315586 208574
rect 315822 208338 351266 208574
rect 351502 208338 351586 208574
rect 351822 208338 387266 208574
rect 387502 208338 387586 208574
rect 387822 208338 423266 208574
rect 423502 208338 423586 208574
rect 423822 208338 459266 208574
rect 459502 208338 459586 208574
rect 459822 208338 495266 208574
rect 495502 208338 495586 208574
rect 495822 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect -6806 208306 590730 208338
rect -4886 205174 588810 205206
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 59546 205174
rect 59782 204938 59866 205174
rect 60102 204938 95546 205174
rect 95782 204938 95866 205174
rect 96102 204938 131546 205174
rect 131782 204938 131866 205174
rect 132102 204938 167546 205174
rect 167782 204938 167866 205174
rect 168102 204938 203546 205174
rect 203782 204938 203866 205174
rect 204102 204938 239546 205174
rect 239782 204938 239866 205174
rect 240102 204938 275546 205174
rect 275782 204938 275866 205174
rect 276102 204938 311546 205174
rect 311782 204938 311866 205174
rect 312102 204938 347546 205174
rect 347782 204938 347866 205174
rect 348102 204938 383546 205174
rect 383782 204938 383866 205174
rect 384102 204938 419546 205174
rect 419782 204938 419866 205174
rect 420102 204938 455546 205174
rect 455782 204938 455866 205174
rect 456102 204938 491546 205174
rect 491782 204938 491866 205174
rect 492102 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect -4886 204854 588810 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 59546 204854
rect 59782 204618 59866 204854
rect 60102 204618 95546 204854
rect 95782 204618 95866 204854
rect 96102 204618 131546 204854
rect 131782 204618 131866 204854
rect 132102 204618 167546 204854
rect 167782 204618 167866 204854
rect 168102 204618 203546 204854
rect 203782 204618 203866 204854
rect 204102 204618 239546 204854
rect 239782 204618 239866 204854
rect 240102 204618 275546 204854
rect 275782 204618 275866 204854
rect 276102 204618 311546 204854
rect 311782 204618 311866 204854
rect 312102 204618 347546 204854
rect 347782 204618 347866 204854
rect 348102 204618 383546 204854
rect 383782 204618 383866 204854
rect 384102 204618 419546 204854
rect 419782 204618 419866 204854
rect 420102 204618 455546 204854
rect 455782 204618 455866 204854
rect 456102 204618 491546 204854
rect 491782 204618 491866 204854
rect 492102 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect -4886 204586 588810 204618
rect -2966 201454 586890 201486
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect -2966 201134 586890 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect -2966 200866 586890 200898
rect -8726 194614 592650 194646
rect -8726 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 84986 194614
rect 85222 194378 85306 194614
rect 85542 194378 120986 194614
rect 121222 194378 121306 194614
rect 121542 194378 156986 194614
rect 157222 194378 157306 194614
rect 157542 194378 192986 194614
rect 193222 194378 193306 194614
rect 193542 194378 228986 194614
rect 229222 194378 229306 194614
rect 229542 194378 264986 194614
rect 265222 194378 265306 194614
rect 265542 194378 300986 194614
rect 301222 194378 301306 194614
rect 301542 194378 336986 194614
rect 337222 194378 337306 194614
rect 337542 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 592650 194614
rect -8726 194294 592650 194378
rect -8726 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 84986 194294
rect 85222 194058 85306 194294
rect 85542 194058 120986 194294
rect 121222 194058 121306 194294
rect 121542 194058 156986 194294
rect 157222 194058 157306 194294
rect 157542 194058 192986 194294
rect 193222 194058 193306 194294
rect 193542 194058 228986 194294
rect 229222 194058 229306 194294
rect 229542 194058 264986 194294
rect 265222 194058 265306 194294
rect 265542 194058 300986 194294
rect 301222 194058 301306 194294
rect 301542 194058 336986 194294
rect 337222 194058 337306 194294
rect 337542 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 592650 194294
rect -8726 194026 592650 194058
rect -6806 190894 590730 190926
rect -6806 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 81266 190894
rect 81502 190658 81586 190894
rect 81822 190658 117266 190894
rect 117502 190658 117586 190894
rect 117822 190658 153266 190894
rect 153502 190658 153586 190894
rect 153822 190658 189266 190894
rect 189502 190658 189586 190894
rect 189822 190658 225266 190894
rect 225502 190658 225586 190894
rect 225822 190658 261266 190894
rect 261502 190658 261586 190894
rect 261822 190658 297266 190894
rect 297502 190658 297586 190894
rect 297822 190658 333266 190894
rect 333502 190658 333586 190894
rect 333822 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 590730 190894
rect -6806 190574 590730 190658
rect -6806 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 81266 190574
rect 81502 190338 81586 190574
rect 81822 190338 117266 190574
rect 117502 190338 117586 190574
rect 117822 190338 153266 190574
rect 153502 190338 153586 190574
rect 153822 190338 189266 190574
rect 189502 190338 189586 190574
rect 189822 190338 225266 190574
rect 225502 190338 225586 190574
rect 225822 190338 261266 190574
rect 261502 190338 261586 190574
rect 261822 190338 297266 190574
rect 297502 190338 297586 190574
rect 297822 190338 333266 190574
rect 333502 190338 333586 190574
rect 333822 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 590730 190574
rect -6806 190306 590730 190338
rect -4886 187174 588810 187206
rect -4886 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 77546 187174
rect 77782 186938 77866 187174
rect 78102 186938 113546 187174
rect 113782 186938 113866 187174
rect 114102 186938 149546 187174
rect 149782 186938 149866 187174
rect 150102 186938 185546 187174
rect 185782 186938 185866 187174
rect 186102 186938 221546 187174
rect 221782 186938 221866 187174
rect 222102 186938 257546 187174
rect 257782 186938 257866 187174
rect 258102 186938 293546 187174
rect 293782 186938 293866 187174
rect 294102 186938 329546 187174
rect 329782 186938 329866 187174
rect 330102 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 588810 187174
rect -4886 186854 588810 186938
rect -4886 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 77546 186854
rect 77782 186618 77866 186854
rect 78102 186618 113546 186854
rect 113782 186618 113866 186854
rect 114102 186618 149546 186854
rect 149782 186618 149866 186854
rect 150102 186618 185546 186854
rect 185782 186618 185866 186854
rect 186102 186618 221546 186854
rect 221782 186618 221866 186854
rect 222102 186618 257546 186854
rect 257782 186618 257866 186854
rect 258102 186618 293546 186854
rect 293782 186618 293866 186854
rect 294102 186618 329546 186854
rect 329782 186618 329866 186854
rect 330102 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 588810 186854
rect -4886 186586 588810 186618
rect -2966 183454 586890 183486
rect -2966 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 586890 183454
rect -2966 183134 586890 183218
rect -2966 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 586890 183134
rect -2966 182866 586890 182898
rect -8726 176614 592650 176646
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 174986 176614
rect 175222 176378 175306 176614
rect 175542 176378 210986 176614
rect 211222 176378 211306 176614
rect 211542 176378 246986 176614
rect 247222 176378 247306 176614
rect 247542 176378 282986 176614
rect 283222 176378 283306 176614
rect 283542 176378 318986 176614
rect 319222 176378 319306 176614
rect 319542 176378 354986 176614
rect 355222 176378 355306 176614
rect 355542 176378 390986 176614
rect 391222 176378 391306 176614
rect 391542 176378 426986 176614
rect 427222 176378 427306 176614
rect 427542 176378 462986 176614
rect 463222 176378 463306 176614
rect 463542 176378 498986 176614
rect 499222 176378 499306 176614
rect 499542 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect -8726 176294 592650 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 174986 176294
rect 175222 176058 175306 176294
rect 175542 176058 210986 176294
rect 211222 176058 211306 176294
rect 211542 176058 246986 176294
rect 247222 176058 247306 176294
rect 247542 176058 282986 176294
rect 283222 176058 283306 176294
rect 283542 176058 318986 176294
rect 319222 176058 319306 176294
rect 319542 176058 354986 176294
rect 355222 176058 355306 176294
rect 355542 176058 390986 176294
rect 391222 176058 391306 176294
rect 391542 176058 426986 176294
rect 427222 176058 427306 176294
rect 427542 176058 462986 176294
rect 463222 176058 463306 176294
rect 463542 176058 498986 176294
rect 499222 176058 499306 176294
rect 499542 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect -8726 176026 592650 176058
rect -6806 172894 590730 172926
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 63266 172894
rect 63502 172658 63586 172894
rect 63822 172658 171266 172894
rect 171502 172658 171586 172894
rect 171822 172658 207266 172894
rect 207502 172658 207586 172894
rect 207822 172658 243266 172894
rect 243502 172658 243586 172894
rect 243822 172658 315266 172894
rect 315502 172658 315586 172894
rect 315822 172658 351266 172894
rect 351502 172658 351586 172894
rect 351822 172658 387266 172894
rect 387502 172658 387586 172894
rect 387822 172658 423266 172894
rect 423502 172658 423586 172894
rect 423822 172658 459266 172894
rect 459502 172658 459586 172894
rect 459822 172658 495266 172894
rect 495502 172658 495586 172894
rect 495822 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect -6806 172574 590730 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 63266 172574
rect 63502 172338 63586 172574
rect 63822 172338 171266 172574
rect 171502 172338 171586 172574
rect 171822 172338 207266 172574
rect 207502 172338 207586 172574
rect 207822 172338 243266 172574
rect 243502 172338 243586 172574
rect 243822 172338 315266 172574
rect 315502 172338 315586 172574
rect 315822 172338 351266 172574
rect 351502 172338 351586 172574
rect 351822 172338 387266 172574
rect 387502 172338 387586 172574
rect 387822 172338 423266 172574
rect 423502 172338 423586 172574
rect 423822 172338 459266 172574
rect 459502 172338 459586 172574
rect 459822 172338 495266 172574
rect 495502 172338 495586 172574
rect 495822 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect -6806 172306 590730 172338
rect -4886 169174 588810 169206
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 59546 169174
rect 59782 168938 59866 169174
rect 60102 168938 167546 169174
rect 167782 168938 167866 169174
rect 168102 168938 203546 169174
rect 203782 168938 203866 169174
rect 204102 168938 239546 169174
rect 239782 168938 239866 169174
rect 240102 168938 311546 169174
rect 311782 168938 311866 169174
rect 312102 168938 347546 169174
rect 347782 168938 347866 169174
rect 348102 168938 383546 169174
rect 383782 168938 383866 169174
rect 384102 168938 419546 169174
rect 419782 168938 419866 169174
rect 420102 168938 455546 169174
rect 455782 168938 455866 169174
rect 456102 168938 491546 169174
rect 491782 168938 491866 169174
rect 492102 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect -4886 168854 588810 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 59546 168854
rect 59782 168618 59866 168854
rect 60102 168618 167546 168854
rect 167782 168618 167866 168854
rect 168102 168618 203546 168854
rect 203782 168618 203866 168854
rect 204102 168618 239546 168854
rect 239782 168618 239866 168854
rect 240102 168618 311546 168854
rect 311782 168618 311866 168854
rect 312102 168618 347546 168854
rect 347782 168618 347866 168854
rect 348102 168618 383546 168854
rect 383782 168618 383866 168854
rect 384102 168618 419546 168854
rect 419782 168618 419866 168854
rect 420102 168618 455546 168854
rect 455782 168618 455866 168854
rect 456102 168618 491546 168854
rect 491782 168618 491866 168854
rect 492102 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect -4886 168586 588810 168618
rect -2966 165454 586890 165486
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 69128 165454
rect 69364 165218 164192 165454
rect 164428 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 221249 165454
rect 221485 165218 224513 165454
rect 224749 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 272249 165454
rect 272485 165218 275513 165454
rect 275749 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect -2966 165134 586890 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 69128 165134
rect 69364 164898 164192 165134
rect 164428 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 221249 165134
rect 221485 164898 224513 165134
rect 224749 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 272249 165134
rect 272485 164898 275513 165134
rect 275749 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect -2966 164866 586890 164898
rect -8726 158614 592650 158646
rect -8726 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 192986 158614
rect 193222 158378 193306 158614
rect 193542 158378 264986 158614
rect 265222 158378 265306 158614
rect 265542 158378 300986 158614
rect 301222 158378 301306 158614
rect 301542 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 592650 158614
rect -8726 158294 592650 158378
rect -8726 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 192986 158294
rect 193222 158058 193306 158294
rect 193542 158058 264986 158294
rect 265222 158058 265306 158294
rect 265542 158058 300986 158294
rect 301222 158058 301306 158294
rect 301542 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 592650 158294
rect -8726 158026 592650 158058
rect -6806 154894 590730 154926
rect -6806 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 189266 154894
rect 189502 154658 189586 154894
rect 189822 154658 261266 154894
rect 261502 154658 261586 154894
rect 261822 154658 297266 154894
rect 297502 154658 297586 154894
rect 297822 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 441266 154894
rect 441502 154658 441586 154894
rect 441822 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 590730 154894
rect -6806 154574 590730 154658
rect -6806 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 189266 154574
rect 189502 154338 189586 154574
rect 189822 154338 261266 154574
rect 261502 154338 261586 154574
rect 261822 154338 297266 154574
rect 297502 154338 297586 154574
rect 297822 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 441266 154574
rect 441502 154338 441586 154574
rect 441822 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 590730 154574
rect -6806 154306 590730 154338
rect -4886 151174 588810 151206
rect -4886 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 257546 151174
rect 257782 150938 257866 151174
rect 258102 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 588810 151174
rect -4886 150854 588810 150938
rect -4886 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 257546 150854
rect 257782 150618 257866 150854
rect 258102 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 588810 150854
rect -4886 150586 588810 150618
rect -2966 147454 586890 147486
rect -2966 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 69808 147454
rect 70044 147218 163512 147454
rect 163748 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 219617 147454
rect 219853 147218 222881 147454
rect 223117 147218 226145 147454
rect 226381 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 270617 147454
rect 270853 147218 273881 147454
rect 274117 147218 277145 147454
rect 277381 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 586890 147454
rect -2966 147134 586890 147218
rect -2966 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 69808 147134
rect 70044 146898 163512 147134
rect 163748 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 219617 147134
rect 219853 146898 222881 147134
rect 223117 146898 226145 147134
rect 226381 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 270617 147134
rect 270853 146898 273881 147134
rect 274117 146898 277145 147134
rect 277381 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 586890 147134
rect -2966 146866 586890 146898
rect -8726 140614 592650 140646
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 174986 140614
rect 175222 140378 175306 140614
rect 175542 140378 210986 140614
rect 211222 140378 211306 140614
rect 211542 140378 246986 140614
rect 247222 140378 247306 140614
rect 247542 140378 282986 140614
rect 283222 140378 283306 140614
rect 283542 140378 318986 140614
rect 319222 140378 319306 140614
rect 319542 140378 354986 140614
rect 355222 140378 355306 140614
rect 355542 140378 390986 140614
rect 391222 140378 391306 140614
rect 391542 140378 426986 140614
rect 427222 140378 427306 140614
rect 427542 140378 462986 140614
rect 463222 140378 463306 140614
rect 463542 140378 498986 140614
rect 499222 140378 499306 140614
rect 499542 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect -8726 140294 592650 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 174986 140294
rect 175222 140058 175306 140294
rect 175542 140058 210986 140294
rect 211222 140058 211306 140294
rect 211542 140058 246986 140294
rect 247222 140058 247306 140294
rect 247542 140058 282986 140294
rect 283222 140058 283306 140294
rect 283542 140058 318986 140294
rect 319222 140058 319306 140294
rect 319542 140058 354986 140294
rect 355222 140058 355306 140294
rect 355542 140058 390986 140294
rect 391222 140058 391306 140294
rect 391542 140058 426986 140294
rect 427222 140058 427306 140294
rect 427542 140058 462986 140294
rect 463222 140058 463306 140294
rect 463542 140058 498986 140294
rect 499222 140058 499306 140294
rect 499542 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect -8726 140026 592650 140058
rect -6806 136894 590730 136926
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 63266 136894
rect 63502 136658 63586 136894
rect 63822 136658 171266 136894
rect 171502 136658 171586 136894
rect 171822 136658 207266 136894
rect 207502 136658 207586 136894
rect 207822 136658 243266 136894
rect 243502 136658 243586 136894
rect 243822 136658 315266 136894
rect 315502 136658 315586 136894
rect 315822 136658 351266 136894
rect 351502 136658 351586 136894
rect 351822 136658 387266 136894
rect 387502 136658 387586 136894
rect 387822 136658 423266 136894
rect 423502 136658 423586 136894
rect 423822 136658 459266 136894
rect 459502 136658 459586 136894
rect 459822 136658 495266 136894
rect 495502 136658 495586 136894
rect 495822 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect -6806 136574 590730 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 63266 136574
rect 63502 136338 63586 136574
rect 63822 136338 171266 136574
rect 171502 136338 171586 136574
rect 171822 136338 207266 136574
rect 207502 136338 207586 136574
rect 207822 136338 243266 136574
rect 243502 136338 243586 136574
rect 243822 136338 315266 136574
rect 315502 136338 315586 136574
rect 315822 136338 351266 136574
rect 351502 136338 351586 136574
rect 351822 136338 387266 136574
rect 387502 136338 387586 136574
rect 387822 136338 423266 136574
rect 423502 136338 423586 136574
rect 423822 136338 459266 136574
rect 459502 136338 459586 136574
rect 459822 136338 495266 136574
rect 495502 136338 495586 136574
rect 495822 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect -6806 136306 590730 136338
rect -4886 133174 588810 133206
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 59546 133174
rect 59782 132938 59866 133174
rect 60102 132938 167546 133174
rect 167782 132938 167866 133174
rect 168102 132938 203546 133174
rect 203782 132938 203866 133174
rect 204102 132938 239546 133174
rect 239782 132938 239866 133174
rect 240102 132938 311546 133174
rect 311782 132938 311866 133174
rect 312102 132938 347546 133174
rect 347782 132938 347866 133174
rect 348102 132938 383546 133174
rect 383782 132938 383866 133174
rect 384102 132938 419546 133174
rect 419782 132938 419866 133174
rect 420102 132938 455546 133174
rect 455782 132938 455866 133174
rect 456102 132938 491546 133174
rect 491782 132938 491866 133174
rect 492102 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect -4886 132854 588810 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 59546 132854
rect 59782 132618 59866 132854
rect 60102 132618 167546 132854
rect 167782 132618 167866 132854
rect 168102 132618 203546 132854
rect 203782 132618 203866 132854
rect 204102 132618 239546 132854
rect 239782 132618 239866 132854
rect 240102 132618 311546 132854
rect 311782 132618 311866 132854
rect 312102 132618 347546 132854
rect 347782 132618 347866 132854
rect 348102 132618 383546 132854
rect 383782 132618 383866 132854
rect 384102 132618 419546 132854
rect 419782 132618 419866 132854
rect 420102 132618 455546 132854
rect 455782 132618 455866 132854
rect 456102 132618 491546 132854
rect 491782 132618 491866 132854
rect 492102 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect -4886 132586 588810 132618
rect -2966 129454 586890 129486
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 69128 129454
rect 69364 129218 164192 129454
rect 164428 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 221249 129454
rect 221485 129218 224513 129454
rect 224749 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 272249 129454
rect 272485 129218 275513 129454
rect 275749 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect -2966 129134 586890 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 69128 129134
rect 69364 128898 164192 129134
rect 164428 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 221249 129134
rect 221485 128898 224513 129134
rect 224749 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 272249 129134
rect 272485 128898 275513 129134
rect 275749 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect -2966 128866 586890 128898
rect -8726 122614 592650 122646
rect -8726 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 192986 122614
rect 193222 122378 193306 122614
rect 193542 122378 264986 122614
rect 265222 122378 265306 122614
rect 265542 122378 300986 122614
rect 301222 122378 301306 122614
rect 301542 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 444986 122614
rect 445222 122378 445306 122614
rect 445542 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 592650 122614
rect -8726 122294 592650 122378
rect -8726 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 192986 122294
rect 193222 122058 193306 122294
rect 193542 122058 264986 122294
rect 265222 122058 265306 122294
rect 265542 122058 300986 122294
rect 301222 122058 301306 122294
rect 301542 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 444986 122294
rect 445222 122058 445306 122294
rect 445542 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 592650 122294
rect -8726 122026 592650 122058
rect -6806 118894 590730 118926
rect -6806 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 189266 118894
rect 189502 118658 189586 118894
rect 189822 118658 261266 118894
rect 261502 118658 261586 118894
rect 261822 118658 297266 118894
rect 297502 118658 297586 118894
rect 297822 118658 333266 118894
rect 333502 118658 333586 118894
rect 333822 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 441266 118894
rect 441502 118658 441586 118894
rect 441822 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 590730 118894
rect -6806 118574 590730 118658
rect -6806 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 189266 118574
rect 189502 118338 189586 118574
rect 189822 118338 261266 118574
rect 261502 118338 261586 118574
rect 261822 118338 297266 118574
rect 297502 118338 297586 118574
rect 297822 118338 333266 118574
rect 333502 118338 333586 118574
rect 333822 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 441266 118574
rect 441502 118338 441586 118574
rect 441822 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 590730 118574
rect -6806 118306 590730 118338
rect -4886 115174 588810 115206
rect -4886 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 185546 115174
rect 185782 114938 185866 115174
rect 186102 114938 257546 115174
rect 257782 114938 257866 115174
rect 258102 114938 293546 115174
rect 293782 114938 293866 115174
rect 294102 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 588810 115174
rect -4886 114854 588810 114938
rect -4886 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 185546 114854
rect 185782 114618 185866 114854
rect 186102 114618 257546 114854
rect 257782 114618 257866 114854
rect 258102 114618 293546 114854
rect 293782 114618 293866 114854
rect 294102 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 588810 114854
rect -4886 114586 588810 114618
rect -2966 111454 586890 111486
rect -2966 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 69808 111454
rect 70044 111218 163512 111454
rect 163748 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 219617 111454
rect 219853 111218 222881 111454
rect 223117 111218 226145 111454
rect 226381 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 270617 111454
rect 270853 111218 273881 111454
rect 274117 111218 277145 111454
rect 277381 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 586890 111454
rect -2966 111134 586890 111218
rect -2966 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 69808 111134
rect 70044 110898 163512 111134
rect 163748 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 219617 111134
rect 219853 110898 222881 111134
rect 223117 110898 226145 111134
rect 226381 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 270617 111134
rect 270853 110898 273881 111134
rect 274117 110898 277145 111134
rect 277381 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 586890 111134
rect -2966 110866 586890 110898
rect -8726 104614 592650 104646
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 174986 104614
rect 175222 104378 175306 104614
rect 175542 104378 210986 104614
rect 211222 104378 211306 104614
rect 211542 104378 246986 104614
rect 247222 104378 247306 104614
rect 247542 104378 282986 104614
rect 283222 104378 283306 104614
rect 283542 104378 318986 104614
rect 319222 104378 319306 104614
rect 319542 104378 354986 104614
rect 355222 104378 355306 104614
rect 355542 104378 390986 104614
rect 391222 104378 391306 104614
rect 391542 104378 426986 104614
rect 427222 104378 427306 104614
rect 427542 104378 462986 104614
rect 463222 104378 463306 104614
rect 463542 104378 498986 104614
rect 499222 104378 499306 104614
rect 499542 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect -8726 104294 592650 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 174986 104294
rect 175222 104058 175306 104294
rect 175542 104058 210986 104294
rect 211222 104058 211306 104294
rect 211542 104058 246986 104294
rect 247222 104058 247306 104294
rect 247542 104058 282986 104294
rect 283222 104058 283306 104294
rect 283542 104058 318986 104294
rect 319222 104058 319306 104294
rect 319542 104058 354986 104294
rect 355222 104058 355306 104294
rect 355542 104058 390986 104294
rect 391222 104058 391306 104294
rect 391542 104058 426986 104294
rect 427222 104058 427306 104294
rect 427542 104058 462986 104294
rect 463222 104058 463306 104294
rect 463542 104058 498986 104294
rect 499222 104058 499306 104294
rect 499542 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect -8726 104026 592650 104058
rect -6806 100894 590730 100926
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 63266 100894
rect 63502 100658 63586 100894
rect 63822 100658 171266 100894
rect 171502 100658 171586 100894
rect 171822 100658 207266 100894
rect 207502 100658 207586 100894
rect 207822 100658 243266 100894
rect 243502 100658 243586 100894
rect 243822 100658 315266 100894
rect 315502 100658 315586 100894
rect 315822 100658 351266 100894
rect 351502 100658 351586 100894
rect 351822 100658 387266 100894
rect 387502 100658 387586 100894
rect 387822 100658 423266 100894
rect 423502 100658 423586 100894
rect 423822 100658 459266 100894
rect 459502 100658 459586 100894
rect 459822 100658 495266 100894
rect 495502 100658 495586 100894
rect 495822 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect -6806 100574 590730 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 63266 100574
rect 63502 100338 63586 100574
rect 63822 100338 171266 100574
rect 171502 100338 171586 100574
rect 171822 100338 207266 100574
rect 207502 100338 207586 100574
rect 207822 100338 243266 100574
rect 243502 100338 243586 100574
rect 243822 100338 315266 100574
rect 315502 100338 315586 100574
rect 315822 100338 351266 100574
rect 351502 100338 351586 100574
rect 351822 100338 387266 100574
rect 387502 100338 387586 100574
rect 387822 100338 423266 100574
rect 423502 100338 423586 100574
rect 423822 100338 459266 100574
rect 459502 100338 459586 100574
rect 459822 100338 495266 100574
rect 495502 100338 495586 100574
rect 495822 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect -6806 100306 590730 100338
rect -4886 97174 588810 97206
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 59546 97174
rect 59782 96938 59866 97174
rect 60102 96938 167546 97174
rect 167782 96938 167866 97174
rect 168102 96938 203546 97174
rect 203782 96938 203866 97174
rect 204102 96938 239546 97174
rect 239782 96938 239866 97174
rect 240102 96938 311546 97174
rect 311782 96938 311866 97174
rect 312102 96938 347546 97174
rect 347782 96938 347866 97174
rect 348102 96938 383546 97174
rect 383782 96938 383866 97174
rect 384102 96938 419546 97174
rect 419782 96938 419866 97174
rect 420102 96938 455546 97174
rect 455782 96938 455866 97174
rect 456102 96938 491546 97174
rect 491782 96938 491866 97174
rect 492102 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect -4886 96854 588810 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 59546 96854
rect 59782 96618 59866 96854
rect 60102 96618 167546 96854
rect 167782 96618 167866 96854
rect 168102 96618 203546 96854
rect 203782 96618 203866 96854
rect 204102 96618 239546 96854
rect 239782 96618 239866 96854
rect 240102 96618 311546 96854
rect 311782 96618 311866 96854
rect 312102 96618 347546 96854
rect 347782 96618 347866 96854
rect 348102 96618 383546 96854
rect 383782 96618 383866 96854
rect 384102 96618 419546 96854
rect 419782 96618 419866 96854
rect 420102 96618 455546 96854
rect 455782 96618 455866 96854
rect 456102 96618 491546 96854
rect 491782 96618 491866 96854
rect 492102 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect -4886 96586 588810 96618
rect -2966 93454 586890 93486
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect -2966 93134 586890 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect -2966 92866 586890 92898
rect -8726 86614 592650 86646
rect -8726 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 84986 86614
rect 85222 86378 85306 86614
rect 85542 86378 120986 86614
rect 121222 86378 121306 86614
rect 121542 86378 156986 86614
rect 157222 86378 157306 86614
rect 157542 86378 192986 86614
rect 193222 86378 193306 86614
rect 193542 86378 228986 86614
rect 229222 86378 229306 86614
rect 229542 86378 264986 86614
rect 265222 86378 265306 86614
rect 265542 86378 300986 86614
rect 301222 86378 301306 86614
rect 301542 86378 336986 86614
rect 337222 86378 337306 86614
rect 337542 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 592650 86614
rect -8726 86294 592650 86378
rect -8726 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 84986 86294
rect 85222 86058 85306 86294
rect 85542 86058 120986 86294
rect 121222 86058 121306 86294
rect 121542 86058 156986 86294
rect 157222 86058 157306 86294
rect 157542 86058 192986 86294
rect 193222 86058 193306 86294
rect 193542 86058 228986 86294
rect 229222 86058 229306 86294
rect 229542 86058 264986 86294
rect 265222 86058 265306 86294
rect 265542 86058 300986 86294
rect 301222 86058 301306 86294
rect 301542 86058 336986 86294
rect 337222 86058 337306 86294
rect 337542 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 592650 86294
rect -8726 86026 592650 86058
rect -6806 82894 590730 82926
rect -6806 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 81266 82894
rect 81502 82658 81586 82894
rect 81822 82658 117266 82894
rect 117502 82658 117586 82894
rect 117822 82658 153266 82894
rect 153502 82658 153586 82894
rect 153822 82658 189266 82894
rect 189502 82658 189586 82894
rect 189822 82658 225266 82894
rect 225502 82658 225586 82894
rect 225822 82658 261266 82894
rect 261502 82658 261586 82894
rect 261822 82658 297266 82894
rect 297502 82658 297586 82894
rect 297822 82658 333266 82894
rect 333502 82658 333586 82894
rect 333822 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 590730 82894
rect -6806 82574 590730 82658
rect -6806 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 81266 82574
rect 81502 82338 81586 82574
rect 81822 82338 117266 82574
rect 117502 82338 117586 82574
rect 117822 82338 153266 82574
rect 153502 82338 153586 82574
rect 153822 82338 189266 82574
rect 189502 82338 189586 82574
rect 189822 82338 225266 82574
rect 225502 82338 225586 82574
rect 225822 82338 261266 82574
rect 261502 82338 261586 82574
rect 261822 82338 297266 82574
rect 297502 82338 297586 82574
rect 297822 82338 333266 82574
rect 333502 82338 333586 82574
rect 333822 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 590730 82574
rect -6806 82306 590730 82338
rect -4886 79174 588810 79206
rect -4886 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 77546 79174
rect 77782 78938 77866 79174
rect 78102 78938 113546 79174
rect 113782 78938 113866 79174
rect 114102 78938 149546 79174
rect 149782 78938 149866 79174
rect 150102 78938 185546 79174
rect 185782 78938 185866 79174
rect 186102 78938 221546 79174
rect 221782 78938 221866 79174
rect 222102 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 588810 79174
rect -4886 78854 588810 78938
rect -4886 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 77546 78854
rect 77782 78618 77866 78854
rect 78102 78618 113546 78854
rect 113782 78618 113866 78854
rect 114102 78618 149546 78854
rect 149782 78618 149866 78854
rect 150102 78618 185546 78854
rect 185782 78618 185866 78854
rect 186102 78618 221546 78854
rect 221782 78618 221866 78854
rect 222102 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 588810 78854
rect -4886 78586 588810 78618
rect -2966 75454 586890 75486
rect -2966 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 586890 75454
rect -2966 75134 586890 75218
rect -2966 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 586890 75134
rect -2966 74866 586890 74898
rect -8726 68614 592650 68646
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 66986 68614
rect 67222 68378 67306 68614
rect 67542 68378 102986 68614
rect 103222 68378 103306 68614
rect 103542 68378 138986 68614
rect 139222 68378 139306 68614
rect 139542 68378 174986 68614
rect 175222 68378 175306 68614
rect 175542 68378 210986 68614
rect 211222 68378 211306 68614
rect 211542 68378 246986 68614
rect 247222 68378 247306 68614
rect 247542 68378 282986 68614
rect 283222 68378 283306 68614
rect 283542 68378 318986 68614
rect 319222 68378 319306 68614
rect 319542 68378 354986 68614
rect 355222 68378 355306 68614
rect 355542 68378 390986 68614
rect 391222 68378 391306 68614
rect 391542 68378 426986 68614
rect 427222 68378 427306 68614
rect 427542 68378 462986 68614
rect 463222 68378 463306 68614
rect 463542 68378 498986 68614
rect 499222 68378 499306 68614
rect 499542 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect -8726 68294 592650 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 66986 68294
rect 67222 68058 67306 68294
rect 67542 68058 102986 68294
rect 103222 68058 103306 68294
rect 103542 68058 138986 68294
rect 139222 68058 139306 68294
rect 139542 68058 174986 68294
rect 175222 68058 175306 68294
rect 175542 68058 210986 68294
rect 211222 68058 211306 68294
rect 211542 68058 246986 68294
rect 247222 68058 247306 68294
rect 247542 68058 282986 68294
rect 283222 68058 283306 68294
rect 283542 68058 318986 68294
rect 319222 68058 319306 68294
rect 319542 68058 354986 68294
rect 355222 68058 355306 68294
rect 355542 68058 390986 68294
rect 391222 68058 391306 68294
rect 391542 68058 426986 68294
rect 427222 68058 427306 68294
rect 427542 68058 462986 68294
rect 463222 68058 463306 68294
rect 463542 68058 498986 68294
rect 499222 68058 499306 68294
rect 499542 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect -8726 68026 592650 68058
rect -6806 64894 590730 64926
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 63266 64894
rect 63502 64658 63586 64894
rect 63822 64658 99266 64894
rect 99502 64658 99586 64894
rect 99822 64658 135266 64894
rect 135502 64658 135586 64894
rect 135822 64658 171266 64894
rect 171502 64658 171586 64894
rect 171822 64658 207266 64894
rect 207502 64658 207586 64894
rect 207822 64658 243266 64894
rect 243502 64658 243586 64894
rect 243822 64658 279266 64894
rect 279502 64658 279586 64894
rect 279822 64658 315266 64894
rect 315502 64658 315586 64894
rect 315822 64658 351266 64894
rect 351502 64658 351586 64894
rect 351822 64658 387266 64894
rect 387502 64658 387586 64894
rect 387822 64658 423266 64894
rect 423502 64658 423586 64894
rect 423822 64658 459266 64894
rect 459502 64658 459586 64894
rect 459822 64658 495266 64894
rect 495502 64658 495586 64894
rect 495822 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect -6806 64574 590730 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 63266 64574
rect 63502 64338 63586 64574
rect 63822 64338 99266 64574
rect 99502 64338 99586 64574
rect 99822 64338 135266 64574
rect 135502 64338 135586 64574
rect 135822 64338 171266 64574
rect 171502 64338 171586 64574
rect 171822 64338 207266 64574
rect 207502 64338 207586 64574
rect 207822 64338 243266 64574
rect 243502 64338 243586 64574
rect 243822 64338 279266 64574
rect 279502 64338 279586 64574
rect 279822 64338 315266 64574
rect 315502 64338 315586 64574
rect 315822 64338 351266 64574
rect 351502 64338 351586 64574
rect 351822 64338 387266 64574
rect 387502 64338 387586 64574
rect 387822 64338 423266 64574
rect 423502 64338 423586 64574
rect 423822 64338 459266 64574
rect 459502 64338 459586 64574
rect 459822 64338 495266 64574
rect 495502 64338 495586 64574
rect 495822 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect -6806 64306 590730 64338
rect -4886 61174 588810 61206
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 59546 61174
rect 59782 60938 59866 61174
rect 60102 60938 95546 61174
rect 95782 60938 95866 61174
rect 96102 60938 131546 61174
rect 131782 60938 131866 61174
rect 132102 60938 167546 61174
rect 167782 60938 167866 61174
rect 168102 60938 203546 61174
rect 203782 60938 203866 61174
rect 204102 60938 239546 61174
rect 239782 60938 239866 61174
rect 240102 60938 275546 61174
rect 275782 60938 275866 61174
rect 276102 60938 311546 61174
rect 311782 60938 311866 61174
rect 312102 60938 347546 61174
rect 347782 60938 347866 61174
rect 348102 60938 383546 61174
rect 383782 60938 383866 61174
rect 384102 60938 419546 61174
rect 419782 60938 419866 61174
rect 420102 60938 455546 61174
rect 455782 60938 455866 61174
rect 456102 60938 491546 61174
rect 491782 60938 491866 61174
rect 492102 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect -4886 60854 588810 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 59546 60854
rect 59782 60618 59866 60854
rect 60102 60618 95546 60854
rect 95782 60618 95866 60854
rect 96102 60618 131546 60854
rect 131782 60618 131866 60854
rect 132102 60618 167546 60854
rect 167782 60618 167866 60854
rect 168102 60618 203546 60854
rect 203782 60618 203866 60854
rect 204102 60618 239546 60854
rect 239782 60618 239866 60854
rect 240102 60618 275546 60854
rect 275782 60618 275866 60854
rect 276102 60618 311546 60854
rect 311782 60618 311866 60854
rect 312102 60618 347546 60854
rect 347782 60618 347866 60854
rect 348102 60618 383546 60854
rect 383782 60618 383866 60854
rect 384102 60618 419546 60854
rect 419782 60618 419866 60854
rect 420102 60618 455546 60854
rect 455782 60618 455866 60854
rect 456102 60618 491546 60854
rect 491782 60618 491866 60854
rect 492102 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect -4886 60586 588810 60618
rect -2966 57454 586890 57486
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect -2966 57134 586890 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect -2966 56866 586890 56898
rect -8726 50614 592650 50646
rect -8726 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 592650 50614
rect -8726 50294 592650 50378
rect -8726 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 592650 50294
rect -8726 50026 592650 50058
rect -6806 46894 590730 46926
rect -6806 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 590730 46894
rect -6806 46574 590730 46658
rect -6806 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 590730 46574
rect -6806 46306 590730 46338
rect -4886 43174 588810 43206
rect -4886 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 588810 43174
rect -4886 42854 588810 42938
rect -4886 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 588810 42854
rect -4886 42586 588810 42618
rect -2966 39454 586890 39486
rect -2966 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 586890 39454
rect -2966 39134 586890 39218
rect -2966 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 586890 39134
rect -2966 38866 586890 38898
rect -8726 32614 592650 32646
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect -8726 32294 592650 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect -8726 32026 592650 32058
rect -6806 28894 590730 28926
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect -6806 28574 590730 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect -6806 28306 590730 28338
rect -4886 25174 588810 25206
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect -4886 24854 588810 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect -4886 24586 588810 24618
rect -2966 21454 586890 21486
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect -2966 21134 586890 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect -2966 20866 586890 20898
rect -8726 14614 592650 14646
rect -8726 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 592650 14614
rect -8726 14294 592650 14378
rect -8726 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 592650 14294
rect -8726 14026 592650 14058
rect -6806 10894 590730 10926
rect -6806 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 590730 10894
rect -6806 10574 590730 10658
rect -6806 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 590730 10574
rect -6806 10306 590730 10338
rect -4886 7174 588810 7206
rect -4886 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 588810 7174
rect -4886 6854 588810 6938
rect -4886 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 588810 6854
rect -4886 6586 588810 6618
rect -2966 3454 586890 3486
rect -2966 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 586890 3454
rect -2966 3134 586890 3218
rect -2966 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 586890 3134
rect -2966 2866 586890 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use wrapped_spell  wrapped_spell_1
timestamp 1640364529
transform 1 0 68770 0 1 241592
box 0 0 88000 88000
use wrapped_silife  wrapped_silife_4
timestamp 1640364529
transform 1 0 200000 0 1 377600
box -10 0 156249 158393
use wrapped_ppm_decoder  wrapped_ppm_decoder_3
timestamp 1640364529
transform 1 0 68770 0 1 539166
box -10 0 20000 50000
use wrapped_ppm_coder  wrapped_ppm_coder_2
timestamp 1640364529
transform 1 0 68770 0 1 390356
box -10 0 51907 54051
use wrapped_function_generator  wrapped_function_generator_0
timestamp 1640364529
transform 1 0 200200 0 1 240182
box 0 0 44000 44000
use wb_openram_wrapper  wb_openram_wrapper
timestamp 1640364529
transform 1 0 217000 0 1 96000
box 0 144 12000 79688
use wb_bridge_2way  wb_bridge_2way
timestamp 1640364529
transform 1 0 268000 0 1 96000
box 0 0 12000 79688
use sky130_sram_1kbyte_1rw1r_32x256_8  openram_1kB
timestamp 1640364529
transform 1 0 68800 0 1 95100
box 0 0 95956 79500
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 30 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 31 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 32 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 33 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 37 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 38 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 39 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 41 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 42 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 44 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 45 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 46 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 47 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 48 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 49 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 50 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 51 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 52 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 53 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 54 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 55 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 56 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 57 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 58 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 59 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 61 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 62 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 63 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 64 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 65 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 66 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 67 nsew signal tristate
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 68 nsew signal tristate
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 69 nsew signal tristate
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 70 nsew signal tristate
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 71 nsew signal tristate
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 72 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 73 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 74 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 75 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 76 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 77 nsew signal tristate
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 78 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 79 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 80 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 81 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 82 nsew signal tristate
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 83 nsew signal tristate
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 84 nsew signal tristate
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 85 nsew signal tristate
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 86 nsew signal tristate
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 87 nsew signal tristate
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 88 nsew signal tristate
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 89 nsew signal tristate
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 90 nsew signal tristate
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 91 nsew signal tristate
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 92 nsew signal tristate
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 93 nsew signal tristate
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 94 nsew signal tristate
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 95 nsew signal tristate
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 96 nsew signal tristate
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 97 nsew signal tristate
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 98 nsew signal tristate
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 99 nsew signal tristate
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 100 nsew signal tristate
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 101 nsew signal tristate
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 102 nsew signal tristate
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 103 nsew signal tristate
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 104 nsew signal tristate
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 105 nsew signal tristate
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 106 nsew signal tristate
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 107 nsew signal tristate
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 108 nsew signal tristate
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 109 nsew signal tristate
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 110 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 111 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 112 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 113 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 114 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 115 nsew signal tristate
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 116 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 117 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 118 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 119 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 120 nsew signal tristate
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 121 nsew signal tristate
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 122 nsew signal tristate
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 123 nsew signal tristate
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 124 nsew signal tristate
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 125 nsew signal tristate
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 126 nsew signal tristate
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 127 nsew signal tristate
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 128 nsew signal tristate
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 129 nsew signal tristate
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 130 nsew signal tristate
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 131 nsew signal tristate
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 132 nsew signal tristate
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 133 nsew signal tristate
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 134 nsew signal tristate
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 135 nsew signal tristate
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 136 nsew signal tristate
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 137 nsew signal tristate
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 138 nsew signal tristate
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 139 nsew signal tristate
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 140 nsew signal tristate
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 141 nsew signal tristate
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 142 nsew signal tristate
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 271 nsew signal tristate
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 274 nsew signal tristate
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 276 nsew signal tristate
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 278 nsew signal tristate
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 279 nsew signal tristate
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 282 nsew signal tristate
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 283 nsew signal tristate
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 284 nsew signal tristate
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 287 nsew signal tristate
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 290 nsew signal tristate
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 292 nsew signal tristate
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 293 nsew signal tristate
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 295 nsew signal tristate
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 296 nsew signal tristate
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 304 nsew signal tristate
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 305 nsew signal tristate
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 306 nsew signal tristate
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 307 nsew signal tristate
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 311 nsew signal tristate
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 312 nsew signal tristate
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 313 nsew signal tristate
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 316 nsew signal tristate
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 322 nsew signal tristate
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 323 nsew signal tristate
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 326 nsew signal tristate
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 330 nsew signal tristate
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 332 nsew signal tristate
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 333 nsew signal tristate
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 335 nsew signal tristate
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 336 nsew signal tristate
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 343 nsew signal tristate
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 345 nsew signal tristate
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 347 nsew signal tristate
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 352 nsew signal tristate
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 356 nsew signal tristate
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 358 nsew signal tristate
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 361 nsew signal tristate
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 362 nsew signal tristate
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 374 nsew signal tristate
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 376 nsew signal tristate
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 378 nsew signal tristate
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 379 nsew signal tristate
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 380 nsew signal tristate
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 383 nsew signal tristate
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 384 nsew signal tristate
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 386 nsew signal tristate
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 387 nsew signal tristate
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 396 nsew signal tristate
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 397 nsew signal tristate
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 404 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 407 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 410 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 411 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 414 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 416 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 421 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 422 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 424 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 428 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 429 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 430 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 432 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 433 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 435 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 436 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 438 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 441 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 442 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 443 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 445 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 449 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 451 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 452 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 454 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 455 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 457 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 458 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 461 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 462 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 463 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 464 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 466 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 468 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 472 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 473 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 476 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 478 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 479 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 482 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 483 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 488 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 493 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 494 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 495 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 496 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 497 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 498 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 499 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 500 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 504 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 505 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 506 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 507 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 508 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 509 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 510 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 512 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 515 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 518 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 520 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 522 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 526 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 527 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 528 nsew signal tristate
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 529 nsew signal tristate
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 530 nsew signal tristate
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 531 nsew power input
rlabel metal5 s -2966 2866 586890 3486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 38866 586890 39486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 74866 586890 75486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 110866 586890 111486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 146866 586890 147486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 182866 586890 183486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 218866 586890 219486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 254866 586890 255486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 290866 586890 291486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 326866 586890 327486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 362866 586890 363486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 398866 586890 399486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 434866 586890 435486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 470866 586890 471486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 506866 586890 507486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 542866 586890 543486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 578866 586890 579486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 614866 586890 615486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 650866 586890 651486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 686866 586890 687486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 -1894 74414 93100 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 -1894 110414 93100 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 -1894 146414 93100 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 -1894 218414 94000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 178000 218414 238182 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 176600 74414 239592 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 176600 110414 239592 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 176600 146414 239592 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 286182 218414 375600 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 -1894 254414 375600 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 -1894 290414 375600 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 -1894 326414 375600 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 331592 74414 388356 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 331592 110414 388356 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 446407 74414 537166 6 vccd1
port 531 nsew power input
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 531 nsew power input
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 1794 -1894 2414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 -1894 38414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 591166 74414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 446407 110414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 331592 146414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 -1894 182414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 537993 218414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 537993 254414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 537993 290414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 537993 326414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 -1894 362414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 -1894 398414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 -1894 434414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 -1894 470414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 -1894 506414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 -1894 542414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 577794 -1894 578414 705830 6 vccd1
port 531 nsew power input
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 532 nsew power input
rlabel metal5 s -4886 6586 588810 7206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 42586 588810 43206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 78586 588810 79206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 114586 588810 115206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 150586 588810 151206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 186586 588810 187206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 222586 588810 223206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 258586 588810 259206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 294586 588810 295206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 330586 588810 331206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 366586 588810 367206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 402586 588810 403206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 438586 588810 439206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 474586 588810 475206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 510586 588810 511206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 546586 588810 547206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 582586 588810 583206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 618586 588810 619206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 654586 588810 655206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 690586 588810 691206 6 vccd2
port 532 nsew power input
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 -3814 78134 93100 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 -3814 114134 93100 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 -3814 150134 93100 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 -3814 222134 94000 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 178000 222134 238182 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 176600 78134 239592 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 176600 114134 239592 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 176600 150134 239592 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 286182 222134 375600 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 -3814 258134 375600 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 -3814 294134 375600 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 -3814 330134 375600 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 331592 78134 388356 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 331592 114134 388356 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 446407 78134 537166 6 vccd2
port 532 nsew power input
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 532 nsew power input
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 5514 -3814 6134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 41514 -3814 42134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 591166 78134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 446407 114134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 331592 150134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 -3814 186134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 537993 222134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 537993 258134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 537993 294134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 537993 330134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 -3814 366134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 -3814 402134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 -3814 438134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 -3814 474134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 -3814 510134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 545514 -3814 546134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 581514 -3814 582134 707750 6 vccd2
port 532 nsew power input
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 533 nsew power input
rlabel metal5 s -6806 10306 590730 10926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 46306 590730 46926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 82306 590730 82926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 118306 590730 118926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 154306 590730 154926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 190306 590730 190926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 226306 590730 226926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 262306 590730 262926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 298306 590730 298926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 334306 590730 334926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 370306 590730 370926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 406306 590730 406926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 442306 590730 442926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 478306 590730 478926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 514306 590730 514926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 550306 590730 550926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 586306 590730 586926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 622306 590730 622926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 658306 590730 658926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 694306 590730 694926 6 vdda1
port 533 nsew power input
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 -5734 81854 93100 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 -5734 117854 93100 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 -5734 153854 93100 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 -5734 225854 94000 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 178000 225854 238182 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 176600 81854 239592 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 176600 117854 239592 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 176600 153854 239592 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 286182 225854 375600 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 -5734 261854 375600 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 -5734 297854 375600 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 -5734 333854 375600 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 331592 81854 388356 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 331592 117854 388356 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 446407 81854 537166 6 vdda1
port 533 nsew power input
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 533 nsew power input
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 9234 -5734 9854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 45234 -5734 45854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 591166 81854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 446407 117854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 331592 153854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 -5734 189854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 537993 225854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 537993 261854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 537993 297854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 537993 333854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 -5734 369854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 -5734 405854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 -5734 441854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 -5734 477854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 -5734 513854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 549234 -5734 549854 709670 6 vdda1
port 533 nsew power input
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 534 nsew power input
rlabel metal5 s -8726 14026 592650 14646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 50026 592650 50646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 86026 592650 86646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 122026 592650 122646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 158026 592650 158646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 194026 592650 194646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 230026 592650 230646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 266026 592650 266646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 302026 592650 302646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 338026 592650 338646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 374026 592650 374646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 410026 592650 410646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 446026 592650 446646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 482026 592650 482646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 518026 592650 518646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 554026 592650 554646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 590026 592650 590646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 626026 592650 626646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 662026 592650 662646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 698026 592650 698646 6 vdda2
port 534 nsew power input
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 -7654 85574 93100 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 -7654 121574 93100 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 -7654 157574 93100 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 -7654 229574 94000 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 178000 229574 238182 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 176600 85574 239592 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 176600 121574 239592 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 176600 157574 239592 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 286182 229574 375600 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 -7654 265574 375600 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 -7654 301574 375600 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 -7654 337574 375600 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 331592 85574 388356 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 331592 121574 388356 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 446407 85574 537166 6 vdda2
port 534 nsew power input
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 534 nsew power input
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 12954 -7654 13574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 48954 -7654 49574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 591166 85574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 446407 121574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 331592 157574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 -7654 193574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 537993 229574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 537993 265574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 537993 301574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 537993 337574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 -7654 373574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 -7654 409574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 -7654 445574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 -7654 481574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 -7654 517574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 552954 -7654 553574 711590 6 vdda2
port 534 nsew power input
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 28306 590730 28926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 64306 590730 64926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 100306 590730 100926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 136306 590730 136926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 172306 590730 172926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 208306 590730 208926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 244306 590730 244926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 280306 590730 280926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 316306 590730 316926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 352306 590730 352926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 388306 590730 388926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 424306 590730 424926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 460306 590730 460926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 496306 590730 496926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 532306 590730 532926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 568306 590730 568926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 604306 590730 604926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 640306 590730 640926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 676306 590730 676926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 -5734 99854 93100 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 -5734 135854 93100 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 -5734 279854 94000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 -5734 207854 238182 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 -5734 243854 238182 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 176600 99854 239592 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 176600 135854 239592 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 286182 207854 375600 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 286182 243854 375600 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 178000 279854 375600 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 -5734 315854 375600 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 -5734 351854 375600 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 331592 99854 388356 6 vssa1
port 535 nsew ground input
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 535 nsew ground input
rlabel metal4 s 27234 -5734 27854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 -5734 63854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 446407 99854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 331592 135854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 -5734 171854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 537993 207854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 537993 243854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 537993 279854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 537993 315854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 537993 351854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 -5734 387854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 -5734 423854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 -5734 459854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 -5734 495854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 -5734 531854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 567234 -5734 567854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 32026 592650 32646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 68026 592650 68646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 104026 592650 104646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 140026 592650 140646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 176026 592650 176646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 212026 592650 212646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 248026 592650 248646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 284026 592650 284646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 320026 592650 320646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 356026 592650 356646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 392026 592650 392646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 428026 592650 428646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 464026 592650 464646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 500026 592650 500646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 536026 592650 536646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 572026 592650 572646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 608026 592650 608646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 644026 592650 644646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 680026 592650 680646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 -7654 67574 93100 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 -7654 103574 93100 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 -7654 139574 93100 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 -7654 211574 238182 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 176600 67574 239592 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 176600 103574 239592 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 176600 139574 239592 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 286182 211574 375600 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 -7654 247574 375600 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 -7654 283574 375600 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 -7654 319574 375600 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 -7654 355574 375600 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 331592 67574 388356 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 331592 103574 388356 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 446407 67574 537166 6 vssa2
port 536 nsew ground input
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 536 nsew ground input
rlabel metal4 s 30954 -7654 31574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 591166 67574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 446407 103574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 331592 139574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 -7654 175574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 537993 211574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 537993 247574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 537993 283574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 537993 319574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 537993 355574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 -7654 391574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 -7654 427574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 -7654 463574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 -7654 499574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 -7654 535574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 570954 -7654 571574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 20866 586890 21486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 56866 586890 57486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 92866 586890 93486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 128866 586890 129486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 164866 586890 165486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 200866 586890 201486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 236866 586890 237486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 272866 586890 273486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 308866 586890 309486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 344866 586890 345486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 380866 586890 381486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 416866 586890 417486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 452866 586890 453486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 488866 586890 489486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 524866 586890 525486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 560866 586890 561486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 596866 586890 597486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 632866 586890 633486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 668866 586890 669486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 -1894 92414 93100 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 -1894 128414 93100 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 -1894 164414 93100 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 -1894 272414 94000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 -1894 200414 238182 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 -1894 236414 238182 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 176600 92414 239592 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 176600 128414 239592 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 286182 200414 375600 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 286182 236414 375600 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 178000 272414 375600 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 -1894 308414 375600 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 -1894 344414 375600 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 331592 92414 388356 6 vssd1
port 537 nsew ground input
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 537 nsew ground input
rlabel metal4 s 19794 -1894 20414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 -1894 56414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 446407 92414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 331592 128414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 176600 164414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 537993 200414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 537993 236414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 537993 272414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 537993 308414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 537993 344414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 -1894 380414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 -1894 416414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 -1894 452414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 -1894 488414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 523794 -1894 524414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 559794 -1894 560414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 24586 588810 25206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 60586 588810 61206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 96586 588810 97206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 132586 588810 133206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 168586 588810 169206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 204586 588810 205206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 240586 588810 241206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 276586 588810 277206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 312586 588810 313206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 348586 588810 349206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 384586 588810 385206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 420586 588810 421206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 456586 588810 457206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 492586 588810 493206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 528586 588810 529206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 564586 588810 565206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 600586 588810 601206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 636586 588810 637206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 672586 588810 673206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 -3814 96134 93100 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 -3814 132134 93100 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 -3814 276134 94000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 -3814 204134 238182 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 -3814 240134 238182 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 176600 96134 239592 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 176600 132134 239592 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 286182 204134 375600 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 286182 240134 375600 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 178000 276134 375600 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 -3814 312134 375600 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 -3814 348134 375600 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 331592 96134 388356 6 vssd2
port 538 nsew ground input
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 538 nsew ground input
rlabel metal4 s 23514 -3814 24134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 -3814 60134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 446407 96134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 331592 132134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 -3814 168134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 537993 204134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 537993 240134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 537993 276134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 537993 312134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 537993 348134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 -3814 384134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 -3814 420134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 -3814 456134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 -3814 492134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 -3814 528134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 563514 -3814 564134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 539 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 540 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 541 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 542 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 543 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 544 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 545 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 546 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 547 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 548 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 549 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 550 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 551 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 552 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 553 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 554 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 555 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 556 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 557 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 558 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 559 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 560 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 561 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 562 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 563 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 564 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 565 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 566 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 567 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 568 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 569 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 570 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 571 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 572 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 573 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 574 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 575 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 576 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 577 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 578 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 579 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 580 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 581 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 582 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 583 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 584 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 585 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 586 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 587 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 588 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 589 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 590 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 591 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 592 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 593 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 594 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 595 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 596 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 597 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 598 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 599 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 600 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 601 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 602 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 603 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 604 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 605 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 606 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 607 nsew signal tristate
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 608 nsew signal tristate
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 609 nsew signal tristate
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 610 nsew signal tristate
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 611 nsew signal tristate
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 612 nsew signal tristate
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 613 nsew signal tristate
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 614 nsew signal tristate
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 615 nsew signal tristate
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 616 nsew signal tristate
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 617 nsew signal tristate
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 618 nsew signal tristate
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 619 nsew signal tristate
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 620 nsew signal tristate
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 621 nsew signal tristate
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 622 nsew signal tristate
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 623 nsew signal tristate
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 624 nsew signal tristate
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 625 nsew signal tristate
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 626 nsew signal tristate
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 627 nsew signal tristate
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 628 nsew signal tristate
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 629 nsew signal tristate
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 630 nsew signal tristate
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 631 nsew signal tristate
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 632 nsew signal tristate
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 633 nsew signal tristate
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 634 nsew signal tristate
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 635 nsew signal tristate
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 636 nsew signal tristate
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 637 nsew signal tristate
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 638 nsew signal tristate
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 639 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 640 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 641 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 642 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 643 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
