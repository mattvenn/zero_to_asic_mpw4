magic
tech sky130A
magscale 1 2
timestamp 1640693535
<< metal1 >>
rect 331214 702992 331220 703044
rect 331272 703032 331278 703044
rect 332502 703032 332508 703044
rect 331272 703004 332508 703032
rect 331272 702992 331278 703004
rect 332502 702992 332508 703004
rect 332560 702992 332566 703044
rect 62022 702924 62028 702976
rect 62080 702964 62086 702976
rect 267642 702964 267648 702976
rect 62080 702936 267648 702964
rect 62080 702924 62086 702936
rect 267642 702924 267648 702936
rect 267700 702924 267706 702976
rect 283834 702924 283840 702976
rect 283892 702964 283898 702976
rect 351914 702964 351920 702976
rect 283892 702936 351920 702964
rect 283892 702924 283898 702936
rect 351914 702924 351920 702936
rect 351972 702924 351978 702976
rect 202782 702856 202788 702908
rect 202840 702896 202846 702908
rect 273254 702896 273260 702908
rect 202840 702868 273260 702896
rect 202840 702856 202846 702868
rect 273254 702856 273260 702868
rect 273312 702856 273318 702908
rect 276658 702856 276664 702908
rect 276716 702896 276722 702908
rect 478506 702896 478512 702908
rect 276716 702868 478512 702896
rect 276716 702856 276722 702868
rect 478506 702856 478512 702868
rect 478564 702856 478570 702908
rect 281534 702828 281540 702840
rect 171106 702800 281540 702828
rect 67634 702652 67640 702704
rect 67692 702692 67698 702704
rect 170306 702692 170312 702704
rect 67692 702664 170312 702692
rect 67692 702652 67698 702664
rect 170306 702652 170312 702664
rect 170364 702692 170370 702704
rect 171106 702692 171134 702800
rect 281534 702788 281540 702800
rect 281592 702788 281598 702840
rect 349798 702788 349804 702840
rect 349856 702828 349862 702840
rect 494790 702828 494796 702840
rect 349856 702800 494796 702828
rect 349856 702788 349862 702800
rect 494790 702788 494796 702800
rect 494848 702788 494854 702840
rect 233878 702720 233884 702772
rect 233936 702760 233942 702772
rect 397362 702760 397368 702772
rect 233936 702732 397368 702760
rect 233936 702720 233942 702732
rect 397362 702720 397368 702732
rect 397420 702720 397426 702772
rect 170364 702664 171134 702692
rect 170364 702652 170370 702664
rect 191742 702652 191748 702704
rect 191800 702692 191806 702704
rect 364978 702692 364984 702704
rect 191800 702664 364984 702692
rect 191800 702652 191806 702664
rect 364978 702652 364984 702664
rect 365036 702652 365042 702704
rect 378778 702652 378784 702704
rect 378836 702692 378842 702704
rect 462314 702692 462320 702704
rect 378836 702664 462320 702692
rect 378836 702652 378842 702664
rect 462314 702652 462320 702664
rect 462372 702652 462378 702704
rect 24302 702584 24308 702636
rect 24360 702624 24366 702636
rect 79318 702624 79324 702636
rect 24360 702596 79324 702624
rect 24360 702584 24366 702596
rect 79318 702584 79324 702596
rect 79376 702584 79382 702636
rect 95142 702584 95148 702636
rect 95200 702624 95206 702636
rect 300118 702624 300124 702636
rect 95200 702596 300124 702624
rect 95200 702584 95206 702596
rect 300118 702584 300124 702596
rect 300176 702624 300182 702636
rect 300762 702624 300768 702636
rect 300176 702596 300768 702624
rect 300176 702584 300182 702596
rect 300762 702584 300768 702596
rect 300820 702584 300826 702636
rect 359458 702584 359464 702636
rect 359516 702624 359522 702636
rect 543458 702624 543464 702636
rect 359516 702596 543464 702624
rect 359516 702584 359522 702596
rect 543458 702584 543464 702596
rect 543516 702584 543522 702636
rect 88242 702516 88248 702568
rect 88300 702556 88306 702568
rect 235166 702556 235172 702568
rect 88300 702528 235172 702556
rect 88300 702516 88306 702528
rect 235166 702516 235172 702528
rect 235224 702516 235230 702568
rect 264238 702516 264244 702568
rect 264296 702556 264302 702568
rect 559650 702556 559656 702568
rect 264296 702528 559656 702556
rect 264296 702516 264302 702528
rect 559650 702516 559656 702528
rect 559708 702516 559714 702568
rect 8110 702448 8116 702500
rect 8168 702488 8174 702500
rect 88794 702488 88800 702500
rect 8168 702460 88800 702488
rect 8168 702448 8174 702460
rect 88794 702448 88800 702460
rect 88852 702448 88858 702500
rect 99282 702448 99288 702500
rect 99340 702488 99346 702500
rect 527174 702488 527180 702500
rect 99340 702460 527180 702488
rect 99340 702448 99346 702460
rect 527174 702448 527180 702460
rect 527232 702448 527238 702500
rect 124858 700340 124864 700392
rect 124916 700380 124922 700392
rect 137830 700380 137836 700392
rect 124916 700352 137836 700380
rect 124916 700340 124922 700352
rect 137830 700340 137836 700352
rect 137888 700340 137894 700392
rect 75178 700272 75184 700324
rect 75236 700312 75242 700324
rect 105446 700312 105452 700324
rect 75236 700284 105452 700312
rect 75236 700272 75242 700284
rect 105446 700272 105452 700284
rect 105504 700272 105510 700324
rect 128998 700272 129004 700324
rect 129056 700312 129062 700324
rect 218974 700312 218980 700324
rect 129056 700284 218980 700312
rect 129056 700272 129062 700284
rect 218974 700272 218980 700284
rect 219032 700272 219038 700324
rect 300762 700272 300768 700324
rect 300820 700312 300826 700324
rect 341518 700312 341524 700324
rect 300820 700284 341524 700312
rect 300820 700272 300826 700284
rect 341518 700272 341524 700284
rect 341576 700272 341582 700324
rect 342898 700272 342904 700324
rect 342956 700312 342962 700324
rect 348786 700312 348792 700324
rect 342956 700284 348792 700312
rect 342956 700272 342962 700284
rect 348786 700272 348792 700284
rect 348844 700272 348850 700324
rect 382918 700272 382924 700324
rect 382976 700312 382982 700324
rect 429838 700312 429844 700324
rect 382976 700284 429844 700312
rect 382976 700272 382982 700284
rect 429838 700272 429844 700284
rect 429896 700272 429902 700324
rect 66162 699660 66168 699712
rect 66220 699700 66226 699712
rect 72970 699700 72976 699712
rect 66220 699672 72976 699700
rect 66220 699660 66226 699672
rect 72970 699660 72976 699672
rect 73028 699660 73034 699712
rect 86218 699660 86224 699712
rect 86276 699700 86282 699712
rect 89162 699700 89168 699712
rect 86276 699672 89168 699700
rect 86276 699660 86282 699672
rect 89162 699660 89168 699672
rect 89220 699660 89226 699712
rect 3418 683136 3424 683188
rect 3476 683176 3482 683188
rect 21358 683176 21364 683188
rect 3476 683148 21364 683176
rect 3476 683136 3482 683148
rect 21358 683136 21364 683148
rect 21416 683136 21422 683188
rect 3510 670692 3516 670744
rect 3568 670732 3574 670744
rect 22738 670732 22744 670744
rect 3568 670704 22744 670732
rect 3568 670692 3574 670704
rect 22738 670692 22744 670704
rect 22796 670692 22802 670744
rect 3510 632068 3516 632120
rect 3568 632108 3574 632120
rect 11698 632108 11704 632120
rect 3568 632080 11704 632108
rect 3568 632068 3574 632080
rect 11698 632068 11704 632080
rect 11756 632068 11762 632120
rect 3510 618264 3516 618316
rect 3568 618304 3574 618316
rect 14458 618304 14464 618316
rect 3568 618276 14464 618304
rect 3568 618264 3574 618276
rect 14458 618264 14464 618276
rect 14516 618264 14522 618316
rect 3510 605820 3516 605872
rect 3568 605860 3574 605872
rect 90358 605860 90364 605872
rect 3568 605832 90364 605860
rect 3568 605820 3574 605832
rect 90358 605820 90364 605832
rect 90416 605820 90422 605872
rect 71774 605072 71780 605124
rect 71832 605112 71838 605124
rect 86218 605112 86224 605124
rect 71832 605084 86224 605112
rect 71832 605072 71838 605084
rect 86218 605072 86224 605084
rect 86276 605072 86282 605124
rect 70302 596164 70308 596216
rect 70360 596204 70366 596216
rect 349798 596204 349804 596216
rect 70360 596176 349804 596204
rect 70360 596164 70366 596176
rect 349798 596164 349804 596176
rect 349856 596164 349862 596216
rect 79318 595620 79324 595672
rect 79376 595660 79382 595672
rect 80330 595660 80336 595672
rect 79376 595632 80336 595660
rect 79376 595620 79382 595632
rect 80330 595620 80336 595632
rect 80388 595620 80394 595672
rect 80330 594872 80336 594924
rect 80388 594912 80394 594924
rect 106918 594912 106924 594924
rect 80388 594884 106924 594912
rect 80388 594872 80394 594884
rect 106918 594872 106924 594884
rect 106976 594872 106982 594924
rect 85942 594804 85948 594856
rect 86000 594844 86006 594856
rect 141418 594844 141424 594856
rect 86000 594816 141424 594844
rect 86000 594804 86006 594816
rect 141418 594804 141424 594816
rect 141476 594804 141482 594856
rect 90358 594260 90364 594312
rect 90416 594300 90422 594312
rect 91094 594300 91100 594312
rect 90416 594272 91100 594300
rect 90416 594260 90422 594272
rect 91094 594260 91100 594272
rect 91152 594260 91158 594312
rect 40034 594056 40040 594108
rect 40092 594096 40098 594108
rect 89806 594096 89812 594108
rect 40092 594068 89812 594096
rect 40092 594056 40098 594068
rect 89806 594056 89812 594068
rect 89864 594056 89870 594108
rect 88242 593376 88248 593428
rect 88300 593416 88306 593428
rect 113174 593416 113180 593428
rect 88300 593388 113180 593416
rect 88300 593376 88306 593388
rect 113174 593376 113180 593388
rect 113232 593376 113238 593428
rect 67358 592696 67364 592748
rect 67416 592736 67422 592748
rect 75178 592736 75184 592748
rect 67416 592708 75184 592736
rect 67416 592696 67422 592708
rect 75178 592696 75184 592708
rect 75236 592696 75242 592748
rect 3418 592628 3424 592680
rect 3476 592668 3482 592680
rect 69106 592668 69112 592680
rect 3476 592640 69112 592668
rect 3476 592628 3482 592640
rect 69106 592628 69112 592640
rect 69164 592628 69170 592680
rect 78582 592084 78588 592136
rect 78640 592124 78646 592136
rect 103514 592124 103520 592136
rect 78640 592096 103520 592124
rect 78640 592084 78646 592096
rect 103514 592084 103520 592096
rect 103572 592084 103578 592136
rect 84102 592016 84108 592068
rect 84160 592056 84166 592068
rect 112438 592056 112444 592068
rect 84160 592028 112444 592056
rect 84160 592016 84166 592028
rect 112438 592016 112444 592028
rect 112496 592016 112502 592068
rect 85022 591948 85028 592000
rect 85080 591988 85086 592000
rect 88242 591988 88248 592000
rect 85080 591960 88248 591988
rect 85080 591948 85086 591960
rect 88242 591948 88248 591960
rect 88300 591948 88306 592000
rect 73062 590792 73068 590844
rect 73120 590832 73126 590844
rect 79318 590832 79324 590844
rect 73120 590804 79324 590832
rect 73120 590792 73126 590804
rect 79318 590792 79324 590804
rect 79376 590792 79382 590844
rect 63310 590724 63316 590776
rect 63368 590764 63374 590776
rect 73890 590764 73896 590776
rect 63368 590736 73896 590764
rect 63368 590724 63374 590736
rect 73890 590724 73896 590736
rect 73948 590724 73954 590776
rect 86862 590656 86868 590708
rect 86920 590696 86926 590708
rect 115290 590696 115296 590708
rect 86920 590668 115296 590696
rect 86920 590656 86926 590668
rect 115290 590656 115296 590668
rect 115348 590656 115354 590708
rect 69106 589364 69112 589416
rect 69164 589404 69170 589416
rect 89070 589404 89076 589416
rect 69164 589376 89076 589404
rect 69164 589364 69170 589376
rect 89070 589364 89076 589376
rect 89128 589364 89134 589416
rect 3418 589296 3424 589348
rect 3476 589336 3482 589348
rect 74902 589336 74908 589348
rect 3476 589308 74908 589336
rect 3476 589296 3482 589308
rect 74902 589296 74908 589308
rect 74960 589296 74966 589348
rect 76742 589296 76748 589348
rect 76800 589336 76806 589348
rect 101398 589336 101404 589348
rect 76800 589308 101404 589336
rect 76800 589296 76806 589308
rect 101398 589296 101404 589308
rect 101456 589296 101462 589348
rect 79318 588616 79324 588668
rect 79376 588656 79382 588668
rect 94498 588656 94504 588668
rect 79376 588628 94504 588656
rect 79376 588616 79382 588628
rect 94498 588616 94504 588628
rect 94556 588616 94562 588668
rect 79778 588548 79784 588600
rect 79836 588588 79842 588600
rect 105538 588588 105544 588600
rect 79836 588560 105544 588588
rect 79836 588548 79842 588560
rect 105538 588548 105544 588560
rect 105596 588548 105602 588600
rect 75914 588412 75920 588464
rect 75972 588412 75978 588464
rect 52270 587868 52276 587920
rect 52328 587908 52334 587920
rect 66806 587908 66812 587920
rect 52328 587880 66812 587908
rect 52328 587868 52334 587880
rect 66806 587868 66812 587880
rect 66864 587868 66870 587920
rect 75932 587840 75960 588412
rect 88886 588344 88892 588396
rect 88944 588344 88950 588396
rect 88904 588192 88932 588344
rect 88886 588140 88892 588192
rect 88944 588140 88950 588192
rect 88978 587840 88984 587852
rect 75932 587812 88984 587840
rect 88978 587800 88984 587812
rect 89036 587800 89042 587852
rect 88978 586576 88984 586628
rect 89036 586616 89042 586628
rect 98638 586616 98644 586628
rect 89036 586588 98644 586616
rect 89036 586576 89042 586588
rect 98638 586576 98644 586588
rect 98696 586576 98702 586628
rect 55122 586508 55128 586560
rect 55180 586548 55186 586560
rect 66254 586548 66260 586560
rect 55180 586520 66260 586548
rect 55180 586508 55186 586520
rect 66254 586508 66260 586520
rect 66312 586508 66318 586560
rect 91738 586508 91744 586560
rect 91796 586548 91802 586560
rect 95234 586548 95240 586560
rect 91796 586520 95240 586548
rect 91796 586508 91802 586520
rect 95234 586508 95240 586520
rect 95292 586508 95298 586560
rect 57790 585148 57796 585200
rect 57848 585188 57854 585200
rect 66806 585188 66812 585200
rect 57848 585160 66812 585188
rect 57848 585148 57854 585160
rect 66806 585148 66812 585160
rect 66864 585148 66870 585200
rect 88886 584468 88892 584520
rect 88944 584508 88950 584520
rect 116578 584508 116584 584520
rect 88944 584480 116584 584508
rect 88944 584468 88950 584480
rect 116578 584468 116584 584480
rect 116636 584468 116642 584520
rect 91370 584400 91376 584452
rect 91428 584440 91434 584452
rect 95142 584440 95148 584452
rect 91428 584412 95148 584440
rect 91428 584400 91434 584412
rect 95142 584400 95148 584412
rect 95200 584440 95206 584452
rect 132494 584440 132500 584452
rect 95200 584412 132500 584440
rect 95200 584400 95206 584412
rect 132494 584400 132500 584412
rect 132552 584400 132558 584452
rect 91186 583652 91192 583704
rect 91244 583692 91250 583704
rect 99282 583692 99288 583704
rect 91244 583664 99288 583692
rect 91244 583652 91250 583664
rect 99282 583652 99288 583664
rect 99340 583652 99346 583704
rect 99282 582972 99288 583024
rect 99340 583012 99346 583024
rect 108298 583012 108304 583024
rect 99340 582984 108304 583012
rect 99340 582972 99346 582984
rect 108298 582972 108304 582984
rect 108356 582972 108362 583024
rect 50982 582360 50988 582412
rect 51040 582400 51046 582412
rect 66806 582400 66812 582412
rect 51040 582372 66812 582400
rect 51040 582360 51046 582372
rect 66806 582360 66812 582372
rect 66864 582360 66870 582412
rect 59262 581000 59268 581052
rect 59320 581040 59326 581052
rect 66714 581040 66720 581052
rect 59320 581012 66720 581040
rect 59320 581000 59326 581012
rect 66714 581000 66720 581012
rect 66772 581000 66778 581052
rect 91738 581000 91744 581052
rect 91796 581040 91802 581052
rect 148410 581040 148416 581052
rect 91796 581012 148416 581040
rect 91796 581000 91802 581012
rect 148410 581000 148416 581012
rect 148468 581000 148474 581052
rect 64782 579640 64788 579692
rect 64840 579680 64846 579692
rect 66806 579680 66812 579692
rect 64840 579652 66812 579680
rect 64840 579640 64846 579652
rect 66806 579640 66812 579652
rect 66864 579640 66870 579692
rect 91738 579640 91744 579692
rect 91796 579680 91802 579692
rect 142798 579680 142804 579692
rect 91796 579652 142804 579680
rect 91796 579640 91802 579652
rect 142798 579640 142804 579652
rect 142856 579640 142862 579692
rect 91738 578212 91744 578264
rect 91796 578252 91802 578264
rect 120718 578252 120724 578264
rect 91796 578224 120724 578252
rect 91796 578212 91802 578224
rect 120718 578212 120724 578224
rect 120776 578212 120782 578264
rect 95878 577464 95884 577516
rect 95936 577504 95942 577516
rect 109034 577504 109040 577516
rect 95936 577476 109040 577504
rect 95936 577464 95942 577476
rect 109034 577464 109040 577476
rect 109092 577464 109098 577516
rect 11698 576104 11704 576156
rect 11756 576144 11762 576156
rect 67450 576144 67456 576156
rect 11756 576116 67456 576144
rect 11756 576104 11762 576116
rect 67450 576104 67456 576116
rect 67508 576104 67514 576156
rect 91094 576104 91100 576156
rect 91152 576144 91158 576156
rect 123110 576144 123116 576156
rect 91152 576116 123116 576144
rect 91152 576104 91158 576116
rect 123110 576104 123116 576116
rect 123168 576104 123174 576156
rect 142798 574744 142804 574796
rect 142856 574784 142862 574796
rect 276014 574784 276020 574796
rect 142856 574756 276020 574784
rect 142856 574744 142862 574756
rect 276014 574744 276020 574756
rect 276072 574744 276078 574796
rect 276014 574404 276020 574456
rect 276072 574444 276078 574456
rect 276658 574444 276664 574456
rect 276072 574416 276664 574444
rect 276072 574404 276078 574416
rect 276658 574404 276664 574416
rect 276716 574404 276722 574456
rect 61930 574064 61936 574116
rect 61988 574104 61994 574116
rect 67358 574104 67364 574116
rect 61988 574076 67364 574104
rect 61988 574064 61994 574076
rect 67358 574064 67364 574076
rect 67416 574064 67422 574116
rect 91094 574064 91100 574116
rect 91152 574104 91158 574116
rect 122190 574104 122196 574116
rect 91152 574076 122196 574104
rect 91152 574064 91158 574076
rect 122190 574064 122196 574076
rect 122248 574064 122254 574116
rect 91094 572704 91100 572756
rect 91152 572744 91158 572756
rect 115198 572744 115204 572756
rect 91152 572716 115204 572744
rect 91152 572704 91158 572716
rect 115198 572704 115204 572716
rect 115256 572704 115262 572756
rect 49602 571344 49608 571396
rect 49660 571384 49666 571396
rect 66806 571384 66812 571396
rect 49660 571356 66812 571384
rect 49660 571344 49666 571356
rect 66806 571344 66812 571356
rect 66864 571344 66870 571396
rect 91094 571344 91100 571396
rect 91152 571384 91158 571396
rect 95142 571384 95148 571396
rect 91152 571356 95148 571384
rect 91152 571344 91158 571356
rect 95142 571344 95148 571356
rect 95200 571344 95206 571396
rect 91186 570596 91192 570648
rect 91244 570636 91250 570648
rect 121546 570636 121552 570648
rect 91244 570608 121552 570636
rect 91244 570596 91250 570608
rect 121546 570596 121552 570608
rect 121604 570596 121610 570648
rect 91094 569916 91100 569968
rect 91152 569956 91158 569968
rect 101490 569956 101496 569968
rect 91152 569928 101496 569956
rect 91152 569916 91158 569928
rect 101490 569916 101496 569928
rect 101548 569916 101554 569968
rect 95142 569168 95148 569220
rect 95200 569208 95206 569220
rect 129734 569208 129740 569220
rect 95200 569180 129740 569208
rect 95200 569168 95206 569180
rect 129734 569168 129740 569180
rect 129792 569168 129798 569220
rect 60642 568556 60648 568608
rect 60700 568596 60706 568608
rect 66806 568596 66812 568608
rect 60700 568568 66812 568596
rect 60700 568556 60706 568568
rect 66806 568556 66812 568568
rect 66864 568556 66870 568608
rect 91094 568556 91100 568608
rect 91152 568596 91158 568608
rect 100018 568596 100024 568608
rect 91152 568568 100024 568596
rect 91152 568556 91158 568568
rect 100018 568556 100024 568568
rect 100076 568556 100082 568608
rect 129734 568556 129740 568608
rect 129792 568596 129798 568608
rect 213914 568596 213920 568608
rect 129792 568568 213920 568596
rect 129792 568556 129798 568568
rect 213914 568556 213920 568568
rect 213972 568556 213978 568608
rect 120718 568488 120724 568540
rect 120776 568528 120782 568540
rect 121362 568528 121368 568540
rect 120776 568500 121368 568528
rect 120776 568488 120782 568500
rect 121362 568488 121368 568500
rect 121420 568488 121426 568540
rect 53650 567196 53656 567248
rect 53708 567236 53714 567248
rect 66806 567236 66812 567248
rect 53708 567208 66812 567236
rect 53708 567196 53714 567208
rect 66806 567196 66812 567208
rect 66864 567196 66870 567248
rect 121362 567196 121368 567248
rect 121420 567236 121426 567248
rect 332594 567236 332600 567248
rect 121420 567208 332600 567236
rect 121420 567196 121426 567208
rect 332594 567196 332600 567208
rect 332652 567196 332658 567248
rect 101490 566448 101496 566500
rect 101548 566488 101554 566500
rect 127434 566488 127440 566500
rect 101548 566460 127440 566488
rect 101548 566448 101554 566460
rect 127434 566448 127440 566460
rect 127492 566448 127498 566500
rect 184198 565904 184204 565956
rect 184256 565944 184262 565956
rect 311894 565944 311900 565956
rect 184256 565916 311900 565944
rect 184256 565904 184262 565916
rect 311894 565904 311900 565916
rect 311952 565904 311958 565956
rect 59078 565836 59084 565888
rect 59136 565876 59142 565888
rect 67634 565876 67640 565888
rect 59136 565848 67640 565876
rect 59136 565836 59142 565848
rect 67634 565836 67640 565848
rect 67692 565836 67698 565888
rect 91370 565836 91376 565888
rect 91428 565876 91434 565888
rect 102778 565876 102784 565888
rect 91428 565848 102784 565876
rect 91428 565836 91434 565848
rect 102778 565836 102784 565848
rect 102836 565836 102842 565888
rect 126974 565836 126980 565888
rect 127032 565876 127038 565888
rect 127434 565876 127440 565888
rect 127032 565848 127440 565876
rect 127032 565836 127038 565848
rect 127434 565836 127440 565848
rect 127492 565876 127498 565888
rect 291194 565876 291200 565888
rect 127492 565848 291200 565876
rect 127492 565836 127498 565848
rect 291194 565836 291200 565848
rect 291252 565836 291258 565888
rect 91462 565088 91468 565140
rect 91520 565128 91526 565140
rect 134518 565128 134524 565140
rect 91520 565100 134524 565128
rect 91520 565088 91526 565100
rect 134518 565088 134524 565100
rect 134576 565088 134582 565140
rect 54478 564408 54484 564460
rect 54536 564448 54542 564460
rect 66806 564448 66812 564460
rect 54536 564420 66812 564448
rect 54536 564408 54542 564420
rect 66806 564408 66812 564420
rect 66864 564408 66870 564460
rect 91370 564408 91376 564460
rect 91428 564448 91434 564460
rect 101490 564448 101496 564460
rect 91428 564420 101496 564448
rect 91428 564408 91434 564420
rect 101490 564408 101496 564420
rect 101548 564408 101554 564460
rect 162762 564408 162768 564460
rect 162820 564448 162826 564460
rect 309134 564448 309140 564460
rect 162820 564420 309140 564448
rect 162820 564408 162826 564420
rect 309134 564408 309140 564420
rect 309192 564408 309198 564460
rect 194594 563156 194600 563168
rect 180766 563128 194600 563156
rect 52362 563048 52368 563100
rect 52420 563088 52426 563100
rect 66806 563088 66812 563100
rect 52420 563060 66812 563088
rect 52420 563048 52426 563060
rect 66806 563048 66812 563060
rect 66864 563048 66870 563100
rect 91370 563048 91376 563100
rect 91428 563088 91434 563100
rect 180766 563088 180794 563128
rect 194594 563116 194600 563128
rect 194652 563156 194658 563168
rect 241514 563156 241520 563168
rect 194652 563128 241520 563156
rect 194652 563116 194658 563128
rect 241514 563116 241520 563128
rect 241572 563116 241578 563168
rect 91428 563060 180794 563088
rect 91428 563048 91434 563060
rect 196618 563048 196624 563100
rect 196676 563088 196682 563100
rect 295978 563088 295984 563100
rect 196676 563060 295984 563088
rect 196676 563048 196682 563060
rect 295978 563048 295984 563060
rect 296036 563048 296042 563100
rect 115290 562504 115296 562556
rect 115348 562544 115354 562556
rect 117958 562544 117964 562556
rect 115348 562516 117964 562544
rect 115348 562504 115354 562516
rect 117958 562504 117964 562516
rect 118016 562504 118022 562556
rect 67450 562300 67456 562352
rect 67508 562340 67514 562352
rect 68278 562340 68284 562352
rect 67508 562312 68284 562340
rect 67508 562300 67514 562312
rect 68278 562300 68284 562312
rect 68336 562300 68342 562352
rect 166350 561756 166356 561808
rect 166408 561796 166414 561808
rect 335354 561796 335360 561808
rect 166408 561768 335360 561796
rect 166408 561756 166414 561768
rect 335354 561756 335360 561768
rect 335412 561756 335418 561808
rect 37182 561688 37188 561740
rect 37240 561728 37246 561740
rect 66806 561728 66812 561740
rect 37240 561700 66812 561728
rect 37240 561688 37246 561700
rect 66806 561688 66812 561700
rect 66864 561688 66870 561740
rect 111058 561688 111064 561740
rect 111116 561728 111122 561740
rect 111702 561728 111708 561740
rect 111116 561700 111708 561728
rect 111116 561688 111122 561700
rect 111702 561688 111708 561700
rect 111760 561728 111766 561740
rect 357526 561728 357532 561740
rect 111760 561700 357532 561728
rect 111760 561688 111766 561700
rect 357526 561688 357532 561700
rect 357584 561688 357590 561740
rect 153102 560328 153108 560380
rect 153160 560368 153166 560380
rect 215294 560368 215300 560380
rect 153160 560340 215300 560368
rect 153160 560328 153166 560340
rect 215294 560328 215300 560340
rect 215352 560328 215358 560380
rect 44082 560260 44088 560312
rect 44140 560300 44146 560312
rect 66806 560300 66812 560312
rect 44140 560272 66812 560300
rect 44140 560260 44146 560272
rect 66806 560260 66812 560272
rect 66864 560260 66870 560312
rect 194502 560260 194508 560312
rect 194560 560300 194566 560312
rect 268378 560300 268384 560312
rect 194560 560272 268384 560300
rect 194560 560260 194566 560272
rect 268378 560260 268384 560272
rect 268436 560260 268442 560312
rect 273254 559648 273260 559700
rect 273312 559688 273318 559700
rect 273898 559688 273904 559700
rect 273312 559660 273904 559688
rect 273312 559648 273318 559660
rect 273898 559648 273904 559660
rect 273956 559648 273962 559700
rect 198458 558968 198464 559020
rect 198516 559008 198522 559020
rect 273898 559008 273904 559020
rect 198516 558980 273904 559008
rect 198516 558968 198522 558980
rect 273898 558968 273904 558980
rect 273956 558968 273962 559020
rect 89622 558900 89628 558952
rect 89680 558940 89686 558952
rect 122098 558940 122104 558952
rect 89680 558912 122104 558940
rect 89680 558900 89686 558912
rect 122098 558900 122104 558912
rect 122156 558900 122162 558952
rect 122190 558900 122196 558952
rect 122248 558940 122254 558952
rect 122926 558940 122932 558952
rect 122248 558912 122932 558940
rect 122248 558900 122254 558912
rect 122926 558900 122932 558912
rect 122984 558900 122990 558952
rect 196710 558900 196716 558952
rect 196768 558940 196774 558952
rect 343634 558940 343640 558952
rect 196768 558912 343640 558940
rect 196768 558900 196774 558912
rect 343634 558900 343640 558912
rect 343692 558900 343698 558952
rect 60734 558628 60740 558680
rect 60792 558668 60798 558680
rect 62022 558668 62028 558680
rect 60792 558640 62028 558668
rect 60792 558628 60798 558640
rect 62022 558628 62028 558640
rect 62080 558668 62086 558680
rect 66254 558668 66260 558680
rect 62080 558640 66260 558668
rect 62080 558628 62086 558640
rect 66254 558628 66260 558640
rect 66312 558628 66318 558680
rect 39942 558152 39948 558204
rect 40000 558192 40006 558204
rect 60734 558192 60740 558204
rect 40000 558164 60740 558192
rect 40000 558152 40006 558164
rect 60734 558152 60740 558164
rect 60792 558152 60798 558204
rect 198642 558152 198648 558204
rect 198700 558192 198706 558204
rect 582926 558192 582932 558204
rect 198700 558164 582932 558192
rect 198700 558152 198706 558164
rect 582926 558152 582932 558164
rect 582984 558152 582990 558204
rect 91186 557540 91192 557592
rect 91244 557580 91250 557592
rect 151814 557580 151820 557592
rect 91244 557552 151820 557580
rect 91244 557540 91250 557552
rect 151814 557540 151820 557552
rect 151872 557540 151878 557592
rect 191098 557540 191104 557592
rect 191156 557580 191162 557592
rect 270494 557580 270500 557592
rect 191156 557552 270500 557580
rect 191156 557540 191162 557552
rect 270494 557540 270500 557552
rect 270552 557540 270558 557592
rect 91278 556248 91284 556300
rect 91336 556288 91342 556300
rect 121454 556288 121460 556300
rect 91336 556260 121460 556288
rect 91336 556248 91342 556260
rect 121454 556248 121460 556260
rect 121512 556248 121518 556300
rect 195882 556248 195888 556300
rect 195940 556288 195946 556300
rect 288434 556288 288440 556300
rect 195940 556260 288440 556288
rect 195940 556248 195946 556260
rect 288434 556248 288440 556260
rect 288492 556248 288498 556300
rect 112438 556180 112444 556232
rect 112496 556220 112502 556232
rect 226978 556220 226984 556232
rect 112496 556192 226984 556220
rect 112496 556180 112502 556192
rect 226978 556180 226984 556192
rect 227036 556180 227042 556232
rect 187050 554820 187056 554872
rect 187108 554860 187114 554872
rect 237374 554860 237380 554872
rect 187108 554832 237380 554860
rect 187108 554820 187114 554832
rect 237374 554820 237380 554832
rect 237432 554820 237438 554872
rect 56502 554752 56508 554804
rect 56560 554792 56566 554804
rect 66806 554792 66812 554804
rect 56560 554764 66812 554792
rect 56560 554752 56566 554764
rect 66806 554752 66812 554764
rect 66864 554752 66870 554804
rect 198090 554752 198096 554804
rect 198148 554792 198154 554804
rect 268286 554792 268292 554804
rect 198148 554764 268292 554792
rect 198148 554752 198154 554764
rect 268286 554752 268292 554764
rect 268344 554752 268350 554804
rect 188614 553460 188620 553512
rect 188672 553500 188678 553512
rect 260098 553500 260104 553512
rect 188672 553472 260104 553500
rect 188672 553460 188678 553472
rect 260098 553460 260104 553472
rect 260156 553460 260162 553512
rect 3326 553392 3332 553444
rect 3384 553432 3390 553444
rect 43438 553432 43444 553444
rect 3384 553404 43444 553432
rect 3384 553392 3390 553404
rect 43438 553392 43444 553404
rect 43496 553392 43502 553444
rect 64690 553392 64696 553444
rect 64748 553432 64754 553444
rect 66438 553432 66444 553444
rect 64748 553404 66444 553432
rect 64748 553392 64754 553404
rect 66438 553392 66444 553404
rect 66496 553392 66502 553444
rect 91094 553392 91100 553444
rect 91152 553432 91158 553444
rect 112530 553432 112536 553444
rect 91152 553404 112536 553432
rect 91152 553392 91158 553404
rect 112530 553392 112536 553404
rect 112588 553392 112594 553444
rect 134518 553392 134524 553444
rect 134576 553432 134582 553444
rect 210418 553432 210424 553444
rect 134576 553404 210424 553432
rect 134576 553392 134582 553404
rect 210418 553392 210424 553404
rect 210476 553392 210482 553444
rect 91094 552100 91100 552152
rect 91152 552140 91158 552152
rect 104250 552140 104256 552152
rect 91152 552112 104256 552140
rect 91152 552100 91158 552112
rect 104250 552100 104256 552112
rect 104308 552100 104314 552152
rect 156598 552100 156604 552152
rect 156656 552140 156662 552152
rect 238754 552140 238760 552152
rect 156656 552112 238760 552140
rect 156656 552100 156662 552112
rect 238754 552100 238760 552112
rect 238812 552100 238818 552152
rect 92106 552032 92112 552084
rect 92164 552072 92170 552084
rect 108390 552072 108396 552084
rect 92164 552044 108396 552072
rect 92164 552032 92170 552044
rect 108390 552032 108396 552044
rect 108448 552032 108454 552084
rect 124950 552032 124956 552084
rect 125008 552072 125014 552084
rect 351914 552072 351920 552084
rect 125008 552044 351920 552072
rect 125008 552032 125014 552044
rect 351914 552032 351920 552044
rect 351972 552032 351978 552084
rect 117958 551964 117964 552016
rect 118016 552004 118022 552016
rect 118602 552004 118608 552016
rect 118016 551976 118608 552004
rect 118016 551964 118022 551976
rect 118602 551964 118608 551976
rect 118660 551964 118666 552016
rect 91094 550672 91100 550724
rect 91152 550712 91158 550724
rect 128354 550712 128360 550724
rect 91152 550684 128360 550712
rect 91152 550672 91158 550684
rect 128354 550672 128360 550684
rect 128412 550712 128418 550724
rect 180242 550712 180248 550724
rect 128412 550684 180248 550712
rect 128412 550672 128418 550684
rect 180242 550672 180248 550684
rect 180300 550672 180306 550724
rect 182082 550672 182088 550724
rect 182140 550712 182146 550724
rect 240226 550712 240232 550724
rect 182140 550684 240232 550712
rect 182140 550672 182146 550684
rect 240226 550672 240232 550684
rect 240284 550672 240290 550724
rect 118602 550604 118608 550656
rect 118660 550644 118666 550656
rect 212534 550644 212540 550656
rect 118660 550616 212540 550644
rect 118660 550604 118666 550616
rect 212534 550604 212540 550616
rect 212592 550604 212598 550656
rect 193950 549312 193956 549364
rect 194008 549352 194014 549364
rect 223666 549352 223672 549364
rect 194008 549324 223672 549352
rect 194008 549312 194014 549324
rect 223666 549312 223672 549324
rect 223724 549312 223730 549364
rect 60550 549244 60556 549296
rect 60608 549284 60614 549296
rect 66806 549284 66812 549296
rect 60608 549256 66812 549284
rect 60608 549244 60614 549256
rect 66806 549244 66812 549256
rect 66864 549244 66870 549296
rect 187602 549244 187608 549296
rect 187660 549284 187666 549296
rect 220814 549284 220820 549296
rect 187660 549256 220820 549284
rect 187660 549244 187666 549256
rect 220814 549244 220820 549256
rect 220872 549244 220878 549296
rect 192478 547952 192484 548004
rect 192536 547992 192542 548004
rect 287054 547992 287060 548004
rect 192536 547964 287060 547992
rect 192536 547952 192542 547964
rect 287054 547952 287060 547964
rect 287112 547952 287118 548004
rect 57698 547884 57704 547936
rect 57756 547924 57762 547936
rect 66806 547924 66812 547936
rect 57756 547896 66812 547924
rect 57756 547884 57762 547896
rect 66806 547884 66812 547896
rect 66864 547884 66870 547936
rect 91370 547884 91376 547936
rect 91428 547924 91434 547936
rect 245654 547924 245660 547936
rect 91428 547896 245660 547924
rect 91428 547884 91434 547896
rect 245654 547884 245660 547896
rect 245712 547884 245718 547936
rect 295334 547884 295340 547936
rect 295392 547924 295398 547936
rect 372614 547924 372620 547936
rect 295392 547896 372620 547924
rect 295392 547884 295398 547896
rect 372614 547884 372620 547896
rect 372672 547884 372678 547936
rect 204898 546524 204904 546576
rect 204956 546564 204962 546576
rect 251818 546564 251824 546576
rect 204956 546536 251824 546564
rect 204956 546524 204962 546536
rect 251818 546524 251824 546536
rect 251876 546524 251882 546576
rect 62022 546456 62028 546508
rect 62080 546496 62086 546508
rect 66898 546496 66904 546508
rect 62080 546468 66904 546496
rect 62080 546456 62086 546468
rect 66898 546456 66904 546468
rect 66956 546456 66962 546508
rect 91554 546456 91560 546508
rect 91612 546496 91618 546508
rect 104158 546496 104164 546508
rect 91612 546468 104164 546496
rect 91612 546456 91618 546468
rect 104158 546456 104164 546468
rect 104216 546456 104222 546508
rect 188430 546456 188436 546508
rect 188488 546496 188494 546508
rect 304994 546496 305000 546508
rect 188488 546468 305000 546496
rect 188488 546456 188494 546468
rect 304994 546456 305000 546468
rect 305052 546456 305058 546508
rect 327074 546456 327080 546508
rect 327132 546496 327138 546508
rect 361850 546496 361856 546508
rect 327132 546468 361856 546496
rect 327132 546456 327138 546468
rect 361850 546456 361856 546468
rect 361908 546456 361914 546508
rect 199378 545164 199384 545216
rect 199436 545204 199442 545216
rect 298370 545204 298376 545216
rect 199436 545176 298376 545204
rect 199436 545164 199442 545176
rect 298370 545164 298376 545176
rect 298428 545164 298434 545216
rect 314930 545164 314936 545216
rect 314988 545204 314994 545216
rect 363046 545204 363052 545216
rect 314988 545176 363052 545204
rect 314988 545164 314994 545176
rect 363046 545164 363052 545176
rect 363104 545164 363110 545216
rect 50890 545096 50896 545148
rect 50948 545136 50954 545148
rect 66898 545136 66904 545148
rect 50948 545108 66904 545136
rect 50948 545096 50954 545108
rect 66898 545096 66904 545108
rect 66956 545096 66962 545148
rect 91094 545096 91100 545148
rect 91152 545136 91158 545148
rect 94590 545136 94596 545148
rect 91152 545108 94596 545136
rect 91152 545096 91158 545108
rect 94590 545096 94596 545108
rect 94648 545096 94654 545148
rect 186958 545096 186964 545148
rect 187016 545136 187022 545148
rect 324314 545136 324320 545148
rect 187016 545108 324320 545136
rect 187016 545096 187022 545108
rect 324314 545096 324320 545108
rect 324372 545096 324378 545148
rect 331674 545096 331680 545148
rect 331732 545136 331738 545148
rect 364426 545136 364432 545148
rect 331732 545108 364432 545136
rect 331732 545096 331738 545108
rect 364426 545096 364432 545108
rect 364484 545096 364490 545148
rect 199470 543804 199476 543856
rect 199528 543844 199534 543856
rect 229094 543844 229100 543856
rect 199528 543816 229100 543844
rect 199528 543804 199534 543816
rect 229094 543804 229100 543816
rect 229152 543804 229158 543856
rect 318242 543804 318248 543856
rect 318300 543844 318306 543856
rect 365714 543844 365720 543856
rect 318300 543816 365720 543844
rect 318300 543804 318306 543816
rect 365714 543804 365720 543816
rect 365772 543804 365778 543856
rect 48222 543736 48228 543788
rect 48280 543776 48286 543788
rect 66898 543776 66904 543788
rect 48280 543748 66904 543776
rect 48280 543736 48286 543748
rect 66898 543736 66904 543748
rect 66956 543736 66962 543788
rect 182818 543736 182824 543788
rect 182876 543776 182882 543788
rect 321554 543776 321560 543788
rect 182876 543748 321560 543776
rect 182876 543736 182882 543748
rect 321554 543736 321560 543748
rect 321612 543736 321618 543788
rect 330018 543736 330024 543788
rect 330076 543776 330082 543788
rect 376846 543776 376852 543788
rect 330076 543748 376852 543776
rect 330076 543736 330082 543748
rect 376846 543736 376852 543748
rect 376904 543736 376910 543788
rect 21358 542988 21364 543040
rect 21416 543028 21422 543040
rect 34514 543028 34520 543040
rect 21416 543000 34520 543028
rect 21416 542988 21422 543000
rect 34514 542988 34520 543000
rect 34572 542988 34578 543040
rect 175918 542444 175924 542496
rect 175976 542484 175982 542496
rect 280154 542484 280160 542496
rect 175976 542456 280160 542484
rect 175976 542444 175982 542456
rect 280154 542444 280160 542456
rect 280212 542444 280218 542496
rect 338298 542444 338304 542496
rect 338356 542484 338362 542496
rect 367278 542484 367284 542496
rect 338356 542456 367284 542484
rect 338356 542444 338362 542456
rect 367278 542444 367284 542456
rect 367336 542444 367342 542496
rect 34514 542376 34520 542428
rect 34572 542416 34578 542428
rect 35802 542416 35808 542428
rect 34572 542388 35808 542416
rect 34572 542376 34578 542388
rect 35802 542376 35808 542388
rect 35860 542416 35866 542428
rect 66898 542416 66904 542428
rect 35860 542388 66904 542416
rect 35860 542376 35866 542388
rect 66898 542376 66904 542388
rect 66956 542376 66962 542428
rect 91094 542376 91100 542428
rect 91152 542416 91158 542428
rect 95878 542416 95884 542428
rect 91152 542388 95884 542416
rect 91152 542376 91158 542388
rect 95878 542376 95884 542388
rect 95936 542376 95942 542428
rect 133138 542376 133144 542428
rect 133196 542416 133202 542428
rect 357434 542416 357440 542428
rect 133196 542388 357440 542416
rect 133196 542376 133202 542388
rect 357434 542376 357440 542388
rect 357492 542376 357498 542428
rect 22738 541628 22744 541680
rect 22796 541668 22802 541680
rect 66990 541668 66996 541680
rect 22796 541640 66996 541668
rect 22796 541628 22802 541640
rect 66990 541628 66996 541640
rect 67048 541668 67054 541680
rect 67266 541668 67272 541680
rect 67048 541640 67272 541668
rect 67048 541628 67054 541640
rect 67266 541628 67272 541640
rect 67324 541628 67330 541680
rect 91094 541628 91100 541680
rect 91152 541668 91158 541680
rect 124858 541668 124864 541680
rect 91152 541640 124864 541668
rect 91152 541628 91158 541640
rect 124858 541628 124864 541640
rect 124916 541668 124922 541680
rect 131574 541668 131580 541680
rect 124916 541640 131580 541668
rect 124916 541628 124922 541640
rect 131574 541628 131580 541640
rect 131632 541628 131638 541680
rect 131114 541016 131120 541068
rect 131172 541056 131178 541068
rect 131574 541056 131580 541068
rect 131172 541028 131580 541056
rect 131172 541016 131178 541028
rect 131574 541016 131580 541028
rect 131632 541056 131638 541068
rect 258442 541056 258448 541068
rect 131632 541028 258448 541056
rect 131632 541016 131638 541028
rect 258442 541016 258448 541028
rect 258500 541016 258506 541068
rect 88886 540948 88892 541000
rect 88944 540988 88950 541000
rect 266354 540988 266360 541000
rect 88944 540960 266360 540988
rect 88944 540948 88950 540960
rect 266354 540948 266360 540960
rect 266412 540948 266418 541000
rect 324314 540880 324320 540932
rect 324372 540920 324378 540932
rect 324958 540920 324964 540932
rect 324372 540892 324964 540920
rect 324372 540880 324378 540892
rect 324958 540880 324964 540892
rect 325016 540920 325022 540932
rect 342898 540920 342904 540932
rect 325016 540892 342904 540920
rect 325016 540880 325022 540892
rect 342898 540880 342904 540892
rect 342956 540880 342962 540932
rect 3418 540200 3424 540252
rect 3476 540240 3482 540252
rect 3476 540212 64874 540240
rect 3476 540200 3482 540212
rect 64846 539696 64874 540212
rect 67542 539724 67548 539776
rect 67600 539764 67606 539776
rect 67600 539736 71912 539764
rect 67600 539724 67606 539736
rect 64846 539668 69428 539696
rect 69400 539640 69428 539668
rect 71884 539640 71912 539736
rect 91094 539656 91100 539708
rect 91152 539696 91158 539708
rect 101582 539696 101588 539708
rect 91152 539668 101588 539696
rect 91152 539656 91158 539668
rect 101582 539656 101588 539668
rect 101640 539656 101646 539708
rect 144822 539656 144828 539708
rect 144880 539696 144886 539708
rect 283926 539696 283932 539708
rect 144880 539668 283932 539696
rect 144880 539656 144886 539668
rect 283926 539656 283932 539668
rect 283984 539656 283990 539708
rect 328822 539656 328828 539708
rect 328880 539696 328886 539708
rect 360470 539696 360476 539708
rect 328880 539668 360476 539696
rect 328880 539656 328886 539668
rect 360470 539656 360476 539668
rect 360528 539656 360534 539708
rect 63402 539588 63408 539640
rect 63460 539628 63466 539640
rect 67542 539628 67548 539640
rect 63460 539600 67548 539628
rect 63460 539588 63466 539600
rect 67542 539588 67548 539600
rect 67600 539588 67606 539640
rect 69382 539588 69388 539640
rect 69440 539588 69446 539640
rect 71866 539588 71872 539640
rect 71924 539588 71930 539640
rect 81158 539588 81164 539640
rect 81216 539628 81222 539640
rect 88794 539628 88800 539640
rect 81216 539600 88800 539628
rect 81216 539588 81222 539600
rect 88794 539588 88800 539600
rect 88852 539588 88858 539640
rect 250622 539628 250628 539640
rect 88904 539600 250628 539628
rect 88150 539520 88156 539572
rect 88208 539560 88214 539572
rect 88904 539560 88932 539600
rect 250622 539588 250628 539600
rect 250680 539588 250686 539640
rect 349982 539588 349988 539640
rect 350040 539628 350046 539640
rect 393958 539628 393964 539640
rect 350040 539600 393964 539628
rect 350040 539588 350046 539600
rect 393958 539588 393964 539600
rect 394016 539588 394022 539640
rect 88208 539532 88932 539560
rect 88208 539520 88214 539532
rect 268378 539520 268384 539572
rect 268436 539560 268442 539572
rect 272334 539560 272340 539572
rect 268436 539532 272340 539560
rect 268436 539520 268442 539532
rect 272334 539520 272340 539532
rect 272392 539520 272398 539572
rect 273898 539520 273904 539572
rect 273956 539560 273962 539572
rect 275646 539560 275652 539572
rect 273956 539532 275652 539560
rect 273956 539520 273962 539532
rect 275646 539520 275652 539532
rect 275704 539520 275710 539572
rect 278038 539520 278044 539572
rect 278096 539560 278102 539572
rect 278958 539560 278964 539572
rect 278096 539532 278964 539560
rect 278096 539520 278102 539532
rect 278958 539520 278964 539532
rect 279016 539520 279022 539572
rect 17218 538840 17224 538892
rect 17276 538880 17282 538892
rect 91186 538880 91192 538892
rect 17276 538852 91192 538880
rect 17276 538840 17282 538852
rect 91186 538840 91192 538852
rect 91244 538840 91250 538892
rect 172422 538840 172428 538892
rect 172480 538880 172486 538892
rect 195238 538880 195244 538892
rect 172480 538852 195244 538880
rect 172480 538840 172486 538852
rect 195238 538840 195244 538852
rect 195296 538840 195302 538892
rect 195790 538296 195796 538348
rect 195848 538336 195854 538348
rect 202782 538336 202788 538348
rect 195848 538308 202788 538336
rect 195848 538296 195854 538308
rect 202782 538296 202788 538308
rect 202840 538296 202846 538348
rect 221090 538296 221096 538348
rect 221148 538336 221154 538348
rect 232406 538336 232412 538348
rect 221148 538308 232412 538336
rect 221148 538296 221154 538308
rect 232406 538296 232412 538308
rect 232464 538296 232470 538348
rect 295978 538296 295984 538348
rect 296036 538336 296042 538348
rect 297174 538336 297180 538348
rect 296036 538308 297180 538336
rect 296036 538296 296042 538308
rect 297174 538296 297180 538308
rect 297232 538296 297238 538348
rect 323670 538296 323676 538348
rect 323728 538336 323734 538348
rect 340782 538336 340788 538348
rect 323728 538308 340788 538336
rect 323728 538296 323734 538308
rect 340782 538296 340788 538308
rect 340840 538296 340846 538348
rect 347038 538296 347044 538348
rect 347096 538336 347102 538348
rect 360194 538336 360200 538348
rect 347096 538308 360200 538336
rect 347096 538296 347102 538308
rect 360194 538296 360200 538308
rect 360252 538296 360258 538348
rect 67818 538228 67824 538280
rect 67876 538268 67882 538280
rect 76558 538268 76564 538280
rect 67876 538240 76564 538268
rect 67876 538228 67882 538240
rect 76558 538228 76564 538240
rect 76616 538228 76622 538280
rect 166258 538228 166264 538280
rect 166316 538268 166322 538280
rect 204162 538268 204168 538280
rect 166316 538240 204168 538268
rect 166316 538228 166322 538240
rect 204162 538228 204168 538240
rect 204220 538228 204226 538280
rect 208394 538228 208400 538280
rect 208452 538268 208458 538280
rect 356330 538268 356336 538280
rect 208452 538240 356336 538268
rect 208452 538228 208458 538240
rect 356330 538228 356336 538240
rect 356388 538228 356394 538280
rect 86862 538160 86868 538212
rect 86920 538200 86926 538212
rect 128998 538200 129004 538212
rect 86920 538172 129004 538200
rect 86920 538160 86926 538172
rect 128998 538160 129004 538172
rect 129056 538160 129062 538212
rect 340782 538160 340788 538212
rect 340840 538200 340846 538212
rect 579890 538200 579896 538212
rect 340840 538172 579896 538200
rect 340840 538160 340846 538172
rect 579890 538160 579896 538172
rect 579948 538160 579954 538212
rect 8202 537480 8208 537532
rect 8260 537520 8266 537532
rect 91278 537520 91284 537532
rect 8260 537492 91284 537520
rect 8260 537480 8266 537492
rect 91278 537480 91284 537492
rect 91336 537480 91342 537532
rect 198734 537480 198740 537532
rect 198792 537520 198798 537532
rect 208394 537520 208400 537532
rect 198792 537492 208400 537520
rect 198792 537480 198798 537492
rect 208394 537480 208400 537492
rect 208452 537480 208458 537532
rect 129642 536800 129648 536852
rect 129700 536840 129706 536852
rect 267182 536840 267188 536852
rect 129700 536812 267188 536840
rect 129700 536800 129706 536812
rect 267182 536800 267188 536812
rect 267240 536800 267246 536852
rect 43438 536732 43444 536784
rect 43496 536772 43502 536784
rect 70486 536772 70492 536784
rect 43496 536744 70492 536772
rect 43496 536732 43502 536744
rect 70486 536732 70492 536744
rect 70544 536732 70550 536784
rect 72326 536732 72332 536784
rect 72384 536772 72390 536784
rect 81158 536772 81164 536784
rect 72384 536744 81164 536772
rect 72384 536732 72390 536744
rect 81158 536732 81164 536744
rect 81216 536732 81222 536784
rect 68646 536664 68652 536716
rect 68704 536704 68710 536716
rect 88150 536704 88156 536716
rect 68704 536676 88156 536704
rect 68704 536664 68710 536676
rect 88150 536664 88156 536676
rect 88208 536664 88214 536716
rect 353938 536052 353944 536104
rect 353996 536092 354002 536104
rect 354582 536092 354588 536104
rect 353996 536064 354588 536092
rect 353996 536052 354002 536064
rect 354582 536052 354588 536064
rect 354640 536092 354646 536104
rect 359458 536092 359464 536104
rect 354640 536064 359464 536092
rect 354640 536052 354646 536064
rect 359458 536052 359464 536064
rect 359516 536052 359522 536104
rect 197998 535576 198004 535628
rect 198056 535616 198062 535628
rect 201310 535616 201316 535628
rect 198056 535588 201316 535616
rect 198056 535576 198062 535588
rect 201310 535576 201316 535588
rect 201368 535576 201374 535628
rect 148318 535508 148324 535560
rect 148376 535548 148382 535560
rect 293494 535548 293500 535560
rect 148376 535520 293500 535548
rect 148376 535508 148382 535520
rect 293494 535508 293500 535520
rect 293552 535508 293558 535560
rect 82722 535440 82728 535492
rect 82780 535480 82786 535492
rect 86218 535480 86224 535492
rect 82780 535452 86224 535480
rect 82780 535440 82786 535452
rect 86218 535440 86224 535452
rect 86276 535440 86282 535492
rect 201402 535440 201408 535492
rect 201460 535480 201466 535492
rect 580258 535480 580264 535492
rect 201460 535452 580264 535480
rect 201460 535440 201466 535452
rect 580258 535440 580264 535452
rect 580316 535440 580322 535492
rect 204898 535276 204904 535288
rect 200086 535248 204904 535276
rect 78306 534760 78312 534812
rect 78364 534800 78370 534812
rect 124214 534800 124220 534812
rect 78364 534772 124220 534800
rect 78364 534760 78370 534772
rect 124214 534760 124220 534772
rect 124272 534800 124278 534812
rect 125042 534800 125048 534812
rect 124272 534772 125048 534800
rect 124272 534760 124278 534772
rect 125042 534760 125048 534772
rect 125100 534760 125106 534812
rect 177298 534760 177304 534812
rect 177356 534800 177362 534812
rect 193950 534800 193956 534812
rect 177356 534772 193956 534800
rect 177356 534760 177362 534772
rect 193950 534760 193956 534772
rect 194008 534760 194014 534812
rect 199838 534760 199844 534812
rect 199896 534800 199902 534812
rect 200086 534800 200114 535248
rect 204898 535236 204904 535248
rect 204956 535236 204962 535288
rect 355594 535236 355600 535288
rect 355652 535276 355658 535288
rect 355652 535248 364334 535276
rect 355652 535236 355658 535248
rect 199896 534772 200114 534800
rect 364306 534800 364334 535248
rect 427814 534800 427820 534812
rect 364306 534772 427820 534800
rect 199896 534760 199902 534772
rect 427814 534760 427820 534772
rect 427872 534760 427878 534812
rect 18598 534692 18604 534744
rect 18656 534732 18662 534744
rect 91186 534732 91192 534744
rect 18656 534704 91192 534732
rect 18656 534692 18662 534704
rect 91186 534692 91192 534704
rect 91244 534692 91250 534744
rect 180058 534692 180064 534744
rect 180116 534732 180122 534744
rect 198734 534732 198740 534744
rect 180116 534704 198740 534732
rect 180116 534692 180122 534704
rect 198734 534692 198740 534704
rect 198792 534692 198798 534744
rect 125042 534080 125048 534132
rect 125100 534120 125106 534132
rect 140774 534120 140780 534132
rect 125100 534092 140780 534120
rect 125100 534080 125106 534092
rect 140774 534080 140780 534092
rect 140832 534080 140838 534132
rect 193858 534080 193864 534132
rect 193916 534120 193922 534132
rect 197354 534120 197360 534132
rect 193916 534092 197360 534120
rect 193916 534080 193922 534092
rect 197354 534080 197360 534092
rect 197412 534080 197418 534132
rect 67358 534012 67364 534064
rect 67416 534052 67422 534064
rect 188614 534052 188620 534064
rect 67416 534024 188620 534052
rect 67416 534012 67422 534024
rect 188614 534012 188620 534024
rect 188672 534012 188678 534064
rect 81066 532652 81072 532704
rect 81124 532692 81130 532704
rect 97994 532692 98000 532704
rect 81124 532664 98000 532692
rect 81124 532652 81130 532664
rect 97994 532652 98000 532664
rect 98052 532652 98058 532704
rect 140774 532652 140780 532704
rect 140832 532692 140838 532704
rect 197354 532692 197360 532704
rect 140832 532664 197360 532692
rect 140832 532652 140838 532664
rect 197354 532652 197360 532664
rect 197412 532652 197418 532704
rect 3418 531972 3424 532024
rect 3476 532012 3482 532024
rect 89714 532012 89720 532024
rect 3476 531984 89720 532012
rect 3476 531972 3482 531984
rect 89714 531972 89720 531984
rect 89772 531972 89778 532024
rect 358722 531972 358728 532024
rect 358780 532012 358786 532024
rect 582926 532012 582932 532024
rect 358780 531984 582932 532012
rect 358780 531972 358786 531984
rect 582926 531972 582932 531984
rect 582984 531972 582990 532024
rect 97994 531292 98000 531344
rect 98052 531332 98058 531344
rect 155218 531332 155224 531344
rect 98052 531304 155224 531332
rect 98052 531292 98058 531304
rect 155218 531292 155224 531304
rect 155276 531292 155282 531344
rect 44082 531224 44088 531276
rect 44140 531264 44146 531276
rect 188522 531264 188528 531276
rect 44140 531236 188528 531264
rect 44140 531224 44146 531236
rect 188522 531224 188528 531236
rect 188580 531224 188586 531276
rect 64782 530544 64788 530596
rect 64840 530584 64846 530596
rect 77938 530584 77944 530596
rect 64840 530556 77944 530584
rect 64840 530544 64846 530556
rect 77938 530544 77944 530556
rect 77996 530544 78002 530596
rect 176010 530544 176016 530596
rect 176068 530584 176074 530596
rect 199470 530584 199476 530596
rect 176068 530556 199476 530584
rect 176068 530544 176074 530556
rect 199470 530544 199476 530556
rect 199528 530544 199534 530596
rect 124858 529864 124864 529916
rect 124916 529904 124922 529916
rect 197354 529904 197360 529916
rect 124916 529876 197360 529904
rect 124916 529864 124922 529876
rect 197354 529864 197360 529876
rect 197412 529864 197418 529916
rect 64690 529796 64696 529848
rect 64748 529836 64754 529848
rect 124950 529836 124956 529848
rect 64748 529808 124956 529836
rect 64748 529796 64754 529808
rect 124950 529796 124956 529808
rect 125008 529796 125014 529848
rect 79318 529728 79324 529780
rect 79376 529768 79382 529780
rect 79962 529768 79968 529780
rect 79376 529740 79968 529768
rect 79376 529728 79382 529740
rect 79962 529728 79968 529740
rect 80020 529728 80026 529780
rect 59262 529184 59268 529236
rect 59320 529224 59326 529236
rect 79318 529224 79324 529236
rect 59320 529196 79324 529224
rect 59320 529184 59326 529196
rect 79318 529184 79324 529196
rect 79376 529184 79382 529236
rect 358722 528572 358728 528624
rect 358780 528612 358786 528624
rect 371234 528612 371240 528624
rect 358780 528584 371240 528612
rect 358780 528572 358786 528584
rect 371234 528572 371240 528584
rect 371292 528572 371298 528624
rect 180242 528504 180248 528556
rect 180300 528544 180306 528556
rect 197354 528544 197360 528556
rect 180300 528516 197360 528544
rect 180300 528504 180306 528516
rect 197354 528504 197360 528516
rect 197412 528504 197418 528556
rect 70394 527484 70400 527536
rect 70452 527524 70458 527536
rect 71038 527524 71044 527536
rect 70452 527496 71044 527524
rect 70452 527484 70458 527496
rect 71038 527484 71044 527496
rect 71096 527484 71102 527536
rect 71038 527144 71044 527196
rect 71096 527184 71102 527196
rect 141510 527184 141516 527196
rect 71096 527156 141516 527184
rect 71096 527144 71102 527156
rect 141510 527144 141516 527156
rect 141568 527144 141574 527196
rect 358722 527144 358728 527196
rect 358780 527184 358786 527196
rect 376754 527184 376760 527196
rect 358780 527156 376760 527184
rect 358780 527144 358786 527156
rect 376754 527144 376760 527156
rect 376812 527144 376818 527196
rect 50890 527076 50896 527128
rect 50948 527116 50954 527128
rect 160830 527116 160836 527128
rect 50948 527088 160836 527116
rect 50948 527076 50954 527088
rect 160830 527076 160836 527088
rect 160888 527076 160894 527128
rect 173158 525036 173164 525088
rect 173216 525076 173222 525088
rect 197998 525076 198004 525088
rect 173216 525048 198004 525076
rect 173216 525036 173222 525048
rect 197998 525036 198004 525048
rect 198056 525036 198062 525088
rect 170398 524424 170404 524476
rect 170456 524464 170462 524476
rect 197354 524464 197360 524476
rect 170456 524436 197360 524464
rect 170456 524424 170462 524436
rect 197354 524424 197360 524436
rect 197412 524424 197418 524476
rect 358722 524424 358728 524476
rect 358780 524464 358786 524476
rect 375466 524464 375472 524476
rect 358780 524436 375472 524464
rect 358780 524424 358786 524436
rect 375466 524424 375472 524436
rect 375524 524424 375530 524476
rect 59170 523676 59176 523728
rect 59228 523716 59234 523728
rect 78766 523716 78772 523728
rect 59228 523688 78772 523716
rect 59228 523676 59234 523688
rect 78766 523676 78772 523688
rect 78824 523676 78830 523728
rect 66898 522248 66904 522300
rect 66956 522288 66962 522300
rect 177390 522288 177396 522300
rect 66956 522260 177396 522288
rect 66956 522248 66962 522260
rect 177390 522248 177396 522260
rect 177448 522248 177454 522300
rect 147582 521636 147588 521688
rect 147640 521676 147646 521688
rect 197354 521676 197360 521688
rect 147640 521648 197360 521676
rect 147640 521636 147646 521648
rect 197354 521636 197360 521648
rect 197412 521636 197418 521688
rect 34422 520888 34428 520940
rect 34480 520928 34486 520940
rect 195238 520928 195244 520940
rect 34480 520900 195244 520928
rect 34480 520888 34486 520900
rect 195238 520888 195244 520900
rect 195296 520888 195302 520940
rect 358722 520888 358728 520940
rect 358780 520928 358786 520940
rect 395982 520928 395988 520940
rect 358780 520900 395988 520928
rect 358780 520888 358786 520900
rect 395982 520888 395988 520900
rect 396040 520888 396046 520940
rect 395982 520276 395988 520328
rect 396040 520316 396046 520328
rect 582466 520316 582472 520328
rect 396040 520288 582472 520316
rect 396040 520276 396046 520288
rect 582466 520276 582472 520288
rect 582524 520276 582530 520328
rect 55122 519528 55128 519580
rect 55180 519568 55186 519580
rect 85574 519568 85580 519580
rect 55180 519540 85580 519568
rect 55180 519528 55186 519540
rect 85574 519528 85580 519540
rect 85632 519528 85638 519580
rect 358722 519528 358728 519580
rect 358780 519568 358786 519580
rect 388438 519568 388444 519580
rect 358780 519540 388444 519568
rect 358780 519528 358786 519540
rect 388438 519528 388444 519540
rect 388496 519528 388502 519580
rect 62022 517420 62028 517472
rect 62080 517460 62086 517472
rect 186958 517460 186964 517472
rect 62080 517432 186964 517460
rect 62080 517420 62086 517432
rect 186958 517420 186964 517432
rect 187016 517420 187022 517472
rect 180242 516128 180248 516180
rect 180300 516168 180306 516180
rect 197354 516168 197360 516180
rect 180300 516140 197360 516168
rect 180300 516128 180306 516140
rect 197354 516128 197360 516140
rect 197412 516128 197418 516180
rect 358722 516128 358728 516180
rect 358780 516168 358786 516180
rect 374730 516168 374736 516180
rect 358780 516140 374736 516168
rect 358780 516128 358786 516140
rect 374730 516128 374736 516140
rect 374788 516128 374794 516180
rect 3510 514768 3516 514820
rect 3568 514808 3574 514820
rect 14458 514808 14464 514820
rect 3568 514780 14464 514808
rect 3568 514768 3574 514780
rect 14458 514768 14464 514780
rect 14516 514768 14522 514820
rect 175182 514768 175188 514820
rect 175240 514808 175246 514820
rect 197354 514808 197360 514820
rect 175240 514780 197360 514808
rect 175240 514768 175246 514780
rect 197354 514768 197360 514780
rect 197412 514768 197418 514820
rect 60550 514700 60556 514752
rect 60608 514740 60614 514752
rect 188430 514740 188436 514752
rect 60608 514712 188436 514740
rect 60608 514700 60614 514712
rect 188430 514700 188436 514712
rect 188488 514700 188494 514752
rect 41322 511232 41328 511284
rect 41380 511272 41386 511284
rect 180150 511272 180156 511284
rect 41380 511244 180156 511272
rect 41380 511232 41386 511244
rect 180150 511232 180156 511244
rect 180208 511232 180214 511284
rect 141510 510552 141516 510604
rect 141568 510592 141574 510604
rect 197354 510592 197360 510604
rect 141568 510564 197360 510592
rect 141568 510552 141574 510564
rect 197354 510552 197360 510564
rect 197412 510552 197418 510604
rect 358722 509668 358728 509720
rect 358780 509708 358786 509720
rect 360286 509708 360292 509720
rect 358780 509680 360292 509708
rect 358780 509668 358786 509680
rect 360286 509668 360292 509680
rect 360344 509668 360350 509720
rect 46842 507084 46848 507136
rect 46900 507124 46906 507136
rect 196802 507124 196808 507136
rect 46900 507096 196808 507124
rect 46900 507084 46906 507096
rect 196802 507084 196808 507096
rect 196860 507084 196866 507136
rect 358722 505112 358728 505164
rect 358780 505152 358786 505164
rect 414658 505152 414664 505164
rect 358780 505124 414664 505152
rect 358780 505112 358786 505124
rect 414658 505112 414664 505124
rect 414716 505112 414722 505164
rect 164878 504364 164884 504416
rect 164936 504404 164942 504416
rect 197354 504404 197360 504416
rect 164936 504376 197360 504404
rect 164936 504364 164942 504376
rect 197354 504364 197360 504376
rect 197412 504364 197418 504416
rect 358722 502324 358728 502376
rect 358780 502364 358786 502376
rect 369854 502364 369860 502376
rect 358780 502336 369860 502364
rect 358780 502324 358786 502336
rect 369854 502324 369860 502336
rect 369912 502324 369918 502376
rect 3510 502256 3516 502308
rect 3568 502296 3574 502308
rect 18598 502296 18604 502308
rect 3568 502268 18604 502296
rect 3568 502256 3574 502268
rect 18598 502256 18604 502268
rect 18656 502256 18662 502308
rect 155218 500896 155224 500948
rect 155276 500936 155282 500948
rect 198274 500936 198280 500948
rect 155276 500908 198280 500936
rect 155276 500896 155282 500908
rect 198274 500896 198280 500908
rect 198332 500896 198338 500948
rect 155862 498788 155868 498840
rect 155920 498828 155926 498840
rect 180242 498828 180248 498840
rect 155920 498800 180248 498828
rect 155920 498788 155926 498800
rect 180242 498788 180248 498800
rect 180300 498788 180306 498840
rect 180150 496816 180156 496868
rect 180208 496856 180214 496868
rect 197354 496856 197360 496868
rect 180208 496828 197360 496856
rect 180208 496816 180214 496828
rect 197354 496816 197360 496828
rect 197412 496816 197418 496868
rect 357158 496748 357164 496800
rect 357216 496788 357222 496800
rect 583018 496788 583024 496800
rect 357216 496760 583024 496788
rect 357216 496748 357222 496760
rect 583018 496748 583024 496760
rect 583076 496748 583082 496800
rect 178678 495456 178684 495508
rect 178736 495496 178742 495508
rect 197354 495496 197360 495508
rect 178736 495468 197360 495496
rect 178736 495456 178742 495468
rect 197354 495456 197360 495468
rect 197412 495456 197418 495508
rect 358630 493960 358636 494012
rect 358688 494000 358694 494012
rect 412634 494000 412640 494012
rect 358688 493972 412640 494000
rect 358688 493960 358694 493972
rect 412634 493960 412640 493972
rect 412692 493960 412698 494012
rect 138658 492668 138664 492720
rect 138716 492708 138722 492720
rect 197354 492708 197360 492720
rect 138716 492680 197360 492708
rect 138716 492668 138722 492680
rect 197354 492668 197360 492680
rect 197412 492668 197418 492720
rect 127618 488520 127624 488572
rect 127676 488560 127682 488572
rect 151814 488560 151820 488572
rect 127676 488532 151820 488560
rect 127676 488520 127682 488532
rect 151786 488520 151820 488532
rect 151872 488520 151878 488572
rect 151786 488492 151814 488520
rect 197354 488492 197360 488504
rect 151786 488464 197360 488492
rect 197354 488452 197360 488464
rect 197412 488452 197418 488504
rect 358722 486412 358728 486464
rect 358780 486452 358786 486464
rect 385034 486452 385040 486464
rect 358780 486424 385040 486452
rect 358780 486412 358786 486424
rect 385034 486412 385040 486424
rect 385092 486412 385098 486464
rect 181622 483624 181628 483676
rect 181680 483664 181686 483676
rect 197354 483664 197360 483676
rect 181680 483636 197360 483664
rect 181680 483624 181686 483636
rect 197354 483624 197360 483636
rect 197412 483624 197418 483676
rect 358722 481652 358728 481704
rect 358780 481692 358786 481704
rect 364334 481692 364340 481704
rect 358780 481664 364340 481692
rect 358780 481652 358786 481664
rect 364334 481652 364340 481664
rect 364392 481652 364398 481704
rect 180242 480224 180248 480276
rect 180300 480264 180306 480276
rect 197354 480264 197360 480276
rect 180300 480236 197360 480264
rect 180300 480224 180306 480236
rect 197354 480224 197360 480236
rect 197412 480224 197418 480276
rect 358722 480224 358728 480276
rect 358780 480264 358786 480276
rect 378134 480264 378140 480276
rect 358780 480236 378140 480264
rect 358780 480224 358786 480236
rect 378134 480224 378140 480236
rect 378192 480224 378198 480276
rect 124858 477504 124864 477556
rect 124916 477544 124922 477556
rect 171042 477544 171048 477556
rect 124916 477516 171048 477544
rect 124916 477504 124922 477516
rect 171042 477504 171048 477516
rect 171100 477544 171106 477556
rect 197354 477544 197360 477556
rect 171100 477516 197360 477544
rect 171100 477504 171106 477516
rect 197354 477504 197360 477516
rect 197412 477504 197418 477556
rect 358722 477504 358728 477556
rect 358780 477544 358786 477556
rect 367186 477544 367192 477556
rect 358780 477516 367192 477544
rect 358780 477504 358786 477516
rect 367186 477504 367192 477516
rect 367244 477504 367250 477556
rect 68278 476076 68284 476128
rect 68336 476116 68342 476128
rect 68922 476116 68928 476128
rect 68336 476088 68928 476116
rect 68336 476076 68342 476088
rect 68922 476076 68928 476088
rect 68980 476116 68986 476128
rect 68980 476088 147168 476116
rect 68980 476076 68986 476088
rect 147140 476048 147168 476088
rect 147490 476048 147496 476060
rect 147140 476020 147496 476048
rect 147490 476008 147496 476020
rect 147548 476048 147554 476060
rect 180058 476048 180064 476060
rect 147548 476020 180064 476048
rect 147548 476008 147554 476020
rect 180058 476008 180064 476020
rect 180116 476008 180122 476060
rect 3326 475328 3332 475380
rect 3384 475368 3390 475380
rect 8202 475368 8208 475380
rect 3384 475340 8208 475368
rect 3384 475328 3390 475340
rect 8202 475328 8208 475340
rect 8260 475368 8266 475380
rect 15838 475368 15844 475380
rect 8260 475340 15844 475368
rect 8260 475328 8266 475340
rect 15838 475328 15844 475340
rect 15896 475328 15902 475380
rect 177390 474716 177396 474768
rect 177448 474756 177454 474768
rect 197354 474756 197360 474768
rect 177448 474728 197360 474756
rect 177448 474716 177454 474728
rect 197354 474716 197360 474728
rect 197412 474716 197418 474768
rect 137278 473356 137284 473408
rect 137336 473396 137342 473408
rect 197354 473396 197360 473408
rect 137336 473368 197360 473396
rect 137336 473356 137342 473368
rect 197354 473356 197360 473368
rect 197412 473356 197418 473408
rect 358538 471996 358544 472048
rect 358596 472036 358602 472048
rect 389174 472036 389180 472048
rect 358596 472008 389180 472036
rect 358596 471996 358602 472008
rect 389174 471996 389180 472008
rect 389232 471996 389238 472048
rect 191190 471248 191196 471300
rect 191248 471288 191254 471300
rect 198090 471288 198096 471300
rect 191248 471260 198096 471288
rect 191248 471248 191254 471260
rect 198090 471248 198096 471260
rect 198148 471248 198154 471300
rect 357894 470568 357900 470620
rect 357952 470608 357958 470620
rect 368566 470608 368572 470620
rect 357952 470580 368572 470608
rect 357952 470568 357958 470580
rect 368566 470568 368572 470580
rect 368624 470568 368630 470620
rect 165522 467848 165528 467900
rect 165580 467888 165586 467900
rect 197354 467888 197360 467900
rect 165580 467860 197360 467888
rect 165580 467848 165586 467860
rect 197354 467848 197360 467860
rect 197412 467848 197418 467900
rect 105538 467780 105544 467832
rect 105596 467820 105602 467832
rect 182082 467820 182088 467832
rect 105596 467792 182088 467820
rect 105596 467780 105602 467792
rect 182082 467780 182088 467792
rect 182140 467820 182146 467832
rect 188430 467820 188436 467832
rect 182140 467792 188436 467820
rect 182140 467780 182146 467792
rect 188430 467780 188436 467792
rect 188488 467780 188494 467832
rect 104894 466420 104900 466472
rect 104952 466460 104958 466472
rect 105538 466460 105544 466472
rect 104952 466432 105544 466460
rect 104952 466420 104958 466432
rect 105538 466420 105544 466432
rect 105596 466420 105602 466472
rect 93762 465672 93768 465724
rect 93820 465712 93826 465724
rect 107654 465712 107660 465724
rect 93820 465684 107660 465712
rect 93820 465672 93826 465684
rect 107654 465672 107660 465684
rect 107712 465672 107718 465724
rect 131758 465060 131764 465112
rect 131816 465100 131822 465112
rect 186958 465100 186964 465112
rect 131816 465072 186964 465100
rect 131816 465060 131822 465072
rect 186958 465060 186964 465072
rect 187016 465100 187022 465112
rect 197354 465100 197360 465112
rect 187016 465072 197360 465100
rect 187016 465060 187022 465072
rect 197354 465060 197360 465072
rect 197412 465060 197418 465112
rect 358722 465060 358728 465112
rect 358780 465100 358786 465112
rect 376938 465100 376944 465112
rect 358780 465072 376944 465100
rect 358780 465060 358786 465072
rect 376938 465060 376944 465072
rect 376996 465100 377002 465112
rect 583018 465100 583024 465112
rect 376996 465072 583024 465100
rect 376996 465060 377002 465072
rect 583018 465060 583024 465072
rect 583076 465060 583082 465112
rect 106182 462952 106188 463004
rect 106240 462992 106246 463004
rect 120810 462992 120816 463004
rect 106240 462964 120816 462992
rect 106240 462952 106246 462964
rect 120810 462952 120816 462964
rect 120868 462952 120874 463004
rect 3510 462340 3516 462392
rect 3568 462380 3574 462392
rect 25498 462380 25504 462392
rect 3568 462352 25504 462380
rect 3568 462340 3574 462352
rect 25498 462340 25504 462352
rect 25556 462340 25562 462392
rect 50982 462340 50988 462392
rect 51040 462380 51046 462392
rect 67726 462380 67732 462392
rect 51040 462352 67732 462380
rect 51040 462340 51046 462352
rect 67726 462340 67732 462352
rect 67784 462380 67790 462392
rect 68830 462380 68836 462392
rect 67784 462352 68836 462380
rect 67784 462340 67790 462352
rect 68830 462340 68836 462352
rect 68888 462340 68894 462392
rect 187142 462340 187148 462392
rect 187200 462380 187206 462392
rect 197354 462380 197360 462392
rect 187200 462352 197360 462380
rect 187200 462340 187206 462352
rect 197354 462340 197360 462352
rect 197412 462340 197418 462392
rect 68830 461592 68836 461644
rect 68888 461632 68894 461644
rect 81434 461632 81440 461644
rect 68888 461604 81440 461632
rect 68888 461592 68894 461604
rect 81434 461592 81440 461604
rect 81492 461592 81498 461644
rect 76006 461456 76012 461508
rect 76064 461496 76070 461508
rect 76558 461496 76564 461508
rect 76064 461468 76564 461496
rect 76064 461456 76070 461468
rect 76558 461456 76564 461468
rect 76616 461456 76622 461508
rect 76558 460912 76564 460964
rect 76616 460952 76622 460964
rect 159358 460952 159364 460964
rect 76616 460924 159364 460952
rect 76616 460912 76622 460924
rect 159358 460912 159364 460924
rect 159416 460912 159422 460964
rect 57882 460164 57888 460216
rect 57940 460204 57946 460216
rect 95234 460204 95240 460216
rect 57940 460176 95240 460204
rect 57940 460164 57946 460176
rect 95234 460164 95240 460176
rect 95292 460164 95298 460216
rect 148962 460164 148968 460216
rect 149020 460204 149026 460216
rect 197354 460204 197360 460216
rect 149020 460176 197360 460204
rect 149020 460164 149026 460176
rect 197354 460164 197360 460176
rect 197412 460164 197418 460216
rect 375282 460164 375288 460216
rect 375340 460204 375346 460216
rect 582558 460204 582564 460216
rect 375340 460176 582564 460204
rect 375340 460164 375346 460176
rect 582558 460164 582564 460176
rect 582616 460164 582622 460216
rect 148410 459552 148416 459604
rect 148468 459592 148474 459604
rect 148962 459592 148968 459604
rect 148468 459564 148968 459592
rect 148468 459552 148474 459564
rect 148962 459552 148968 459564
rect 149020 459552 149026 459604
rect 358446 459552 358452 459604
rect 358504 459592 358510 459604
rect 374086 459592 374092 459604
rect 358504 459564 374092 459592
rect 358504 459552 358510 459564
rect 374086 459552 374092 459564
rect 374144 459592 374150 459604
rect 375282 459592 375288 459604
rect 374144 459564 375288 459592
rect 374144 459552 374150 459564
rect 375282 459552 375288 459564
rect 375340 459552 375346 459604
rect 14458 459484 14464 459536
rect 14516 459524 14522 459536
rect 112438 459524 112444 459536
rect 14516 459496 112444 459524
rect 14516 459484 14522 459496
rect 112438 459484 112444 459496
rect 112496 459484 112502 459536
rect 127710 458192 127716 458244
rect 127768 458232 127774 458244
rect 197354 458232 197360 458244
rect 127768 458204 197360 458232
rect 127768 458192 127774 458204
rect 197354 458192 197360 458204
rect 197412 458192 197418 458244
rect 52270 457444 52276 457496
rect 52328 457484 52334 457496
rect 87046 457484 87052 457496
rect 52328 457456 87052 457484
rect 52328 457444 52334 457456
rect 87046 457444 87052 457456
rect 87104 457444 87110 457496
rect 60642 456696 60648 456748
rect 60700 456736 60706 456748
rect 65610 456736 65616 456748
rect 60700 456708 65616 456736
rect 60700 456696 60706 456708
rect 65610 456696 65616 456708
rect 65668 456696 65674 456748
rect 57790 456016 57796 456068
rect 57848 456056 57854 456068
rect 82814 456056 82820 456068
rect 57848 456028 82820 456056
rect 57848 456016 57854 456028
rect 82814 456016 82820 456028
rect 82872 456016 82878 456068
rect 65610 455404 65616 455456
rect 65668 455444 65674 455456
rect 65886 455444 65892 455456
rect 65668 455416 65892 455444
rect 65668 455404 65674 455416
rect 65886 455404 65892 455416
rect 65944 455444 65950 455456
rect 195238 455444 195244 455456
rect 65944 455416 195244 455444
rect 65944 455404 65950 455416
rect 195238 455404 195244 455416
rect 195296 455404 195302 455456
rect 358722 455404 358728 455456
rect 358780 455444 358786 455456
rect 363230 455444 363236 455456
rect 358780 455416 363236 455444
rect 358780 455404 358786 455416
rect 363230 455404 363236 455416
rect 363288 455444 363294 455456
rect 582466 455444 582472 455456
rect 363288 455416 582472 455444
rect 363288 455404 363294 455416
rect 582466 455404 582472 455416
rect 582524 455404 582530 455456
rect 172238 455336 172244 455388
rect 172296 455376 172302 455388
rect 172422 455376 172428 455388
rect 172296 455348 172428 455376
rect 172296 455336 172302 455348
rect 172422 455336 172428 455348
rect 172480 455376 172486 455388
rect 173250 455376 173256 455388
rect 172480 455348 173256 455376
rect 172480 455336 172486 455348
rect 173250 455336 173256 455348
rect 173308 455336 173314 455388
rect 88334 454792 88340 454844
rect 88392 454832 88398 454844
rect 88978 454832 88984 454844
rect 88392 454804 88984 454832
rect 88392 454792 88398 454804
rect 88978 454792 88984 454804
rect 89036 454792 89042 454844
rect 63310 454656 63316 454708
rect 63368 454696 63374 454708
rect 95878 454696 95884 454708
rect 63368 454668 95884 454696
rect 63368 454656 63374 454668
rect 95878 454656 95884 454668
rect 95936 454656 95942 454708
rect 88334 454044 88340 454096
rect 88392 454084 88398 454096
rect 133874 454084 133880 454096
rect 88392 454056 133880 454084
rect 88392 454044 88398 454056
rect 133874 454044 133880 454056
rect 133932 454044 133938 454096
rect 65978 453976 65984 454028
rect 66036 454016 66042 454028
rect 71038 454016 71044 454028
rect 66036 453988 71044 454016
rect 66036 453976 66042 453988
rect 71038 453976 71044 453988
rect 71096 453976 71102 454028
rect 97258 453976 97264 454028
rect 97316 454016 97322 454028
rect 102134 454016 102140 454028
rect 97316 453988 102140 454016
rect 97316 453976 97322 453988
rect 102134 453976 102140 453988
rect 102192 453976 102198 454028
rect 57606 453296 57612 453348
rect 57664 453336 57670 453348
rect 73154 453336 73160 453348
rect 57664 453308 73160 453336
rect 57664 453296 57670 453308
rect 73154 453296 73160 453308
rect 73212 453296 73218 453348
rect 102778 453296 102784 453348
rect 102836 453336 102842 453348
rect 125594 453336 125600 453348
rect 102836 453308 125600 453336
rect 102836 453296 102842 453308
rect 125594 453296 125600 453308
rect 125652 453296 125658 453348
rect 77938 452616 77944 452668
rect 77996 452656 78002 452668
rect 128446 452656 128452 452668
rect 77996 452628 128452 452656
rect 77996 452616 78002 452628
rect 128446 452616 128452 452628
rect 128504 452616 128510 452668
rect 358722 452616 358728 452668
rect 358780 452656 358786 452668
rect 398834 452656 398840 452668
rect 358780 452628 398840 452656
rect 358780 452616 358786 452628
rect 398834 452616 398840 452628
rect 398892 452616 398898 452668
rect 116578 451936 116584 451988
rect 116636 451976 116642 451988
rect 124306 451976 124312 451988
rect 116636 451948 124312 451976
rect 116636 451936 116642 451948
rect 124306 451936 124312 451948
rect 124364 451936 124370 451988
rect 3418 451868 3424 451920
rect 3476 451908 3482 451920
rect 121638 451908 121644 451920
rect 3476 451880 121644 451908
rect 3476 451868 3482 451880
rect 121638 451868 121644 451880
rect 121696 451868 121702 451920
rect 95878 451188 95884 451240
rect 95936 451228 95942 451240
rect 124858 451228 124864 451240
rect 95936 451200 124864 451228
rect 95936 451188 95942 451200
rect 124858 451188 124864 451200
rect 124916 451188 124922 451240
rect 106918 451120 106924 451172
rect 106976 451160 106982 451172
rect 127710 451160 127716 451172
rect 106976 451132 127716 451160
rect 106976 451120 106982 451132
rect 127710 451120 127716 451132
rect 127768 451120 127774 451172
rect 63218 450508 63224 450560
rect 63276 450548 63282 450560
rect 75914 450548 75920 450560
rect 63276 450520 75920 450548
rect 63276 450508 63282 450520
rect 75914 450508 75920 450520
rect 75972 450508 75978 450560
rect 358722 449896 358728 449948
rect 358780 449936 358786 449948
rect 375374 449936 375380 449948
rect 358780 449908 375380 449936
rect 358780 449896 358786 449908
rect 375374 449896 375380 449908
rect 375432 449896 375438 449948
rect 25498 449828 25504 449880
rect 25556 449868 25562 449880
rect 71774 449868 71780 449880
rect 25556 449840 71780 449868
rect 25556 449828 25562 449840
rect 71774 449828 71780 449840
rect 71832 449828 71838 449880
rect 64690 449216 64696 449268
rect 64748 449256 64754 449268
rect 78674 449256 78680 449268
rect 64748 449228 78680 449256
rect 64748 449216 64754 449228
rect 78674 449216 78680 449228
rect 78732 449216 78738 449268
rect 100018 449216 100024 449268
rect 100076 449256 100082 449268
rect 123570 449256 123576 449268
rect 100076 449228 123576 449256
rect 100076 449216 100082 449228
rect 123570 449216 123576 449228
rect 123628 449216 123634 449268
rect 71774 449148 71780 449200
rect 71832 449188 71838 449200
rect 72694 449188 72700 449200
rect 71832 449160 72700 449188
rect 71832 449148 71838 449160
rect 72694 449148 72700 449160
rect 72752 449188 72758 449200
rect 103514 449188 103520 449200
rect 72752 449160 103520 449188
rect 72752 449148 72758 449160
rect 103514 449148 103520 449160
rect 103572 449188 103578 449200
rect 103698 449188 103704 449200
rect 103572 449160 103704 449188
rect 103572 449148 103578 449160
rect 103698 449148 103704 449160
rect 103756 449148 103762 449200
rect 358722 449148 358728 449200
rect 358780 449188 358786 449200
rect 365898 449188 365904 449200
rect 358780 449160 365904 449188
rect 358780 449148 358786 449160
rect 365898 449148 365904 449160
rect 365956 449188 365962 449200
rect 582650 449188 582656 449200
rect 365956 449160 582656 449188
rect 365956 449148 365962 449160
rect 582650 449148 582656 449160
rect 582708 449148 582714 449200
rect 3142 448536 3148 448588
rect 3200 448576 3206 448588
rect 18598 448576 18604 448588
rect 3200 448548 18604 448576
rect 3200 448536 3206 448548
rect 18598 448536 18604 448548
rect 18656 448536 18662 448588
rect 119338 448536 119344 448588
rect 119396 448576 119402 448588
rect 137370 448576 137376 448588
rect 119396 448548 137376 448576
rect 119396 448536 119402 448548
rect 137370 448536 137376 448548
rect 137428 448536 137434 448588
rect 184750 448536 184756 448588
rect 184808 448576 184814 448588
rect 197354 448576 197360 448588
rect 184808 448548 197360 448576
rect 184808 448536 184814 448548
rect 197354 448536 197360 448548
rect 197412 448536 197418 448588
rect 94498 448468 94504 448520
rect 94556 448508 94562 448520
rect 187142 448508 187148 448520
rect 94556 448480 187148 448508
rect 94556 448468 94562 448480
rect 187142 448468 187148 448480
rect 187200 448468 187206 448520
rect 61930 447788 61936 447840
rect 61988 447828 61994 447840
rect 71774 447828 71780 447840
rect 61988 447800 71780 447828
rect 61988 447788 61994 447800
rect 71774 447788 71780 447800
rect 71832 447788 71838 447840
rect 68278 447176 68284 447228
rect 68336 447216 68342 447228
rect 71866 447216 71872 447228
rect 68336 447188 71872 447216
rect 68336 447176 68342 447188
rect 71866 447176 71872 447188
rect 71924 447176 71930 447228
rect 71774 447108 71780 447160
rect 71832 447148 71838 447160
rect 124858 447148 124864 447160
rect 71832 447120 124864 447148
rect 71832 447108 71838 447120
rect 124858 447108 124864 447120
rect 124916 447108 124922 447160
rect 68922 447040 68928 447092
rect 68980 447080 68986 447092
rect 73154 447080 73160 447092
rect 68980 447052 73160 447080
rect 68980 447040 68986 447052
rect 73154 447040 73160 447052
rect 73212 447040 73218 447092
rect 109034 447040 109040 447092
rect 109092 447080 109098 447092
rect 109770 447080 109776 447092
rect 109092 447052 109776 447080
rect 109092 447040 109098 447052
rect 109770 447040 109776 447052
rect 109828 447080 109834 447092
rect 148318 447080 148324 447092
rect 109828 447052 148324 447080
rect 109828 447040 109834 447052
rect 148318 447040 148324 447052
rect 148376 447040 148382 447092
rect 140774 446768 140780 446820
rect 140832 446808 140838 446820
rect 142062 446808 142068 446820
rect 140832 446780 142068 446808
rect 140832 446768 140838 446780
rect 142062 446768 142068 446780
rect 142120 446808 142126 446820
rect 142982 446808 142988 446820
rect 142120 446780 142988 446808
rect 142120 446768 142126 446780
rect 142982 446768 142988 446780
rect 143040 446768 143046 446820
rect 71866 446700 71872 446752
rect 71924 446740 71930 446752
rect 74810 446740 74816 446752
rect 71924 446712 74816 446740
rect 71924 446700 71930 446712
rect 74810 446700 74816 446712
rect 74868 446700 74874 446752
rect 49602 446360 49608 446412
rect 49660 446400 49666 446412
rect 67818 446400 67824 446412
rect 49660 446372 67824 446400
rect 49660 446360 49666 446372
rect 67818 446360 67824 446372
rect 67876 446400 67882 446412
rect 68738 446400 68744 446412
rect 67876 446372 68744 446400
rect 67876 446360 67882 446372
rect 68738 446360 68744 446372
rect 68796 446360 68802 446412
rect 112438 445748 112444 445800
rect 112496 445788 112502 445800
rect 112898 445788 112904 445800
rect 112496 445760 112904 445788
rect 112496 445748 112502 445760
rect 112898 445748 112904 445760
rect 112956 445788 112962 445800
rect 124950 445788 124956 445800
rect 112956 445760 124956 445788
rect 112956 445748 112962 445760
rect 124950 445748 124956 445760
rect 125008 445748 125014 445800
rect 195330 445748 195336 445800
rect 195388 445788 195394 445800
rect 197354 445788 197360 445800
rect 195388 445760 197360 445788
rect 195388 445748 195394 445760
rect 197354 445748 197360 445760
rect 197412 445748 197418 445800
rect 358722 445748 358728 445800
rect 358780 445788 358786 445800
rect 368474 445788 368480 445800
rect 358780 445760 368480 445788
rect 358780 445748 358786 445760
rect 368474 445748 368480 445760
rect 368532 445748 368538 445800
rect 130378 445000 130384 445052
rect 130436 445040 130442 445052
rect 195330 445040 195336 445052
rect 130436 445012 195336 445040
rect 130436 445000 130442 445012
rect 195330 445000 195336 445012
rect 195388 445000 195394 445052
rect 59262 444456 59268 444508
rect 59320 444496 59326 444508
rect 79410 444496 79416 444508
rect 59320 444468 79416 444496
rect 59320 444456 59326 444468
rect 79410 444456 79416 444468
rect 79468 444456 79474 444508
rect 101398 444456 101404 444508
rect 101456 444496 101462 444508
rect 127710 444496 127716 444508
rect 101456 444468 127716 444496
rect 101456 444456 101462 444468
rect 127710 444456 127716 444468
rect 127768 444456 127774 444508
rect 4798 444388 4804 444440
rect 4856 444428 4862 444440
rect 118694 444428 118700 444440
rect 4856 444400 118700 444428
rect 4856 444388 4862 444400
rect 118694 444388 118700 444400
rect 118752 444388 118758 444440
rect 120074 444388 120080 444440
rect 120132 444428 120138 444440
rect 120718 444428 120724 444440
rect 120132 444400 120724 444428
rect 120132 444388 120138 444400
rect 120718 444388 120724 444400
rect 120776 444428 120782 444440
rect 130470 444428 130476 444440
rect 120776 444400 130476 444428
rect 120776 444388 120782 444400
rect 130470 444388 130476 444400
rect 130528 444388 130534 444440
rect 124122 444320 124128 444372
rect 124180 444360 124186 444372
rect 124306 444360 124312 444372
rect 124180 444332 124312 444360
rect 124180 444320 124186 444332
rect 124306 444320 124312 444332
rect 124364 444360 124370 444372
rect 166350 444360 166356 444372
rect 124364 444332 166356 444360
rect 124364 444320 124370 444332
rect 166350 444320 166356 444332
rect 166408 444320 166414 444372
rect 147490 444252 147496 444304
rect 147548 444292 147554 444304
rect 148318 444292 148324 444304
rect 147548 444264 148324 444292
rect 147548 444252 147554 444264
rect 148318 444252 148324 444264
rect 148376 444252 148382 444304
rect 191282 443980 191288 444032
rect 191340 444020 191346 444032
rect 191742 444020 191748 444032
rect 191340 443992 191748 444020
rect 191340 443980 191346 443992
rect 191742 443980 191748 443992
rect 191800 444020 191806 444032
rect 197354 444020 197360 444032
rect 191800 443992 197360 444020
rect 191800 443980 191806 443992
rect 197354 443980 197360 443992
rect 197412 443980 197418 444032
rect 358722 442960 358728 443012
rect 358780 443000 358786 443012
rect 372706 443000 372712 443012
rect 358780 442972 372712 443000
rect 358780 442960 358786 442972
rect 372706 442960 372712 442972
rect 372764 442960 372770 443012
rect 124122 441600 124128 441652
rect 124180 441640 124186 441652
rect 163498 441640 163504 441652
rect 124180 441612 163504 441640
rect 124180 441600 124186 441612
rect 163498 441600 163504 441612
rect 163556 441600 163562 441652
rect 195238 441396 195244 441448
rect 195296 441436 195302 441448
rect 197722 441436 197728 441448
rect 195296 441408 197728 441436
rect 195296 441396 195302 441408
rect 197722 441396 197728 441408
rect 197780 441396 197786 441448
rect 49602 440852 49608 440904
rect 49660 440892 49666 440904
rect 68278 440892 68284 440904
rect 49660 440864 68284 440892
rect 49660 440852 49666 440864
rect 68278 440852 68284 440864
rect 68336 440852 68342 440904
rect 358722 440240 358728 440292
rect 358780 440280 358786 440292
rect 367094 440280 367100 440292
rect 358780 440252 367100 440280
rect 358780 440240 358786 440252
rect 367094 440240 367100 440252
rect 367152 440240 367158 440292
rect 121638 440172 121644 440224
rect 121696 440212 121702 440224
rect 131758 440212 131764 440224
rect 121696 440184 131764 440212
rect 121696 440172 121702 440184
rect 131758 440172 131764 440184
rect 131816 440172 131822 440224
rect 65886 439628 65892 439680
rect 65944 439668 65950 439680
rect 66346 439668 66352 439680
rect 65944 439640 66352 439668
rect 65944 439628 65950 439640
rect 66346 439628 66352 439640
rect 66404 439628 66410 439680
rect 133138 439492 133144 439544
rect 133196 439532 133202 439544
rect 169018 439532 169024 439544
rect 133196 439504 169024 439532
rect 133196 439492 133202 439504
rect 169018 439492 169024 439504
rect 169076 439492 169082 439544
rect 180058 438880 180064 438932
rect 180116 438920 180122 438932
rect 197354 438920 197360 438932
rect 180116 438892 197360 438920
rect 180116 438880 180122 438892
rect 197354 438880 197360 438892
rect 197412 438880 197418 438932
rect 358722 438880 358728 438932
rect 358780 438920 358786 438932
rect 392578 438920 392584 438932
rect 358780 438892 392584 438920
rect 358780 438880 358786 438892
rect 392578 438880 392584 438892
rect 392636 438880 392642 438932
rect 124122 438812 124128 438864
rect 124180 438852 124186 438864
rect 132494 438852 132500 438864
rect 124180 438824 132500 438852
rect 124180 438812 124186 438824
rect 132494 438812 132500 438824
rect 132552 438852 132558 438864
rect 133782 438852 133788 438864
rect 132552 438824 133788 438852
rect 132552 438812 132558 438824
rect 133782 438812 133788 438824
rect 133840 438812 133846 438864
rect 53650 438132 53656 438184
rect 53708 438172 53714 438184
rect 60734 438172 60740 438184
rect 53708 438144 60740 438172
rect 53708 438132 53714 438144
rect 60734 438132 60740 438144
rect 60792 438132 60798 438184
rect 133782 438132 133788 438184
rect 133840 438172 133846 438184
rect 151078 438172 151084 438184
rect 133840 438144 151084 438172
rect 133840 438132 133846 438144
rect 151078 438132 151084 438144
rect 151136 438132 151142 438184
rect 60734 437452 60740 437504
rect 60792 437492 60798 437504
rect 61930 437492 61936 437504
rect 60792 437464 61936 437492
rect 60792 437452 60798 437464
rect 61930 437452 61936 437464
rect 61988 437492 61994 437504
rect 66806 437492 66812 437504
rect 61988 437464 66812 437492
rect 61988 437452 61994 437464
rect 66806 437452 66812 437464
rect 66864 437452 66870 437504
rect 124950 436704 124956 436756
rect 125008 436744 125014 436756
rect 157978 436744 157984 436756
rect 125008 436716 157984 436744
rect 125008 436704 125014 436716
rect 157978 436704 157984 436716
rect 158036 436704 158042 436756
rect 162210 436092 162216 436144
rect 162268 436132 162274 436144
rect 197354 436132 197360 436144
rect 162268 436104 197360 436132
rect 162268 436092 162274 436104
rect 197354 436092 197360 436104
rect 197412 436092 197418 436144
rect 357894 436092 357900 436144
rect 357952 436132 357958 436144
rect 360378 436132 360384 436144
rect 357952 436104 360384 436132
rect 357952 436092 357958 436104
rect 360378 436092 360384 436104
rect 360436 436092 360442 436144
rect 41230 435344 41236 435396
rect 41288 435384 41294 435396
rect 59078 435384 59084 435396
rect 41288 435356 59084 435384
rect 41288 435344 41294 435356
rect 59078 435344 59084 435356
rect 59136 435384 59142 435396
rect 66254 435384 66260 435396
rect 59136 435356 66260 435384
rect 59136 435344 59142 435356
rect 66254 435344 66260 435356
rect 66312 435344 66318 435396
rect 147490 434664 147496 434716
rect 147548 434704 147554 434716
rect 148410 434704 148416 434716
rect 147548 434676 148416 434704
rect 147548 434664 147554 434676
rect 148410 434664 148416 434676
rect 148468 434664 148474 434716
rect 44082 433304 44088 433356
rect 44140 433344 44146 433356
rect 54478 433344 54484 433356
rect 44140 433316 54484 433344
rect 44140 433304 44146 433316
rect 54478 433304 54484 433316
rect 54536 433344 54542 433356
rect 54536 433316 55214 433344
rect 54536 433304 54542 433316
rect 55186 433276 55214 433316
rect 124122 433304 124128 433356
rect 124180 433344 124186 433356
rect 147490 433344 147496 433356
rect 124180 433316 147496 433344
rect 124180 433304 124186 433316
rect 147490 433304 147496 433316
rect 147548 433304 147554 433356
rect 358722 433304 358728 433356
rect 358780 433344 358786 433356
rect 370038 433344 370044 433356
rect 358780 433316 370044 433344
rect 358780 433304 358786 433316
rect 370038 433304 370044 433316
rect 370096 433304 370102 433356
rect 66254 433276 66260 433288
rect 55186 433248 66260 433276
rect 66254 433236 66260 433248
rect 66312 433236 66318 433288
rect 124030 431876 124036 431928
rect 124088 431916 124094 431928
rect 142798 431916 142804 431928
rect 124088 431888 142804 431916
rect 124088 431876 124094 431888
rect 142798 431876 142804 431888
rect 142856 431876 142862 431928
rect 52362 431196 52368 431248
rect 52420 431236 52426 431248
rect 65886 431236 65892 431248
rect 52420 431208 65892 431236
rect 52420 431196 52426 431208
rect 65886 431196 65892 431208
rect 65944 431236 65950 431248
rect 66530 431236 66536 431248
rect 65944 431208 66536 431236
rect 65944 431196 65950 431208
rect 66530 431196 66536 431208
rect 66588 431196 66594 431248
rect 183462 430584 183468 430636
rect 183520 430624 183526 430636
rect 197354 430624 197360 430636
rect 183520 430596 197360 430624
rect 183520 430584 183526 430596
rect 197354 430584 197360 430596
rect 197412 430584 197418 430636
rect 358722 430584 358728 430636
rect 358780 430624 358786 430636
rect 371326 430624 371332 430636
rect 358780 430596 371332 430624
rect 358780 430584 358786 430596
rect 371326 430584 371332 430596
rect 371384 430584 371390 430636
rect 121362 429156 121368 429208
rect 121420 429196 121426 429208
rect 121638 429196 121644 429208
rect 121420 429168 121644 429196
rect 121420 429156 121426 429168
rect 121638 429156 121644 429168
rect 121696 429156 121702 429208
rect 36722 429088 36728 429140
rect 36780 429128 36786 429140
rect 37182 429128 37188 429140
rect 36780 429100 37188 429128
rect 36780 429088 36786 429100
rect 37182 429088 37188 429100
rect 37240 429128 37246 429140
rect 66806 429128 66812 429140
rect 37240 429100 66812 429128
rect 37240 429088 37246 429100
rect 66806 429088 66812 429100
rect 66864 429088 66870 429140
rect 14458 428408 14464 428460
rect 14516 428448 14522 428460
rect 36722 428448 36728 428460
rect 14516 428420 36728 428448
rect 14516 428408 14522 428420
rect 36722 428408 36728 428420
rect 36780 428408 36786 428460
rect 169018 427796 169024 427848
rect 169076 427836 169082 427848
rect 197354 427836 197360 427848
rect 169076 427808 197360 427836
rect 169076 427796 169082 427808
rect 197354 427796 197360 427808
rect 197412 427796 197418 427848
rect 358722 427796 358728 427848
rect 358780 427836 358786 427848
rect 382274 427836 382280 427848
rect 358780 427808 382280 427836
rect 358780 427796 358786 427808
rect 382274 427796 382280 427808
rect 382332 427796 382338 427848
rect 43990 427048 43996 427100
rect 44048 427088 44054 427100
rect 52454 427088 52460 427100
rect 44048 427060 52460 427088
rect 44048 427048 44054 427060
rect 52454 427048 52460 427060
rect 52512 427048 52518 427100
rect 140038 426436 140044 426488
rect 140096 426476 140102 426488
rect 197354 426476 197360 426488
rect 140096 426448 197360 426476
rect 140096 426436 140102 426448
rect 197354 426436 197360 426448
rect 197412 426436 197418 426488
rect 358722 426436 358728 426488
rect 358780 426476 358786 426488
rect 369946 426476 369952 426488
rect 358780 426448 369952 426476
rect 358780 426436 358786 426448
rect 369946 426436 369952 426448
rect 370004 426436 370010 426488
rect 52454 425688 52460 425740
rect 52512 425728 52518 425740
rect 53650 425728 53656 425740
rect 52512 425700 53656 425728
rect 52512 425688 52518 425700
rect 53650 425688 53656 425700
rect 53708 425728 53714 425740
rect 66806 425728 66812 425740
rect 53708 425700 66812 425728
rect 53708 425688 53714 425700
rect 66806 425688 66812 425700
rect 66864 425688 66870 425740
rect 59078 423648 59084 423700
rect 59136 423688 59142 423700
rect 66070 423688 66076 423700
rect 59136 423660 66076 423688
rect 59136 423648 59142 423660
rect 66070 423648 66076 423660
rect 66128 423648 66134 423700
rect 167638 423648 167644 423700
rect 167696 423688 167702 423700
rect 197354 423688 197360 423700
rect 167696 423660 197360 423688
rect 167696 423648 167702 423660
rect 197354 423648 197360 423660
rect 197412 423648 197418 423700
rect 3142 422900 3148 422952
rect 3200 422940 3206 422952
rect 17218 422940 17224 422952
rect 3200 422912 17224 422940
rect 3200 422900 3206 422912
rect 17218 422900 17224 422912
rect 17276 422900 17282 422952
rect 39942 421540 39948 421592
rect 40000 421580 40006 421592
rect 66070 421580 66076 421592
rect 40000 421552 66076 421580
rect 40000 421540 40006 421552
rect 66070 421540 66076 421552
rect 66128 421580 66134 421592
rect 66622 421580 66628 421592
rect 66128 421552 66628 421580
rect 66128 421540 66134 421552
rect 66622 421540 66628 421552
rect 66680 421540 66686 421592
rect 122926 421540 122932 421592
rect 122984 421580 122990 421592
rect 143442 421580 143448 421592
rect 122984 421552 143448 421580
rect 122984 421540 122990 421552
rect 143442 421540 143448 421552
rect 143500 421580 143506 421592
rect 178770 421580 178776 421592
rect 143500 421552 178776 421580
rect 143500 421540 143506 421552
rect 178770 421540 178776 421552
rect 178828 421540 178834 421592
rect 358722 420928 358728 420980
rect 358780 420968 358786 420980
rect 371418 420968 371424 420980
rect 358780 420940 371424 420968
rect 358780 420928 358786 420940
rect 371418 420928 371424 420940
rect 371476 420928 371482 420980
rect 124306 420860 124312 420912
rect 124364 420900 124370 420912
rect 160738 420900 160744 420912
rect 124364 420872 160744 420900
rect 124364 420860 124370 420872
rect 160738 420860 160744 420872
rect 160796 420860 160802 420912
rect 358078 420180 358084 420232
rect 358136 420220 358142 420232
rect 379514 420220 379520 420232
rect 358136 420192 379520 420220
rect 358136 420180 358142 420192
rect 379514 420180 379520 420192
rect 379572 420180 379578 420232
rect 181438 418140 181444 418192
rect 181496 418180 181502 418192
rect 197354 418180 197360 418192
rect 181496 418152 197360 418180
rect 181496 418140 181502 418152
rect 197354 418140 197360 418152
rect 197412 418140 197418 418192
rect 358722 418140 358728 418192
rect 358780 418180 358786 418192
rect 361666 418180 361672 418192
rect 358780 418152 361672 418180
rect 358780 418140 358786 418152
rect 361666 418140 361672 418152
rect 361724 418140 361730 418192
rect 195790 416780 195796 416832
rect 195848 416820 195854 416832
rect 197354 416820 197360 416832
rect 195848 416792 197360 416820
rect 195848 416780 195854 416792
rect 197354 416780 197360 416792
rect 197412 416780 197418 416832
rect 358722 416780 358728 416832
rect 358780 416820 358786 416832
rect 365806 416820 365812 416832
rect 358780 416792 365812 416820
rect 358780 416780 358786 416792
rect 365806 416780 365812 416792
rect 365864 416780 365870 416832
rect 122926 415148 122932 415200
rect 122984 415188 122990 415200
rect 129734 415188 129740 415200
rect 122984 415160 129740 415188
rect 122984 415148 122990 415160
rect 129734 415148 129740 415160
rect 129792 415148 129798 415200
rect 57790 414672 57796 414724
rect 57848 414712 57854 414724
rect 64782 414712 64788 414724
rect 57848 414684 64788 414712
rect 57848 414672 57854 414684
rect 64782 414672 64788 414684
rect 64840 414712 64846 414724
rect 66806 414712 66812 414724
rect 64840 414684 66812 414712
rect 64840 414672 64846 414684
rect 66806 414672 66812 414684
rect 66864 414672 66870 414724
rect 193950 413992 193956 414044
rect 194008 414032 194014 414044
rect 197354 414032 197360 414044
rect 194008 414004 197360 414032
rect 194008 413992 194014 414004
rect 197354 413992 197360 414004
rect 197412 413992 197418 414044
rect 358722 413992 358728 414044
rect 358780 414032 358786 414044
rect 365990 414032 365996 414044
rect 358780 414004 365996 414032
rect 358780 413992 358786 414004
rect 365990 413992 365996 414004
rect 366048 413992 366054 414044
rect 125686 413924 125692 413976
rect 125744 413964 125750 413976
rect 126974 413964 126980 413976
rect 125744 413936 126980 413964
rect 125744 413924 125750 413936
rect 126974 413924 126980 413936
rect 127032 413924 127038 413976
rect 124122 412700 124128 412752
rect 124180 412740 124186 412752
rect 125686 412740 125692 412752
rect 124180 412712 125692 412740
rect 124180 412700 124186 412712
rect 125686 412700 125692 412712
rect 125744 412700 125750 412752
rect 56410 411272 56416 411324
rect 56468 411312 56474 411324
rect 66714 411312 66720 411324
rect 56468 411284 66720 411312
rect 56468 411272 56474 411284
rect 66714 411272 66720 411284
rect 66772 411272 66778 411324
rect 164142 411272 164148 411324
rect 164200 411312 164206 411324
rect 197354 411312 197360 411324
rect 164200 411284 197360 411312
rect 164200 411272 164206 411284
rect 197354 411272 197360 411284
rect 197412 411272 197418 411324
rect 358722 411272 358728 411324
rect 358780 411312 358786 411324
rect 373994 411312 374000 411324
rect 358780 411284 374000 411312
rect 358780 411272 358786 411284
rect 373994 411272 374000 411284
rect 374052 411272 374058 411324
rect 130470 409776 130476 409828
rect 130528 409816 130534 409828
rect 197354 409816 197360 409828
rect 130528 409788 197360 409816
rect 130528 409776 130534 409788
rect 197354 409776 197360 409788
rect 197412 409776 197418 409828
rect 358722 408484 358728 408536
rect 358780 408524 358786 408536
rect 367370 408524 367376 408536
rect 358780 408496 367376 408524
rect 358780 408484 358786 408496
rect 367370 408484 367376 408496
rect 367428 408484 367434 408536
rect 124122 407736 124128 407788
rect 124180 407776 124186 407788
rect 134518 407776 134524 407788
rect 124180 407748 134524 407776
rect 124180 407736 124186 407748
rect 134518 407736 134524 407748
rect 134576 407736 134582 407788
rect 124122 406172 124128 406224
rect 124180 406212 124186 406224
rect 125502 406212 125508 406224
rect 124180 406184 125508 406212
rect 124180 406172 124186 406184
rect 125502 406172 125508 406184
rect 125560 406172 125566 406224
rect 57698 405764 57704 405816
rect 57756 405804 57762 405816
rect 64782 405804 64788 405816
rect 57756 405776 64788 405804
rect 57756 405764 57762 405776
rect 64782 405764 64788 405776
rect 64840 405804 64846 405816
rect 66346 405804 66352 405816
rect 64840 405776 66352 405804
rect 64840 405764 64846 405776
rect 66346 405764 66352 405776
rect 66404 405764 66410 405816
rect 189718 405696 189724 405748
rect 189776 405736 189782 405748
rect 197354 405736 197360 405748
rect 189776 405708 197360 405736
rect 189776 405696 189782 405708
rect 197354 405696 197360 405708
rect 197412 405696 197418 405748
rect 358722 405696 358728 405748
rect 358780 405736 358786 405748
rect 364518 405736 364524 405748
rect 358780 405708 364524 405736
rect 358780 405696 358786 405708
rect 364518 405696 364524 405708
rect 364576 405696 364582 405748
rect 48130 403588 48136 403640
rect 48188 403628 48194 403640
rect 62022 403628 62028 403640
rect 48188 403600 62028 403628
rect 48188 403588 48194 403600
rect 62022 403588 62028 403600
rect 62080 403628 62086 403640
rect 66346 403628 66352 403640
rect 62080 403600 66352 403628
rect 62080 403588 62086 403600
rect 66346 403588 66352 403600
rect 66404 403588 66410 403640
rect 358722 403452 358728 403504
rect 358780 403492 358786 403504
rect 363138 403492 363144 403504
rect 358780 403464 363144 403492
rect 358780 403452 358786 403464
rect 363138 403452 363144 403464
rect 363196 403452 363202 403504
rect 123846 403316 123852 403368
rect 123904 403356 123910 403368
rect 124950 403356 124956 403368
rect 123904 403328 124956 403356
rect 123904 403316 123910 403328
rect 124950 403316 124956 403328
rect 125008 403316 125014 403368
rect 125502 402296 125508 402348
rect 125560 402336 125566 402348
rect 127802 402336 127808 402348
rect 125560 402308 127808 402336
rect 125560 402296 125566 402308
rect 127802 402296 127808 402308
rect 127860 402296 127866 402348
rect 358722 401616 358728 401668
rect 358780 401656 358786 401668
rect 406378 401656 406384 401668
rect 358780 401628 406384 401656
rect 358780 401616 358786 401628
rect 406378 401616 406384 401628
rect 406436 401616 406442 401668
rect 123938 400868 123944 400920
rect 123996 400908 124002 400920
rect 194594 400908 194600 400920
rect 123996 400880 194600 400908
rect 123996 400868 124002 400880
rect 194594 400868 194600 400880
rect 194652 400868 194658 400920
rect 188982 400392 188988 400444
rect 189040 400432 189046 400444
rect 191282 400432 191288 400444
rect 189040 400404 191288 400432
rect 189040 400392 189046 400404
rect 191282 400392 191288 400404
rect 191340 400392 191346 400444
rect 50890 400188 50896 400240
rect 50948 400228 50954 400240
rect 55030 400228 55036 400240
rect 50948 400200 55036 400228
rect 50948 400188 50954 400200
rect 55030 400188 55036 400200
rect 55088 400228 55094 400240
rect 66346 400228 66352 400240
rect 55088 400200 66352 400228
rect 55088 400188 55094 400200
rect 66346 400188 66352 400200
rect 66404 400188 66410 400240
rect 194594 400188 194600 400240
rect 194652 400228 194658 400240
rect 195238 400228 195244 400240
rect 194652 400200 195244 400228
rect 194652 400188 194658 400200
rect 195238 400188 195244 400200
rect 195296 400188 195302 400240
rect 191742 398896 191748 398948
rect 191800 398936 191806 398948
rect 197354 398936 197360 398948
rect 191800 398908 197360 398936
rect 191800 398896 191806 398908
rect 197354 398896 197360 398908
rect 197412 398896 197418 398948
rect 48222 398828 48228 398880
rect 48280 398868 48286 398880
rect 50890 398868 50896 398880
rect 48280 398840 50896 398868
rect 48280 398828 48286 398840
rect 50890 398828 50896 398840
rect 50948 398868 50954 398880
rect 66346 398868 66352 398880
rect 50948 398840 66352 398868
rect 50948 398828 50954 398840
rect 66346 398828 66352 398840
rect 66404 398828 66410 398880
rect 124122 398828 124128 398880
rect 124180 398868 124186 398880
rect 125594 398868 125600 398880
rect 124180 398840 125600 398868
rect 124180 398828 124186 398840
rect 125594 398828 125600 398840
rect 125652 398868 125658 398880
rect 192570 398868 192576 398880
rect 125652 398840 192576 398868
rect 125652 398828 125658 398840
rect 192570 398828 192576 398840
rect 192628 398828 192634 398880
rect 358630 398828 358636 398880
rect 358688 398868 358694 398880
rect 361758 398868 361764 398880
rect 358688 398840 361764 398868
rect 358688 398828 358694 398840
rect 361758 398828 361764 398840
rect 361816 398828 361822 398880
rect 2774 398692 2780 398744
rect 2832 398732 2838 398744
rect 4798 398732 4804 398744
rect 2832 398704 4804 398732
rect 2832 398692 2838 398704
rect 4798 398692 4804 398704
rect 4856 398692 4862 398744
rect 125042 397468 125048 397520
rect 125100 397508 125106 397520
rect 191282 397508 191288 397520
rect 125100 397480 191288 397508
rect 125100 397468 125106 397480
rect 191282 397468 191288 397480
rect 191340 397508 191346 397520
rect 191742 397508 191748 397520
rect 191340 397480 191748 397508
rect 191340 397468 191346 397480
rect 191742 397468 191748 397480
rect 191800 397468 191806 397520
rect 35802 396720 35808 396772
rect 35860 396760 35866 396772
rect 66990 396760 66996 396772
rect 35860 396732 66996 396760
rect 35860 396720 35866 396732
rect 66990 396720 66996 396732
rect 67048 396720 67054 396772
rect 177850 396040 177856 396092
rect 177908 396080 177914 396092
rect 197354 396080 197360 396092
rect 177908 396052 197360 396080
rect 177908 396040 177914 396052
rect 197354 396040 197360 396052
rect 197412 396040 197418 396092
rect 121546 395972 121552 396024
rect 121604 396012 121610 396024
rect 127618 396012 127624 396024
rect 121604 395984 127624 396012
rect 121604 395972 121610 395984
rect 127618 395972 127624 395984
rect 127676 395972 127682 396024
rect 143350 394680 143356 394732
rect 143408 394720 143414 394732
rect 197354 394720 197360 394732
rect 143408 394692 197360 394720
rect 143408 394680 143414 394692
rect 197354 394680 197360 394692
rect 197412 394680 197418 394732
rect 123754 393932 123760 393984
rect 123812 393972 123818 393984
rect 160738 393972 160744 393984
rect 123812 393944 160744 393972
rect 123812 393932 123818 393944
rect 160738 393932 160744 393944
rect 160796 393932 160802 393984
rect 358722 393320 358728 393372
rect 358780 393360 358786 393372
rect 368658 393360 368664 393372
rect 358780 393332 368664 393360
rect 358780 393320 358786 393332
rect 368658 393320 368664 393332
rect 368716 393320 368722 393372
rect 63310 391960 63316 392012
rect 63368 392000 63374 392012
rect 66806 392000 66812 392012
rect 63368 391972 66812 392000
rect 63368 391960 63374 391972
rect 66806 391960 66812 391972
rect 66864 391960 66870 392012
rect 121454 391960 121460 392012
rect 121512 392000 121518 392012
rect 153930 392000 153936 392012
rect 121512 391972 153936 392000
rect 121512 391960 121518 391972
rect 153930 391960 153936 391972
rect 153988 391960 153994 392012
rect 3418 391212 3424 391264
rect 3476 391252 3482 391264
rect 131114 391252 131120 391264
rect 3476 391224 64874 391252
rect 3476 391212 3482 391224
rect 64846 391048 64874 391224
rect 113146 391224 131120 391252
rect 73338 391048 73344 391060
rect 64846 391020 73344 391048
rect 73338 391008 73344 391020
rect 73396 391008 73402 391060
rect 104066 391008 104072 391060
rect 104124 391048 104130 391060
rect 113146 391048 113174 391224
rect 131114 391212 131120 391224
rect 131172 391212 131178 391264
rect 104124 391020 113174 391048
rect 104124 391008 104130 391020
rect 120442 390260 120448 390312
rect 120500 390300 120506 390312
rect 120810 390300 120816 390312
rect 120500 390272 120816 390300
rect 120500 390260 120506 390272
rect 120810 390260 120816 390272
rect 120868 390260 120874 390312
rect 113082 389784 113088 389836
rect 113140 389824 113146 389836
rect 120626 389824 120632 389836
rect 113140 389796 120632 389824
rect 113140 389784 113146 389796
rect 120626 389784 120632 389796
rect 120684 389784 120690 389836
rect 59170 389240 59176 389292
rect 59228 389280 59234 389292
rect 87046 389280 87052 389292
rect 59228 389252 87052 389280
rect 59228 389240 59234 389252
rect 87046 389240 87052 389252
rect 87104 389240 87110 389292
rect 15838 389172 15844 389224
rect 15896 389212 15902 389224
rect 111426 389212 111432 389224
rect 15896 389184 111432 389212
rect 15896 389172 15902 389184
rect 111426 389172 111432 389184
rect 111484 389172 111490 389224
rect 67634 389104 67640 389156
rect 67692 389144 67698 389156
rect 68462 389144 68468 389156
rect 67692 389116 68468 389144
rect 67692 389104 67698 389116
rect 68462 389104 68468 389116
rect 68520 389104 68526 389156
rect 96154 389104 96160 389156
rect 96212 389144 96218 389156
rect 125042 389144 125048 389156
rect 96212 389116 125048 389144
rect 96212 389104 96218 389116
rect 125042 389104 125048 389116
rect 125100 389104 125106 389156
rect 65978 389036 65984 389088
rect 66036 389076 66042 389088
rect 73154 389076 73160 389088
rect 66036 389048 73160 389076
rect 66036 389036 66042 389048
rect 73154 389036 73160 389048
rect 73212 389076 73218 389088
rect 73798 389076 73804 389088
rect 73212 389048 73804 389076
rect 73212 389036 73218 389048
rect 73798 389036 73804 389048
rect 73856 389036 73862 389088
rect 101398 389036 101404 389088
rect 101456 389076 101462 389088
rect 103790 389076 103796 389088
rect 101456 389048 103796 389076
rect 101456 389036 101462 389048
rect 103790 389036 103796 389048
rect 103848 389036 103854 389088
rect 57606 388968 57612 389020
rect 57664 389008 57670 389020
rect 77846 389008 77852 389020
rect 57664 388980 77852 389008
rect 57664 388968 57670 388980
rect 77846 388968 77852 388980
rect 77904 388968 77910 389020
rect 88518 388628 88524 388680
rect 88576 388668 88582 388680
rect 92474 388668 92480 388680
rect 88576 388640 92480 388668
rect 88576 388628 88582 388640
rect 92474 388628 92480 388640
rect 92532 388628 92538 388680
rect 79502 388492 79508 388544
rect 79560 388532 79566 388544
rect 86218 388532 86224 388544
rect 79560 388504 86224 388532
rect 79560 388492 79566 388504
rect 86218 388492 86224 388504
rect 86276 388492 86282 388544
rect 93026 388424 93032 388476
rect 93084 388464 93090 388476
rect 98638 388464 98644 388476
rect 93084 388436 98644 388464
rect 93084 388424 93090 388436
rect 98638 388424 98644 388436
rect 98696 388424 98702 388476
rect 118970 388424 118976 388476
rect 119028 388464 119034 388476
rect 148410 388464 148416 388476
rect 119028 388436 148416 388464
rect 119028 388424 119034 388436
rect 148410 388424 148416 388436
rect 148468 388424 148474 388476
rect 167178 388424 167184 388476
rect 167236 388464 167242 388476
rect 168282 388464 168288 388476
rect 167236 388436 168288 388464
rect 167236 388424 167242 388436
rect 168282 388424 168288 388436
rect 168340 388464 168346 388476
rect 180242 388464 180248 388476
rect 168340 388436 180248 388464
rect 168340 388424 168346 388436
rect 180242 388424 180248 388436
rect 180300 388424 180306 388476
rect 66162 387744 66168 387796
rect 66220 387784 66226 387796
rect 82078 387784 82084 387796
rect 66220 387756 82084 387784
rect 66220 387744 66226 387756
rect 82078 387744 82084 387756
rect 82136 387744 82142 387796
rect 114462 387744 114468 387796
rect 114520 387784 114526 387796
rect 128354 387784 128360 387796
rect 114520 387756 128360 387784
rect 114520 387744 114526 387756
rect 128354 387744 128360 387756
rect 128412 387744 128418 387796
rect 171870 387132 171876 387184
rect 171928 387172 171934 387184
rect 181622 387172 181628 387184
rect 171928 387144 181628 387172
rect 171928 387132 171934 387144
rect 181622 387132 181628 387144
rect 181680 387132 181686 387184
rect 67818 387064 67824 387116
rect 67876 387104 67882 387116
rect 146938 387104 146944 387116
rect 67876 387076 146944 387104
rect 67876 387064 67882 387076
rect 146938 387064 146944 387076
rect 146996 387064 147002 387116
rect 147490 387064 147496 387116
rect 147548 387104 147554 387116
rect 178034 387104 178040 387116
rect 147548 387076 178040 387104
rect 147548 387064 147554 387076
rect 178034 387064 178040 387076
rect 178092 387064 178098 387116
rect 180334 387064 180340 387116
rect 180392 387104 180398 387116
rect 196710 387104 196716 387116
rect 180392 387076 196716 387104
rect 180392 387064 180398 387076
rect 196710 387064 196716 387076
rect 196768 387064 196774 387116
rect 181530 386384 181536 386436
rect 181588 386424 181594 386436
rect 197354 386424 197360 386436
rect 181588 386396 197360 386424
rect 181588 386384 181594 386396
rect 197354 386384 197360 386396
rect 197412 386384 197418 386436
rect 358722 386384 358728 386436
rect 358780 386424 358786 386436
rect 385126 386424 385132 386436
rect 358780 386396 385132 386424
rect 358780 386384 358786 386396
rect 385126 386384 385132 386396
rect 385184 386384 385190 386436
rect 63218 386316 63224 386368
rect 63276 386356 63282 386368
rect 80054 386356 80060 386368
rect 63276 386328 80060 386356
rect 63276 386316 63282 386328
rect 80054 386316 80060 386328
rect 80112 386356 80118 386368
rect 80882 386356 80888 386368
rect 80112 386328 80888 386356
rect 80112 386316 80118 386328
rect 80882 386316 80888 386328
rect 80940 386316 80946 386368
rect 99190 385704 99196 385756
rect 99248 385744 99254 385756
rect 122926 385744 122932 385756
rect 99248 385716 122932 385744
rect 99248 385704 99254 385716
rect 122926 385704 122932 385716
rect 122984 385704 122990 385756
rect 111426 385636 111432 385688
rect 111484 385676 111490 385688
rect 156690 385676 156696 385688
rect 111484 385648 156696 385676
rect 111484 385636 111490 385648
rect 156690 385636 156696 385648
rect 156748 385636 156754 385688
rect 123478 385024 123484 385076
rect 123536 385064 123542 385076
rect 189074 385064 189080 385076
rect 123536 385036 189080 385064
rect 123536 385024 123542 385036
rect 189074 385024 189080 385036
rect 189132 385024 189138 385076
rect 45462 384956 45468 385008
rect 45520 384996 45526 385008
rect 76558 384996 76564 385008
rect 45520 384968 76564 384996
rect 45520 384956 45526 384968
rect 76558 384956 76564 384968
rect 76616 384956 76622 385008
rect 73798 383664 73804 383716
rect 73856 383704 73862 383716
rect 184290 383704 184296 383716
rect 73856 383676 184296 383704
rect 73856 383664 73862 383676
rect 184290 383664 184296 383676
rect 184348 383664 184354 383716
rect 358722 383664 358728 383716
rect 358780 383704 358786 383716
rect 403618 383704 403624 383716
rect 358780 383676 403624 383704
rect 358780 383664 358786 383676
rect 403618 383664 403624 383676
rect 403676 383664 403682 383716
rect 17218 383596 17224 383648
rect 17276 383636 17282 383648
rect 125594 383636 125600 383648
rect 17276 383608 125600 383636
rect 17276 383596 17282 383608
rect 125594 383596 125600 383608
rect 125652 383596 125658 383648
rect 118602 382916 118608 382968
rect 118660 382956 118666 382968
rect 195974 382956 195980 382968
rect 118660 382928 195980 382956
rect 118660 382916 118666 382928
rect 195974 382916 195980 382928
rect 196032 382916 196038 382968
rect 80054 381488 80060 381540
rect 80112 381528 80118 381540
rect 166994 381528 167000 381540
rect 80112 381500 167000 381528
rect 80112 381488 80118 381500
rect 166994 381488 167000 381500
rect 167052 381488 167058 381540
rect 166994 380944 167000 380996
rect 167052 380984 167058 380996
rect 194502 380984 194508 380996
rect 167052 380956 194508 380984
rect 167052 380944 167058 380956
rect 194502 380944 194508 380956
rect 194560 380944 194566 380996
rect 3510 380876 3516 380928
rect 3568 380916 3574 380928
rect 104986 380916 104992 380928
rect 3568 380888 104992 380916
rect 3568 380876 3574 380888
rect 104986 380876 104992 380888
rect 105044 380916 105050 380928
rect 105538 380916 105544 380928
rect 105044 380888 105544 380916
rect 105044 380876 105050 380888
rect 105538 380876 105544 380888
rect 105596 380876 105602 380928
rect 109678 380876 109684 380928
rect 109736 380916 109742 380928
rect 171134 380916 171140 380928
rect 109736 380888 171140 380916
rect 109736 380876 109742 380888
rect 171134 380876 171140 380888
rect 171192 380916 171198 380928
rect 171870 380916 171876 380928
rect 171192 380888 171876 380916
rect 171192 380876 171198 380888
rect 171870 380876 171876 380888
rect 171928 380876 171934 380928
rect 39298 380128 39304 380180
rect 39356 380168 39362 380180
rect 125686 380168 125692 380180
rect 39356 380140 125692 380168
rect 39356 380128 39362 380140
rect 125686 380128 125692 380140
rect 125744 380128 125750 380180
rect 160738 380128 160744 380180
rect 160796 380168 160802 380180
rect 178126 380168 178132 380180
rect 160796 380140 178132 380168
rect 160796 380128 160802 380140
rect 178126 380128 178132 380140
rect 178184 380128 178190 380180
rect 178126 379584 178132 379636
rect 178184 379624 178190 379636
rect 178770 379624 178776 379636
rect 178184 379596 178776 379624
rect 178184 379584 178190 379596
rect 178770 379584 178776 379596
rect 178828 379624 178834 379636
rect 197354 379624 197360 379636
rect 178828 379596 197360 379624
rect 178828 379584 178834 379596
rect 197354 379584 197360 379596
rect 197412 379584 197418 379636
rect 48222 379516 48228 379568
rect 48280 379556 48286 379568
rect 188522 379556 188528 379568
rect 48280 379528 188528 379556
rect 48280 379516 48286 379528
rect 188522 379516 188528 379528
rect 188580 379516 188586 379568
rect 358630 379516 358636 379568
rect 358688 379556 358694 379568
rect 361574 379556 361580 379568
rect 358688 379528 361580 379556
rect 358688 379516 358694 379528
rect 361574 379516 361580 379528
rect 361632 379516 361638 379568
rect 110230 378768 110236 378820
rect 110288 378808 110294 378820
rect 160830 378808 160836 378820
rect 110288 378780 160836 378808
rect 110288 378768 110294 378780
rect 160830 378768 160836 378780
rect 160888 378768 160894 378820
rect 131298 378156 131304 378208
rect 131356 378196 131362 378208
rect 184198 378196 184204 378208
rect 131356 378168 184204 378196
rect 131356 378156 131362 378168
rect 184198 378156 184204 378168
rect 184256 378156 184262 378208
rect 50890 378088 50896 378140
rect 50948 378128 50954 378140
rect 187694 378128 187700 378140
rect 50948 378100 187700 378128
rect 50948 378088 50954 378100
rect 187694 378088 187700 378100
rect 187752 378088 187758 378140
rect 41230 378020 41236 378072
rect 41288 378060 41294 378072
rect 124398 378060 124404 378072
rect 41288 378032 124404 378060
rect 41288 378020 41294 378032
rect 124398 378020 124404 378032
rect 124456 378020 124462 378072
rect 124950 378020 124956 378072
rect 125008 378060 125014 378072
rect 130470 378060 130476 378072
rect 125008 378032 130476 378060
rect 125008 378020 125014 378032
rect 130470 378020 130476 378032
rect 130528 378020 130534 378072
rect 194410 377476 194416 377528
rect 194468 377516 194474 377528
rect 201586 377516 201592 377528
rect 194468 377488 201592 377516
rect 194468 377476 194474 377488
rect 201586 377476 201592 377488
rect 201644 377476 201650 377528
rect 189074 377408 189080 377460
rect 189132 377448 189138 377460
rect 194134 377448 194140 377460
rect 189132 377420 194140 377448
rect 189132 377408 189138 377420
rect 194134 377408 194140 377420
rect 194192 377408 194198 377460
rect 345658 377408 345664 377460
rect 345716 377448 345722 377460
rect 357710 377448 357716 377460
rect 345716 377420 357716 377448
rect 345716 377408 345722 377420
rect 357710 377408 357716 377420
rect 357768 377408 357774 377460
rect 198734 377272 198740 377324
rect 198792 377312 198798 377324
rect 199654 377312 199660 377324
rect 198792 377284 199660 377312
rect 198792 377272 198798 377284
rect 199654 377272 199660 377284
rect 199712 377272 199718 377324
rect 140682 376728 140688 376780
rect 140740 376768 140746 376780
rect 198734 376768 198740 376780
rect 140740 376740 198740 376768
rect 140740 376728 140746 376740
rect 198734 376728 198740 376740
rect 198792 376728 198798 376780
rect 192570 376660 192576 376712
rect 192628 376700 192634 376712
rect 215202 376700 215208 376712
rect 192628 376672 215208 376700
rect 192628 376660 192634 376672
rect 215202 376660 215208 376672
rect 215260 376660 215266 376712
rect 342898 376048 342904 376100
rect 342956 376088 342962 376100
rect 357618 376088 357624 376100
rect 342956 376060 357624 376088
rect 342956 376048 342962 376060
rect 357618 376048 357624 376060
rect 357676 376048 357682 376100
rect 81342 375980 81348 376032
rect 81400 376020 81406 376032
rect 95234 376020 95240 376032
rect 81400 375992 95240 376020
rect 81400 375980 81406 375992
rect 95234 375980 95240 375992
rect 95292 375980 95298 376032
rect 198826 375980 198832 376032
rect 198884 376020 198890 376032
rect 204346 376020 204352 376032
rect 198884 375992 204352 376020
rect 198884 375980 198890 375992
rect 204346 375980 204352 375992
rect 204404 375980 204410 376032
rect 247034 375980 247040 376032
rect 247092 376020 247098 376032
rect 248046 376020 248052 376032
rect 247092 375992 248052 376020
rect 247092 375980 247098 375992
rect 248046 375980 248052 375992
rect 248104 376020 248110 376032
rect 382918 376020 382924 376032
rect 248104 375992 382924 376020
rect 248104 375980 248110 375992
rect 382918 375980 382924 375992
rect 382976 375980 382982 376032
rect 104158 375436 104164 375488
rect 104216 375476 104222 375488
rect 195422 375476 195428 375488
rect 104216 375448 195428 375476
rect 104216 375436 104222 375448
rect 195422 375436 195428 375448
rect 195480 375436 195486 375488
rect 67542 375368 67548 375420
rect 67600 375408 67606 375420
rect 192662 375408 192668 375420
rect 67600 375380 192668 375408
rect 67600 375368 67606 375380
rect 192662 375368 192668 375380
rect 192720 375368 192726 375420
rect 195974 375300 195980 375352
rect 196032 375340 196038 375352
rect 196032 375312 200114 375340
rect 196032 375300 196038 375312
rect 200086 375272 200114 375312
rect 201678 375300 201684 375352
rect 201736 375340 201742 375352
rect 202782 375340 202788 375352
rect 201736 375312 202788 375340
rect 201736 375300 201742 375312
rect 202782 375300 202788 375312
rect 202840 375300 202846 375352
rect 205634 375300 205640 375352
rect 205692 375340 205698 375352
rect 206646 375340 206652 375352
rect 205692 375312 206652 375340
rect 205692 375300 205698 375312
rect 206646 375300 206652 375312
rect 206704 375300 206710 375352
rect 215202 375300 215208 375352
rect 215260 375340 215266 375352
rect 218238 375340 218244 375352
rect 215260 375312 218244 375340
rect 215260 375300 215266 375312
rect 218238 375300 218244 375312
rect 218296 375300 218302 375352
rect 258718 375300 258724 375352
rect 258776 375340 258782 375352
rect 261478 375340 261484 375352
rect 258776 375312 261484 375340
rect 258776 375300 258782 375312
rect 261478 375300 261484 375312
rect 261536 375300 261542 375352
rect 278130 375300 278136 375352
rect 278188 375340 278194 375352
rect 279694 375340 279700 375352
rect 278188 375312 279700 375340
rect 278188 375300 278194 375312
rect 279694 375300 279700 375312
rect 279752 375300 279758 375352
rect 298830 375300 298836 375352
rect 298888 375340 298894 375352
rect 301222 375340 301228 375352
rect 298888 375312 301228 375340
rect 298888 375300 298894 375312
rect 301222 375300 301228 375312
rect 301280 375300 301286 375352
rect 335998 375300 336004 375352
rect 336056 375340 336062 375352
rect 337838 375340 337844 375352
rect 336056 375312 337844 375340
rect 336056 375300 336062 375312
rect 337838 375300 337844 375312
rect 337896 375300 337902 375352
rect 339494 375300 339500 375352
rect 339552 375340 339558 375352
rect 378778 375340 378784 375352
rect 339552 375312 378784 375340
rect 339552 375300 339558 375312
rect 378778 375300 378784 375312
rect 378836 375300 378842 375352
rect 205652 375272 205680 375300
rect 200086 375244 205680 375272
rect 311894 375164 311900 375216
rect 311952 375204 311958 375216
rect 312814 375204 312820 375216
rect 311952 375176 312820 375204
rect 311952 375164 311958 375176
rect 312814 375164 312820 375176
rect 312872 375164 312878 375216
rect 233878 375028 233884 375080
rect 233936 375068 233942 375080
rect 238110 375068 238116 375080
rect 233936 375040 238116 375068
rect 233936 375028 233942 375040
rect 238110 375028 238116 375040
rect 238168 375028 238174 375080
rect 254670 374756 254676 374808
rect 254728 374796 254734 374808
rect 255406 374796 255412 374808
rect 254728 374768 255412 374796
rect 254728 374756 254734 374768
rect 255406 374756 255412 374768
rect 255464 374756 255470 374808
rect 250438 374688 250444 374740
rect 250496 374728 250502 374740
rect 251358 374728 251364 374740
rect 250496 374700 251364 374728
rect 250496 374688 250502 374700
rect 251358 374688 251364 374700
rect 251416 374688 251422 374740
rect 261478 374688 261484 374740
rect 261536 374728 261542 374740
rect 274726 374728 274732 374740
rect 261536 374700 274732 374728
rect 261536 374688 261542 374700
rect 274726 374688 274732 374700
rect 274784 374688 274790 374740
rect 295242 374688 295248 374740
rect 295300 374728 295306 374740
rect 296254 374728 296260 374740
rect 295300 374700 296260 374728
rect 295300 374688 295306 374700
rect 296254 374688 296260 374700
rect 296312 374688 296318 374740
rect 77938 374620 77944 374672
rect 77996 374660 78002 374672
rect 138658 374660 138664 374672
rect 77996 374632 138664 374660
rect 77996 374620 78002 374632
rect 138658 374620 138664 374632
rect 138716 374620 138722 374672
rect 209682 374620 209688 374672
rect 209740 374660 209746 374672
rect 216582 374660 216588 374672
rect 209740 374632 216588 374660
rect 209740 374620 209746 374632
rect 216582 374620 216588 374632
rect 216640 374620 216646 374672
rect 228358 374620 228364 374672
rect 228416 374660 228422 374672
rect 233142 374660 233148 374672
rect 228416 374632 233148 374660
rect 228416 374620 228422 374632
rect 233142 374620 233148 374632
rect 233200 374620 233206 374672
rect 262858 374620 262864 374672
rect 262916 374660 262922 374672
rect 294598 374660 294604 374672
rect 262916 374632 294604 374660
rect 262916 374620 262922 374632
rect 294598 374620 294604 374632
rect 294656 374620 294662 374672
rect 322198 374620 322204 374672
rect 322256 374660 322262 374672
rect 334526 374660 334532 374672
rect 322256 374632 334532 374660
rect 322256 374620 322262 374632
rect 334526 374620 334532 374632
rect 334584 374620 334590 374672
rect 334710 374620 334716 374672
rect 334768 374660 334774 374672
rect 339494 374660 339500 374672
rect 334768 374632 339500 374660
rect 334768 374620 334774 374632
rect 339494 374620 339500 374632
rect 339552 374620 339558 374672
rect 143534 374076 143540 374128
rect 143592 374116 143598 374128
rect 164878 374116 164884 374128
rect 143592 374088 164884 374116
rect 143592 374076 143598 374088
rect 164878 374076 164884 374088
rect 164936 374076 164942 374128
rect 200022 374076 200028 374128
rect 200080 374116 200086 374128
rect 201678 374116 201684 374128
rect 200080 374088 201684 374116
rect 200080 374076 200086 374088
rect 201678 374076 201684 374088
rect 201736 374076 201742 374128
rect 234614 374076 234620 374128
rect 234672 374116 234678 374128
rect 238018 374116 238024 374128
rect 234672 374088 238024 374116
rect 234672 374076 234678 374088
rect 238018 374076 238024 374088
rect 238076 374076 238082 374128
rect 246390 374076 246396 374128
rect 246448 374116 246454 374128
rect 255958 374116 255964 374128
rect 246448 374088 255964 374116
rect 246448 374076 246454 374088
rect 255958 374076 255964 374088
rect 256016 374076 256022 374128
rect 300210 374076 300216 374128
rect 300268 374116 300274 374128
rect 311894 374116 311900 374128
rect 300268 374088 311900 374116
rect 300268 374076 300274 374088
rect 311894 374076 311900 374088
rect 311952 374076 311958 374128
rect 119982 374008 119988 374060
rect 120040 374048 120046 374060
rect 120040 374020 195652 374048
rect 120040 374008 120046 374020
rect 195624 373980 195652 374020
rect 295978 374008 295984 374060
rect 296036 374048 296042 374060
rect 297910 374048 297916 374060
rect 296036 374020 297916 374048
rect 296036 374008 296042 374020
rect 297910 374008 297916 374020
rect 297968 374008 297974 374060
rect 307754 374008 307760 374060
rect 307812 374048 307818 374060
rect 313918 374048 313924 374060
rect 307812 374020 313924 374048
rect 307812 374008 307818 374020
rect 313918 374008 313924 374020
rect 313976 374008 313982 374060
rect 326338 374008 326344 374060
rect 326396 374048 326402 374060
rect 329098 374048 329104 374060
rect 326396 374020 329104 374048
rect 326396 374008 326402 374020
rect 329098 374008 329104 374020
rect 329156 374008 329162 374060
rect 354030 374008 354036 374060
rect 354088 374048 354094 374060
rect 356054 374048 356060 374060
rect 354088 374020 356060 374048
rect 354088 374008 354094 374020
rect 356054 374008 356060 374020
rect 356112 374008 356118 374060
rect 234614 373980 234620 373992
rect 195624 373952 234620 373980
rect 234614 373940 234620 373952
rect 234672 373940 234678 373992
rect 70302 373260 70308 373312
rect 70360 373300 70366 373312
rect 158714 373300 158720 373312
rect 70360 373272 158720 373300
rect 70360 373260 70366 373272
rect 158714 373260 158720 373272
rect 158772 373260 158778 373312
rect 350534 373260 350540 373312
rect 350592 373300 350598 373312
rect 452654 373300 452660 373312
rect 350592 373272 452660 373300
rect 350592 373260 350598 373272
rect 452654 373260 452660 373272
rect 452712 373260 452718 373312
rect 153930 372580 153936 372632
rect 153988 372620 153994 372632
rect 208394 372620 208400 372632
rect 153988 372592 208400 372620
rect 153988 372580 153994 372592
rect 208394 372580 208400 372592
rect 208452 372580 208458 372632
rect 184290 371832 184296 371884
rect 184348 371872 184354 371884
rect 206370 371872 206376 371884
rect 184348 371844 206376 371872
rect 184348 371832 184354 371844
rect 206370 371832 206376 371844
rect 206428 371832 206434 371884
rect 235258 371696 235264 371748
rect 235316 371736 235322 371748
rect 238754 371736 238760 371748
rect 235316 371708 238760 371736
rect 235316 371696 235322 371708
rect 238754 371696 238760 371708
rect 238812 371696 238818 371748
rect 134518 371492 134524 371544
rect 134576 371532 134582 371544
rect 135162 371532 135168 371544
rect 134576 371504 135168 371532
rect 134576 371492 134582 371504
rect 135162 371492 135168 371504
rect 135220 371492 135226 371544
rect 3234 371356 3240 371408
rect 3292 371396 3298 371408
rect 4798 371396 4804 371408
rect 3292 371368 4804 371396
rect 3292 371356 3298 371368
rect 4798 371356 4804 371368
rect 4856 371356 4862 371408
rect 117958 371288 117964 371340
rect 118016 371328 118022 371340
rect 169110 371328 169116 371340
rect 118016 371300 169116 371328
rect 118016 371288 118022 371300
rect 169110 371288 169116 371300
rect 169168 371288 169174 371340
rect 71682 371220 71688 371272
rect 71740 371260 71746 371272
rect 73798 371260 73804 371272
rect 71740 371232 73804 371260
rect 71740 371220 71746 371232
rect 73798 371220 73804 371232
rect 73856 371220 73862 371272
rect 135162 371220 135168 371272
rect 135220 371260 135226 371272
rect 196802 371260 196808 371272
rect 135220 371232 196808 371260
rect 135220 371220 135226 371232
rect 196802 371220 196808 371232
rect 196860 371220 196866 371272
rect 358170 371220 358176 371272
rect 358228 371260 358234 371272
rect 360470 371260 360476 371272
rect 358228 371232 360476 371260
rect 358228 371220 358234 371232
rect 360470 371220 360476 371232
rect 360528 371220 360534 371272
rect 86310 371152 86316 371204
rect 86368 371192 86374 371204
rect 148502 371192 148508 371204
rect 86368 371164 148508 371192
rect 86368 371152 86374 371164
rect 148502 371152 148508 371164
rect 148560 371152 148566 371204
rect 85574 370676 85580 370728
rect 85632 370716 85638 370728
rect 86310 370716 86316 370728
rect 85632 370688 86316 370716
rect 85632 370676 85638 370688
rect 86310 370676 86316 370688
rect 86368 370676 86374 370728
rect 53466 370472 53472 370524
rect 53524 370512 53530 370524
rect 143534 370512 143540 370524
rect 53524 370484 143540 370512
rect 53524 370472 53530 370484
rect 143534 370472 143540 370484
rect 143592 370472 143598 370524
rect 188522 370472 188528 370524
rect 188580 370512 188586 370524
rect 199562 370512 199568 370524
rect 188580 370484 199568 370512
rect 188580 370472 188586 370484
rect 199562 370472 199568 370484
rect 199620 370472 199626 370524
rect 199654 370472 199660 370524
rect 199712 370512 199718 370524
rect 242158 370512 242164 370524
rect 199712 370484 242164 370512
rect 199712 370472 199718 370484
rect 242158 370472 242164 370484
rect 242216 370472 242222 370524
rect 345014 370472 345020 370524
rect 345072 370512 345078 370524
rect 420914 370512 420920 370524
rect 345072 370484 420920 370512
rect 345072 370472 345078 370484
rect 420914 370472 420920 370484
rect 420972 370472 420978 370524
rect 146202 369860 146208 369912
rect 146260 369900 146266 369912
rect 207014 369900 207020 369912
rect 146260 369872 207020 369900
rect 146260 369860 146266 369872
rect 207014 369860 207020 369872
rect 207072 369900 207078 369912
rect 207658 369900 207664 369912
rect 207072 369872 207664 369900
rect 207072 369860 207078 369872
rect 207658 369860 207664 369872
rect 207716 369860 207722 369912
rect 343634 369792 343640 369844
rect 343692 369832 343698 369844
rect 344278 369832 344284 369844
rect 343692 369804 344284 369832
rect 343692 369792 343698 369804
rect 344278 369792 344284 369804
rect 344336 369832 344342 369844
rect 580350 369832 580356 369844
rect 344336 369804 580356 369832
rect 344336 369792 344342 369804
rect 580350 369792 580356 369804
rect 580408 369792 580414 369844
rect 98638 369180 98644 369232
rect 98696 369220 98702 369232
rect 151814 369220 151820 369232
rect 98696 369192 151820 369220
rect 98696 369180 98702 369192
rect 151814 369180 151820 369192
rect 151872 369180 151878 369232
rect 153838 369180 153844 369232
rect 153896 369220 153902 369232
rect 169202 369220 169208 369232
rect 153896 369192 169208 369220
rect 153896 369180 153902 369192
rect 169202 369180 169208 369192
rect 169260 369180 169266 369232
rect 191282 369180 191288 369232
rect 191340 369220 191346 369232
rect 267826 369220 267832 369232
rect 191340 369192 267832 369220
rect 191340 369180 191346 369192
rect 267826 369180 267832 369192
rect 267884 369180 267890 369232
rect 67726 369112 67732 369164
rect 67784 369152 67790 369164
rect 123478 369152 123484 369164
rect 67784 369124 123484 369152
rect 67784 369112 67790 369124
rect 123478 369112 123484 369124
rect 123536 369112 123542 369164
rect 145558 369112 145564 369164
rect 145616 369152 145622 369164
rect 202874 369152 202880 369164
rect 145616 369124 202880 369152
rect 145616 369112 145622 369124
rect 202874 369112 202880 369124
rect 202932 369152 202938 369164
rect 206278 369152 206284 369164
rect 202932 369124 206284 369152
rect 202932 369112 202938 369124
rect 206278 369112 206284 369124
rect 206336 369112 206342 369164
rect 232498 369112 232504 369164
rect 232556 369152 232562 369164
rect 361666 369152 361672 369164
rect 232556 369124 361672 369152
rect 232556 369112 232562 369124
rect 361666 369112 361672 369124
rect 361724 369112 361730 369164
rect 66162 368976 66168 369028
rect 66220 369016 66226 369028
rect 67634 369016 67640 369028
rect 66220 368988 67640 369016
rect 66220 368976 66226 368988
rect 67634 368976 67640 368988
rect 67692 368976 67698 369028
rect 197262 368432 197268 368484
rect 197320 368472 197326 368484
rect 200206 368472 200212 368484
rect 197320 368444 200212 368472
rect 197320 368432 197326 368444
rect 200206 368432 200212 368444
rect 200264 368432 200270 368484
rect 113818 367888 113824 367940
rect 113876 367928 113882 367940
rect 114462 367928 114468 367940
rect 113876 367900 114468 367928
rect 113876 367888 113882 367900
rect 114462 367888 114468 367900
rect 114520 367888 114526 367940
rect 348418 367820 348424 367872
rect 348476 367860 348482 367872
rect 364426 367860 364432 367872
rect 348476 367832 364432 367860
rect 348476 367820 348482 367832
rect 364426 367820 364432 367832
rect 364484 367820 364490 367872
rect 79962 367752 79968 367804
rect 80020 367792 80026 367804
rect 133138 367792 133144 367804
rect 80020 367764 133144 367792
rect 80020 367752 80026 367764
rect 133138 367752 133144 367764
rect 133196 367752 133202 367804
rect 345750 367752 345756 367804
rect 345808 367792 345814 367804
rect 365714 367792 365720 367804
rect 345808 367764 365720 367792
rect 345808 367752 345814 367764
rect 365714 367752 365720 367764
rect 365772 367752 365778 367804
rect 113818 367072 113824 367124
rect 113876 367112 113882 367124
rect 271874 367112 271880 367124
rect 113876 367084 271880 367112
rect 113876 367072 113882 367084
rect 271874 367072 271880 367084
rect 271932 367072 271938 367124
rect 340138 366392 340144 366444
rect 340196 366432 340202 366444
rect 356238 366432 356244 366444
rect 340196 366404 356244 366432
rect 340196 366392 340202 366404
rect 356238 366392 356244 366404
rect 356296 366392 356302 366444
rect 64782 366324 64788 366376
rect 64840 366364 64846 366376
rect 107746 366364 107752 366376
rect 64840 366336 107752 366364
rect 64840 366324 64846 366336
rect 107746 366324 107752 366336
rect 107804 366324 107810 366376
rect 341610 366324 341616 366376
rect 341668 366364 341674 366376
rect 367278 366364 367284 366376
rect 341668 366336 367284 366364
rect 341668 366324 341674 366336
rect 367278 366324 367284 366336
rect 367336 366324 367342 366376
rect 126238 365780 126244 365832
rect 126296 365820 126302 365832
rect 199378 365820 199384 365832
rect 126296 365792 199384 365820
rect 126296 365780 126302 365792
rect 199378 365780 199384 365792
rect 199436 365780 199442 365832
rect 144730 365712 144736 365764
rect 144788 365752 144794 365764
rect 340138 365752 340144 365764
rect 144788 365724 340144 365752
rect 144788 365712 144794 365724
rect 340138 365712 340144 365724
rect 340196 365712 340202 365764
rect 66898 365644 66904 365696
rect 66956 365684 66962 365696
rect 67358 365684 67364 365696
rect 66956 365656 67364 365684
rect 66956 365644 66962 365656
rect 67358 365644 67364 365656
rect 67416 365684 67422 365696
rect 359090 365684 359096 365696
rect 67416 365656 359096 365684
rect 67416 365644 67422 365656
rect 359090 365644 359096 365656
rect 359148 365644 359154 365696
rect 192754 364964 192760 365016
rect 192812 365004 192818 365016
rect 213822 365004 213828 365016
rect 192812 364976 213828 365004
rect 192812 364964 192818 364976
rect 213822 364964 213828 364976
rect 213880 364964 213886 365016
rect 358722 364964 358728 365016
rect 358780 365004 358786 365016
rect 370038 365004 370044 365016
rect 358780 364976 370044 365004
rect 358780 364964 358786 364976
rect 370038 364964 370044 364976
rect 370096 364964 370102 365016
rect 104894 364352 104900 364404
rect 104952 364392 104958 364404
rect 191282 364392 191288 364404
rect 104952 364364 191288 364392
rect 104952 364352 104958 364364
rect 191282 364352 191288 364364
rect 191340 364352 191346 364404
rect 281442 363672 281448 363724
rect 281500 363712 281506 363724
rect 413278 363712 413284 363724
rect 281500 363684 413284 363712
rect 281500 363672 281506 363684
rect 413278 363672 413284 363684
rect 413336 363672 413342 363724
rect 59078 363604 59084 363656
rect 59136 363644 59142 363656
rect 130378 363644 130384 363656
rect 59136 363616 130384 363644
rect 59136 363604 59142 363616
rect 130378 363604 130384 363616
rect 130436 363604 130442 363656
rect 166902 363604 166908 363656
rect 166960 363644 166966 363656
rect 309134 363644 309140 363656
rect 166960 363616 309140 363644
rect 166960 363604 166966 363616
rect 309134 363604 309140 363616
rect 309192 363604 309198 363656
rect 139302 362992 139308 363044
rect 139360 363032 139366 363044
rect 143350 363032 143356 363044
rect 139360 363004 143356 363032
rect 139360 362992 139366 363004
rect 143350 362992 143356 363004
rect 143408 362992 143414 363044
rect 110322 362924 110328 362976
rect 110380 362964 110386 362976
rect 196618 362964 196624 362976
rect 110380 362936 196624 362964
rect 110380 362924 110386 362936
rect 196618 362924 196624 362936
rect 196676 362924 196682 362976
rect 354582 362244 354588 362296
rect 354640 362284 354646 362296
rect 363046 362284 363052 362296
rect 354640 362256 363052 362284
rect 354640 362244 354646 362256
rect 363046 362244 363052 362256
rect 363104 362244 363110 362296
rect 70302 362176 70308 362228
rect 70360 362216 70366 362228
rect 175090 362216 175096 362228
rect 70360 362188 175096 362216
rect 70360 362176 70366 362188
rect 175090 362176 175096 362188
rect 175148 362216 175154 362228
rect 200758 362216 200764 362228
rect 175148 362188 200764 362216
rect 175148 362176 175154 362188
rect 200758 362176 200764 362188
rect 200816 362176 200822 362228
rect 338758 362176 338764 362228
rect 338816 362216 338822 362228
rect 361574 362216 361580 362228
rect 338816 362188 361580 362216
rect 338816 362176 338822 362188
rect 361574 362176 361580 362188
rect 361632 362176 361638 362228
rect 111794 361564 111800 361616
rect 111852 361604 111858 361616
rect 113082 361604 113088 361616
rect 111852 361576 113088 361604
rect 111852 361564 111858 361576
rect 113082 361564 113088 361576
rect 113140 361604 113146 361616
rect 232590 361604 232596 361616
rect 113140 361576 232596 361604
rect 113140 361564 113146 361576
rect 232590 361564 232596 361576
rect 232648 361564 232654 361616
rect 92198 360884 92204 360936
rect 92256 360924 92262 360936
rect 120810 360924 120816 360936
rect 92256 360896 120816 360924
rect 92256 360884 92262 360896
rect 120810 360884 120816 360896
rect 120868 360884 120874 360936
rect 81618 360816 81624 360868
rect 81676 360856 81682 360868
rect 82078 360856 82084 360868
rect 81676 360828 82084 360856
rect 81676 360816 81682 360828
rect 82078 360816 82084 360828
rect 82136 360856 82142 360868
rect 258166 360856 258172 360868
rect 82136 360828 258172 360856
rect 82136 360816 82142 360828
rect 258166 360816 258172 360828
rect 258224 360856 258230 360868
rect 258718 360856 258724 360868
rect 258224 360828 258724 360856
rect 258224 360816 258230 360828
rect 258718 360816 258724 360828
rect 258776 360816 258782 360868
rect 146110 360204 146116 360256
rect 146168 360244 146174 360256
rect 187050 360244 187056 360256
rect 146168 360216 187056 360244
rect 146168 360204 146174 360216
rect 187050 360204 187056 360216
rect 187108 360204 187114 360256
rect 101122 359524 101128 359576
rect 101180 359564 101186 359576
rect 177390 359564 177396 359576
rect 101180 359536 177396 359564
rect 101180 359524 101186 359536
rect 177390 359524 177396 359536
rect 177448 359524 177454 359576
rect 126974 359456 126980 359508
rect 127032 359496 127038 359508
rect 127710 359496 127716 359508
rect 127032 359468 127716 359496
rect 127032 359456 127038 359468
rect 127710 359456 127716 359468
rect 127768 359496 127774 359508
rect 259454 359496 259460 359508
rect 127768 359468 259460 359496
rect 127768 359456 127774 359468
rect 259454 359456 259460 359468
rect 259512 359456 259518 359508
rect 146938 358708 146944 358760
rect 146996 358748 147002 358760
rect 147582 358748 147588 358760
rect 146996 358720 147588 358748
rect 146996 358708 147002 358720
rect 147582 358708 147588 358720
rect 147640 358708 147646 358760
rect 3418 358572 3424 358624
rect 3476 358612 3482 358624
rect 7558 358612 7564 358624
rect 3476 358584 7564 358612
rect 3476 358572 3482 358584
rect 7558 358572 7564 358584
rect 7616 358572 7622 358624
rect 167730 358096 167736 358148
rect 167788 358136 167794 358148
rect 232498 358136 232504 358148
rect 167788 358108 232504 358136
rect 167788 358096 167794 358108
rect 232498 358096 232504 358108
rect 232556 358096 232562 358148
rect 56318 358028 56324 358080
rect 56376 358068 56382 358080
rect 109678 358068 109684 358080
rect 56376 358040 109684 358068
rect 56376 358028 56382 358040
rect 109678 358028 109684 358040
rect 109736 358028 109742 358080
rect 147582 358028 147588 358080
rect 147640 358068 147646 358080
rect 167086 358068 167092 358080
rect 147640 358040 167092 358068
rect 147640 358028 147646 358040
rect 167086 358028 167092 358040
rect 167144 358068 167150 358080
rect 167638 358068 167644 358080
rect 167144 358040 167644 358068
rect 167144 358028 167150 358040
rect 167638 358028 167644 358040
rect 167696 358028 167702 358080
rect 207658 358028 207664 358080
rect 207716 358068 207722 358080
rect 307018 358068 307024 358080
rect 207716 358040 307024 358068
rect 207716 358028 207722 358040
rect 307018 358028 307024 358040
rect 307076 358028 307082 358080
rect 107746 357416 107752 357468
rect 107804 357456 107810 357468
rect 206462 357456 206468 357468
rect 107804 357428 206468 357456
rect 107804 357416 107810 357428
rect 206462 357416 206468 357428
rect 206520 357416 206526 357468
rect 93762 357348 93768 357400
rect 93820 357388 93826 357400
rect 131022 357388 131028 357400
rect 93820 357360 131028 357388
rect 93820 357348 93826 357360
rect 131022 357348 131028 357360
rect 131080 357348 131086 357400
rect 229094 357348 229100 357400
rect 229152 357388 229158 357400
rect 238110 357388 238116 357400
rect 229152 357360 238116 357388
rect 229152 357348 229158 357360
rect 238110 357348 238116 357360
rect 238168 357348 238174 357400
rect 167086 356804 167092 356856
rect 167144 356844 167150 356856
rect 191190 356844 191196 356856
rect 167144 356816 191196 356844
rect 167144 356804 167150 356816
rect 191190 356804 191196 356816
rect 191248 356804 191254 356856
rect 140774 356736 140780 356788
rect 140832 356776 140838 356788
rect 141418 356776 141424 356788
rect 140832 356748 141424 356776
rect 140832 356736 140838 356748
rect 141418 356736 141424 356748
rect 141476 356776 141482 356788
rect 167730 356776 167736 356788
rect 141476 356748 167736 356776
rect 141476 356736 141482 356748
rect 167730 356736 167736 356748
rect 167788 356736 167794 356788
rect 194134 356736 194140 356788
rect 194192 356776 194198 356788
rect 227070 356776 227076 356788
rect 194192 356748 227076 356776
rect 194192 356736 194198 356748
rect 227070 356736 227076 356748
rect 227128 356736 227134 356788
rect 252554 356776 252560 356788
rect 238726 356748 252560 356776
rect 76558 356668 76564 356720
rect 76616 356708 76622 356720
rect 123018 356708 123024 356720
rect 76616 356680 123024 356708
rect 76616 356668 76622 356680
rect 123018 356668 123024 356680
rect 123076 356708 123082 356720
rect 124030 356708 124036 356720
rect 123076 356680 124036 356708
rect 123076 356668 123082 356680
rect 124030 356668 124036 356680
rect 124088 356668 124094 356720
rect 160738 356668 160744 356720
rect 160796 356708 160802 356720
rect 238726 356708 238754 356748
rect 252554 356736 252560 356748
rect 252612 356776 252618 356788
rect 300118 356776 300124 356788
rect 252612 356748 300124 356776
rect 252612 356736 252618 356748
rect 300118 356736 300124 356748
rect 300176 356736 300182 356788
rect 160796 356680 238754 356708
rect 160796 356668 160802 356680
rect 282178 356668 282184 356720
rect 282236 356708 282242 356720
rect 376938 356708 376944 356720
rect 282236 356680 376944 356708
rect 282236 356668 282242 356680
rect 376938 356668 376944 356680
rect 376996 356668 377002 356720
rect 96522 355376 96528 355428
rect 96580 355416 96586 355428
rect 99190 355416 99196 355428
rect 96580 355388 99196 355416
rect 96580 355376 96586 355388
rect 99190 355376 99196 355388
rect 99248 355376 99254 355428
rect 245654 355376 245660 355428
rect 245712 355416 245718 355428
rect 263594 355416 263600 355428
rect 245712 355388 263600 355416
rect 245712 355376 245718 355388
rect 263594 355376 263600 355388
rect 263652 355376 263658 355428
rect 84102 355308 84108 355360
rect 84160 355348 84166 355360
rect 108758 355348 108764 355360
rect 84160 355320 108764 355348
rect 84160 355308 84166 355320
rect 108758 355308 108764 355320
rect 108816 355308 108822 355360
rect 111702 355308 111708 355360
rect 111760 355348 111766 355360
rect 300210 355348 300216 355360
rect 111760 355320 300216 355348
rect 111760 355308 111766 355320
rect 300210 355308 300216 355320
rect 300268 355308 300274 355360
rect 309870 355308 309876 355360
rect 309928 355348 309934 355360
rect 358998 355348 359004 355360
rect 309928 355320 359004 355348
rect 309928 355308 309934 355320
rect 358998 355308 359004 355320
rect 359056 355308 359062 355360
rect 201586 355172 201592 355224
rect 201644 355212 201650 355224
rect 202138 355212 202144 355224
rect 201644 355184 202144 355212
rect 201644 355172 201650 355184
rect 202138 355172 202144 355184
rect 202196 355172 202202 355224
rect 102042 354696 102048 354748
rect 102100 354736 102106 354748
rect 201586 354736 201592 354748
rect 102100 354708 201592 354736
rect 102100 354696 102106 354708
rect 201586 354696 201592 354708
rect 201644 354696 201650 354748
rect 72418 354016 72424 354068
rect 72476 354056 72482 354068
rect 87046 354056 87052 354068
rect 72476 354028 87052 354056
rect 72476 354016 72482 354028
rect 87046 354016 87052 354028
rect 87104 354016 87110 354068
rect 273898 354016 273904 354068
rect 273956 354056 273962 354068
rect 295978 354056 295984 354068
rect 273956 354028 295984 354056
rect 273956 354016 273962 354028
rect 295978 354016 295984 354028
rect 296036 354016 296042 354068
rect 67726 353948 67732 354000
rect 67784 353988 67790 354000
rect 117958 353988 117964 354000
rect 67784 353960 117964 353988
rect 67784 353948 67790 353960
rect 117958 353948 117964 353960
rect 118016 353948 118022 354000
rect 195238 353948 195244 354000
rect 195296 353988 195302 354000
rect 211154 353988 211160 354000
rect 195296 353960 211160 353988
rect 195296 353948 195302 353960
rect 211154 353948 211160 353960
rect 211212 353948 211218 354000
rect 226978 353948 226984 354000
rect 227036 353988 227042 354000
rect 364518 353988 364524 354000
rect 227036 353960 364524 353988
rect 227036 353948 227042 353960
rect 364518 353948 364524 353960
rect 364576 353948 364582 354000
rect 121454 353336 121460 353388
rect 121512 353376 121518 353388
rect 177298 353376 177304 353388
rect 121512 353348 177304 353376
rect 121512 353336 121518 353348
rect 177298 353336 177304 353348
rect 177356 353336 177362 353388
rect 114462 353268 114468 353320
rect 114520 353308 114526 353320
rect 153838 353308 153844 353320
rect 114520 353280 153844 353308
rect 114520 353268 114526 353280
rect 153838 353268 153844 353280
rect 153896 353268 153902 353320
rect 154666 353268 154672 353320
rect 154724 353308 154730 353320
rect 155310 353308 155316 353320
rect 154724 353280 155316 353308
rect 154724 353268 154730 353280
rect 155310 353268 155316 353280
rect 155368 353308 155374 353320
rect 234522 353308 234528 353320
rect 155368 353280 234528 353308
rect 155368 353268 155374 353280
rect 234522 353268 234528 353280
rect 234580 353308 234586 353320
rect 240134 353308 240140 353320
rect 234580 353280 240140 353308
rect 234580 353268 234586 353280
rect 240134 353268 240140 353280
rect 240192 353268 240198 353320
rect 77202 352588 77208 352640
rect 77260 352628 77266 352640
rect 152458 352628 152464 352640
rect 77260 352600 152464 352628
rect 77260 352588 77266 352600
rect 152458 352588 152464 352600
rect 152516 352588 152522 352640
rect 152642 352588 152648 352640
rect 152700 352628 152706 352640
rect 223574 352628 223580 352640
rect 152700 352600 223580 352628
rect 152700 352588 152706 352600
rect 223574 352588 223580 352600
rect 223632 352588 223638 352640
rect 86862 352520 86868 352572
rect 86920 352560 86926 352572
rect 99374 352560 99380 352572
rect 86920 352532 99380 352560
rect 86920 352520 86926 352532
rect 99374 352520 99380 352532
rect 99432 352520 99438 352572
rect 105538 352520 105544 352572
rect 105596 352560 105602 352572
rect 181622 352560 181628 352572
rect 105596 352532 181628 352560
rect 105596 352520 105602 352532
rect 181622 352520 181628 352532
rect 181680 352520 181686 352572
rect 152642 351908 152648 351960
rect 152700 351948 152706 351960
rect 153102 351948 153108 351960
rect 152700 351920 153108 351948
rect 152700 351908 152706 351920
rect 153102 351908 153108 351920
rect 153160 351908 153166 351960
rect 223574 351908 223580 351960
rect 223632 351948 223638 351960
rect 224310 351948 224316 351960
rect 223632 351920 224316 351948
rect 223632 351908 223638 351920
rect 224310 351908 224316 351920
rect 224368 351908 224374 351960
rect 74442 351228 74448 351280
rect 74500 351268 74506 351280
rect 113818 351268 113824 351280
rect 74500 351240 113824 351268
rect 74500 351228 74506 351240
rect 113818 351228 113824 351240
rect 113876 351228 113882 351280
rect 90450 351160 90456 351212
rect 90508 351200 90514 351212
rect 195238 351200 195244 351212
rect 90508 351172 195244 351200
rect 90508 351160 90514 351172
rect 195238 351160 195244 351172
rect 195296 351160 195302 351212
rect 195330 351160 195336 351212
rect 195388 351200 195394 351212
rect 224218 351200 224224 351212
rect 195388 351172 224224 351200
rect 195388 351160 195394 351172
rect 224218 351160 224224 351172
rect 224276 351160 224282 351212
rect 120074 350548 120080 350600
rect 120132 350588 120138 350600
rect 120810 350588 120816 350600
rect 120132 350560 120816 350588
rect 120132 350548 120138 350560
rect 120810 350548 120816 350560
rect 120868 350588 120874 350600
rect 156782 350588 156788 350600
rect 120868 350560 156788 350588
rect 120868 350548 120874 350560
rect 156782 350548 156788 350560
rect 156840 350548 156846 350600
rect 121546 349868 121552 349920
rect 121604 349908 121610 349920
rect 126238 349908 126244 349920
rect 121604 349880 126244 349908
rect 121604 349868 121610 349880
rect 126238 349868 126244 349880
rect 126296 349868 126302 349920
rect 71590 349800 71596 349852
rect 71648 349840 71654 349852
rect 121454 349840 121460 349852
rect 71648 349812 121460 349840
rect 71648 349800 71654 349812
rect 121454 349800 121460 349812
rect 121512 349800 121518 349852
rect 192662 349800 192668 349852
rect 192720 349840 192726 349852
rect 202782 349840 202788 349852
rect 192720 349812 202788 349840
rect 192720 349800 192726 349812
rect 202782 349800 202788 349812
rect 202840 349840 202846 349852
rect 335354 349840 335360 349852
rect 202840 349812 335360 349840
rect 202840 349800 202846 349812
rect 335354 349800 335360 349812
rect 335412 349800 335418 349852
rect 126790 349188 126796 349240
rect 126848 349228 126854 349240
rect 176194 349228 176200 349240
rect 126848 349200 176200 349228
rect 126848 349188 126854 349200
rect 176194 349188 176200 349200
rect 176252 349188 176258 349240
rect 63218 349120 63224 349172
rect 63276 349160 63282 349172
rect 66898 349160 66904 349172
rect 63276 349132 66904 349160
rect 63276 349120 63282 349132
rect 66898 349120 66904 349132
rect 66956 349160 66962 349172
rect 67358 349160 67364 349172
rect 66956 349132 67364 349160
rect 66956 349120 66962 349132
rect 67358 349120 67364 349132
rect 67416 349120 67422 349172
rect 80146 349120 80152 349172
rect 80204 349160 80210 349172
rect 81342 349160 81348 349172
rect 80204 349132 81348 349160
rect 80204 349120 80210 349132
rect 81342 349120 81348 349132
rect 81400 349160 81406 349172
rect 195330 349160 195336 349172
rect 81400 349132 195336 349160
rect 81400 349120 81406 349132
rect 195330 349120 195336 349132
rect 195388 349120 195394 349172
rect 356698 349120 356704 349172
rect 356756 349160 356762 349172
rect 357342 349160 357348 349172
rect 356756 349132 357348 349160
rect 356756 349120 356762 349132
rect 357342 349120 357348 349132
rect 357400 349160 357406 349172
rect 400214 349160 400220 349172
rect 357400 349132 400220 349160
rect 357400 349120 357406 349132
rect 400214 349120 400220 349132
rect 400272 349120 400278 349172
rect 208486 349052 208492 349104
rect 208544 349092 208550 349104
rect 209038 349092 209044 349104
rect 208544 349064 209044 349092
rect 208544 349052 208550 349064
rect 209038 349052 209044 349064
rect 209096 349052 209102 349104
rect 241422 348440 241428 348492
rect 241480 348480 241486 348492
rect 357342 348480 357348 348492
rect 241480 348452 357348 348480
rect 241480 348440 241486 348452
rect 357342 348440 357348 348452
rect 357400 348440 357406 348492
rect 121730 348372 121736 348424
rect 121788 348412 121794 348424
rect 246390 348412 246396 348424
rect 121788 348384 246396 348412
rect 121788 348372 121794 348384
rect 246390 348372 246396 348384
rect 246448 348372 246454 348424
rect 90358 347760 90364 347812
rect 90416 347800 90422 347812
rect 209038 347800 209044 347812
rect 90416 347772 209044 347800
rect 90416 347760 90422 347772
rect 209038 347760 209044 347772
rect 209096 347760 209102 347812
rect 134978 347692 134984 347744
rect 135036 347732 135042 347744
rect 244274 347732 244280 347744
rect 135036 347704 244280 347732
rect 135036 347692 135042 347704
rect 244274 347692 244280 347704
rect 244332 347732 244338 347744
rect 244918 347732 244924 347744
rect 244332 347704 244924 347732
rect 244332 347692 244338 347704
rect 244918 347692 244924 347704
rect 244976 347692 244982 347744
rect 108298 347080 108304 347132
rect 108356 347120 108362 347132
rect 122098 347120 122104 347132
rect 108356 347092 122104 347120
rect 108356 347080 108362 347092
rect 122098 347080 122104 347092
rect 122156 347080 122162 347132
rect 81342 347012 81348 347064
rect 81400 347052 81406 347064
rect 133874 347052 133880 347064
rect 81400 347024 133880 347052
rect 81400 347012 81406 347024
rect 133874 347012 133880 347024
rect 133932 347052 133938 347064
rect 134978 347052 134984 347064
rect 133932 347024 134984 347052
rect 133932 347012 133938 347024
rect 134978 347012 134984 347024
rect 135036 347012 135042 347064
rect 185578 347012 185584 347064
rect 185636 347052 185642 347064
rect 204438 347052 204444 347064
rect 185636 347024 204444 347052
rect 185636 347012 185642 347024
rect 204438 347012 204444 347024
rect 204496 347012 204502 347064
rect 240870 347012 240876 347064
rect 240928 347052 240934 347064
rect 582926 347052 582932 347064
rect 240928 347024 582932 347052
rect 240928 347012 240934 347024
rect 582926 347012 582932 347024
rect 582984 347012 582990 347064
rect 140130 346400 140136 346452
rect 140188 346440 140194 346452
rect 162946 346440 162952 346452
rect 140188 346412 162952 346440
rect 140188 346400 140194 346412
rect 162946 346400 162952 346412
rect 163004 346400 163010 346452
rect 206462 346332 206468 346384
rect 206520 346372 206526 346384
rect 240134 346372 240140 346384
rect 206520 346344 240140 346372
rect 206520 346332 206526 346344
rect 240134 346332 240140 346344
rect 240192 346372 240198 346384
rect 241422 346372 241428 346384
rect 240192 346344 241428 346372
rect 240192 346332 240198 346344
rect 241422 346332 241428 346344
rect 241480 346332 241486 346384
rect 249610 346332 249616 346384
rect 249668 346372 249674 346384
rect 261478 346372 261484 346384
rect 249668 346344 261484 346372
rect 249668 346332 249674 346344
rect 261478 346332 261484 346344
rect 261536 346332 261542 346384
rect 124858 345652 124864 345704
rect 124916 345692 124922 345704
rect 248506 345692 248512 345704
rect 124916 345664 248512 345692
rect 124916 345652 124922 345664
rect 248506 345652 248512 345664
rect 248564 345692 248570 345704
rect 249610 345692 249616 345704
rect 248564 345664 249616 345692
rect 248564 345652 248570 345664
rect 249610 345652 249616 345664
rect 249668 345652 249674 345704
rect 59078 345040 59084 345092
rect 59136 345080 59142 345092
rect 197354 345080 197360 345092
rect 59136 345052 197360 345080
rect 59136 345040 59142 345052
rect 197354 345040 197360 345052
rect 197412 345040 197418 345092
rect 227622 344972 227628 345024
rect 227680 345012 227686 345024
rect 332594 345012 332600 345024
rect 227680 344984 332600 345012
rect 227680 344972 227686 344984
rect 332594 344972 332600 344984
rect 332652 344972 332658 345024
rect 227070 344428 227076 344480
rect 227128 344468 227134 344480
rect 227622 344468 227628 344480
rect 227128 344440 227628 344468
rect 227128 344428 227134 344440
rect 227622 344428 227628 344440
rect 227680 344428 227686 344480
rect 301314 344292 301320 344344
rect 301372 344332 301378 344344
rect 355318 344332 355324 344344
rect 301372 344304 355324 344332
rect 301372 344292 301378 344304
rect 355318 344292 355324 344304
rect 355376 344292 355382 344344
rect 67266 343680 67272 343732
rect 67324 343720 67330 343732
rect 156506 343720 156512 343732
rect 67324 343692 156512 343720
rect 67324 343680 67330 343692
rect 156506 343680 156512 343692
rect 156564 343680 156570 343732
rect 156690 343680 156696 343732
rect 156748 343720 156754 343732
rect 161474 343720 161480 343732
rect 156748 343692 161480 343720
rect 156748 343680 156754 343692
rect 161474 343680 161480 343692
rect 161532 343720 161538 343732
rect 221550 343720 221556 343732
rect 161532 343692 221556 343720
rect 161532 343680 161538 343692
rect 221550 343680 221556 343692
rect 221608 343680 221614 343732
rect 54938 343612 54944 343664
rect 54996 343652 55002 343664
rect 134794 343652 134800 343664
rect 54996 343624 134800 343652
rect 54996 343612 55002 343624
rect 134794 343612 134800 343624
rect 134852 343612 134858 343664
rect 137278 343612 137284 343664
rect 137336 343652 137342 343664
rect 228358 343652 228364 343664
rect 137336 343624 228364 343652
rect 137336 343612 137342 343624
rect 228358 343612 228364 343624
rect 228416 343612 228422 343664
rect 240778 343612 240784 343664
rect 240836 343652 240842 343664
rect 300946 343652 300952 343664
rect 240836 343624 300952 343652
rect 240836 343612 240842 343624
rect 300946 343612 300952 343624
rect 301004 343652 301010 343664
rect 301314 343652 301320 343664
rect 301004 343624 301320 343652
rect 301004 343612 301010 343624
rect 301314 343612 301320 343624
rect 301372 343612 301378 343664
rect 107562 343000 107568 343052
rect 107620 343040 107626 343052
rect 157334 343040 157340 343052
rect 107620 343012 157340 343040
rect 107620 343000 107626 343012
rect 157334 343000 157340 343012
rect 157392 343000 157398 343052
rect 199562 342932 199568 342984
rect 199620 342972 199626 342984
rect 215938 342972 215944 342984
rect 199620 342944 215944 342972
rect 199620 342932 199626 342944
rect 215938 342932 215944 342944
rect 215996 342932 216002 342984
rect 107470 342864 107476 342916
rect 107528 342904 107534 342916
rect 202230 342904 202236 342916
rect 107528 342876 202236 342904
rect 107528 342864 107534 342876
rect 202230 342864 202236 342876
rect 202288 342864 202294 342916
rect 232590 342864 232596 342916
rect 232648 342904 232654 342916
rect 260098 342904 260104 342916
rect 232648 342876 260104 342904
rect 232648 342864 232654 342876
rect 260098 342864 260104 342876
rect 260156 342864 260162 342916
rect 289722 342864 289728 342916
rect 289780 342904 289786 342916
rect 375466 342904 375472 342916
rect 289780 342876 375472 342904
rect 289780 342864 289786 342876
rect 375466 342864 375472 342876
rect 375524 342864 375530 342916
rect 61746 342252 61752 342304
rect 61804 342292 61810 342304
rect 66254 342292 66260 342304
rect 61804 342264 66260 342292
rect 61804 342252 61810 342264
rect 66254 342252 66260 342264
rect 66312 342292 66318 342304
rect 67358 342292 67364 342304
rect 66312 342264 67364 342292
rect 66312 342252 66318 342264
rect 67358 342252 67364 342264
rect 67416 342252 67422 342304
rect 77110 341504 77116 341556
rect 77168 341544 77174 341556
rect 87598 341544 87604 341556
rect 77168 341516 87604 341544
rect 77168 341504 77174 341516
rect 87598 341504 87604 341516
rect 87656 341504 87662 341556
rect 206370 341504 206376 341556
rect 206428 341544 206434 341556
rect 245102 341544 245108 341556
rect 206428 341516 245108 341544
rect 206428 341504 206434 341516
rect 245102 341504 245108 341516
rect 245160 341504 245166 341556
rect 117222 340960 117228 341012
rect 117280 341000 117286 341012
rect 183002 341000 183008 341012
rect 117280 340972 183008 341000
rect 117280 340960 117286 340972
rect 183002 340960 183008 340972
rect 183060 340960 183066 341012
rect 85574 340892 85580 340944
rect 85632 340932 85638 340944
rect 249886 340932 249892 340944
rect 85632 340904 249892 340932
rect 85632 340892 85638 340904
rect 249886 340892 249892 340904
rect 249944 340892 249950 340944
rect 78582 340212 78588 340264
rect 78640 340252 78646 340264
rect 95142 340252 95148 340264
rect 78640 340224 95148 340252
rect 78640 340212 78646 340224
rect 95142 340212 95148 340224
rect 95200 340212 95206 340264
rect 93486 340144 93492 340196
rect 93544 340184 93550 340196
rect 122190 340184 122196 340196
rect 93544 340156 122196 340184
rect 93544 340144 93550 340156
rect 122190 340144 122196 340156
rect 122248 340144 122254 340196
rect 135162 340144 135168 340196
rect 135220 340184 135226 340196
rect 139486 340184 139492 340196
rect 135220 340156 139492 340184
rect 135220 340144 135226 340156
rect 139486 340144 139492 340156
rect 139544 340144 139550 340196
rect 162946 340144 162952 340196
rect 163004 340184 163010 340196
rect 216674 340184 216680 340196
rect 163004 340156 216680 340184
rect 163004 340144 163010 340156
rect 216674 340144 216680 340156
rect 216732 340144 216738 340196
rect 156506 339872 156512 339924
rect 156564 339912 156570 339924
rect 158806 339912 158812 339924
rect 156564 339884 158812 339912
rect 156564 339872 156570 339884
rect 158806 339872 158812 339884
rect 158864 339872 158870 339924
rect 139394 339532 139400 339584
rect 139452 339572 139458 339584
rect 152458 339572 152464 339584
rect 139452 339544 152464 339572
rect 139452 339532 139458 339544
rect 152458 339532 152464 339544
rect 152516 339532 152522 339584
rect 95142 339464 95148 339516
rect 95200 339504 95206 339516
rect 248414 339504 248420 339516
rect 95200 339476 248420 339504
rect 95200 339464 95206 339476
rect 248414 339464 248420 339476
rect 248472 339464 248478 339516
rect 216122 338716 216128 338768
rect 216180 338756 216186 338768
rect 235994 338756 236000 338768
rect 216180 338728 236000 338756
rect 216180 338716 216186 338728
rect 235994 338716 236000 338728
rect 236052 338716 236058 338768
rect 236638 338716 236644 338768
rect 236696 338756 236702 338768
rect 263778 338756 263784 338768
rect 236696 338728 263784 338756
rect 236696 338716 236702 338728
rect 263778 338716 263784 338728
rect 263836 338716 263842 338768
rect 280798 338716 280804 338768
rect 280856 338756 280862 338768
rect 353938 338756 353944 338768
rect 280856 338728 353944 338756
rect 280856 338716 280862 338728
rect 353938 338716 353944 338728
rect 353996 338716 354002 338768
rect 85390 338376 85396 338428
rect 85448 338416 85454 338428
rect 90450 338416 90456 338428
rect 85448 338388 90456 338416
rect 85448 338376 85454 338388
rect 90450 338376 90456 338388
rect 90508 338376 90514 338428
rect 112346 338172 112352 338224
rect 112404 338212 112410 338224
rect 162302 338212 162308 338224
rect 112404 338184 162308 338212
rect 112404 338172 112410 338184
rect 162302 338172 162308 338184
rect 162360 338172 162366 338224
rect 106274 338104 106280 338156
rect 106332 338144 106338 338156
rect 229186 338144 229192 338156
rect 106332 338116 229192 338144
rect 106332 338104 106338 338116
rect 229186 338104 229192 338116
rect 229244 338104 229250 338156
rect 58618 337356 58624 337408
rect 58676 337396 58682 337408
rect 72418 337396 72424 337408
rect 58676 337368 72424 337396
rect 58676 337356 58682 337368
rect 72418 337356 72424 337368
rect 72476 337356 72482 337408
rect 97074 337356 97080 337408
rect 97132 337396 97138 337408
rect 128446 337396 128452 337408
rect 97132 337368 128452 337396
rect 97132 337356 97138 337368
rect 128446 337356 128452 337368
rect 128504 337396 128510 337408
rect 149238 337396 149244 337408
rect 128504 337368 149244 337396
rect 128504 337356 128510 337368
rect 149238 337356 149244 337368
rect 149296 337356 149302 337408
rect 196802 337356 196808 337408
rect 196860 337396 196866 337408
rect 260926 337396 260932 337408
rect 196860 337368 260932 337396
rect 196860 337356 196866 337368
rect 260926 337356 260932 337368
rect 260984 337356 260990 337408
rect 307110 337356 307116 337408
rect 307168 337396 307174 337408
rect 358170 337396 358176 337408
rect 307168 337368 358176 337396
rect 307168 337356 307174 337368
rect 358170 337356 358176 337368
rect 358228 337356 358234 337408
rect 150342 336812 150348 336864
rect 150400 336852 150406 336864
rect 199654 336852 199660 336864
rect 150400 336824 199660 336852
rect 150400 336812 150406 336824
rect 199654 336812 199660 336824
rect 199712 336812 199718 336864
rect 107838 336744 107844 336796
rect 107896 336784 107902 336796
rect 176102 336784 176108 336796
rect 107896 336756 176108 336784
rect 107896 336744 107902 336756
rect 176102 336744 176108 336756
rect 176160 336744 176166 336796
rect 134794 336676 134800 336728
rect 134852 336716 134858 336728
rect 154206 336716 154212 336728
rect 134852 336688 154212 336716
rect 134852 336676 134858 336688
rect 154206 336676 154212 336688
rect 154264 336676 154270 336728
rect 162946 336104 162952 336116
rect 142126 336076 162952 336104
rect 14 335996 20 336048
rect 72 336036 78 336048
rect 50982 336036 50988 336048
rect 72 336008 50988 336036
rect 72 335996 78 336008
rect 50982 335996 50988 336008
rect 51040 336036 51046 336048
rect 94222 336036 94228 336048
rect 51040 336008 94228 336036
rect 51040 335996 51046 336008
rect 94222 335996 94228 336008
rect 94280 335996 94286 336048
rect 118234 335996 118240 336048
rect 118292 336036 118298 336048
rect 133966 336036 133972 336048
rect 118292 336008 133972 336036
rect 118292 335996 118298 336008
rect 133966 335996 133972 336008
rect 134024 335996 134030 336048
rect 140038 335996 140044 336048
rect 140096 336036 140102 336048
rect 142126 336036 142154 336076
rect 162946 336064 162952 336076
rect 163004 336064 163010 336116
rect 140096 336008 142154 336036
rect 140096 335996 140102 336008
rect 153838 335996 153844 336048
rect 153896 336036 153902 336048
rect 224310 336036 224316 336048
rect 153896 336008 224316 336036
rect 153896 335996 153902 336008
rect 224310 335996 224316 336008
rect 224368 335996 224374 336048
rect 228450 335996 228456 336048
rect 228508 336036 228514 336048
rect 300854 336036 300860 336048
rect 228508 336008 300860 336036
rect 228508 335996 228514 336008
rect 300854 335996 300860 336008
rect 300912 335996 300918 336048
rect 154666 335724 154672 335776
rect 154724 335764 154730 335776
rect 155862 335764 155868 335776
rect 154724 335736 155868 335764
rect 154724 335724 154730 335736
rect 155862 335724 155868 335736
rect 155920 335764 155926 335776
rect 158898 335764 158904 335776
rect 155920 335736 158904 335764
rect 155920 335724 155926 335736
rect 158898 335724 158904 335736
rect 158956 335724 158962 335776
rect 61930 335316 61936 335368
rect 61988 335356 61994 335368
rect 132494 335356 132500 335368
rect 61988 335328 132500 335356
rect 61988 335316 61994 335328
rect 132494 335316 132500 335328
rect 132552 335316 132558 335368
rect 64506 334568 64512 334620
rect 64564 334608 64570 334620
rect 108298 334608 108304 334620
rect 64564 334580 108304 334608
rect 64564 334568 64570 334580
rect 108298 334568 108304 334580
rect 108356 334568 108362 334620
rect 135162 334024 135168 334076
rect 135220 334064 135226 334076
rect 158898 334064 158904 334076
rect 135220 334036 158904 334064
rect 135220 334024 135226 334036
rect 158898 334024 158904 334036
rect 158956 334024 158962 334076
rect 104434 333956 104440 334008
rect 104492 333996 104498 334008
rect 170582 333996 170588 334008
rect 104492 333968 170588 333996
rect 104492 333956 104498 333968
rect 170582 333956 170588 333968
rect 170640 333956 170646 334008
rect 154758 333276 154764 333328
rect 154816 333316 154822 333328
rect 217318 333316 217324 333328
rect 154816 333288 217324 333316
rect 154816 333276 154822 333288
rect 217318 333276 217324 333288
rect 217376 333276 217382 333328
rect 75638 333208 75644 333260
rect 75696 333248 75702 333260
rect 140130 333248 140136 333260
rect 75696 333220 140136 333248
rect 75696 333208 75702 333220
rect 140130 333208 140136 333220
rect 140188 333208 140194 333260
rect 195974 333208 195980 333260
rect 196032 333248 196038 333260
rect 582374 333248 582380 333260
rect 196032 333220 582380 333248
rect 196032 333208 196038 333220
rect 582374 333208 582380 333220
rect 582432 333208 582438 333260
rect 67818 332596 67824 332648
rect 67876 332636 67882 332648
rect 71774 332636 71780 332648
rect 67876 332608 71780 332636
rect 67876 332596 67882 332608
rect 71774 332596 71780 332608
rect 71832 332596 71838 332648
rect 148134 332596 148140 332648
rect 148192 332636 148198 332648
rect 158254 332636 158260 332648
rect 148192 332608 158260 332636
rect 148192 332596 148198 332608
rect 158254 332596 158260 332608
rect 158312 332596 158318 332648
rect 260098 332528 260104 332580
rect 260156 332568 260162 332580
rect 344278 332568 344284 332580
rect 260156 332540 344284 332568
rect 260156 332528 260162 332540
rect 344278 332528 344284 332540
rect 344336 332528 344342 332580
rect 166350 332188 166356 332240
rect 166408 332228 166414 332240
rect 168374 332228 168380 332240
rect 166408 332200 168380 332228
rect 166408 332188 166414 332200
rect 168374 332188 168380 332200
rect 168432 332188 168438 332240
rect 76650 332120 76656 332172
rect 76708 332160 76714 332172
rect 77110 332160 77116 332172
rect 76708 332132 77116 332160
rect 76708 332120 76714 332132
rect 77110 332120 77116 332132
rect 77168 332120 77174 332172
rect 83090 332120 83096 332172
rect 83148 332160 83154 332172
rect 84102 332160 84108 332172
rect 83148 332132 84108 332160
rect 83148 332120 83154 332132
rect 84102 332120 84108 332132
rect 84160 332120 84166 332172
rect 91922 332120 91928 332172
rect 91980 332160 91986 332172
rect 92382 332160 92388 332172
rect 91980 332132 92388 332160
rect 91980 332120 91986 332132
rect 92382 332120 92388 332132
rect 92440 332120 92446 332172
rect 95602 332120 95608 332172
rect 95660 332160 95666 332172
rect 96338 332160 96344 332172
rect 95660 332132 96344 332160
rect 95660 332120 95666 332132
rect 96338 332120 96344 332132
rect 96396 332120 96402 332172
rect 100018 332120 100024 332172
rect 100076 332160 100082 332172
rect 100570 332160 100576 332172
rect 100076 332132 100576 332160
rect 100076 332120 100082 332132
rect 100570 332120 100576 332132
rect 100628 332120 100634 332172
rect 102962 332120 102968 332172
rect 103020 332160 103026 332172
rect 103422 332160 103428 332172
rect 103020 332132 103428 332160
rect 103020 332120 103026 332132
rect 103422 332120 103428 332132
rect 103480 332120 103486 332172
rect 113818 332120 113824 332172
rect 113876 332160 113882 332172
rect 114370 332160 114376 332172
rect 113876 332132 114376 332160
rect 113876 332120 113882 332132
rect 114370 332120 114376 332132
rect 114428 332120 114434 332172
rect 116762 332120 116768 332172
rect 116820 332160 116826 332172
rect 117222 332160 117228 332172
rect 116820 332132 117228 332160
rect 116820 332120 116826 332132
rect 117222 332120 117228 332132
rect 117280 332120 117286 332172
rect 177390 331916 177396 331968
rect 177448 331956 177454 331968
rect 200850 331956 200856 331968
rect 177448 331928 200856 331956
rect 177448 331916 177454 331928
rect 200850 331916 200856 331928
rect 200908 331916 200914 331968
rect 70762 331848 70768 331900
rect 70820 331888 70826 331900
rect 71498 331888 71504 331900
rect 70820 331860 71504 331888
rect 70820 331848 70826 331860
rect 71498 331848 71504 331860
rect 71556 331848 71562 331900
rect 156598 331848 156604 331900
rect 156656 331888 156662 331900
rect 166258 331888 166264 331900
rect 156656 331860 166264 331888
rect 156656 331848 156662 331860
rect 166258 331848 166264 331860
rect 166316 331848 166322 331900
rect 167638 331848 167644 331900
rect 167696 331888 167702 331900
rect 195422 331888 195428 331900
rect 167696 331860 195428 331888
rect 167696 331848 167702 331860
rect 195422 331848 195428 331860
rect 195480 331848 195486 331900
rect 195514 331848 195520 331900
rect 195572 331888 195578 331900
rect 261018 331888 261024 331900
rect 195572 331860 261024 331888
rect 195572 331848 195578 331860
rect 261018 331848 261024 331860
rect 261076 331848 261082 331900
rect 146754 331780 146760 331832
rect 146812 331820 146818 331832
rect 150342 331820 150348 331832
rect 146812 331792 150348 331820
rect 146812 331780 146818 331792
rect 150342 331780 150348 331792
rect 150400 331780 150406 331832
rect 79962 331712 79968 331764
rect 80020 331752 80026 331764
rect 84378 331752 84384 331764
rect 80020 331724 84384 331752
rect 80020 331712 80026 331724
rect 84378 331712 84384 331724
rect 84436 331712 84442 331764
rect 88242 331712 88248 331764
rect 88300 331752 88306 331764
rect 90358 331752 90364 331764
rect 88300 331724 90364 331752
rect 88300 331712 88306 331724
rect 90358 331712 90364 331724
rect 90416 331712 90422 331764
rect 132770 331644 132776 331696
rect 132828 331684 132834 331696
rect 133782 331684 133788 331696
rect 132828 331656 133788 331684
rect 132828 331644 132834 331656
rect 133782 331644 133788 331656
rect 133840 331644 133846 331696
rect 80238 331576 80244 331628
rect 80296 331616 80302 331628
rect 81342 331616 81348 331628
rect 80296 331588 81348 331616
rect 80296 331576 80302 331588
rect 81342 331576 81348 331588
rect 81400 331576 81406 331628
rect 118878 331576 118884 331628
rect 118936 331616 118942 331628
rect 119890 331616 119896 331628
rect 118936 331588 119896 331616
rect 118936 331576 118942 331588
rect 119890 331576 119896 331588
rect 119948 331576 119954 331628
rect 123386 331576 123392 331628
rect 123444 331616 123450 331628
rect 124122 331616 124128 331628
rect 123444 331588 124128 331616
rect 123444 331576 123450 331588
rect 124122 331576 124128 331588
rect 124180 331576 124186 331628
rect 109402 331508 109408 331560
rect 109460 331548 109466 331560
rect 110322 331548 110328 331560
rect 109460 331520 110328 331548
rect 109460 331508 109466 331520
rect 110322 331508 110328 331520
rect 110380 331508 110386 331560
rect 129274 331508 129280 331560
rect 129332 331548 129338 331560
rect 135162 331548 135168 331560
rect 129332 331520 135168 331548
rect 129332 331508 129338 331520
rect 135162 331508 135168 331520
rect 135220 331508 135226 331560
rect 88978 331440 88984 331492
rect 89036 331480 89042 331492
rect 89622 331480 89628 331492
rect 89036 331452 89628 331480
rect 89036 331440 89042 331452
rect 89622 331440 89628 331452
rect 89680 331440 89686 331492
rect 90450 331440 90456 331492
rect 90508 331480 90514 331492
rect 93118 331480 93124 331492
rect 90508 331452 93124 331480
rect 90508 331440 90514 331452
rect 93118 331440 93124 331452
rect 93176 331440 93182 331492
rect 94130 331440 94136 331492
rect 94188 331480 94194 331492
rect 95142 331480 95148 331492
rect 94188 331452 95148 331480
rect 94188 331440 94194 331452
rect 95142 331440 95148 331452
rect 95200 331440 95206 331492
rect 98546 331440 98552 331492
rect 98604 331480 98610 331492
rect 99282 331480 99288 331492
rect 98604 331452 99288 331480
rect 98604 331440 98610 331452
rect 99282 331440 99288 331452
rect 99340 331440 99346 331492
rect 124122 331440 124128 331492
rect 124180 331480 124186 331492
rect 124858 331480 124864 331492
rect 124180 331452 124864 331480
rect 124180 331440 124186 331452
rect 124858 331440 124864 331452
rect 124916 331440 124922 331492
rect 130010 331440 130016 331492
rect 130068 331480 130074 331492
rect 131022 331480 131028 331492
rect 130068 331452 131028 331480
rect 130068 331440 130074 331452
rect 131022 331440 131028 331452
rect 131080 331440 131086 331492
rect 138658 331440 138664 331492
rect 138716 331480 138722 331492
rect 139302 331480 139308 331492
rect 138716 331452 139308 331480
rect 138716 331440 138722 331452
rect 139302 331440 139308 331452
rect 139360 331440 139366 331492
rect 143074 331372 143080 331424
rect 143132 331412 143138 331424
rect 144914 331412 144920 331424
rect 143132 331384 144920 331412
rect 143132 331372 143138 331384
rect 144914 331372 144920 331384
rect 144972 331372 144978 331424
rect 153028 331384 153240 331412
rect 50982 331304 50988 331356
rect 51040 331344 51046 331356
rect 69290 331344 69296 331356
rect 51040 331316 69296 331344
rect 51040 331304 51046 331316
rect 69290 331304 69296 331316
rect 69348 331304 69354 331356
rect 72234 331304 72240 331356
rect 72292 331344 72298 331356
rect 75638 331344 75644 331356
rect 72292 331316 75644 331344
rect 72292 331304 72298 331316
rect 75638 331304 75644 331316
rect 75696 331304 75702 331356
rect 110874 331304 110880 331356
rect 110932 331344 110938 331356
rect 111702 331344 111708 331356
rect 110932 331316 111708 331344
rect 110932 331304 110938 331316
rect 111702 331304 111708 331316
rect 111760 331304 111766 331356
rect 119982 331304 119988 331356
rect 120040 331344 120046 331356
rect 120534 331344 120540 331356
rect 120040 331316 120540 331344
rect 120040 331304 120046 331316
rect 120534 331304 120540 331316
rect 120592 331304 120598 331356
rect 143810 331304 143816 331356
rect 143868 331344 143874 331356
rect 144730 331344 144736 331356
rect 143868 331316 144736 331344
rect 143868 331304 143874 331316
rect 144730 331304 144736 331316
rect 144788 331304 144794 331356
rect 151170 331304 151176 331356
rect 151228 331344 151234 331356
rect 152918 331344 152924 331356
rect 151228 331316 152924 331344
rect 151228 331304 151234 331316
rect 152918 331304 152924 331316
rect 152976 331304 152982 331356
rect 67358 331236 67364 331288
rect 67416 331276 67422 331288
rect 153028 331276 153056 331384
rect 67416 331248 153056 331276
rect 153212 331276 153240 331384
rect 154114 331304 154120 331356
rect 154172 331344 154178 331356
rect 158990 331344 158996 331356
rect 154172 331316 158996 331344
rect 154172 331304 154178 331316
rect 158990 331304 158996 331316
rect 159048 331304 159054 331356
rect 153212 331248 156644 331276
rect 67416 331236 67422 331248
rect 49602 331168 49608 331220
rect 49660 331208 49666 331220
rect 137002 331208 137008 331220
rect 49660 331180 137008 331208
rect 49660 331168 49666 331180
rect 137002 331168 137008 331180
rect 137060 331208 137066 331220
rect 137278 331208 137284 331220
rect 137060 331180 137284 331208
rect 137060 331168 137066 331180
rect 137278 331168 137284 331180
rect 137336 331168 137342 331220
rect 144914 331168 144920 331220
rect 144972 331208 144978 331220
rect 153010 331208 153016 331220
rect 144972 331180 153016 331208
rect 144972 331168 144978 331180
rect 153010 331168 153016 331180
rect 153068 331168 153074 331220
rect 156616 331208 156644 331248
rect 260098 331236 260104 331288
rect 260156 331276 260162 331288
rect 260742 331276 260748 331288
rect 260156 331248 260748 331276
rect 260156 331236 260162 331248
rect 260742 331236 260748 331248
rect 260800 331236 260806 331288
rect 157426 331208 157432 331220
rect 156616 331180 157432 331208
rect 157426 331168 157432 331180
rect 157484 331168 157490 331220
rect 298002 331168 298008 331220
rect 298060 331208 298066 331220
rect 371234 331208 371240 331220
rect 298060 331180 371240 331208
rect 298060 331168 298066 331180
rect 371234 331168 371240 331180
rect 371292 331168 371298 331220
rect 152918 331100 152924 331152
rect 152976 331140 152982 331152
rect 156046 331140 156052 331152
rect 152976 331112 156052 331140
rect 152976 331100 152982 331112
rect 156046 331100 156052 331112
rect 156104 331100 156110 331152
rect 167730 330964 167736 331016
rect 167788 331004 167794 331016
rect 169110 331004 169116 331016
rect 167788 330976 169116 331004
rect 167788 330964 167794 330976
rect 169110 330964 169116 330976
rect 169168 330964 169174 331016
rect 162946 330828 162952 330880
rect 163004 330868 163010 330880
rect 165614 330868 165620 330880
rect 163004 330840 165620 330868
rect 163004 330828 163010 330840
rect 165614 330828 165620 330840
rect 165672 330828 165678 330880
rect 150342 330556 150348 330608
rect 150400 330596 150406 330608
rect 155862 330596 155868 330608
rect 150400 330568 155868 330596
rect 150400 330556 150406 330568
rect 155862 330556 155868 330568
rect 155920 330556 155926 330608
rect 165890 330556 165896 330608
rect 165948 330596 165954 330608
rect 199562 330596 199568 330608
rect 165948 330568 199568 330596
rect 165948 330556 165954 330568
rect 199562 330556 199568 330568
rect 199620 330556 199626 330608
rect 245010 330556 245016 330608
rect 245068 330596 245074 330608
rect 305730 330596 305736 330608
rect 245068 330568 305736 330596
rect 245068 330556 245074 330568
rect 305730 330556 305736 330568
rect 305788 330556 305794 330608
rect 36538 330488 36544 330540
rect 36596 330528 36602 330540
rect 49602 330528 49608 330540
rect 36596 330500 49608 330528
rect 36596 330488 36602 330500
rect 49602 330488 49608 330500
rect 49660 330488 49666 330540
rect 195330 330488 195336 330540
rect 195388 330528 195394 330540
rect 266446 330528 266452 330540
rect 195388 330500 266452 330528
rect 195388 330488 195394 330500
rect 266446 330488 266452 330500
rect 266504 330488 266510 330540
rect 7558 329808 7564 329860
rect 7616 329848 7622 329860
rect 125594 329848 125600 329860
rect 7616 329820 125600 329848
rect 7616 329808 7622 329820
rect 125594 329808 125600 329820
rect 125652 329808 125658 329860
rect 155862 329808 155868 329860
rect 155920 329848 155926 329860
rect 167638 329848 167644 329860
rect 155920 329820 167644 329848
rect 155920 329808 155926 329820
rect 167638 329808 167644 329820
rect 167696 329808 167702 329860
rect 149238 329740 149244 329792
rect 149296 329780 149302 329792
rect 155954 329780 155960 329792
rect 149296 329752 155960 329780
rect 149296 329740 149302 329752
rect 155954 329740 155960 329752
rect 156012 329740 156018 329792
rect 156046 329740 156052 329792
rect 156104 329780 156110 329792
rect 159450 329780 159456 329792
rect 156104 329752 159456 329780
rect 156104 329740 156110 329752
rect 159450 329740 159456 329752
rect 159508 329740 159514 329792
rect 169202 329740 169208 329792
rect 169260 329780 169266 329792
rect 172606 329780 172612 329792
rect 169260 329752 172612 329780
rect 169260 329740 169266 329752
rect 172606 329740 172612 329752
rect 172664 329740 172670 329792
rect 173250 329740 173256 329792
rect 173308 329780 173314 329792
rect 175274 329780 175280 329792
rect 173308 329752 175280 329780
rect 173308 329740 173314 329752
rect 175274 329740 175280 329752
rect 175332 329740 175338 329792
rect 194042 329740 194048 329792
rect 194100 329780 194106 329792
rect 259546 329780 259552 329792
rect 194100 329752 259552 329780
rect 194100 329740 194106 329752
rect 259546 329740 259552 329752
rect 259604 329780 259610 329792
rect 374086 329780 374092 329792
rect 259604 329752 374092 329780
rect 259604 329740 259610 329752
rect 374086 329740 374092 329752
rect 374144 329740 374150 329792
rect 114646 329672 114652 329724
rect 114704 329712 114710 329724
rect 115704 329712 115710 329724
rect 114704 329684 115710 329712
rect 114704 329672 114710 329684
rect 115704 329672 115710 329684
rect 115762 329672 115768 329724
rect 150434 329672 150440 329724
rect 150492 329712 150498 329724
rect 156690 329712 156696 329724
rect 150492 329684 156696 329712
rect 150492 329672 150498 329684
rect 156690 329672 156696 329684
rect 156748 329672 156754 329724
rect 69382 329536 69388 329588
rect 69440 329576 69446 329588
rect 76558 329576 76564 329588
rect 69440 329548 76564 329576
rect 69440 329536 69446 329548
rect 76558 329536 76564 329548
rect 76616 329536 76622 329588
rect 158898 329128 158904 329180
rect 158956 329168 158962 329180
rect 166442 329168 166448 329180
rect 158956 329140 166448 329168
rect 158956 329128 158962 329140
rect 166442 329128 166448 329140
rect 166500 329128 166506 329180
rect 176194 329128 176200 329180
rect 176252 329168 176258 329180
rect 184474 329168 184480 329180
rect 176252 329140 184480 329168
rect 176252 329128 176258 329140
rect 184474 329128 184480 329140
rect 184532 329128 184538 329180
rect 115382 329100 115388 329112
rect 103486 329072 115388 329100
rect 11698 328448 11704 328500
rect 11756 328488 11762 328500
rect 103486 328488 103514 329072
rect 115382 329060 115388 329072
rect 115440 329060 115446 329112
rect 124306 329060 124312 329112
rect 124364 329060 124370 329112
rect 139302 329060 139308 329112
rect 139360 329100 139366 329112
rect 139360 329072 151814 329100
rect 139360 329060 139366 329072
rect 11756 328460 103514 328488
rect 11756 328448 11762 328460
rect 124324 328420 124352 329060
rect 103486 328392 124352 328420
rect 22738 327700 22744 327752
rect 22796 327740 22802 327752
rect 103486 327740 103514 328392
rect 151786 328284 151814 329072
rect 152642 329060 152648 329112
rect 152700 329060 152706 329112
rect 156322 329060 156328 329112
rect 156380 329100 156386 329112
rect 156380 329072 156736 329100
rect 156380 329060 156386 329072
rect 152660 328352 152688 329060
rect 156708 328840 156736 329072
rect 165154 329060 165160 329112
rect 165212 329100 165218 329112
rect 235258 329100 235264 329112
rect 165212 329072 235264 329100
rect 165212 329060 165218 329072
rect 235258 329060 235264 329072
rect 235316 329060 235322 329112
rect 374730 329060 374736 329112
rect 374788 329100 374794 329112
rect 409874 329100 409880 329112
rect 374788 329072 409880 329100
rect 374788 329060 374794 329072
rect 409874 329060 409880 329072
rect 409932 329060 409938 329112
rect 156690 328788 156696 328840
rect 156748 328788 156754 328840
rect 156874 328448 156880 328500
rect 156932 328488 156938 328500
rect 165154 328488 165160 328500
rect 156932 328460 165160 328488
rect 156932 328448 156938 328460
rect 165154 328448 165160 328460
rect 165212 328448 165218 328500
rect 266446 328380 266452 328432
rect 266504 328420 266510 328432
rect 267642 328420 267648 328432
rect 266504 328392 267648 328420
rect 266504 328380 266510 328392
rect 267642 328380 267648 328392
rect 267700 328420 267706 328432
rect 349154 328420 349160 328432
rect 267700 328392 349160 328420
rect 267700 328380 267706 328392
rect 349154 328380 349160 328392
rect 349212 328380 349218 328432
rect 156874 328352 156880 328364
rect 152660 328324 156880 328352
rect 156874 328312 156880 328324
rect 156932 328312 156938 328364
rect 156782 328284 156788 328296
rect 151786 328256 156788 328284
rect 156782 328244 156788 328256
rect 156840 328244 156846 328296
rect 158898 327836 158904 327888
rect 158956 327876 158962 327888
rect 161474 327876 161480 327888
rect 158956 327848 161480 327876
rect 158956 327836 158962 327848
rect 161474 327836 161480 327848
rect 161532 327836 161538 327888
rect 189810 327768 189816 327820
rect 189868 327808 189874 327820
rect 211890 327808 211896 327820
rect 189868 327780 211896 327808
rect 189868 327768 189874 327780
rect 211890 327768 211896 327780
rect 211948 327768 211954 327820
rect 22796 327712 103514 327740
rect 22796 327700 22802 327712
rect 168098 327700 168104 327752
rect 168156 327740 168162 327752
rect 195974 327740 195980 327752
rect 168156 327712 195980 327740
rect 168156 327700 168162 327712
rect 195974 327700 195980 327712
rect 196032 327700 196038 327752
rect 239122 327700 239128 327752
rect 239180 327740 239186 327752
rect 259362 327740 259368 327752
rect 239180 327712 259368 327740
rect 239180 327700 239186 327712
rect 259362 327700 259368 327712
rect 259420 327700 259426 327752
rect 156966 327292 156972 327344
rect 157024 327332 157030 327344
rect 161474 327332 161480 327344
rect 157024 327304 161480 327332
rect 157024 327292 157030 327304
rect 161474 327292 161480 327304
rect 161532 327292 161538 327344
rect 216030 327088 216036 327140
rect 216088 327128 216094 327140
rect 275278 327128 275284 327140
rect 216088 327100 275284 327128
rect 216088 327088 216094 327100
rect 275278 327088 275284 327100
rect 275336 327088 275342 327140
rect 259362 327020 259368 327072
rect 259420 327060 259426 327072
rect 358078 327060 358084 327072
rect 259420 327032 358084 327060
rect 259420 327020 259426 327032
rect 358078 327020 358084 327032
rect 358136 327020 358142 327072
rect 199654 326408 199660 326460
rect 199712 326448 199718 326460
rect 221458 326448 221464 326460
rect 199712 326420 221464 326448
rect 199712 326408 199718 326420
rect 221458 326408 221464 326420
rect 221516 326408 221522 326460
rect 165614 326340 165620 326392
rect 165672 326380 165678 326392
rect 201586 326380 201592 326392
rect 165672 326352 201592 326380
rect 165672 326340 165678 326352
rect 201586 326340 201592 326352
rect 201644 326340 201650 326392
rect 207750 326340 207756 326392
rect 207808 326380 207814 326392
rect 212626 326380 212632 326392
rect 207808 326352 212632 326380
rect 207808 326340 207814 326352
rect 212626 326340 212632 326352
rect 212684 326340 212690 326392
rect 214650 326340 214656 326392
rect 214708 326380 214714 326392
rect 255406 326380 255412 326392
rect 214708 326352 255412 326380
rect 214708 326340 214714 326352
rect 255406 326340 255412 326352
rect 255464 326340 255470 326392
rect 326982 326340 326988 326392
rect 327040 326380 327046 326392
rect 348418 326380 348424 326392
rect 327040 326352 348424 326380
rect 327040 326340 327046 326352
rect 348418 326340 348424 326352
rect 348476 326340 348482 326392
rect 55122 325660 55128 325712
rect 55180 325700 55186 325712
rect 66898 325700 66904 325712
rect 55180 325672 66904 325700
rect 55180 325660 55186 325672
rect 66898 325660 66904 325672
rect 66956 325660 66962 325712
rect 158898 325660 158904 325712
rect 158956 325700 158962 325712
rect 191374 325700 191380 325712
rect 158956 325672 191380 325700
rect 158956 325660 158962 325672
rect 191374 325660 191380 325672
rect 191432 325660 191438 325712
rect 238662 325660 238668 325712
rect 238720 325700 238726 325712
rect 325694 325700 325700 325712
rect 238720 325672 325700 325700
rect 238720 325660 238726 325672
rect 325694 325660 325700 325672
rect 325752 325700 325758 325712
rect 326982 325700 326988 325712
rect 325752 325672 326988 325700
rect 325752 325660 325758 325672
rect 326982 325660 326988 325672
rect 327040 325660 327046 325712
rect 158254 325388 158260 325440
rect 158312 325428 158318 325440
rect 163590 325428 163596 325440
rect 158312 325400 163596 325428
rect 158312 325388 158318 325400
rect 163590 325388 163596 325400
rect 163648 325388 163654 325440
rect 188522 325048 188528 325100
rect 188580 325088 188586 325100
rect 206554 325088 206560 325100
rect 188580 325060 206560 325088
rect 188580 325048 188586 325060
rect 206554 325048 206560 325060
rect 206612 325048 206618 325100
rect 196618 324980 196624 325032
rect 196676 325020 196682 325032
rect 228450 325020 228456 325032
rect 196676 324992 228456 325020
rect 196676 324980 196682 324992
rect 228450 324980 228456 324992
rect 228508 324980 228514 325032
rect 161474 324912 161480 324964
rect 161532 324952 161538 324964
rect 195146 324952 195152 324964
rect 161532 324924 195152 324952
rect 161532 324912 161538 324924
rect 195146 324912 195152 324924
rect 195204 324912 195210 324964
rect 214558 324912 214564 324964
rect 214616 324952 214622 324964
rect 341518 324952 341524 324964
rect 214616 324924 341524 324952
rect 214616 324912 214622 324924
rect 341518 324912 341524 324924
rect 341576 324912 341582 324964
rect 162946 324844 162952 324896
rect 163004 324884 163010 324896
rect 165062 324884 165068 324896
rect 163004 324856 165068 324884
rect 163004 324844 163010 324856
rect 165062 324844 165068 324856
rect 165120 324844 165126 324896
rect 158898 324164 158904 324216
rect 158956 324204 158962 324216
rect 160738 324204 160744 324216
rect 158956 324176 160744 324204
rect 158956 324164 158962 324176
rect 160738 324164 160744 324176
rect 160796 324164 160802 324216
rect 187050 323552 187056 323604
rect 187108 323592 187114 323604
rect 220078 323592 220084 323604
rect 187108 323564 220084 323592
rect 187108 323552 187114 323564
rect 220078 323552 220084 323564
rect 220136 323552 220142 323604
rect 254578 323552 254584 323604
rect 254636 323592 254642 323604
rect 282270 323592 282276 323604
rect 254636 323564 282276 323592
rect 254636 323552 254642 323564
rect 282270 323552 282276 323564
rect 282328 323552 282334 323604
rect 330294 323552 330300 323604
rect 330352 323592 330358 323604
rect 351178 323592 351184 323604
rect 330352 323564 351184 323592
rect 330352 323552 330358 323564
rect 351178 323552 351184 323564
rect 351236 323552 351242 323604
rect 158714 323008 158720 323060
rect 158772 323048 158778 323060
rect 243630 323048 243636 323060
rect 158772 323020 243636 323048
rect 158772 323008 158778 323020
rect 243630 323008 243636 323020
rect 243688 323008 243694 323060
rect 236638 322940 236644 322992
rect 236696 322980 236702 322992
rect 237282 322980 237288 322992
rect 236696 322952 237288 322980
rect 236696 322940 236702 322952
rect 237282 322940 237288 322952
rect 237340 322980 237346 322992
rect 329834 322980 329840 322992
rect 237340 322952 329840 322980
rect 237340 322940 237346 322952
rect 329834 322940 329840 322952
rect 329892 322980 329898 322992
rect 330294 322980 330300 322992
rect 329892 322952 330300 322980
rect 329892 322940 329898 322952
rect 330294 322940 330300 322952
rect 330352 322940 330358 322992
rect 191282 322260 191288 322312
rect 191340 322300 191346 322312
rect 220170 322300 220176 322312
rect 191340 322272 220176 322300
rect 191340 322260 191346 322272
rect 220170 322260 220176 322272
rect 220228 322260 220234 322312
rect 195146 322192 195152 322244
rect 195204 322232 195210 322244
rect 234062 322232 234068 322244
rect 195204 322204 234068 322232
rect 195204 322192 195210 322204
rect 234062 322192 234068 322204
rect 234120 322192 234126 322244
rect 289722 322192 289728 322244
rect 289780 322232 289786 322244
rect 313274 322232 313280 322244
rect 289780 322204 313280 322232
rect 289780 322192 289786 322204
rect 313274 322192 313280 322204
rect 313332 322192 313338 322244
rect 158714 321580 158720 321632
rect 158772 321620 158778 321632
rect 166350 321620 166356 321632
rect 158772 321592 166356 321620
rect 158772 321580 158778 321592
rect 166350 321580 166356 321592
rect 166408 321580 166414 321632
rect 233970 321580 233976 321632
rect 234028 321620 234034 321632
rect 259454 321620 259460 321632
rect 234028 321592 259460 321620
rect 234028 321580 234034 321592
rect 259454 321580 259460 321592
rect 259512 321620 259518 321632
rect 260098 321620 260104 321632
rect 259512 321592 260104 321620
rect 259512 321580 259518 321592
rect 260098 321580 260104 321592
rect 260156 321580 260162 321632
rect 4798 321512 4804 321564
rect 4856 321552 4862 321564
rect 66898 321552 66904 321564
rect 4856 321524 66904 321552
rect 4856 321512 4862 321524
rect 66898 321512 66904 321524
rect 66956 321512 66962 321564
rect 184198 320900 184204 320952
rect 184256 320940 184262 320952
rect 232590 320940 232596 320952
rect 184256 320912 232596 320940
rect 184256 320900 184262 320912
rect 232590 320900 232596 320912
rect 232648 320900 232654 320952
rect 166442 320832 166448 320884
rect 166500 320872 166506 320884
rect 196618 320872 196624 320884
rect 166500 320844 196624 320872
rect 166500 320832 166506 320844
rect 196618 320832 196624 320844
rect 196676 320832 196682 320884
rect 214558 320832 214564 320884
rect 214616 320872 214622 320884
rect 277394 320872 277400 320884
rect 214616 320844 277400 320872
rect 214616 320832 214622 320844
rect 277394 320832 277400 320844
rect 277452 320832 277458 320884
rect 285766 320832 285772 320884
rect 285824 320872 285830 320884
rect 286962 320872 286968 320884
rect 285824 320844 286968 320872
rect 285824 320832 285830 320844
rect 286962 320832 286968 320844
rect 287020 320872 287026 320884
rect 360194 320872 360200 320884
rect 287020 320844 360200 320872
rect 287020 320832 287026 320844
rect 360194 320832 360200 320844
rect 360252 320832 360258 320884
rect 52362 320152 52368 320204
rect 52420 320192 52426 320204
rect 66806 320192 66812 320204
rect 52420 320164 66812 320192
rect 52420 320152 52426 320164
rect 66806 320152 66812 320164
rect 66864 320152 66870 320204
rect 158714 320152 158720 320204
rect 158772 320192 158778 320204
rect 164970 320192 164976 320204
rect 158772 320164 164976 320192
rect 158772 320152 158778 320164
rect 164970 320152 164976 320164
rect 165028 320152 165034 320204
rect 241974 320152 241980 320204
rect 242032 320192 242038 320204
rect 285766 320192 285772 320204
rect 242032 320164 285772 320192
rect 242032 320152 242038 320164
rect 285766 320152 285772 320164
rect 285824 320152 285830 320204
rect 176010 319472 176016 319524
rect 176068 319512 176074 319524
rect 209130 319512 209136 319524
rect 176068 319484 209136 319512
rect 176068 319472 176074 319484
rect 209130 319472 209136 319484
rect 209188 319472 209194 319524
rect 245102 319472 245108 319524
rect 245160 319512 245166 319524
rect 255314 319512 255320 319524
rect 245160 319484 255320 319512
rect 245160 319472 245166 319484
rect 255314 319472 255320 319484
rect 255372 319472 255378 319524
rect 53650 319404 53656 319456
rect 53708 319444 53714 319456
rect 66990 319444 66996 319456
rect 53708 319416 66996 319444
rect 53708 319404 53714 319416
rect 66990 319404 66996 319416
rect 67048 319444 67054 319456
rect 67266 319444 67272 319456
rect 67048 319416 67272 319444
rect 67048 319404 67054 319416
rect 67266 319404 67272 319416
rect 67324 319404 67330 319456
rect 158714 319404 158720 319456
rect 158772 319444 158778 319456
rect 166994 319444 167000 319456
rect 158772 319416 167000 319444
rect 158772 319404 158778 319416
rect 166994 319404 167000 319416
rect 167052 319404 167058 319456
rect 170582 319404 170588 319456
rect 170640 319444 170646 319456
rect 206278 319444 206284 319456
rect 170640 319416 206284 319444
rect 170640 319404 170646 319416
rect 206278 319404 206284 319416
rect 206336 319404 206342 319456
rect 253198 319404 253204 319456
rect 253256 319444 253262 319456
rect 264974 319444 264980 319456
rect 253256 319416 264980 319444
rect 253256 319404 253262 319416
rect 264974 319404 264980 319416
rect 265032 319404 265038 319456
rect 4062 318724 4068 318776
rect 4120 318764 4126 318776
rect 39298 318764 39304 318776
rect 4120 318736 39304 318764
rect 4120 318724 4126 318736
rect 39298 318724 39304 318736
rect 39356 318724 39362 318776
rect 63218 318520 63224 318572
rect 63276 318560 63282 318572
rect 66806 318560 66812 318572
rect 63276 318532 66812 318560
rect 63276 318520 63282 318532
rect 66806 318520 66812 318532
rect 66864 318520 66870 318572
rect 252462 318044 252468 318096
rect 252520 318084 252526 318096
rect 342254 318084 342260 318096
rect 252520 318056 342260 318084
rect 252520 318044 252526 318056
rect 342254 318044 342260 318056
rect 342312 318044 342318 318096
rect 169662 317500 169668 317552
rect 169720 317540 169726 317552
rect 173158 317540 173164 317552
rect 169720 317512 173164 317540
rect 169720 317500 169726 317512
rect 173158 317500 173164 317512
rect 173216 317500 173222 317552
rect 205910 317500 205916 317552
rect 205968 317540 205974 317552
rect 259454 317540 259460 317552
rect 205968 317512 259460 317540
rect 205968 317500 205974 317512
rect 259454 317500 259460 317512
rect 259512 317500 259518 317552
rect 61930 317432 61936 317484
rect 61988 317472 61994 317484
rect 66714 317472 66720 317484
rect 61988 317444 66720 317472
rect 61988 317432 61994 317444
rect 66714 317432 66720 317444
rect 66772 317432 66778 317484
rect 158714 317432 158720 317484
rect 158772 317472 158778 317484
rect 240962 317472 240968 317484
rect 158772 317444 240968 317472
rect 158772 317432 158778 317444
rect 240962 317432 240968 317444
rect 241020 317432 241026 317484
rect 158806 317364 158812 317416
rect 158864 317404 158870 317416
rect 166442 317404 166448 317416
rect 158864 317376 166448 317404
rect 158864 317364 158870 317376
rect 166442 317364 166448 317376
rect 166500 317404 166506 317416
rect 166718 317404 166724 317416
rect 166500 317376 166724 317404
rect 166500 317364 166506 317376
rect 166718 317364 166724 317376
rect 166776 317364 166782 317416
rect 351914 316752 351920 316804
rect 351972 316792 351978 316804
rect 352558 316792 352564 316804
rect 351972 316764 352564 316792
rect 351972 316752 351978 316764
rect 352558 316752 352564 316764
rect 352616 316752 352622 316804
rect 29638 316684 29644 316736
rect 29696 316724 29702 316736
rect 64506 316724 64512 316736
rect 29696 316696 64512 316724
rect 29696 316684 29702 316696
rect 64506 316684 64512 316696
rect 64564 316724 64570 316736
rect 66806 316724 66812 316736
rect 64564 316696 66812 316724
rect 64564 316684 64570 316696
rect 66806 316684 66812 316696
rect 66864 316684 66870 316736
rect 166442 316684 166448 316736
rect 166500 316724 166506 316736
rect 184290 316724 184296 316736
rect 166500 316696 184296 316724
rect 166500 316684 166506 316696
rect 184290 316684 184296 316696
rect 184348 316684 184354 316736
rect 211062 316684 211068 316736
rect 211120 316724 211126 316736
rect 240870 316724 240876 316736
rect 211120 316696 240876 316724
rect 211120 316684 211126 316696
rect 240870 316684 240876 316696
rect 240928 316684 240934 316736
rect 320174 316684 320180 316736
rect 320232 316724 320238 316736
rect 360286 316724 360292 316736
rect 320232 316696 360292 316724
rect 320232 316684 320238 316696
rect 360286 316684 360292 316696
rect 360344 316684 360350 316736
rect 245654 316072 245660 316124
rect 245712 316112 245718 316124
rect 320174 316112 320180 316124
rect 245712 316084 320180 316112
rect 245712 316072 245718 316084
rect 320174 316072 320180 316084
rect 320232 316072 320238 316124
rect 61930 316004 61936 316056
rect 61988 316044 61994 316056
rect 65518 316044 65524 316056
rect 61988 316016 65524 316044
rect 61988 316004 61994 316016
rect 65518 316004 65524 316016
rect 65576 316044 65582 316056
rect 65576 316016 66208 316044
rect 65576 316004 65582 316016
rect 66180 315976 66208 316016
rect 188430 316004 188436 316056
rect 188488 316044 188494 316056
rect 209958 316044 209964 316056
rect 188488 316016 209964 316044
rect 188488 316004 188494 316016
rect 209958 316004 209964 316016
rect 210016 316044 210022 316056
rect 211062 316044 211068 316056
rect 210016 316016 211068 316044
rect 210016 316004 210022 316016
rect 211062 316004 211068 316016
rect 211120 316004 211126 316056
rect 223022 316004 223028 316056
rect 223080 316044 223086 316056
rect 352558 316044 352564 316056
rect 223080 316016 352564 316044
rect 223080 316004 223086 316016
rect 352558 316004 352564 316016
rect 352616 316004 352622 316056
rect 66622 315976 66628 315988
rect 66180 315948 66628 315976
rect 66622 315936 66628 315948
rect 66680 315936 66686 315988
rect 209038 315256 209044 315308
rect 209096 315296 209102 315308
rect 215846 315296 215852 315308
rect 209096 315268 215852 315296
rect 209096 315256 209102 315268
rect 215846 315256 215852 315268
rect 215904 315256 215910 315308
rect 63310 314916 63316 314968
rect 63368 314956 63374 314968
rect 66162 314956 66168 314968
rect 63368 314928 66168 314956
rect 63368 314916 63374 314928
rect 66162 314916 66168 314928
rect 66220 314956 66226 314968
rect 66530 314956 66536 314968
rect 66220 314928 66536 314956
rect 66220 314916 66226 314928
rect 66530 314916 66536 314928
rect 66588 314916 66594 314968
rect 158714 314712 158720 314764
rect 158772 314752 158778 314764
rect 175090 314752 175096 314764
rect 158772 314724 175096 314752
rect 158772 314712 158778 314724
rect 175090 314712 175096 314724
rect 175148 314752 175154 314764
rect 178678 314752 178684 314764
rect 175148 314724 178684 314752
rect 175148 314712 175154 314724
rect 178678 314712 178684 314724
rect 178736 314712 178742 314764
rect 164142 314644 164148 314696
rect 164200 314684 164206 314696
rect 262306 314684 262312 314696
rect 164200 314656 262312 314684
rect 164200 314644 164206 314656
rect 262306 314644 262312 314656
rect 262364 314644 262370 314696
rect 60458 314576 60464 314628
rect 60516 314616 60522 314628
rect 66898 314616 66904 314628
rect 60516 314588 66904 314616
rect 60516 314576 60522 314588
rect 66898 314576 66904 314588
rect 66956 314576 66962 314628
rect 158714 314576 158720 314628
rect 158772 314616 158778 314628
rect 164160 314616 164188 314644
rect 158772 314588 164188 314616
rect 158772 314576 158778 314588
rect 178678 313896 178684 313948
rect 178736 313936 178742 313948
rect 188430 313936 188436 313948
rect 178736 313908 188436 313936
rect 178736 313896 178742 313908
rect 188430 313896 188436 313908
rect 188488 313896 188494 313948
rect 195422 313896 195428 313948
rect 195480 313936 195486 313948
rect 212902 313936 212908 313948
rect 195480 313908 212908 313936
rect 195480 313896 195486 313908
rect 212902 313896 212908 313908
rect 212960 313896 212966 313948
rect 217318 313896 217324 313948
rect 217376 313936 217382 313948
rect 235994 313936 236000 313948
rect 217376 313908 236000 313936
rect 217376 313896 217382 313908
rect 235994 313896 236000 313908
rect 236052 313896 236058 313948
rect 238018 313896 238024 313948
rect 238076 313936 238082 313948
rect 251266 313936 251272 313948
rect 238076 313908 251272 313936
rect 238076 313896 238082 313908
rect 251266 313896 251272 313908
rect 251324 313896 251330 313948
rect 158714 313284 158720 313336
rect 158772 313324 158778 313336
rect 180150 313324 180156 313336
rect 158772 313296 180156 313324
rect 158772 313284 158778 313296
rect 180150 313284 180156 313296
rect 180208 313284 180214 313336
rect 226242 313284 226248 313336
rect 226300 313324 226306 313336
rect 269206 313324 269212 313336
rect 226300 313296 269212 313324
rect 226300 313284 226306 313296
rect 269206 313284 269212 313296
rect 269264 313284 269270 313336
rect 54938 313216 54944 313268
rect 54996 313256 55002 313268
rect 66898 313256 66904 313268
rect 54996 313228 66904 313256
rect 54996 313216 55002 313228
rect 66898 313216 66904 313228
rect 66956 313216 66962 313268
rect 191098 312672 191104 312724
rect 191156 312712 191162 312724
rect 221642 312712 221648 312724
rect 191156 312684 221648 312712
rect 191156 312672 191162 312684
rect 221642 312672 221648 312684
rect 221700 312672 221706 312724
rect 188522 312536 188528 312588
rect 188580 312576 188586 312588
rect 205910 312576 205916 312588
rect 188580 312548 205916 312576
rect 188580 312536 188586 312548
rect 205910 312536 205916 312548
rect 205968 312536 205974 312588
rect 221550 312536 221556 312588
rect 221608 312576 221614 312588
rect 252830 312576 252836 312588
rect 221608 312548 252836 312576
rect 221608 312536 221614 312548
rect 252830 312536 252836 312548
rect 252888 312536 252894 312588
rect 260098 312536 260104 312588
rect 260156 312576 260162 312588
rect 460934 312576 460940 312588
rect 260156 312548 460940 312576
rect 260156 312536 260162 312548
rect 460934 312536 460940 312548
rect 460992 312536 460998 312588
rect 212902 311856 212908 311908
rect 212960 311896 212966 311908
rect 327718 311896 327724 311908
rect 212960 311868 327724 311896
rect 212960 311856 212966 311868
rect 327718 311856 327724 311868
rect 327776 311856 327782 311908
rect 164970 311788 164976 311840
rect 165028 311828 165034 311840
rect 245654 311828 245660 311840
rect 165028 311800 245660 311828
rect 165028 311788 165034 311800
rect 245654 311788 245660 311800
rect 245712 311788 245718 311840
rect 39942 311108 39948 311160
rect 40000 311148 40006 311160
rect 67082 311148 67088 311160
rect 40000 311120 67088 311148
rect 40000 311108 40006 311120
rect 67082 311108 67088 311120
rect 67140 311148 67146 311160
rect 67450 311148 67456 311160
rect 67140 311120 67456 311148
rect 67140 311108 67146 311120
rect 67450 311108 67456 311120
rect 67508 311108 67514 311160
rect 246298 311108 246304 311160
rect 246356 311148 246362 311160
rect 256694 311148 256700 311160
rect 246356 311120 256700 311148
rect 246356 311108 246362 311120
rect 256694 311108 256700 311120
rect 256752 311108 256758 311160
rect 4798 310496 4804 310548
rect 4856 310536 4862 310548
rect 39942 310536 39948 310548
rect 4856 310508 39948 310536
rect 4856 310496 4862 310508
rect 39942 310496 39948 310508
rect 40000 310496 40006 310548
rect 206554 310496 206560 310548
rect 206612 310536 206618 310548
rect 206830 310536 206836 310548
rect 206612 310508 206836 310536
rect 206612 310496 206618 310508
rect 206830 310496 206836 310508
rect 206888 310536 206894 310548
rect 276750 310536 276756 310548
rect 206888 310508 276756 310536
rect 206888 310496 206894 310508
rect 276750 310496 276756 310508
rect 276808 310496 276814 310548
rect 292574 310224 292580 310276
rect 292632 310264 292638 310276
rect 293218 310264 293224 310276
rect 292632 310236 293224 310264
rect 292632 310224 292638 310236
rect 293218 310224 293224 310236
rect 293276 310224 293282 310276
rect 193030 309884 193036 309936
rect 193088 309924 193094 309936
rect 216122 309924 216128 309936
rect 193088 309896 216128 309924
rect 193088 309884 193094 309896
rect 216122 309884 216128 309896
rect 216180 309884 216186 309936
rect 196710 309816 196716 309868
rect 196768 309856 196774 309868
rect 239030 309856 239036 309868
rect 196768 309828 239036 309856
rect 196768 309816 196774 309828
rect 239030 309816 239036 309828
rect 239088 309856 239094 309868
rect 240042 309856 240048 309868
rect 239088 309828 240048 309856
rect 239088 309816 239094 309828
rect 240042 309816 240048 309828
rect 240100 309816 240106 309868
rect 32398 309748 32404 309800
rect 32456 309788 32462 309800
rect 61746 309788 61752 309800
rect 32456 309760 61752 309788
rect 32456 309748 32462 309760
rect 61746 309748 61752 309760
rect 61804 309788 61810 309800
rect 66898 309788 66904 309800
rect 61804 309760 66904 309788
rect 61804 309748 61810 309760
rect 66898 309748 66904 309760
rect 66956 309748 66962 309800
rect 177298 309748 177304 309800
rect 177356 309788 177362 309800
rect 188338 309788 188344 309800
rect 177356 309760 188344 309788
rect 177356 309748 177362 309760
rect 188338 309748 188344 309760
rect 188396 309748 188402 309800
rect 216030 309748 216036 309800
rect 216088 309788 216094 309800
rect 292574 309788 292580 309800
rect 216088 309760 292580 309788
rect 216088 309748 216094 309760
rect 292574 309748 292580 309760
rect 292632 309748 292638 309800
rect 240042 309136 240048 309188
rect 240100 309176 240106 309188
rect 358078 309176 358084 309188
rect 240100 309148 358084 309176
rect 240100 309136 240106 309148
rect 358078 309136 358084 309148
rect 358136 309136 358142 309188
rect 192570 309068 192576 309120
rect 192628 309108 192634 309120
rect 226242 309108 226248 309120
rect 192628 309080 226248 309108
rect 192628 309068 192634 309080
rect 226242 309068 226248 309080
rect 226300 309108 226306 309120
rect 226886 309108 226892 309120
rect 226300 309080 226892 309108
rect 226300 309068 226306 309080
rect 226886 309068 226892 309080
rect 226944 309068 226950 309120
rect 228358 308388 228364 308440
rect 228416 308428 228422 308440
rect 244274 308428 244280 308440
rect 228416 308400 244280 308428
rect 228416 308388 228422 308400
rect 244274 308388 244280 308400
rect 244332 308388 244338 308440
rect 63310 307776 63316 307828
rect 63368 307816 63374 307828
rect 67818 307816 67824 307828
rect 63368 307788 67824 307816
rect 63368 307776 63374 307788
rect 67818 307776 67824 307788
rect 67876 307776 67882 307828
rect 197998 307776 198004 307828
rect 198056 307816 198062 307828
rect 276658 307816 276664 307828
rect 198056 307788 276664 307816
rect 198056 307776 198062 307788
rect 276658 307776 276664 307788
rect 276716 307776 276722 307828
rect 64598 307708 64604 307760
rect 64656 307748 64662 307760
rect 66898 307748 66904 307760
rect 64656 307720 66904 307748
rect 64656 307708 64662 307720
rect 66898 307708 66904 307720
rect 66956 307708 66962 307760
rect 199562 307096 199568 307148
rect 199620 307136 199626 307148
rect 214558 307136 214564 307148
rect 199620 307108 214564 307136
rect 199620 307096 199626 307108
rect 214558 307096 214564 307108
rect 214616 307096 214622 307148
rect 170398 307028 170404 307080
rect 170456 307068 170462 307080
rect 187602 307068 187608 307080
rect 170456 307040 187608 307068
rect 170456 307028 170462 307040
rect 187602 307028 187608 307040
rect 187660 307028 187666 307080
rect 200022 307028 200028 307080
rect 200080 307068 200086 307080
rect 240778 307068 240784 307080
rect 200080 307040 240784 307068
rect 200080 307028 200086 307040
rect 240778 307028 240784 307040
rect 240836 307028 240842 307080
rect 298738 307028 298744 307080
rect 298796 307068 298802 307080
rect 345750 307068 345756 307080
rect 298796 307040 345756 307068
rect 298796 307028 298802 307040
rect 345750 307028 345756 307040
rect 345808 307028 345814 307080
rect 158714 306348 158720 306400
rect 158772 306388 158778 306400
rect 195330 306388 195336 306400
rect 158772 306360 195336 306388
rect 158772 306348 158778 306360
rect 195330 306348 195336 306360
rect 195388 306348 195394 306400
rect 215846 306348 215852 306400
rect 215904 306388 215910 306400
rect 289814 306388 289820 306400
rect 215904 306360 289820 306388
rect 215904 306348 215910 306360
rect 289814 306348 289820 306360
rect 289872 306348 289878 306400
rect 3510 306280 3516 306332
rect 3568 306320 3574 306332
rect 36538 306320 36544 306332
rect 3568 306292 36544 306320
rect 3568 306280 3574 306292
rect 36538 306280 36544 306292
rect 36596 306280 36602 306332
rect 223022 306320 223028 306332
rect 209746 306292 223028 306320
rect 208394 306212 208400 306264
rect 208452 306252 208458 306264
rect 209746 306252 209774 306292
rect 223022 306280 223028 306292
rect 223080 306280 223086 306332
rect 208452 306224 209774 306252
rect 208452 306212 208458 306224
rect 223206 305056 223212 305108
rect 223264 305096 223270 305108
rect 360838 305096 360844 305108
rect 223264 305068 360844 305096
rect 223264 305056 223270 305068
rect 360838 305056 360844 305068
rect 360896 305056 360902 305108
rect 53558 304988 53564 305040
rect 53616 305028 53622 305040
rect 66898 305028 66904 305040
rect 53616 305000 66904 305028
rect 53616 304988 53622 305000
rect 66898 304988 66904 305000
rect 66956 304988 66962 305040
rect 158806 304988 158812 305040
rect 158864 305028 158870 305040
rect 194042 305028 194048 305040
rect 158864 305000 194048 305028
rect 158864 304988 158870 305000
rect 194042 304988 194048 305000
rect 194100 304988 194106 305040
rect 198550 304988 198556 305040
rect 198608 305028 198614 305040
rect 233142 305028 233148 305040
rect 198608 305000 233148 305028
rect 198608 304988 198614 305000
rect 233142 304988 233148 305000
rect 233200 304988 233206 305040
rect 233694 304988 233700 305040
rect 233752 305028 233758 305040
rect 234522 305028 234528 305040
rect 233752 305000 234528 305028
rect 233752 304988 233758 305000
rect 234522 304988 234528 305000
rect 234580 305028 234586 305040
rect 447134 305028 447140 305040
rect 234580 305000 447140 305028
rect 234580 304988 234586 305000
rect 447134 304988 447140 305000
rect 447192 304988 447198 305040
rect 63126 304920 63132 304972
rect 63184 304960 63190 304972
rect 66622 304960 66628 304972
rect 63184 304932 66628 304960
rect 63184 304920 63190 304932
rect 66622 304920 66628 304932
rect 66680 304920 66686 304972
rect 218054 304444 218060 304496
rect 218112 304484 218118 304496
rect 219342 304484 219348 304496
rect 218112 304456 219348 304484
rect 218112 304444 218118 304456
rect 219342 304444 219348 304456
rect 219400 304484 219406 304496
rect 221182 304484 221188 304496
rect 219400 304456 221188 304484
rect 219400 304444 219406 304456
rect 221182 304444 221188 304456
rect 221240 304444 221246 304496
rect 191282 304308 191288 304360
rect 191340 304348 191346 304360
rect 207750 304348 207756 304360
rect 191340 304320 207756 304348
rect 191340 304308 191346 304320
rect 207750 304308 207756 304320
rect 207808 304308 207814 304360
rect 222838 304308 222844 304360
rect 222896 304348 222902 304360
rect 234614 304348 234620 304360
rect 222896 304320 234620 304348
rect 222896 304308 222902 304320
rect 234614 304308 234620 304320
rect 234672 304308 234678 304360
rect 159450 304240 159456 304292
rect 159508 304280 159514 304292
rect 164970 304280 164976 304292
rect 159508 304252 164976 304280
rect 159508 304240 159514 304252
rect 164970 304240 164976 304252
rect 165028 304240 165034 304292
rect 183002 304240 183008 304292
rect 183060 304280 183066 304292
rect 195422 304280 195428 304292
rect 183060 304252 195428 304280
rect 183060 304240 183066 304252
rect 195422 304240 195428 304252
rect 195480 304240 195486 304292
rect 206278 304240 206284 304292
rect 206336 304280 206342 304292
rect 247126 304280 247132 304292
rect 206336 304252 247132 304280
rect 206336 304240 206342 304252
rect 247126 304240 247132 304252
rect 247184 304240 247190 304292
rect 234614 303628 234620 303680
rect 234672 303668 234678 303680
rect 435358 303668 435364 303680
rect 234672 303640 435364 303668
rect 234672 303628 234678 303640
rect 435358 303628 435364 303640
rect 435416 303628 435422 303680
rect 160094 302880 160100 302932
rect 160152 302920 160158 302932
rect 169202 302920 169208 302932
rect 160152 302892 169208 302920
rect 160152 302880 160158 302892
rect 169202 302880 169208 302892
rect 169260 302880 169266 302932
rect 247678 302880 247684 302932
rect 247736 302920 247742 302932
rect 251174 302920 251180 302932
rect 247736 302892 251180 302920
rect 247736 302880 247742 302892
rect 251174 302880 251180 302892
rect 251232 302880 251238 302932
rect 188430 302268 188436 302320
rect 188488 302308 188494 302320
rect 189074 302308 189080 302320
rect 188488 302280 189080 302308
rect 188488 302268 188494 302280
rect 189074 302268 189080 302280
rect 189132 302268 189138 302320
rect 159450 302200 159456 302252
rect 159508 302240 159514 302252
rect 258258 302240 258264 302252
rect 159508 302212 258264 302240
rect 159508 302200 159514 302212
rect 258258 302200 258264 302212
rect 258316 302200 258322 302252
rect 53466 302132 53472 302184
rect 53524 302172 53530 302184
rect 66714 302172 66720 302184
rect 53524 302144 66720 302172
rect 53524 302132 53530 302144
rect 66714 302132 66720 302144
rect 66772 302132 66778 302184
rect 158254 301452 158260 301504
rect 158312 301492 158318 301504
rect 188522 301492 188528 301504
rect 158312 301464 188528 301492
rect 158312 301452 158318 301464
rect 188522 301452 188528 301464
rect 188580 301452 188586 301504
rect 201402 301452 201408 301504
rect 201460 301492 201466 301504
rect 274174 301492 274180 301504
rect 201460 301464 274180 301492
rect 201460 301452 201466 301464
rect 274174 301452 274180 301464
rect 274232 301452 274238 301504
rect 60458 300840 60464 300892
rect 60516 300880 60522 300892
rect 66898 300880 66904 300892
rect 60516 300852 66904 300880
rect 60516 300840 60522 300852
rect 66898 300840 66904 300852
rect 66956 300840 66962 300892
rect 185762 300840 185768 300892
rect 185820 300880 185826 300892
rect 186222 300880 186228 300892
rect 185820 300852 186228 300880
rect 185820 300840 185826 300852
rect 186222 300840 186228 300852
rect 186280 300880 186286 300892
rect 214006 300880 214012 300892
rect 186280 300852 214012 300880
rect 186280 300840 186286 300852
rect 214006 300840 214012 300852
rect 214064 300840 214070 300892
rect 216030 300840 216036 300892
rect 216088 300880 216094 300892
rect 411898 300880 411904 300892
rect 216088 300852 411904 300880
rect 216088 300840 216094 300852
rect 411898 300840 411904 300852
rect 411956 300840 411962 300892
rect 244918 300772 244924 300824
rect 244976 300812 244982 300824
rect 247034 300812 247040 300824
rect 244976 300784 247040 300812
rect 244976 300772 244982 300784
rect 247034 300772 247040 300784
rect 247092 300772 247098 300824
rect 48130 300092 48136 300144
rect 48188 300132 48194 300144
rect 66990 300132 66996 300144
rect 48188 300104 66996 300132
rect 48188 300092 48194 300104
rect 66990 300092 66996 300104
rect 67048 300092 67054 300144
rect 189902 299548 189908 299600
rect 189960 299588 189966 299600
rect 244366 299588 244372 299600
rect 189960 299560 244372 299588
rect 189960 299548 189966 299560
rect 244366 299548 244372 299560
rect 244424 299548 244430 299600
rect 198642 299480 198648 299532
rect 198700 299520 198706 299532
rect 284938 299520 284944 299532
rect 198700 299492 284944 299520
rect 198700 299480 198706 299492
rect 284938 299480 284944 299492
rect 284996 299480 285002 299532
rect 204990 299412 204996 299464
rect 205048 299452 205054 299464
rect 223206 299452 223212 299464
rect 205048 299424 223212 299452
rect 205048 299412 205054 299424
rect 223206 299412 223212 299424
rect 223264 299412 223270 299464
rect 64690 298800 64696 298852
rect 64748 298840 64754 298852
rect 66898 298840 66904 298852
rect 64748 298812 66904 298840
rect 64748 298800 64754 298812
rect 66898 298800 66904 298812
rect 66956 298800 66962 298852
rect 188338 298800 188344 298852
rect 188396 298840 188402 298852
rect 201678 298840 201684 298852
rect 188396 298812 201684 298840
rect 188396 298800 188402 298812
rect 201678 298800 201684 298812
rect 201736 298800 201742 298852
rect 158714 298732 158720 298784
rect 158772 298772 158778 298784
rect 158772 298744 238754 298772
rect 158772 298732 158778 298744
rect 238726 298704 238754 298744
rect 244366 298732 244372 298784
rect 244424 298772 244430 298784
rect 265158 298772 265164 298784
rect 244424 298744 265164 298772
rect 244424 298732 244430 298744
rect 265158 298732 265164 298744
rect 265216 298732 265222 298784
rect 324314 298732 324320 298784
rect 324372 298772 324378 298784
rect 341610 298772 341616 298784
rect 324372 298744 341616 298772
rect 324372 298732 324378 298744
rect 341610 298732 341616 298744
rect 341668 298732 341674 298784
rect 244458 298704 244464 298716
rect 238726 298676 244464 298704
rect 244458 298664 244464 298676
rect 244516 298664 244522 298716
rect 228358 298188 228364 298240
rect 228416 298228 228422 298240
rect 279510 298228 279516 298240
rect 228416 298200 279516 298228
rect 228416 298188 228422 298200
rect 279510 298188 279516 298200
rect 279568 298188 279574 298240
rect 267090 298120 267096 298172
rect 267148 298160 267154 298172
rect 324314 298160 324320 298172
rect 267148 298132 324320 298160
rect 267148 298120 267154 298132
rect 324314 298120 324320 298132
rect 324372 298120 324378 298172
rect 41230 298052 41236 298104
rect 41288 298092 41294 298104
rect 66898 298092 66904 298104
rect 41288 298064 66904 298092
rect 41288 298052 41294 298064
rect 66898 298052 66904 298064
rect 66956 298052 66962 298104
rect 233142 297440 233148 297492
rect 233200 297480 233206 297492
rect 309134 297480 309140 297492
rect 233200 297452 309140 297480
rect 233200 297440 233206 297452
rect 309134 297440 309140 297452
rect 309192 297440 309198 297492
rect 158714 297372 158720 297424
rect 158772 297412 158778 297424
rect 175274 297412 175280 297424
rect 158772 297384 175280 297412
rect 158772 297372 158778 297384
rect 175274 297372 175280 297384
rect 175332 297372 175338 297424
rect 177942 297372 177948 297424
rect 178000 297412 178006 297424
rect 204254 297412 204260 297424
rect 178000 297384 204260 297412
rect 178000 297372 178006 297384
rect 204254 297372 204260 297384
rect 204312 297372 204318 297424
rect 209038 297372 209044 297424
rect 209096 297412 209102 297424
rect 215202 297412 215208 297424
rect 209096 297384 215208 297412
rect 209096 297372 209102 297384
rect 215202 297372 215208 297384
rect 215260 297412 215266 297424
rect 389910 297412 389916 297424
rect 215260 297384 389916 297412
rect 215260 297372 215266 297384
rect 389910 297372 389916 297384
rect 389968 297372 389974 297424
rect 175274 297168 175280 297220
rect 175332 297208 175338 297220
rect 176010 297208 176016 297220
rect 175332 297180 176016 297208
rect 175332 297168 175338 297180
rect 176010 297168 176016 297180
rect 176068 297168 176074 297220
rect 160002 296692 160008 296744
rect 160060 296732 160066 296744
rect 209038 296732 209044 296744
rect 160060 296704 209044 296732
rect 160060 296692 160066 296704
rect 209038 296692 209044 296704
rect 209096 296692 209102 296744
rect 191190 296012 191196 296064
rect 191248 296052 191254 296064
rect 206646 296052 206652 296064
rect 191248 296024 206652 296052
rect 191248 296012 191254 296024
rect 206646 296012 206652 296024
rect 206704 296052 206710 296064
rect 216030 296052 216036 296064
rect 206704 296024 216036 296052
rect 206704 296012 206710 296024
rect 216030 296012 216036 296024
rect 216088 296012 216094 296064
rect 194042 295944 194048 295996
rect 194100 295984 194106 295996
rect 236086 295984 236092 295996
rect 194100 295956 236092 295984
rect 194100 295944 194106 295956
rect 236086 295944 236092 295956
rect 236144 295944 236150 295996
rect 304258 295944 304264 295996
rect 304316 295984 304322 295996
rect 358814 295984 358820 295996
rect 304316 295956 358820 295984
rect 304316 295944 304322 295956
rect 358814 295944 358820 295956
rect 358872 295944 358878 295996
rect 242250 295876 242256 295928
rect 242308 295916 242314 295928
rect 243446 295916 243452 295928
rect 242308 295888 243452 295916
rect 242308 295876 242314 295888
rect 243446 295876 243452 295888
rect 243504 295876 243510 295928
rect 49602 295400 49608 295452
rect 49660 295440 49666 295452
rect 66898 295440 66904 295452
rect 49660 295412 66904 295440
rect 49660 295400 49666 295412
rect 66898 295400 66904 295412
rect 66956 295400 66962 295452
rect 243446 295400 243452 295452
rect 243504 295440 243510 295452
rect 303706 295440 303712 295452
rect 243504 295412 303712 295440
rect 243504 295400 243510 295412
rect 303706 295400 303712 295412
rect 303764 295440 303770 295452
rect 304258 295440 304264 295452
rect 303764 295412 304264 295440
rect 303764 295400 303770 295412
rect 304258 295400 304264 295412
rect 304316 295400 304322 295452
rect 17862 295332 17868 295384
rect 17920 295372 17926 295384
rect 67174 295372 67180 295384
rect 17920 295344 67180 295372
rect 17920 295332 17926 295344
rect 67174 295332 67180 295344
rect 67232 295332 67238 295384
rect 226978 295332 226984 295384
rect 227036 295372 227042 295384
rect 227622 295372 227628 295384
rect 227036 295344 227628 295372
rect 227036 295332 227042 295344
rect 227622 295332 227628 295344
rect 227680 295372 227686 295384
rect 308398 295372 308404 295384
rect 227680 295344 308404 295372
rect 227680 295332 227686 295344
rect 308398 295332 308404 295344
rect 308456 295332 308462 295384
rect 59078 295264 59084 295316
rect 59136 295304 59142 295316
rect 66254 295304 66260 295316
rect 59136 295276 66260 295304
rect 59136 295264 59142 295276
rect 66254 295264 66260 295276
rect 66312 295264 66318 295316
rect 158714 295264 158720 295316
rect 158772 295304 158778 295316
rect 187142 295304 187148 295316
rect 158772 295276 187148 295304
rect 158772 295264 158778 295276
rect 187142 295264 187148 295276
rect 187200 295264 187206 295316
rect 159542 294584 159548 294636
rect 159600 294624 159606 294636
rect 178034 294624 178040 294636
rect 159600 294596 178040 294624
rect 159600 294584 159606 294596
rect 178034 294584 178040 294596
rect 178092 294584 178098 294636
rect 295334 294584 295340 294636
rect 295392 294624 295398 294636
rect 382274 294624 382280 294636
rect 295392 294596 382280 294624
rect 295392 294584 295398 294596
rect 382274 294584 382280 294596
rect 382332 294584 382338 294636
rect 266998 294108 267004 294160
rect 267056 294148 267062 294160
rect 269114 294148 269120 294160
rect 267056 294120 269120 294148
rect 267056 294108 267062 294120
rect 269114 294108 269120 294120
rect 269172 294108 269178 294160
rect 222470 294040 222476 294092
rect 222528 294080 222534 294092
rect 222930 294080 222936 294092
rect 222528 294052 222936 294080
rect 222528 294040 222534 294052
rect 222930 294040 222936 294052
rect 222988 294080 222994 294092
rect 252554 294080 252560 294092
rect 222988 294052 252560 294080
rect 222988 294040 222994 294052
rect 252554 294040 252560 294052
rect 252612 294040 252618 294092
rect 187234 293972 187240 294024
rect 187292 294012 187298 294024
rect 262398 294012 262404 294024
rect 187292 293984 262404 294012
rect 187292 293972 187298 293984
rect 262398 293972 262404 293984
rect 262456 293972 262462 294024
rect 19242 293904 19248 293956
rect 19300 293944 19306 293956
rect 66898 293944 66904 293956
rect 19300 293916 66904 293944
rect 19300 293904 19306 293916
rect 66898 293904 66904 293916
rect 66956 293904 66962 293956
rect 194410 293224 194416 293276
rect 194468 293264 194474 293276
rect 204346 293264 204352 293276
rect 194468 293236 204352 293264
rect 194468 293224 194474 293236
rect 204346 293224 204352 293236
rect 204404 293224 204410 293276
rect 270402 293224 270408 293276
rect 270460 293264 270466 293276
rect 278130 293264 278136 293276
rect 270460 293236 278136 293264
rect 270460 293224 270466 293236
rect 278130 293224 278136 293236
rect 278188 293224 278194 293276
rect 315114 293224 315120 293276
rect 315172 293264 315178 293276
rect 362954 293264 362960 293276
rect 315172 293236 362960 293264
rect 315172 293224 315178 293236
rect 362954 293224 362960 293236
rect 363012 293224 363018 293276
rect 158714 292612 158720 292664
rect 158772 292652 158778 292664
rect 194042 292652 194048 292664
rect 158772 292624 194048 292652
rect 158772 292612 158778 292624
rect 194042 292612 194048 292624
rect 194100 292612 194106 292664
rect 204898 292612 204904 292664
rect 204956 292652 204962 292664
rect 262950 292652 262956 292664
rect 204956 292624 262956 292652
rect 204956 292612 204962 292624
rect 262950 292612 262956 292624
rect 263008 292612 263014 292664
rect 3510 292544 3516 292596
rect 3568 292584 3574 292596
rect 18598 292584 18604 292596
rect 3568 292556 18604 292584
rect 3568 292544 3574 292556
rect 18598 292544 18604 292556
rect 18656 292544 18662 292596
rect 158806 292544 158812 292596
rect 158864 292584 158870 292596
rect 220630 292584 220636 292596
rect 158864 292556 220636 292584
rect 158864 292544 158870 292556
rect 220630 292544 220636 292556
rect 220688 292544 220694 292596
rect 234246 292544 234252 292596
rect 234304 292584 234310 292596
rect 268378 292584 268384 292596
rect 234304 292556 268384 292584
rect 234304 292544 234310 292556
rect 268378 292544 268384 292556
rect 268436 292544 268442 292596
rect 60550 292476 60556 292528
rect 60608 292516 60614 292528
rect 66898 292516 66904 292528
rect 60608 292488 66904 292516
rect 60608 292476 60614 292488
rect 66898 292476 66904 292488
rect 66956 292476 66962 292528
rect 283558 291796 283564 291848
rect 283616 291836 283622 291848
rect 322198 291836 322204 291848
rect 283616 291808 322204 291836
rect 283616 291796 283622 291808
rect 322198 291796 322204 291808
rect 322256 291796 322262 291848
rect 389174 291796 389180 291848
rect 389232 291836 389238 291848
rect 407114 291836 407120 291848
rect 389232 291808 407120 291836
rect 389232 291796 389238 291808
rect 407114 291796 407120 291808
rect 407172 291796 407178 291848
rect 158714 291252 158720 291304
rect 158772 291292 158778 291304
rect 248690 291292 248696 291304
rect 158772 291264 248696 291292
rect 158772 291252 158778 291264
rect 248690 291252 248696 291264
rect 248748 291252 248754 291304
rect 174630 291184 174636 291236
rect 174688 291224 174694 291236
rect 204898 291224 204904 291236
rect 174688 291196 204904 291224
rect 174688 291184 174694 291196
rect 204898 291184 204904 291196
rect 204956 291184 204962 291236
rect 241422 291184 241428 291236
rect 241480 291224 241486 291236
rect 401594 291224 401600 291236
rect 241480 291196 401600 291224
rect 241480 291184 241486 291196
rect 401594 291184 401600 291196
rect 401652 291184 401658 291236
rect 52178 291116 52184 291168
rect 52236 291156 52242 291168
rect 56410 291156 56416 291168
rect 52236 291128 56416 291156
rect 52236 291116 52242 291128
rect 56410 291116 56416 291128
rect 56468 291116 56474 291168
rect 220078 291116 220084 291168
rect 220136 291156 220142 291168
rect 222102 291156 222108 291168
rect 220136 291128 222108 291156
rect 220136 291116 220142 291128
rect 222102 291116 222108 291128
rect 222160 291116 222166 291168
rect 166258 290436 166264 290488
rect 166316 290476 166322 290488
rect 211430 290476 211436 290488
rect 166316 290448 211436 290476
rect 166316 290436 166322 290448
rect 211430 290436 211436 290448
rect 211488 290436 211494 290488
rect 159266 290164 159272 290216
rect 159324 290204 159330 290216
rect 162210 290204 162216 290216
rect 159324 290176 162216 290204
rect 159324 290164 159330 290176
rect 162210 290164 162216 290176
rect 162268 290164 162274 290216
rect 224218 289960 224224 290012
rect 224276 290000 224282 290012
rect 445754 290000 445760 290012
rect 224276 289972 445760 290000
rect 224276 289960 224282 289972
rect 445754 289960 445760 289972
rect 445812 289960 445818 290012
rect 211430 289892 211436 289944
rect 211488 289932 211494 289944
rect 218054 289932 218060 289944
rect 211488 289904 218060 289932
rect 211488 289892 211494 289904
rect 218054 289892 218060 289904
rect 218112 289892 218118 289944
rect 222102 289892 222108 289944
rect 222160 289932 222166 289944
rect 254578 289932 254584 289944
rect 222160 289904 254584 289932
rect 222160 289892 222166 289904
rect 254578 289892 254584 289904
rect 254636 289892 254642 289944
rect 56410 289824 56416 289876
rect 56468 289864 56474 289876
rect 66898 289864 66904 289876
rect 56468 289836 66904 289864
rect 56468 289824 56474 289836
rect 66898 289824 66904 289836
rect 66956 289824 66962 289876
rect 158714 289824 158720 289876
rect 158772 289864 158778 289876
rect 224402 289864 224408 289876
rect 158772 289836 224408 289864
rect 158772 289824 158778 289836
rect 224402 289824 224408 289836
rect 224460 289824 224466 289876
rect 56318 289756 56324 289808
rect 56376 289796 56382 289808
rect 66622 289796 66628 289808
rect 56376 289768 66628 289796
rect 56376 289756 56382 289768
rect 66622 289756 66628 289768
rect 66680 289756 66686 289808
rect 165430 289756 165436 289808
rect 165488 289796 165494 289808
rect 166350 289796 166356 289808
rect 165488 289768 166356 289796
rect 165488 289756 165494 289768
rect 166350 289756 166356 289768
rect 166408 289756 166414 289808
rect 191374 289076 191380 289128
rect 191432 289116 191438 289128
rect 210970 289116 210976 289128
rect 191432 289088 210976 289116
rect 191432 289076 191438 289088
rect 210970 289076 210976 289088
rect 211028 289076 211034 289128
rect 240502 289076 240508 289128
rect 240560 289116 240566 289128
rect 258166 289116 258172 289128
rect 240560 289088 258172 289116
rect 240560 289076 240566 289088
rect 258166 289076 258172 289088
rect 258224 289116 258230 289128
rect 280890 289116 280896 289128
rect 258224 289088 280896 289116
rect 258224 289076 258230 289088
rect 280890 289076 280896 289088
rect 280948 289076 280954 289128
rect 291286 289076 291292 289128
rect 291344 289116 291350 289128
rect 369854 289116 369860 289128
rect 291344 289088 369860 289116
rect 291344 289076 291350 289088
rect 369854 289076 369860 289088
rect 369912 289076 369918 289128
rect 235166 288872 235172 288924
rect 235224 288912 235230 288924
rect 235994 288912 236000 288924
rect 235224 288884 236000 288912
rect 235224 288872 235230 288884
rect 235994 288872 236000 288884
rect 236052 288872 236058 288924
rect 210510 288464 210516 288516
rect 210568 288504 210574 288516
rect 210970 288504 210976 288516
rect 210568 288476 210976 288504
rect 210568 288464 210574 288476
rect 210970 288464 210976 288476
rect 211028 288504 211034 288516
rect 247402 288504 247408 288516
rect 211028 288476 247408 288504
rect 211028 288464 211034 288476
rect 247402 288464 247408 288476
rect 247460 288464 247466 288516
rect 158806 288396 158812 288448
rect 158864 288436 158870 288448
rect 231302 288436 231308 288448
rect 158864 288408 231308 288436
rect 158864 288396 158870 288408
rect 231302 288396 231308 288408
rect 231360 288396 231366 288448
rect 165062 287648 165068 287700
rect 165120 287688 165126 287700
rect 182910 287688 182916 287700
rect 165120 287660 182916 287688
rect 165120 287648 165126 287660
rect 182910 287648 182916 287660
rect 182968 287648 182974 287700
rect 247034 287648 247040 287700
rect 247092 287688 247098 287700
rect 260098 287688 260104 287700
rect 247092 287660 260104 287688
rect 247092 287648 247098 287660
rect 260098 287648 260104 287660
rect 260156 287648 260162 287700
rect 287698 287648 287704 287700
rect 287756 287688 287762 287700
rect 347774 287688 347780 287700
rect 287756 287660 347780 287688
rect 287756 287648 287762 287660
rect 347774 287648 347780 287660
rect 347832 287648 347838 287700
rect 189994 287104 190000 287156
rect 190052 287144 190058 287156
rect 216766 287144 216772 287156
rect 190052 287116 216772 287144
rect 190052 287104 190058 287116
rect 216766 287104 216772 287116
rect 216824 287104 216830 287156
rect 220630 287104 220636 287156
rect 220688 287144 220694 287156
rect 248506 287144 248512 287156
rect 220688 287116 248512 287144
rect 220688 287104 220694 287116
rect 248506 287104 248512 287116
rect 248564 287104 248570 287156
rect 158714 287036 158720 287088
rect 158772 287076 158778 287088
rect 166258 287076 166264 287088
rect 158772 287048 166264 287076
rect 158772 287036 158778 287048
rect 166258 287036 166264 287048
rect 166316 287036 166322 287088
rect 187050 287036 187056 287088
rect 187108 287076 187114 287088
rect 223574 287076 223580 287088
rect 187108 287048 223580 287076
rect 187108 287036 187114 287048
rect 223574 287036 223580 287048
rect 223632 287036 223638 287088
rect 224402 287036 224408 287088
rect 224460 287076 224466 287088
rect 245470 287076 245476 287088
rect 224460 287048 245476 287076
rect 224460 287036 224466 287048
rect 245470 287036 245476 287048
rect 245528 287036 245534 287088
rect 158806 286968 158812 287020
rect 158864 287008 158870 287020
rect 189902 287008 189908 287020
rect 158864 286980 189908 287008
rect 158864 286968 158870 286980
rect 189902 286968 189908 286980
rect 189960 286968 189966 287020
rect 158714 286288 158720 286340
rect 158772 286328 158778 286340
rect 164878 286328 164884 286340
rect 158772 286300 164884 286328
rect 158772 286288 158778 286300
rect 164878 286288 164884 286300
rect 164936 286288 164942 286340
rect 214558 286288 214564 286340
rect 214616 286328 214622 286340
rect 225046 286328 225052 286340
rect 214616 286300 225052 286328
rect 214616 286288 214622 286300
rect 225046 286288 225052 286300
rect 225104 286288 225110 286340
rect 255498 286288 255504 286340
rect 255556 286328 255562 286340
rect 273254 286328 273260 286340
rect 255556 286300 273260 286328
rect 255556 286288 255562 286300
rect 273254 286288 273260 286300
rect 273312 286288 273318 286340
rect 194502 285812 194508 285864
rect 194560 285852 194566 285864
rect 200758 285852 200764 285864
rect 194560 285824 200764 285852
rect 194560 285812 194566 285824
rect 200758 285812 200764 285824
rect 200816 285812 200822 285864
rect 204622 285852 204628 285864
rect 201144 285824 204628 285852
rect 191098 285744 191104 285796
rect 191156 285784 191162 285796
rect 201144 285784 201172 285824
rect 204622 285812 204628 285824
rect 204680 285812 204686 285864
rect 230750 285852 230756 285864
rect 219406 285824 230756 285852
rect 191156 285756 201172 285784
rect 191156 285744 191162 285756
rect 201218 285744 201224 285796
rect 201276 285784 201282 285796
rect 201276 285756 209774 285784
rect 201276 285744 201282 285756
rect 62758 285716 62764 285728
rect 62132 285688 62764 285716
rect 46842 285608 46848 285660
rect 46900 285648 46906 285660
rect 62132 285648 62160 285688
rect 62758 285676 62764 285688
rect 62816 285716 62822 285728
rect 66806 285716 66812 285728
rect 62816 285688 66812 285716
rect 62816 285676 62822 285688
rect 66806 285676 66812 285688
rect 66864 285676 66870 285728
rect 182910 285676 182916 285728
rect 182968 285716 182974 285728
rect 187234 285716 187240 285728
rect 182968 285688 187240 285716
rect 182968 285676 182974 285688
rect 187234 285676 187240 285688
rect 187292 285676 187298 285728
rect 203150 285676 203156 285728
rect 203208 285716 203214 285728
rect 204162 285716 204168 285728
rect 203208 285688 204168 285716
rect 203208 285676 203214 285688
rect 204162 285676 204168 285688
rect 204220 285676 204226 285728
rect 204898 285676 204904 285728
rect 204956 285716 204962 285728
rect 206094 285716 206100 285728
rect 204956 285688 206100 285716
rect 204956 285676 204962 285688
rect 206094 285676 206100 285688
rect 206152 285676 206158 285728
rect 209746 285716 209774 285756
rect 213454 285744 213460 285796
rect 213512 285784 213518 285796
rect 213914 285784 213920 285796
rect 213512 285756 213920 285784
rect 213512 285744 213518 285756
rect 213914 285744 213920 285756
rect 213972 285744 213978 285796
rect 215294 285744 215300 285796
rect 215352 285784 215358 285796
rect 216582 285784 216588 285796
rect 215352 285756 216588 285784
rect 215352 285744 215358 285756
rect 216582 285744 216588 285756
rect 216640 285744 216646 285796
rect 219406 285716 219434 285824
rect 230750 285812 230756 285824
rect 230808 285852 230814 285864
rect 230808 285824 237512 285852
rect 230808 285812 230814 285824
rect 235442 285744 235448 285796
rect 235500 285784 235506 285796
rect 237484 285784 237512 285824
rect 237558 285812 237564 285864
rect 237616 285852 237622 285864
rect 238662 285852 238668 285864
rect 237616 285824 238668 285852
rect 237616 285812 237622 285824
rect 238662 285812 238668 285824
rect 238720 285812 238726 285864
rect 244182 285784 244188 285796
rect 235500 285756 237420 285784
rect 237484 285756 244188 285784
rect 235500 285744 235506 285756
rect 209746 285688 219434 285716
rect 225414 285676 225420 285728
rect 225472 285716 225478 285728
rect 226978 285716 226984 285728
rect 225472 285688 226984 285716
rect 225472 285676 225478 285688
rect 226978 285676 226984 285688
rect 227036 285676 227042 285728
rect 233142 285676 233148 285728
rect 233200 285716 233206 285728
rect 233970 285716 233976 285728
rect 233200 285688 233976 285716
rect 233200 285676 233206 285688
rect 233970 285676 233976 285688
rect 234028 285676 234034 285728
rect 236086 285676 236092 285728
rect 236144 285716 236150 285728
rect 237282 285716 237288 285728
rect 236144 285688 237288 285716
rect 236144 285676 236150 285688
rect 237282 285676 237288 285688
rect 237340 285676 237346 285728
rect 237392 285716 237420 285756
rect 244182 285744 244188 285756
rect 244240 285744 244246 285796
rect 238478 285716 238484 285728
rect 237392 285688 238484 285716
rect 238478 285676 238484 285688
rect 238536 285716 238542 285728
rect 251818 285716 251824 285728
rect 238536 285688 251824 285716
rect 238536 285676 238542 285688
rect 251818 285676 251824 285688
rect 251876 285676 251882 285728
rect 46900 285620 62160 285648
rect 46900 285608 46906 285620
rect 218054 285608 218060 285660
rect 218112 285648 218118 285660
rect 218606 285648 218612 285660
rect 218112 285620 218612 285648
rect 218112 285608 218118 285620
rect 218606 285608 218612 285620
rect 218664 285648 218670 285660
rect 237374 285648 237380 285660
rect 218664 285620 237380 285648
rect 218664 285608 218670 285620
rect 237374 285608 237380 285620
rect 237432 285608 237438 285660
rect 238938 285608 238944 285660
rect 238996 285648 239002 285660
rect 239582 285648 239588 285660
rect 238996 285620 239588 285648
rect 238996 285608 239002 285620
rect 239582 285608 239588 285620
rect 239640 285648 239646 285660
rect 267090 285648 267096 285660
rect 239640 285620 267096 285648
rect 239640 285608 239646 285620
rect 267090 285608 267096 285620
rect 267148 285608 267154 285660
rect 181622 284996 181628 285048
rect 181680 285036 181686 285048
rect 190454 285036 190460 285048
rect 181680 285008 190460 285036
rect 181680 284996 181686 285008
rect 190454 284996 190460 285008
rect 190512 285036 190518 285048
rect 191742 285036 191748 285048
rect 190512 285008 191748 285036
rect 190512 284996 190518 285008
rect 191742 284996 191748 285008
rect 191800 284996 191806 285048
rect 234706 284996 234712 285048
rect 234764 285036 234770 285048
rect 244550 285036 244556 285048
rect 234764 285008 244556 285036
rect 234764 284996 234770 285008
rect 244550 284996 244556 285008
rect 244608 284996 244614 285048
rect 164878 284928 164884 284980
rect 164936 284968 164942 284980
rect 185670 284968 185676 284980
rect 164936 284940 185676 284968
rect 164936 284928 164942 284940
rect 185670 284928 185676 284940
rect 185728 284928 185734 284980
rect 195974 284928 195980 284980
rect 196032 284968 196038 284980
rect 235442 284968 235448 284980
rect 196032 284940 235448 284968
rect 196032 284928 196038 284940
rect 235442 284928 235448 284940
rect 235500 284928 235506 284980
rect 245470 284928 245476 284980
rect 245528 284968 245534 284980
rect 258166 284968 258172 284980
rect 245528 284940 258172 284968
rect 245528 284928 245534 284940
rect 258166 284928 258172 284940
rect 258224 284928 258230 284980
rect 63402 284316 63408 284368
rect 63460 284356 63466 284368
rect 66254 284356 66260 284368
rect 63460 284328 66260 284356
rect 63460 284316 63466 284328
rect 66254 284316 66260 284328
rect 66312 284316 66318 284368
rect 158714 284316 158720 284368
rect 158772 284356 158778 284368
rect 162762 284356 162768 284368
rect 158772 284328 162768 284356
rect 158772 284316 158778 284328
rect 162762 284316 162768 284328
rect 162820 284316 162826 284368
rect 166718 284316 166724 284368
rect 166776 284356 166782 284368
rect 169018 284356 169024 284368
rect 166776 284328 169024 284356
rect 166776 284316 166782 284328
rect 169018 284316 169024 284328
rect 169076 284316 169082 284368
rect 199470 284316 199476 284368
rect 199528 284356 199534 284368
rect 210878 284356 210884 284368
rect 199528 284328 210884 284356
rect 199528 284316 199534 284328
rect 210878 284316 210884 284328
rect 210936 284316 210942 284368
rect 61838 284248 61844 284300
rect 61896 284288 61902 284300
rect 66990 284288 66996 284300
rect 61896 284260 66996 284288
rect 61896 284248 61902 284260
rect 66990 284248 66996 284260
rect 67048 284248 67054 284300
rect 181622 283908 181628 283960
rect 181680 283948 181686 283960
rect 201126 283948 201132 283960
rect 181680 283920 201132 283948
rect 181680 283908 181686 283920
rect 201126 283908 201132 283920
rect 201184 283908 201190 283960
rect 201218 283908 201224 283960
rect 201276 283908 201282 283960
rect 162210 283840 162216 283892
rect 162268 283880 162274 283892
rect 201236 283880 201264 283908
rect 162268 283852 201264 283880
rect 162268 283840 162274 283852
rect 244182 283568 244188 283620
rect 244240 283608 244246 283620
rect 260834 283608 260840 283620
rect 244240 283580 260840 283608
rect 244240 283568 244246 283580
rect 260834 283568 260840 283580
rect 260892 283568 260898 283620
rect 282362 283568 282368 283620
rect 282420 283608 282426 283620
rect 352558 283608 352564 283620
rect 282420 283580 352564 283608
rect 282420 283568 282426 283580
rect 352558 283568 352564 283580
rect 352616 283568 352622 283620
rect 246850 283160 246856 283212
rect 246908 283200 246914 283212
rect 247218 283200 247224 283212
rect 246908 283172 247224 283200
rect 246908 283160 246914 283172
rect 247218 283160 247224 283172
rect 247276 283200 247282 283212
rect 249794 283200 249800 283212
rect 247276 283172 249800 283200
rect 247276 283160 247282 283172
rect 249794 283160 249800 283172
rect 249852 283160 249858 283212
rect 260742 282928 260748 282940
rect 260655 282900 260748 282928
rect 260742 282888 260748 282900
rect 260800 282928 260806 282940
rect 319438 282928 319444 282940
rect 260800 282900 319444 282928
rect 260800 282888 260806 282900
rect 319438 282888 319444 282900
rect 319496 282888 319502 282940
rect 245930 282820 245936 282872
rect 245988 282860 245994 282872
rect 260760 282860 260788 282888
rect 245988 282832 260788 282860
rect 245988 282820 245994 282832
rect 278774 282820 278780 282872
rect 278832 282860 278838 282872
rect 298094 282860 298100 282872
rect 278832 282832 298100 282860
rect 278832 282820 278838 282832
rect 298094 282820 298100 282832
rect 298152 282860 298158 282872
rect 298738 282860 298744 282872
rect 298152 282832 298744 282860
rect 298152 282820 298158 282832
rect 298738 282820 298744 282832
rect 298796 282820 298802 282872
rect 158714 282548 158720 282600
rect 158772 282588 158778 282600
rect 162946 282588 162952 282600
rect 158772 282560 162952 282588
rect 158772 282548 158778 282560
rect 162946 282548 162952 282560
rect 163004 282548 163010 282600
rect 163590 282208 163596 282260
rect 163648 282248 163654 282260
rect 189902 282248 189908 282260
rect 163648 282220 189908 282248
rect 163648 282208 163654 282220
rect 189902 282208 189908 282220
rect 189960 282208 189966 282260
rect 249702 282208 249708 282260
rect 249760 282248 249766 282260
rect 254118 282248 254124 282260
rect 249760 282220 254124 282248
rect 249760 282208 249766 282220
rect 254118 282208 254124 282220
rect 254176 282208 254182 282260
rect 414658 282208 414664 282260
rect 414716 282248 414722 282260
rect 431954 282248 431960 282260
rect 414716 282220 431960 282248
rect 414716 282208 414722 282220
rect 431954 282208 431960 282220
rect 432012 282208 432018 282260
rect 162762 282140 162768 282192
rect 162820 282180 162826 282192
rect 193122 282180 193128 282192
rect 162820 282152 193128 282180
rect 162820 282140 162826 282152
rect 193122 282140 193128 282152
rect 193180 282180 193186 282192
rect 197354 282180 197360 282192
rect 193180 282152 197360 282180
rect 193180 282140 193186 282152
rect 197354 282140 197360 282152
rect 197412 282140 197418 282192
rect 254578 282140 254584 282192
rect 254636 282180 254642 282192
rect 279418 282180 279424 282192
rect 254636 282152 279424 282180
rect 254636 282140 254642 282152
rect 279418 282140 279424 282152
rect 279476 282140 279482 282192
rect 302878 282140 302884 282192
rect 302936 282180 302942 282192
rect 414750 282180 414756 282192
rect 302936 282152 414756 282180
rect 302936 282140 302942 282152
rect 414750 282140 414756 282152
rect 414808 282140 414814 282192
rect 64598 281528 64604 281580
rect 64656 281568 64662 281580
rect 66806 281568 66812 281580
rect 64656 281540 66812 281568
rect 64656 281528 64662 281540
rect 66806 281528 66812 281540
rect 66864 281528 66870 281580
rect 281442 281460 281448 281512
rect 281500 281500 281506 281512
rect 297358 281500 297364 281512
rect 281500 281472 297364 281500
rect 281500 281460 281506 281472
rect 297358 281460 297364 281472
rect 297416 281460 297422 281512
rect 245930 280780 245936 280832
rect 245988 280820 245994 280832
rect 280338 280820 280344 280832
rect 245988 280792 280344 280820
rect 245988 280780 245994 280792
rect 280338 280780 280344 280792
rect 280396 280820 280402 280832
rect 281442 280820 281448 280832
rect 280396 280792 281448 280820
rect 280396 280780 280402 280792
rect 281442 280780 281448 280792
rect 281500 280780 281506 280832
rect 293218 280780 293224 280832
rect 293276 280820 293282 280832
rect 421558 280820 421564 280832
rect 293276 280792 421564 280820
rect 293276 280780 293282 280792
rect 421558 280780 421564 280792
rect 421616 280780 421622 280832
rect 158714 280236 158720 280288
rect 158772 280276 158778 280288
rect 169018 280276 169024 280288
rect 158772 280248 169024 280276
rect 158772 280236 158778 280248
rect 169018 280236 169024 280248
rect 169076 280236 169082 280288
rect 34330 280168 34336 280220
rect 34388 280208 34394 280220
rect 67174 280208 67180 280220
rect 34388 280180 67180 280208
rect 34388 280168 34394 280180
rect 67174 280168 67180 280180
rect 67232 280168 67238 280220
rect 163682 280168 163688 280220
rect 163740 280208 163746 280220
rect 197354 280208 197360 280220
rect 163740 280180 197360 280208
rect 163740 280168 163746 280180
rect 197354 280168 197360 280180
rect 197412 280168 197418 280220
rect 158714 280100 158720 280152
rect 158772 280140 158778 280152
rect 171778 280140 171784 280152
rect 158772 280112 171784 280140
rect 158772 280100 158778 280112
rect 171778 280100 171784 280112
rect 171836 280100 171842 280152
rect 245930 280100 245936 280152
rect 245988 280140 245994 280152
rect 255498 280140 255504 280152
rect 245988 280112 255504 280140
rect 245988 280100 245994 280112
rect 255498 280100 255504 280112
rect 255556 280100 255562 280152
rect 162302 279420 162308 279472
rect 162360 279460 162366 279472
rect 176194 279460 176200 279472
rect 162360 279432 176200 279460
rect 162360 279420 162366 279432
rect 176194 279420 176200 279432
rect 176252 279420 176258 279472
rect 181714 279420 181720 279472
rect 181772 279460 181778 279472
rect 196710 279460 196716 279472
rect 181772 279432 196716 279460
rect 181772 279420 181778 279432
rect 196710 279420 196716 279432
rect 196768 279420 196774 279472
rect 195330 279352 195336 279404
rect 195388 279392 195394 279404
rect 197354 279392 197360 279404
rect 195388 279364 197360 279392
rect 195388 279352 195394 279364
rect 197354 279352 197360 279364
rect 197412 279352 197418 279404
rect 158714 278808 158720 278860
rect 158772 278848 158778 278860
rect 162394 278848 162400 278860
rect 158772 278820 162400 278848
rect 158772 278808 158778 278820
rect 162394 278808 162400 278820
rect 162452 278808 162458 278860
rect 64690 278740 64696 278792
rect 64748 278780 64754 278792
rect 66806 278780 66812 278792
rect 64748 278752 66812 278780
rect 64748 278740 64754 278752
rect 66806 278740 66812 278752
rect 66864 278740 66870 278792
rect 249702 278740 249708 278792
rect 249760 278780 249766 278792
rect 309778 278780 309784 278792
rect 249760 278752 309784 278780
rect 249760 278740 249766 278752
rect 309778 278740 309784 278752
rect 309836 278740 309842 278792
rect 195422 278604 195428 278656
rect 195480 278644 195486 278656
rect 197354 278644 197360 278656
rect 195480 278616 197360 278644
rect 195480 278604 195486 278616
rect 197354 278604 197360 278616
rect 197412 278604 197418 278656
rect 180150 278060 180156 278112
rect 180208 278100 180214 278112
rect 185670 278100 185676 278112
rect 180208 278072 185676 278100
rect 180208 278060 180214 278072
rect 185670 278060 185676 278072
rect 185728 278060 185734 278112
rect 156874 277992 156880 278044
rect 156932 278032 156938 278044
rect 195974 278032 195980 278044
rect 156932 278004 195980 278032
rect 156932 277992 156938 278004
rect 195974 277992 195980 278004
rect 196032 277992 196038 278044
rect 254026 277992 254032 278044
rect 254084 278032 254090 278044
rect 373994 278032 374000 278044
rect 254084 278004 374000 278032
rect 254084 277992 254090 278004
rect 373994 277992 374000 278004
rect 374052 278032 374058 278044
rect 376018 278032 376024 278044
rect 374052 278004 376024 278032
rect 374052 277992 374058 278004
rect 376018 277992 376024 278004
rect 376076 277992 376082 278044
rect 245930 277380 245936 277432
rect 245988 277420 245994 277432
rect 254026 277420 254032 277432
rect 245988 277392 254032 277420
rect 245988 277380 245994 277392
rect 254026 277380 254032 277392
rect 254084 277380 254090 277432
rect 169018 277312 169024 277364
rect 169076 277352 169082 277364
rect 197354 277352 197360 277364
rect 169076 277324 197360 277352
rect 169076 277312 169082 277324
rect 197354 277312 197360 277324
rect 197412 277312 197418 277364
rect 158714 277244 158720 277296
rect 158772 277284 158778 277296
rect 182910 277284 182916 277296
rect 158772 277256 182916 277284
rect 158772 277244 158778 277256
rect 182910 277244 182916 277256
rect 182968 277244 182974 277296
rect 281442 276740 281448 276752
rect 277366 276712 281448 276740
rect 4062 276632 4068 276684
rect 4120 276672 4126 276684
rect 43438 276672 43444 276684
rect 4120 276644 43444 276672
rect 4120 276632 4126 276644
rect 43438 276632 43444 276644
rect 43496 276632 43502 276684
rect 183370 276632 183376 276684
rect 183428 276672 183434 276684
rect 191282 276672 191288 276684
rect 183428 276644 191288 276672
rect 183428 276632 183434 276644
rect 191282 276632 191288 276644
rect 191340 276632 191346 276684
rect 268378 276632 268384 276684
rect 268436 276672 268442 276684
rect 277366 276672 277394 276712
rect 281442 276700 281448 276712
rect 281500 276740 281506 276752
rect 322290 276740 322296 276752
rect 281500 276712 322296 276740
rect 281500 276700 281506 276712
rect 322290 276700 322296 276712
rect 322348 276700 322354 276752
rect 268436 276644 277394 276672
rect 268436 276632 268442 276644
rect 282270 276632 282276 276684
rect 282328 276672 282334 276684
rect 296714 276672 296720 276684
rect 282328 276644 296720 276672
rect 282328 276632 282334 276644
rect 296714 276632 296720 276644
rect 296772 276632 296778 276684
rect 308398 276632 308404 276684
rect 308456 276672 308462 276684
rect 395338 276672 395344 276684
rect 308456 276644 395344 276672
rect 308456 276632 308462 276644
rect 395338 276632 395344 276644
rect 395396 276632 395402 276684
rect 52178 276020 52184 276072
rect 52236 276060 52242 276072
rect 66346 276060 66352 276072
rect 52236 276032 66352 276060
rect 52236 276020 52242 276032
rect 66346 276020 66352 276032
rect 66404 276020 66410 276072
rect 245746 275952 245752 276004
rect 245804 275992 245810 276004
rect 263778 275992 263784 276004
rect 245804 275964 263784 275992
rect 245804 275952 245810 275964
rect 263778 275952 263784 275964
rect 263836 275952 263842 276004
rect 245930 275884 245936 275936
rect 245988 275924 245994 275936
rect 253934 275924 253940 275936
rect 245988 275896 253940 275924
rect 245988 275884 245994 275896
rect 253934 275884 253940 275896
rect 253992 275884 253998 275936
rect 169662 275544 169668 275596
rect 169720 275584 169726 275596
rect 172514 275584 172520 275596
rect 169720 275556 172520 275584
rect 169720 275544 169726 275556
rect 172514 275544 172520 275556
rect 172572 275544 172578 275596
rect 263778 275340 263784 275392
rect 263836 275380 263842 275392
rect 353938 275380 353944 275392
rect 263836 275352 353944 275380
rect 263836 275340 263842 275352
rect 353938 275340 353944 275352
rect 353996 275340 354002 275392
rect 163590 275272 163596 275324
rect 163648 275312 163654 275324
rect 185762 275312 185768 275324
rect 163648 275284 185768 275312
rect 163648 275272 163654 275284
rect 185762 275272 185768 275284
rect 185820 275272 185826 275324
rect 253934 275272 253940 275324
rect 253992 275312 253998 275324
rect 417418 275312 417424 275324
rect 253992 275284 417424 275312
rect 253992 275272 253998 275284
rect 417418 275272 417424 275284
rect 417476 275272 417482 275324
rect 158714 274864 158720 274916
rect 158772 274904 158778 274916
rect 161014 274904 161020 274916
rect 158772 274876 161020 274904
rect 158772 274864 158778 274876
rect 161014 274864 161020 274876
rect 161072 274864 161078 274916
rect 191558 274728 191564 274780
rect 191616 274768 191622 274780
rect 195422 274768 195428 274780
rect 191616 274740 195428 274768
rect 191616 274728 191622 274740
rect 195422 274728 195428 274740
rect 195480 274728 195486 274780
rect 180150 274660 180156 274712
rect 180208 274700 180214 274712
rect 197354 274700 197360 274712
rect 180208 274672 197360 274700
rect 180208 274660 180214 274672
rect 197354 274660 197360 274672
rect 197412 274660 197418 274712
rect 34422 274592 34428 274644
rect 34480 274632 34486 274644
rect 65978 274632 65984 274644
rect 34480 274604 65984 274632
rect 34480 274592 34486 274604
rect 65978 274592 65984 274604
rect 66036 274592 66042 274644
rect 158714 274592 158720 274644
rect 158772 274632 158778 274644
rect 170398 274632 170404 274644
rect 158772 274604 170404 274632
rect 158772 274592 158778 274604
rect 170398 274592 170404 274604
rect 170456 274592 170462 274644
rect 279510 274592 279516 274644
rect 279568 274632 279574 274644
rect 358722 274632 358728 274644
rect 279568 274604 358728 274632
rect 279568 274592 279574 274604
rect 358722 274592 358728 274604
rect 358780 274592 358786 274644
rect 167638 273980 167644 274032
rect 167696 274020 167702 274032
rect 182082 274020 182088 274032
rect 167696 273992 182088 274020
rect 167696 273980 167702 273992
rect 182082 273980 182088 273992
rect 182140 273980 182146 274032
rect 176102 273912 176108 273964
rect 176160 273952 176166 273964
rect 195974 273952 195980 273964
rect 176160 273924 195980 273952
rect 176160 273912 176166 273924
rect 195974 273912 195980 273924
rect 196032 273912 196038 273964
rect 262950 273912 262956 273964
rect 263008 273952 263014 273964
rect 370498 273952 370504 273964
rect 263008 273924 370504 273952
rect 263008 273912 263014 273924
rect 370498 273912 370504 273924
rect 370556 273912 370562 273964
rect 63218 273232 63224 273284
rect 63276 273272 63282 273284
rect 66806 273272 66812 273284
rect 63276 273244 66812 273272
rect 63276 273232 63282 273244
rect 66806 273232 66812 273244
rect 66864 273232 66870 273284
rect 182082 273232 182088 273284
rect 182140 273272 182146 273284
rect 197446 273272 197452 273284
rect 182140 273244 197452 273272
rect 182140 273232 182146 273244
rect 197446 273232 197452 273244
rect 197504 273232 197510 273284
rect 245838 273232 245844 273284
rect 245896 273272 245902 273284
rect 253934 273272 253940 273284
rect 245896 273244 253940 273272
rect 245896 273232 245902 273244
rect 253934 273232 253940 273244
rect 253992 273232 253998 273284
rect 358722 273232 358728 273284
rect 358780 273272 358786 273284
rect 363598 273272 363604 273284
rect 358780 273244 363604 273272
rect 358780 273232 358786 273244
rect 363598 273232 363604 273244
rect 363656 273232 363662 273284
rect 180702 273164 180708 273216
rect 180760 273204 180766 273216
rect 197354 273204 197360 273216
rect 180760 273176 197360 273204
rect 180760 273164 180766 273176
rect 197354 273164 197360 273176
rect 197412 273164 197418 273216
rect 245930 273164 245936 273216
rect 245988 273204 245994 273216
rect 254210 273204 254216 273216
rect 245988 273176 254216 273204
rect 245988 273164 245994 273176
rect 254210 273164 254216 273176
rect 254268 273164 254274 273216
rect 276842 273164 276848 273216
rect 276900 273204 276906 273216
rect 277394 273204 277400 273216
rect 276900 273176 277400 273204
rect 276900 273164 276906 273176
rect 277394 273164 277400 273176
rect 277452 273204 277458 273216
rect 376846 273204 376852 273216
rect 277452 273176 376852 273204
rect 277452 273164 277458 273176
rect 376846 273164 376852 273176
rect 376904 273164 376910 273216
rect 251818 272552 251824 272604
rect 251876 272592 251882 272604
rect 262214 272592 262220 272604
rect 251876 272564 262220 272592
rect 251876 272552 251882 272564
rect 262214 272552 262220 272564
rect 262272 272552 262278 272604
rect 188430 272484 188436 272536
rect 188488 272524 188494 272536
rect 199470 272524 199476 272536
rect 188488 272496 199476 272524
rect 188488 272484 188494 272496
rect 199470 272484 199476 272496
rect 199528 272484 199534 272536
rect 245746 272484 245752 272536
rect 245804 272524 245810 272536
rect 251174 272524 251180 272536
rect 245804 272496 251180 272524
rect 245804 272484 245810 272496
rect 251174 272484 251180 272496
rect 251232 272484 251238 272536
rect 254210 272484 254216 272536
rect 254268 272524 254274 272536
rect 313366 272524 313372 272536
rect 254268 272496 313372 272524
rect 254268 272484 254274 272496
rect 313366 272484 313372 272496
rect 313424 272524 313430 272536
rect 358906 272524 358912 272536
rect 313424 272496 358912 272524
rect 313424 272484 313430 272496
rect 358906 272484 358912 272496
rect 358964 272484 358970 272536
rect 50798 271872 50804 271924
rect 50856 271912 50862 271924
rect 66714 271912 66720 271924
rect 50856 271884 66720 271912
rect 50856 271872 50862 271884
rect 66714 271872 66720 271884
rect 66772 271872 66778 271924
rect 56502 271804 56508 271856
rect 56560 271844 56566 271856
rect 66806 271844 66812 271856
rect 56560 271816 66812 271844
rect 56560 271804 56566 271816
rect 66806 271804 66812 271816
rect 66864 271804 66870 271856
rect 282270 271804 282276 271856
rect 282328 271844 282334 271856
rect 385034 271844 385040 271856
rect 282328 271816 385040 271844
rect 282328 271804 282334 271816
rect 385034 271804 385040 271816
rect 385092 271804 385098 271856
rect 245930 271396 245936 271448
rect 245988 271436 245994 271448
rect 248598 271436 248604 271448
rect 245988 271408 248604 271436
rect 245988 271396 245994 271408
rect 248598 271396 248604 271408
rect 248656 271396 248662 271448
rect 158806 271124 158812 271176
rect 158864 271164 158870 271176
rect 167730 271164 167736 271176
rect 158864 271136 167736 271164
rect 158864 271124 158870 271136
rect 167730 271124 167736 271136
rect 167788 271124 167794 271176
rect 274174 271124 274180 271176
rect 274232 271164 274238 271176
rect 293954 271164 293960 271176
rect 274232 271136 293960 271164
rect 274232 271124 274238 271136
rect 293954 271124 293960 271136
rect 294012 271124 294018 271176
rect 168190 270580 168196 270632
rect 168248 270620 168254 270632
rect 197354 270620 197360 270632
rect 168248 270592 197360 270620
rect 168248 270580 168254 270592
rect 197354 270580 197360 270592
rect 197412 270580 197418 270632
rect 158714 270512 158720 270564
rect 158772 270552 158778 270564
rect 196802 270552 196808 270564
rect 158772 270524 196808 270552
rect 158772 270512 158778 270524
rect 196802 270512 196808 270524
rect 196860 270512 196866 270564
rect 245838 270444 245844 270496
rect 245896 270484 245902 270496
rect 262306 270484 262312 270496
rect 245896 270456 262312 270484
rect 245896 270444 245902 270456
rect 262306 270444 262312 270456
rect 262364 270484 262370 270496
rect 262674 270484 262680 270496
rect 262364 270456 262680 270484
rect 262364 270444 262370 270456
rect 262674 270444 262680 270456
rect 262732 270444 262738 270496
rect 244274 270172 244280 270224
rect 244332 270212 244338 270224
rect 248414 270212 248420 270224
rect 244332 270184 248420 270212
rect 244332 270172 244338 270184
rect 248414 270172 248420 270184
rect 248472 270172 248478 270224
rect 169110 269832 169116 269884
rect 169168 269872 169174 269884
rect 178678 269872 178684 269884
rect 169168 269844 178684 269872
rect 169168 269832 169174 269844
rect 178678 269832 178684 269844
rect 178736 269832 178742 269884
rect 159634 269764 159640 269816
rect 159692 269804 159698 269816
rect 170398 269804 170404 269816
rect 159692 269776 170404 269804
rect 159692 269764 159698 269776
rect 170398 269764 170404 269776
rect 170456 269764 170462 269816
rect 172422 269764 172428 269816
rect 172480 269804 172486 269816
rect 191190 269804 191196 269816
rect 172480 269776 191196 269804
rect 172480 269764 172486 269776
rect 191190 269764 191196 269776
rect 191248 269764 191254 269816
rect 262674 269764 262680 269816
rect 262732 269804 262738 269816
rect 291194 269804 291200 269816
rect 262732 269776 291200 269804
rect 262732 269764 262738 269776
rect 291194 269764 291200 269776
rect 291252 269764 291258 269816
rect 178678 269084 178684 269136
rect 178736 269124 178742 269136
rect 197354 269124 197360 269136
rect 178736 269096 197360 269124
rect 178736 269084 178742 269096
rect 197354 269084 197360 269096
rect 197412 269084 197418 269136
rect 158714 269016 158720 269068
rect 158772 269056 158778 269068
rect 187050 269056 187056 269068
rect 158772 269028 187056 269056
rect 158772 269016 158778 269028
rect 187050 269016 187056 269028
rect 187108 269016 187114 269068
rect 178034 268948 178040 269000
rect 178092 268988 178098 269000
rect 178770 268988 178776 269000
rect 178092 268960 178776 268988
rect 178092 268948 178098 268960
rect 178770 268948 178776 268960
rect 178828 268988 178834 269000
rect 197354 268988 197360 269000
rect 178828 268960 197360 268988
rect 178828 268948 178834 268960
rect 197354 268948 197360 268960
rect 197412 268948 197418 269000
rect 253198 268404 253204 268456
rect 253256 268444 253262 268456
rect 264330 268444 264336 268456
rect 253256 268416 264336 268444
rect 253256 268404 253262 268416
rect 264330 268404 264336 268416
rect 264388 268404 264394 268456
rect 167638 268336 167644 268388
rect 167696 268376 167702 268388
rect 178034 268376 178040 268388
rect 167696 268348 178040 268376
rect 167696 268336 167702 268348
rect 178034 268336 178040 268348
rect 178092 268336 178098 268388
rect 246298 268336 246304 268388
rect 246356 268376 246362 268388
rect 323578 268376 323584 268388
rect 246356 268348 323584 268376
rect 246356 268336 246362 268348
rect 323578 268336 323584 268348
rect 323636 268336 323642 268388
rect 355318 268336 355324 268388
rect 355376 268376 355382 268388
rect 580166 268376 580172 268388
rect 355376 268348 580172 268376
rect 355376 268336 355382 268348
rect 580166 268336 580172 268348
rect 580224 268336 580230 268388
rect 191742 268132 191748 268184
rect 191800 268172 191806 268184
rect 197446 268172 197452 268184
rect 191800 268144 197452 268172
rect 191800 268132 191806 268144
rect 197446 268132 197452 268144
rect 197504 268132 197510 268184
rect 64782 267792 64788 267844
rect 64840 267832 64846 267844
rect 66806 267832 66812 267844
rect 64840 267804 66812 267832
rect 64840 267792 64846 267804
rect 66806 267792 66812 267804
rect 66864 267792 66870 267844
rect 245746 267656 245752 267708
rect 245804 267696 245810 267708
rect 265066 267696 265072 267708
rect 245804 267668 265072 267696
rect 245804 267656 245810 267668
rect 265066 267656 265072 267668
rect 265124 267656 265130 267708
rect 166442 267044 166448 267096
rect 166500 267084 166506 267096
rect 175918 267084 175924 267096
rect 166500 267056 175924 267084
rect 166500 267044 166506 267056
rect 175918 267044 175924 267056
rect 175976 267044 175982 267096
rect 179322 267044 179328 267096
rect 179380 267084 179386 267096
rect 188338 267084 188344 267096
rect 179380 267056 188344 267084
rect 179380 267044 179386 267056
rect 188338 267044 188344 267056
rect 188396 267044 188402 267096
rect 3510 266976 3516 267028
rect 3568 267016 3574 267028
rect 14458 267016 14464 267028
rect 3568 266988 14464 267016
rect 3568 266976 3574 266988
rect 14458 266976 14464 266988
rect 14516 266976 14522 267028
rect 57606 266976 57612 267028
rect 57664 267016 57670 267028
rect 66898 267016 66904 267028
rect 57664 266988 66904 267016
rect 57664 266976 57670 266988
rect 66898 266976 66904 266988
rect 66956 266976 66962 267028
rect 173342 266976 173348 267028
rect 173400 267016 173406 267028
rect 184842 267016 184848 267028
rect 173400 266988 184848 267016
rect 173400 266976 173406 266988
rect 184842 266976 184848 266988
rect 184900 266976 184906 267028
rect 265066 266976 265072 267028
rect 265124 267016 265130 267028
rect 302878 267016 302884 267028
rect 265124 266988 302884 267016
rect 265124 266976 265130 266988
rect 302878 266976 302884 266988
rect 302936 266976 302942 267028
rect 304442 266976 304448 267028
rect 304500 267016 304506 267028
rect 367186 267016 367192 267028
rect 304500 266988 367192 267016
rect 304500 266976 304506 266988
rect 367186 266976 367192 266988
rect 367244 266976 367250 267028
rect 188706 266432 188712 266484
rect 188764 266472 188770 266484
rect 195974 266472 195980 266484
rect 188764 266444 195980 266472
rect 188764 266432 188770 266444
rect 195974 266432 195980 266444
rect 196032 266432 196038 266484
rect 184842 266364 184848 266416
rect 184900 266404 184906 266416
rect 197354 266404 197360 266416
rect 184900 266376 197360 266404
rect 184900 266364 184906 266376
rect 197354 266364 197360 266376
rect 197412 266364 197418 266416
rect 245654 265820 245660 265872
rect 245712 265860 245718 265872
rect 249886 265860 249892 265872
rect 245712 265832 249892 265860
rect 245712 265820 245718 265832
rect 249886 265820 249892 265832
rect 249944 265820 249950 265872
rect 173342 265616 173348 265668
rect 173400 265656 173406 265668
rect 181622 265656 181628 265668
rect 173400 265628 181628 265656
rect 173400 265616 173406 265628
rect 181622 265616 181628 265628
rect 181680 265616 181686 265668
rect 255314 265616 255320 265668
rect 255372 265656 255378 265668
rect 371878 265656 371884 265668
rect 255372 265628 371884 265656
rect 255372 265616 255378 265628
rect 371878 265616 371884 265628
rect 371936 265616 371942 265668
rect 53466 264936 53472 264988
rect 53524 264976 53530 264988
rect 66898 264976 66904 264988
rect 53524 264948 66904 264976
rect 53524 264936 53530 264948
rect 66898 264936 66904 264948
rect 66956 264936 66962 264988
rect 158714 264936 158720 264988
rect 158772 264976 158778 264988
rect 180334 264976 180340 264988
rect 158772 264948 180340 264976
rect 158772 264936 158778 264948
rect 180334 264936 180340 264948
rect 180392 264936 180398 264988
rect 245838 264868 245844 264920
rect 245896 264908 245902 264920
rect 266354 264908 266360 264920
rect 245896 264880 266360 264908
rect 245896 264868 245902 264880
rect 266354 264868 266360 264880
rect 266412 264868 266418 264920
rect 268378 264256 268384 264308
rect 268436 264296 268442 264308
rect 316034 264296 316040 264308
rect 268436 264268 316040 264296
rect 268436 264256 268442 264268
rect 316034 264256 316040 264268
rect 316092 264256 316098 264308
rect 266354 264188 266360 264240
rect 266412 264228 266418 264240
rect 267642 264228 267648 264240
rect 266412 264200 267648 264228
rect 266412 264188 266418 264200
rect 267642 264188 267648 264200
rect 267700 264228 267706 264240
rect 298738 264228 298744 264240
rect 267700 264200 298744 264228
rect 267700 264188 267706 264200
rect 298738 264188 298744 264200
rect 298796 264188 298802 264240
rect 304258 264188 304264 264240
rect 304316 264228 304322 264240
rect 450538 264228 450544 264240
rect 304316 264200 450544 264228
rect 304316 264188 304322 264200
rect 450538 264188 450544 264200
rect 450596 264188 450602 264240
rect 188614 263644 188620 263696
rect 188672 263684 188678 263696
rect 197446 263684 197452 263696
rect 188672 263656 197452 263684
rect 188672 263644 188678 263656
rect 197446 263644 197452 263656
rect 197504 263644 197510 263696
rect 59078 263576 59084 263628
rect 59136 263616 59142 263628
rect 59262 263616 59268 263628
rect 59136 263588 59268 263616
rect 59136 263576 59142 263588
rect 59262 263576 59268 263588
rect 59320 263616 59326 263628
rect 66438 263616 66444 263628
rect 59320 263588 66444 263616
rect 59320 263576 59326 263588
rect 66438 263576 66444 263588
rect 66496 263576 66502 263628
rect 187050 263576 187056 263628
rect 187108 263616 187114 263628
rect 197354 263616 197360 263628
rect 187108 263588 197360 263616
rect 187108 263576 187114 263588
rect 197354 263576 197360 263588
rect 197412 263576 197418 263628
rect 244090 263372 244096 263424
rect 244148 263412 244154 263424
rect 245654 263412 245660 263424
rect 244148 263384 245660 263412
rect 244148 263372 244154 263384
rect 245654 263372 245660 263384
rect 245712 263372 245718 263424
rect 67542 262896 67548 262948
rect 67600 262936 67606 262948
rect 68278 262936 68284 262948
rect 67600 262908 68284 262936
rect 67600 262896 67606 262908
rect 68278 262896 68284 262908
rect 68336 262896 68342 262948
rect 280890 262896 280896 262948
rect 280948 262936 280954 262948
rect 308398 262936 308404 262948
rect 280948 262908 308404 262936
rect 280948 262896 280954 262908
rect 308398 262896 308404 262908
rect 308456 262896 308462 262948
rect 160922 262828 160928 262880
rect 160980 262868 160986 262880
rect 165062 262868 165068 262880
rect 160980 262840 165068 262868
rect 160980 262828 160986 262840
rect 165062 262828 165068 262840
rect 165120 262828 165126 262880
rect 165430 262828 165436 262880
rect 165488 262868 165494 262880
rect 180150 262868 180156 262880
rect 165488 262840 180156 262868
rect 165488 262828 165494 262840
rect 180150 262828 180156 262840
rect 180208 262828 180214 262880
rect 262766 262828 262772 262880
rect 262824 262868 262830 262880
rect 378778 262868 378784 262880
rect 262824 262840 378784 262868
rect 262824 262828 262830 262840
rect 378778 262828 378784 262840
rect 378836 262828 378842 262880
rect 57698 262624 57704 262676
rect 57756 262664 57762 262676
rect 59262 262664 59268 262676
rect 57756 262636 59268 262664
rect 57756 262624 57762 262636
rect 59262 262624 59268 262636
rect 59320 262624 59326 262676
rect 158714 262624 158720 262676
rect 158772 262664 158778 262676
rect 160830 262664 160836 262676
rect 158772 262636 160836 262664
rect 158772 262624 158778 262636
rect 160830 262624 160836 262636
rect 160888 262624 160894 262676
rect 181622 262624 181628 262676
rect 181680 262664 181686 262676
rect 184382 262664 184388 262676
rect 181680 262636 184388 262664
rect 181680 262624 181686 262636
rect 184382 262624 184388 262636
rect 184440 262624 184446 262676
rect 59262 262216 59268 262268
rect 59320 262256 59326 262268
rect 66898 262256 66904 262268
rect 59320 262228 66904 262256
rect 59320 262216 59326 262228
rect 66898 262216 66904 262228
rect 66956 262216 66962 262268
rect 195330 262216 195336 262268
rect 195388 262256 195394 262268
rect 197998 262256 198004 262268
rect 195388 262228 198004 262256
rect 195388 262216 195394 262228
rect 197998 262216 198004 262228
rect 198056 262216 198062 262268
rect 245930 262216 245936 262268
rect 245988 262256 245994 262268
rect 255314 262256 255320 262268
rect 245988 262228 255320 262256
rect 245988 262216 245994 262228
rect 255314 262216 255320 262228
rect 255372 262216 255378 262268
rect 186314 262148 186320 262200
rect 186372 262188 186378 262200
rect 186958 262188 186964 262200
rect 186372 262160 186964 262188
rect 186372 262148 186378 262160
rect 186958 262148 186964 262160
rect 187016 262188 187022 262200
rect 197354 262188 197360 262200
rect 187016 262160 197360 262188
rect 187016 262148 187022 262160
rect 197354 262148 197360 262160
rect 197412 262148 197418 262200
rect 185762 262080 185768 262132
rect 185820 262120 185826 262132
rect 195422 262120 195428 262132
rect 185820 262092 195428 262120
rect 185820 262080 185826 262092
rect 195422 262080 195428 262092
rect 195480 262080 195486 262132
rect 158990 261536 158996 261588
rect 159048 261576 159054 261588
rect 159450 261576 159456 261588
rect 159048 261548 159456 261576
rect 159048 261536 159054 261548
rect 159450 261536 159456 261548
rect 159508 261576 159514 261588
rect 170490 261576 170496 261588
rect 159508 261548 170496 261576
rect 159508 261536 159514 261548
rect 170490 261536 170496 261548
rect 170548 261536 170554 261588
rect 265618 261536 265624 261588
rect 265676 261576 265682 261588
rect 302234 261576 302240 261588
rect 265676 261548 302240 261576
rect 265676 261536 265682 261548
rect 302234 261536 302240 261548
rect 302292 261536 302298 261588
rect 43438 261468 43444 261520
rect 43496 261508 43502 261520
rect 65886 261508 65892 261520
rect 43496 261480 65892 261508
rect 43496 261468 43502 261480
rect 65886 261468 65892 261480
rect 65944 261508 65950 261520
rect 66530 261508 66536 261520
rect 65944 261480 66536 261508
rect 65944 261468 65950 261480
rect 66530 261468 66536 261480
rect 66588 261468 66594 261520
rect 161014 261468 161020 261520
rect 161072 261508 161078 261520
rect 175918 261508 175924 261520
rect 161072 261480 175924 261508
rect 161072 261468 161078 261480
rect 175918 261468 175924 261480
rect 175976 261468 175982 261520
rect 299566 261468 299572 261520
rect 299624 261508 299630 261520
rect 354030 261508 354036 261520
rect 299624 261480 354036 261508
rect 299624 261468 299630 261480
rect 354030 261468 354036 261480
rect 354088 261468 354094 261520
rect 245838 260924 245844 260976
rect 245896 260964 245902 260976
rect 248414 260964 248420 260976
rect 245896 260936 248420 260964
rect 245896 260924 245902 260936
rect 248414 260924 248420 260936
rect 248472 260964 248478 260976
rect 248690 260964 248696 260976
rect 248472 260936 248696 260964
rect 248472 260924 248478 260936
rect 248690 260924 248696 260936
rect 248748 260924 248754 260976
rect 56502 260856 56508 260908
rect 56560 260896 56566 260908
rect 66346 260896 66352 260908
rect 56560 260868 66352 260896
rect 56560 260856 56566 260868
rect 66346 260856 66352 260868
rect 66404 260856 66410 260908
rect 162762 260788 162768 260840
rect 162820 260828 162826 260840
rect 162820 260800 180794 260828
rect 162820 260788 162826 260800
rect 180766 260760 180794 260800
rect 182082 260788 182088 260840
rect 182140 260828 182146 260840
rect 182910 260828 182916 260840
rect 182140 260800 182916 260828
rect 182140 260788 182146 260800
rect 182910 260788 182916 260800
rect 182968 260788 182974 260840
rect 182818 260760 182824 260772
rect 180766 260732 182824 260760
rect 182818 260720 182824 260732
rect 182876 260720 182882 260772
rect 288342 260108 288348 260160
rect 288400 260148 288406 260160
rect 375374 260148 375380 260160
rect 288400 260120 375380 260148
rect 288400 260108 288406 260120
rect 375374 260108 375380 260120
rect 375432 260108 375438 260160
rect 245746 259836 245752 259888
rect 245804 259876 245810 259888
rect 249886 259876 249892 259888
rect 245804 259848 249892 259876
rect 245804 259836 245810 259848
rect 249886 259836 249892 259848
rect 249944 259836 249950 259888
rect 194502 259768 194508 259820
rect 194560 259808 194566 259820
rect 196066 259808 196072 259820
rect 194560 259780 196072 259808
rect 194560 259768 194566 259780
rect 196066 259768 196072 259780
rect 196124 259808 196130 259820
rect 197262 259808 197268 259820
rect 196124 259780 197268 259808
rect 196124 259768 196130 259780
rect 197262 259768 197268 259780
rect 197320 259768 197326 259820
rect 170950 259428 170956 259480
rect 171008 259468 171014 259480
rect 171134 259468 171140 259480
rect 171008 259440 171140 259468
rect 171008 259428 171014 259440
rect 171134 259428 171140 259440
rect 171192 259428 171198 259480
rect 183002 259428 183008 259480
rect 183060 259468 183066 259480
rect 197354 259468 197360 259480
rect 183060 259440 197360 259468
rect 183060 259428 183066 259440
rect 197354 259428 197360 259440
rect 197412 259428 197418 259480
rect 246390 259428 246396 259480
rect 246448 259468 246454 259480
rect 287146 259468 287152 259480
rect 246448 259440 287152 259468
rect 246448 259428 246454 259440
rect 287146 259428 287152 259440
rect 287204 259468 287210 259480
rect 288342 259468 288348 259480
rect 287204 259440 288348 259468
rect 287204 259428 287210 259440
rect 288342 259428 288348 259440
rect 288400 259428 288406 259480
rect 186222 259360 186228 259412
rect 186280 259400 186286 259412
rect 187418 259400 187424 259412
rect 186280 259372 187424 259400
rect 186280 259360 186286 259372
rect 187418 259360 187424 259372
rect 187476 259360 187482 259412
rect 245746 259360 245752 259412
rect 245804 259400 245810 259412
rect 265066 259400 265072 259412
rect 245804 259372 265072 259400
rect 245804 259360 245810 259372
rect 265066 259360 265072 259372
rect 265124 259360 265130 259412
rect 186222 259224 186228 259276
rect 186280 259264 186286 259276
rect 189994 259264 190000 259276
rect 186280 259236 190000 259264
rect 186280 259224 186286 259236
rect 189994 259224 190000 259236
rect 190052 259224 190058 259276
rect 265066 258748 265072 258800
rect 265124 258788 265130 258800
rect 292574 258788 292580 258800
rect 265124 258760 292580 258788
rect 265124 258748 265130 258760
rect 292574 258748 292580 258760
rect 292632 258788 292638 258800
rect 368474 258788 368480 258800
rect 292632 258760 368480 258788
rect 292632 258748 292638 258760
rect 368474 258748 368480 258760
rect 368532 258748 368538 258800
rect 164970 258680 164976 258732
rect 165028 258720 165034 258732
rect 181714 258720 181720 258732
rect 165028 258692 181720 258720
rect 165028 258680 165034 258692
rect 181714 258680 181720 258692
rect 181772 258680 181778 258732
rect 288618 258680 288624 258732
rect 288676 258720 288682 258732
rect 372706 258720 372712 258732
rect 288676 258692 372712 258720
rect 288676 258680 288682 258692
rect 372706 258680 372712 258692
rect 372764 258680 372770 258732
rect 187418 258136 187424 258188
rect 187476 258176 187482 258188
rect 197354 258176 197360 258188
rect 187476 258148 197360 258176
rect 187476 258136 187482 258148
rect 197354 258136 197360 258148
rect 197412 258136 197418 258188
rect 66254 258108 66260 258120
rect 57946 258080 66260 258108
rect 53742 258000 53748 258052
rect 53800 258040 53806 258052
rect 57238 258040 57244 258052
rect 53800 258012 57244 258040
rect 53800 258000 53806 258012
rect 57238 258000 57244 258012
rect 57296 258040 57302 258052
rect 57946 258040 57974 258080
rect 66254 258068 66260 258080
rect 66312 258068 66318 258120
rect 158806 258068 158812 258120
rect 158864 258108 158870 258120
rect 186222 258108 186228 258120
rect 158864 258080 186228 258108
rect 158864 258068 158870 258080
rect 186222 258068 186228 258080
rect 186280 258068 186286 258120
rect 244550 258068 244556 258120
rect 244608 258108 244614 258120
rect 288618 258108 288624 258120
rect 244608 258080 288624 258108
rect 244608 258068 244614 258080
rect 288618 258068 288624 258080
rect 288676 258068 288682 258120
rect 57296 258012 57974 258040
rect 57296 258000 57302 258012
rect 158714 258000 158720 258052
rect 158772 258040 158778 258052
rect 163682 258040 163688 258052
rect 158772 258012 163688 258040
rect 158772 258000 158778 258012
rect 163682 258000 163688 258012
rect 163740 258000 163746 258052
rect 172330 258000 172336 258052
rect 172388 258040 172394 258052
rect 173434 258040 173440 258052
rect 172388 258012 173440 258040
rect 172388 258000 172394 258012
rect 173434 258000 173440 258012
rect 173492 258000 173498 258052
rect 245746 258000 245752 258052
rect 245804 258040 245810 258052
rect 256786 258040 256792 258052
rect 245804 258012 256792 258040
rect 245804 258000 245810 258012
rect 256786 258000 256792 258012
rect 256844 258000 256850 258052
rect 184290 257320 184296 257372
rect 184348 257360 184354 257372
rect 199378 257360 199384 257372
rect 184348 257332 199384 257360
rect 184348 257320 184354 257332
rect 199378 257320 199384 257332
rect 199436 257320 199442 257372
rect 256786 257320 256792 257372
rect 256844 257360 256850 257372
rect 295426 257360 295432 257372
rect 256844 257332 295432 257360
rect 256844 257320 256850 257332
rect 295426 257320 295432 257332
rect 295484 257320 295490 257372
rect 308398 257320 308404 257372
rect 308456 257360 308462 257372
rect 383010 257360 383016 257372
rect 308456 257332 383016 257360
rect 308456 257320 308462 257332
rect 383010 257320 383016 257332
rect 383068 257320 383074 257372
rect 272518 256844 272524 256896
rect 272576 256884 272582 256896
rect 279510 256884 279516 256896
rect 272576 256856 279516 256884
rect 272576 256844 272582 256856
rect 279510 256844 279516 256856
rect 279568 256844 279574 256896
rect 61838 256708 61844 256760
rect 61896 256748 61902 256760
rect 66806 256748 66812 256760
rect 61896 256720 66812 256748
rect 61896 256708 61902 256720
rect 66806 256708 66812 256720
rect 66864 256708 66870 256760
rect 164142 256708 164148 256760
rect 164200 256748 164206 256760
rect 189074 256748 189080 256760
rect 164200 256720 189080 256748
rect 164200 256708 164206 256720
rect 189074 256708 189080 256720
rect 189132 256708 189138 256760
rect 196802 256708 196808 256760
rect 196860 256748 196866 256760
rect 197262 256748 197268 256760
rect 196860 256720 197268 256748
rect 196860 256708 196866 256720
rect 197262 256708 197268 256720
rect 197320 256708 197326 256760
rect 194410 256640 194416 256692
rect 194468 256680 194474 256692
rect 197354 256680 197360 256692
rect 194468 256652 197360 256680
rect 194468 256640 194474 256652
rect 197354 256640 197360 256652
rect 197412 256640 197418 256692
rect 169018 255960 169024 256012
rect 169076 256000 169082 256012
rect 194410 256000 194416 256012
rect 169076 255972 194416 256000
rect 169076 255960 169082 255972
rect 194410 255960 194416 255972
rect 194468 255960 194474 256012
rect 245654 255960 245660 256012
rect 245712 256000 245718 256012
rect 302234 256000 302240 256012
rect 245712 255972 302240 256000
rect 245712 255960 245718 255972
rect 302234 255960 302240 255972
rect 302292 256000 302298 256012
rect 360378 256000 360384 256012
rect 302292 255972 360384 256000
rect 302292 255960 302298 255972
rect 360378 255960 360384 255972
rect 360436 255960 360442 256012
rect 245746 255348 245752 255400
rect 245804 255388 245810 255400
rect 249978 255388 249984 255400
rect 245804 255360 249984 255388
rect 245804 255348 245810 255360
rect 249978 255348 249984 255360
rect 250036 255388 250042 255400
rect 251082 255388 251088 255400
rect 250036 255360 251088 255388
rect 250036 255348 250042 255360
rect 251082 255348 251088 255360
rect 251140 255348 251146 255400
rect 158530 255280 158536 255332
rect 158588 255320 158594 255332
rect 177390 255320 177396 255332
rect 158588 255292 177396 255320
rect 158588 255280 158594 255292
rect 177390 255280 177396 255292
rect 177448 255280 177454 255332
rect 245838 255212 245844 255264
rect 245896 255252 245902 255264
rect 252830 255252 252836 255264
rect 245896 255224 252836 255252
rect 245896 255212 245902 255224
rect 252830 255212 252836 255224
rect 252888 255212 252894 255264
rect 156690 254600 156696 254652
rect 156748 254640 156754 254652
rect 170582 254640 170588 254652
rect 156748 254612 170588 254640
rect 156748 254600 156754 254612
rect 170582 254600 170588 254612
rect 170640 254600 170646 254652
rect 180334 254600 180340 254652
rect 180392 254640 180398 254652
rect 196802 254640 196808 254652
rect 180392 254612 196808 254640
rect 180392 254600 180398 254612
rect 196802 254600 196808 254612
rect 196860 254600 196866 254652
rect 252830 254600 252836 254652
rect 252888 254640 252894 254652
rect 334618 254640 334624 254652
rect 252888 254612 334624 254640
rect 252888 254600 252894 254612
rect 334618 254600 334624 254612
rect 334676 254600 334682 254652
rect 158254 254532 158260 254584
rect 158312 254572 158318 254584
rect 191098 254572 191104 254584
rect 158312 254544 191104 254572
rect 158312 254532 158318 254544
rect 191098 254532 191104 254544
rect 191156 254532 191162 254584
rect 251082 254532 251088 254584
rect 251140 254572 251146 254584
rect 358170 254572 358176 254584
rect 251140 254544 358176 254572
rect 251140 254532 251146 254544
rect 358170 254532 358176 254544
rect 358228 254532 358234 254584
rect 2774 254192 2780 254244
rect 2832 254232 2838 254244
rect 4798 254232 4804 254244
rect 2832 254204 4804 254232
rect 2832 254192 2838 254204
rect 4798 254192 4804 254204
rect 4856 254192 4862 254244
rect 54938 253920 54944 253972
rect 54996 253960 55002 253972
rect 66622 253960 66628 253972
rect 54996 253932 66628 253960
rect 54996 253920 55002 253932
rect 66622 253920 66628 253932
rect 66680 253920 66686 253972
rect 194410 253920 194416 253972
rect 194468 253960 194474 253972
rect 197354 253960 197360 253972
rect 194468 253932 197360 253960
rect 194468 253920 194474 253932
rect 197354 253920 197360 253932
rect 197412 253920 197418 253972
rect 246022 253852 246028 253904
rect 246080 253892 246086 253904
rect 262398 253892 262404 253904
rect 246080 253864 262404 253892
rect 246080 253852 246086 253864
rect 262398 253852 262404 253864
rect 262456 253892 262462 253904
rect 262674 253892 262680 253904
rect 262456 253864 262680 253892
rect 262456 253852 262462 253864
rect 262674 253852 262680 253864
rect 262732 253852 262738 253904
rect 245930 253784 245936 253836
rect 245988 253824 245994 253836
rect 258258 253824 258264 253836
rect 245988 253796 258264 253824
rect 245988 253784 245994 253796
rect 258258 253784 258264 253796
rect 258316 253824 258322 253836
rect 259270 253824 259276 253836
rect 258316 253796 259276 253824
rect 258316 253784 258322 253796
rect 259270 253784 259276 253796
rect 259328 253784 259334 253836
rect 259270 253240 259276 253292
rect 259328 253280 259334 253292
rect 307754 253280 307760 253292
rect 259328 253252 307760 253280
rect 259328 253240 259334 253252
rect 307754 253240 307760 253252
rect 307812 253280 307818 253292
rect 371326 253280 371332 253292
rect 307812 253252 371332 253280
rect 307812 253240 307818 253252
rect 371326 253240 371332 253252
rect 371384 253240 371390 253292
rect 52270 253172 52276 253224
rect 52328 253212 52334 253224
rect 60182 253212 60188 253224
rect 52328 253184 60188 253212
rect 52328 253172 52334 253184
rect 60182 253172 60188 253184
rect 60240 253172 60246 253224
rect 67542 253172 67548 253224
rect 67600 253212 67606 253224
rect 68370 253212 68376 253224
rect 67600 253184 68376 253212
rect 67600 253172 67606 253184
rect 68370 253172 68376 253184
rect 68428 253172 68434 253224
rect 158714 253172 158720 253224
rect 158772 253212 158778 253224
rect 179414 253212 179420 253224
rect 158772 253184 179420 253212
rect 158772 253172 158778 253184
rect 179414 253172 179420 253184
rect 179472 253172 179478 253224
rect 185578 253172 185584 253224
rect 185636 253212 185642 253224
rect 186130 253212 186136 253224
rect 185636 253184 186136 253212
rect 185636 253172 185642 253184
rect 186130 253172 186136 253184
rect 186188 253212 186194 253224
rect 197354 253212 197360 253224
rect 186188 253184 197360 253212
rect 186188 253172 186194 253184
rect 197354 253172 197360 253184
rect 197412 253172 197418 253224
rect 262674 253172 262680 253224
rect 262732 253212 262738 253224
rect 306374 253212 306380 253224
rect 262732 253184 306380 253212
rect 262732 253172 262738 253184
rect 306374 253172 306380 253184
rect 306432 253212 306438 253224
rect 369946 253212 369952 253224
rect 306432 253184 369952 253212
rect 306432 253172 306438 253184
rect 369946 253172 369952 253184
rect 370004 253172 370010 253224
rect 60182 252560 60188 252612
rect 60240 252600 60246 252612
rect 60550 252600 60556 252612
rect 60240 252572 60556 252600
rect 60240 252560 60246 252572
rect 60550 252560 60556 252572
rect 60608 252600 60614 252612
rect 66806 252600 66812 252612
rect 60608 252572 66812 252600
rect 60608 252560 60614 252572
rect 66806 252560 66812 252572
rect 66864 252560 66870 252612
rect 158714 252560 158720 252612
rect 158772 252600 158778 252612
rect 166350 252600 166356 252612
rect 158772 252572 166356 252600
rect 158772 252560 158778 252572
rect 166350 252560 166356 252572
rect 166408 252560 166414 252612
rect 192938 252560 192944 252612
rect 192996 252600 193002 252612
rect 197354 252600 197360 252612
rect 192996 252572 197360 252600
rect 192996 252560 193002 252572
rect 197354 252560 197360 252572
rect 197412 252560 197418 252612
rect 179414 252492 179420 252544
rect 179472 252532 179478 252544
rect 195790 252532 195796 252544
rect 179472 252504 195796 252532
rect 179472 252492 179478 252504
rect 195790 252492 195796 252504
rect 195848 252492 195854 252544
rect 245930 252492 245936 252544
rect 245988 252532 245994 252544
rect 261018 252532 261024 252544
rect 245988 252504 261024 252532
rect 245988 252492 245994 252504
rect 261018 252492 261024 252504
rect 261076 252532 261082 252544
rect 262122 252532 262128 252544
rect 261076 252504 262128 252532
rect 261076 252492 261082 252504
rect 262122 252492 262128 252504
rect 262180 252492 262186 252544
rect 156782 252424 156788 252476
rect 156840 252464 156846 252476
rect 163774 252464 163780 252476
rect 156840 252436 163780 252464
rect 156840 252424 156846 252436
rect 163774 252424 163780 252436
rect 163832 252424 163838 252476
rect 180334 251812 180340 251864
rect 180392 251852 180398 251864
rect 187050 251852 187056 251864
rect 180392 251824 187056 251852
rect 180392 251812 180398 251824
rect 187050 251812 187056 251824
rect 187108 251812 187114 251864
rect 245930 251812 245936 251864
rect 245988 251852 245994 251864
rect 251358 251852 251364 251864
rect 245988 251824 251364 251852
rect 245988 251812 245994 251824
rect 251358 251812 251364 251824
rect 251416 251852 251422 251864
rect 252370 251852 252376 251864
rect 251416 251824 252376 251852
rect 251416 251812 251422 251824
rect 252370 251812 252376 251824
rect 252428 251812 252434 251864
rect 262122 251812 262128 251864
rect 262180 251852 262186 251864
rect 322198 251852 322204 251864
rect 262180 251824 322204 251852
rect 262180 251812 262186 251824
rect 322198 251812 322204 251824
rect 322256 251812 322262 251864
rect 195790 251608 195796 251660
rect 195848 251648 195854 251660
rect 197354 251648 197360 251660
rect 195848 251620 197360 251648
rect 195848 251608 195854 251620
rect 197354 251608 197360 251620
rect 197412 251608 197418 251660
rect 158898 251200 158904 251252
rect 158956 251240 158962 251252
rect 180334 251240 180340 251252
rect 158956 251212 180340 251240
rect 158956 251200 158962 251212
rect 180334 251200 180340 251212
rect 180392 251240 180398 251252
rect 180702 251240 180708 251252
rect 180392 251212 180708 251240
rect 180392 251200 180398 251212
rect 180702 251200 180708 251212
rect 180760 251200 180766 251252
rect 252370 251200 252376 251252
rect 252428 251240 252434 251252
rect 356698 251240 356704 251252
rect 252428 251212 356704 251240
rect 252428 251200 252434 251212
rect 356698 251200 356704 251212
rect 356756 251200 356762 251252
rect 245838 251132 245844 251184
rect 245896 251172 245902 251184
rect 259454 251172 259460 251184
rect 245896 251144 259460 251172
rect 245896 251132 245902 251144
rect 259454 251132 259460 251144
rect 259512 251172 259518 251184
rect 260742 251172 260748 251184
rect 259512 251144 260748 251172
rect 259512 251132 259518 251144
rect 260742 251132 260748 251144
rect 260800 251132 260806 251184
rect 331950 251132 331956 251184
rect 332008 251172 332014 251184
rect 334710 251172 334716 251184
rect 332008 251144 334716 251172
rect 332008 251132 332014 251144
rect 334710 251132 334716 251144
rect 334768 251132 334774 251184
rect 177298 250928 177304 250980
rect 177356 250968 177362 250980
rect 180058 250968 180064 250980
rect 177356 250940 180064 250968
rect 177356 250928 177362 250940
rect 180058 250928 180064 250940
rect 180116 250928 180122 250980
rect 278222 250520 278228 250572
rect 278280 250560 278286 250572
rect 301038 250560 301044 250572
rect 278280 250532 301044 250560
rect 278280 250520 278286 250532
rect 301038 250520 301044 250532
rect 301096 250520 301102 250572
rect 63402 250452 63408 250504
rect 63460 250492 63466 250504
rect 67726 250492 67732 250504
rect 63460 250464 67732 250492
rect 63460 250452 63466 250464
rect 67726 250452 67732 250464
rect 67784 250452 67790 250504
rect 162486 250452 162492 250504
rect 162544 250492 162550 250504
rect 173250 250492 173256 250504
rect 162544 250464 173256 250492
rect 162544 250452 162550 250464
rect 173250 250452 173256 250464
rect 173308 250452 173314 250504
rect 260742 250452 260748 250504
rect 260800 250492 260806 250504
rect 310606 250492 310612 250504
rect 260800 250464 310612 250492
rect 260800 250452 260806 250464
rect 310606 250452 310612 250464
rect 310664 250492 310670 250504
rect 365806 250492 365812 250504
rect 310664 250464 365812 250492
rect 310664 250452 310670 250464
rect 365806 250452 365812 250464
rect 365864 250452 365870 250504
rect 180150 249908 180156 249960
rect 180208 249948 180214 249960
rect 180208 249920 180794 249948
rect 180208 249908 180214 249920
rect 180766 249880 180794 249920
rect 197354 249880 197360 249892
rect 180766 249852 197360 249880
rect 197354 249840 197360 249852
rect 197412 249840 197418 249892
rect 64506 249772 64512 249824
rect 64564 249812 64570 249824
rect 66806 249812 66812 249824
rect 64564 249784 66812 249812
rect 64564 249772 64570 249784
rect 66806 249772 66812 249784
rect 66864 249772 66870 249824
rect 158714 249772 158720 249824
rect 158772 249812 158778 249824
rect 173434 249812 173440 249824
rect 158772 249784 173440 249812
rect 158772 249772 158778 249784
rect 173434 249772 173440 249784
rect 173492 249772 173498 249824
rect 178770 249772 178776 249824
rect 178828 249812 178834 249824
rect 197446 249812 197452 249824
rect 178828 249784 197452 249812
rect 178828 249772 178834 249784
rect 197446 249772 197452 249784
rect 197504 249772 197510 249824
rect 186222 249704 186228 249756
rect 186280 249744 186286 249756
rect 188522 249744 188528 249756
rect 186280 249716 188528 249744
rect 186280 249704 186286 249716
rect 188522 249704 188528 249716
rect 188580 249704 188586 249756
rect 245930 249704 245936 249756
rect 245988 249744 245994 249756
rect 248690 249744 248696 249756
rect 245988 249716 248696 249744
rect 245988 249704 245994 249716
rect 248690 249704 248696 249716
rect 248748 249704 248754 249756
rect 264238 249092 264244 249144
rect 264296 249132 264302 249144
rect 348418 249132 348424 249144
rect 264296 249104 348424 249132
rect 264296 249092 264302 249104
rect 348418 249092 348424 249104
rect 348476 249092 348482 249144
rect 167730 249024 167736 249076
rect 167788 249064 167794 249076
rect 187602 249064 187608 249076
rect 167788 249036 187608 249064
rect 167788 249024 167794 249036
rect 187602 249024 187608 249036
rect 187660 249024 187666 249076
rect 299382 249024 299388 249076
rect 299440 249064 299446 249076
rect 582834 249064 582840 249076
rect 299440 249036 582840 249064
rect 299440 249024 299446 249036
rect 582834 249024 582840 249036
rect 582892 249024 582898 249076
rect 196710 248684 196716 248736
rect 196768 248724 196774 248736
rect 197814 248724 197820 248736
rect 196768 248696 197820 248724
rect 196768 248684 196774 248696
rect 197814 248684 197820 248696
rect 197872 248684 197878 248736
rect 158806 248412 158812 248464
rect 158864 248452 158870 248464
rect 182818 248452 182824 248464
rect 158864 248424 182824 248452
rect 158864 248412 158870 248424
rect 182818 248412 182824 248424
rect 182876 248412 182882 248464
rect 187602 248412 187608 248464
rect 187660 248452 187666 248464
rect 197354 248452 197360 248464
rect 187660 248424 197360 248452
rect 187660 248412 187666 248424
rect 197354 248412 197360 248424
rect 197412 248412 197418 248464
rect 299382 248344 299388 248396
rect 299440 248384 299446 248396
rect 300210 248384 300216 248396
rect 299440 248356 300216 248384
rect 299440 248344 299446 248356
rect 300210 248344 300216 248356
rect 300268 248344 300274 248396
rect 162394 247732 162400 247784
rect 162452 247772 162458 247784
rect 179414 247772 179420 247784
rect 162452 247744 179420 247772
rect 162452 247732 162458 247744
rect 179414 247732 179420 247744
rect 179472 247732 179478 247784
rect 168466 247664 168472 247716
rect 168524 247704 168530 247716
rect 188706 247704 188712 247716
rect 168524 247676 188712 247704
rect 168524 247664 168530 247676
rect 188706 247664 188712 247676
rect 188764 247664 188770 247716
rect 245654 247664 245660 247716
rect 245712 247704 245718 247716
rect 300210 247704 300216 247716
rect 245712 247676 300216 247704
rect 245712 247664 245718 247676
rect 300210 247664 300216 247676
rect 300268 247664 300274 247716
rect 195606 247120 195612 247172
rect 195664 247160 195670 247172
rect 196710 247160 196716 247172
rect 195664 247132 196716 247160
rect 195664 247120 195670 247132
rect 196710 247120 196716 247132
rect 196768 247120 196774 247172
rect 185578 247052 185584 247104
rect 185636 247092 185642 247104
rect 197354 247092 197360 247104
rect 185636 247064 197360 247092
rect 185636 247052 185642 247064
rect 197354 247052 197360 247064
rect 197412 247052 197418 247104
rect 245930 247052 245936 247104
rect 245988 247092 245994 247104
rect 251266 247092 251272 247104
rect 245988 247064 251272 247092
rect 245988 247052 245994 247064
rect 251266 247052 251272 247064
rect 251324 247092 251330 247104
rect 377398 247092 377404 247104
rect 251324 247064 377404 247092
rect 251324 247052 251330 247064
rect 377398 247052 377404 247064
rect 377456 247052 377462 247104
rect 62022 246984 62028 247036
rect 62080 247024 62086 247036
rect 66806 247024 66812 247036
rect 62080 246996 66812 247024
rect 62080 246984 62086 246996
rect 66806 246984 66812 246996
rect 66864 246984 66870 247036
rect 179414 246304 179420 246356
rect 179472 246344 179478 246356
rect 196710 246344 196716 246356
rect 179472 246316 196716 246344
rect 179472 246304 179478 246316
rect 196710 246304 196716 246316
rect 196768 246304 196774 246356
rect 317230 246304 317236 246356
rect 317288 246344 317294 246356
rect 331214 246344 331220 246356
rect 317288 246316 331220 246344
rect 317288 246304 317294 246316
rect 331214 246304 331220 246316
rect 331272 246304 331278 246356
rect 244550 245692 244556 245744
rect 244608 245732 244614 245744
rect 281534 245732 281540 245744
rect 244608 245704 281540 245732
rect 244608 245692 244614 245704
rect 281534 245692 281540 245704
rect 281592 245732 281598 245744
rect 283558 245732 283564 245744
rect 281592 245704 283564 245732
rect 281592 245692 281598 245704
rect 283558 245692 283564 245704
rect 283616 245692 283622 245744
rect 181438 245624 181444 245676
rect 181496 245664 181502 245676
rect 184290 245664 184296 245676
rect 181496 245636 184296 245664
rect 181496 245624 181502 245636
rect 184290 245624 184296 245636
rect 184348 245624 184354 245676
rect 184750 245624 184756 245676
rect 184808 245664 184814 245676
rect 191834 245664 191840 245676
rect 184808 245636 191840 245664
rect 184808 245624 184814 245636
rect 191834 245624 191840 245636
rect 191892 245664 191898 245676
rect 198826 245664 198832 245676
rect 191892 245636 198832 245664
rect 191892 245624 191898 245636
rect 198826 245624 198832 245636
rect 198884 245624 198890 245676
rect 245838 245624 245844 245676
rect 245896 245664 245902 245676
rect 255406 245664 255412 245676
rect 245896 245636 255412 245664
rect 245896 245624 245902 245636
rect 255406 245624 255412 245636
rect 255464 245624 255470 245676
rect 260098 245624 260104 245676
rect 260156 245664 260162 245676
rect 316034 245664 316040 245676
rect 260156 245636 316040 245664
rect 260156 245624 260162 245636
rect 316034 245624 316040 245636
rect 316092 245664 316098 245676
rect 317230 245664 317236 245676
rect 316092 245636 317236 245664
rect 316092 245624 316098 245636
rect 317230 245624 317236 245636
rect 317288 245624 317294 245676
rect 48222 245556 48228 245608
rect 48280 245596 48286 245608
rect 66806 245596 66812 245608
rect 48280 245568 66812 245596
rect 48280 245556 48286 245568
rect 66806 245556 66812 245568
rect 66864 245556 66870 245608
rect 328362 244944 328368 244996
rect 328420 244984 328426 244996
rect 363138 244984 363144 244996
rect 328420 244956 363144 244984
rect 328420 244944 328426 244956
rect 363138 244944 363144 244956
rect 363196 244944 363202 244996
rect 161566 244876 161572 244928
rect 161624 244916 161630 244928
rect 189810 244916 189816 244928
rect 161624 244888 189816 244916
rect 161624 244876 161630 244888
rect 189810 244876 189816 244888
rect 189868 244876 189874 244928
rect 189902 244876 189908 244928
rect 189960 244916 189966 244928
rect 197722 244916 197728 244928
rect 189960 244888 197728 244916
rect 189960 244876 189966 244888
rect 197722 244876 197728 244888
rect 197780 244876 197786 244928
rect 252370 244876 252376 244928
rect 252428 244916 252434 244928
rect 340230 244916 340236 244928
rect 252428 244888 340236 244916
rect 252428 244876 252434 244888
rect 340230 244876 340236 244888
rect 340288 244876 340294 244928
rect 356790 244876 356796 244928
rect 356848 244916 356854 244928
rect 436278 244916 436284 244928
rect 356848 244888 436284 244916
rect 356848 244876 356854 244888
rect 436278 244876 436284 244888
rect 436336 244876 436342 244928
rect 158714 244264 158720 244316
rect 158772 244304 158778 244316
rect 193858 244304 193864 244316
rect 158772 244276 193864 244304
rect 158772 244264 158778 244276
rect 193858 244264 193864 244276
rect 193916 244264 193922 244316
rect 245930 244264 245936 244316
rect 245988 244304 245994 244316
rect 327166 244304 327172 244316
rect 245988 244276 327172 244304
rect 245988 244264 245994 244276
rect 327166 244264 327172 244276
rect 327224 244304 327230 244316
rect 328362 244304 328368 244316
rect 327224 244276 328368 244304
rect 327224 244264 327230 244276
rect 328362 244264 328368 244276
rect 328420 244264 328426 244316
rect 59170 244196 59176 244248
rect 59228 244236 59234 244248
rect 66806 244236 66812 244248
rect 59228 244208 66812 244236
rect 59228 244196 59234 244208
rect 66806 244196 66812 244208
rect 66864 244196 66870 244248
rect 189810 244196 189816 244248
rect 189868 244236 189874 244248
rect 193030 244236 193036 244248
rect 189868 244208 193036 244236
rect 189868 244196 189874 244208
rect 193030 244196 193036 244208
rect 193088 244236 193094 244248
rect 197354 244236 197360 244248
rect 193088 244208 197360 244236
rect 193088 244196 193094 244208
rect 197354 244196 197360 244208
rect 197412 244196 197418 244248
rect 157978 243516 157984 243568
rect 158036 243556 158042 243568
rect 171318 243556 171324 243568
rect 158036 243528 171324 243556
rect 158036 243516 158042 243528
rect 171318 243516 171324 243528
rect 171376 243556 171382 243568
rect 171686 243556 171692 243568
rect 171376 243528 171692 243556
rect 171376 243516 171382 243528
rect 171686 243516 171692 243528
rect 171744 243516 171750 243568
rect 171778 243516 171784 243568
rect 171836 243556 171842 243568
rect 173342 243556 173348 243568
rect 171836 243528 173348 243556
rect 171836 243516 171842 243528
rect 173342 243516 173348 243528
rect 173400 243516 173406 243568
rect 177482 243516 177488 243568
rect 177540 243556 177546 243568
rect 192662 243556 192668 243568
rect 177540 243528 192668 243556
rect 177540 243516 177546 243528
rect 192662 243516 192668 243528
rect 192720 243516 192726 243568
rect 259270 243516 259276 243568
rect 259328 243556 259334 243568
rect 342898 243556 342904 243568
rect 259328 243528 342904 243556
rect 259328 243516 259334 243528
rect 342898 243516 342904 243528
rect 342956 243516 342962 243568
rect 158714 242904 158720 242956
rect 158772 242944 158778 242956
rect 184290 242944 184296 242956
rect 158772 242916 184296 242944
rect 158772 242904 158778 242916
rect 184290 242904 184296 242916
rect 184348 242904 184354 242956
rect 245838 242904 245844 242956
rect 245896 242944 245902 242956
rect 258258 242944 258264 242956
rect 245896 242916 258264 242944
rect 245896 242904 245902 242916
rect 258258 242904 258264 242916
rect 258316 242944 258322 242956
rect 259270 242944 259276 242956
rect 258316 242916 259276 242944
rect 258316 242904 258322 242916
rect 259270 242904 259276 242916
rect 259328 242904 259334 242956
rect 260742 242904 260748 242956
rect 260800 242944 260806 242956
rect 302970 242944 302976 242956
rect 260800 242916 302976 242944
rect 260800 242904 260806 242916
rect 302970 242904 302976 242916
rect 303028 242904 303034 242956
rect 183094 242196 183100 242208
rect 161446 242168 183100 242196
rect 155310 242020 155316 242072
rect 155368 242060 155374 242072
rect 161446 242060 161474 242168
rect 183094 242156 183100 242168
rect 183152 242156 183158 242208
rect 311986 242156 311992 242208
rect 312044 242196 312050 242208
rect 345658 242196 345664 242208
rect 312044 242168 345664 242196
rect 312044 242156 312050 242168
rect 345658 242156 345664 242168
rect 345716 242156 345722 242208
rect 155368 242032 161474 242060
rect 155368 242020 155374 242032
rect 246390 241544 246396 241596
rect 246448 241584 246454 241596
rect 247218 241584 247224 241596
rect 246448 241556 247224 241584
rect 246448 241544 246454 241556
rect 247218 241544 247224 241556
rect 247276 241584 247282 241596
rect 311986 241584 311992 241596
rect 247276 241556 311992 241584
rect 247276 241544 247282 241556
rect 311986 241544 311992 241556
rect 312044 241544 312050 241596
rect 156966 241476 156972 241528
rect 157024 241516 157030 241528
rect 186222 241516 186228 241528
rect 157024 241488 186228 241516
rect 157024 241476 157030 241488
rect 186222 241476 186228 241488
rect 186280 241516 186286 241528
rect 197354 241516 197360 241528
rect 186280 241488 197360 241516
rect 186280 241476 186286 241488
rect 197354 241476 197360 241488
rect 197412 241476 197418 241528
rect 245746 241476 245752 241528
rect 245804 241516 245810 241528
rect 463694 241516 463700 241528
rect 245804 241488 463700 241516
rect 245804 241476 245810 241488
rect 463694 241476 463700 241488
rect 463752 241476 463758 241528
rect 57790 241408 57796 241460
rect 57848 241448 57854 241460
rect 58618 241448 58624 241460
rect 57848 241420 58624 241448
rect 57848 241408 57854 241420
rect 58618 241408 58624 241420
rect 58676 241408 58682 241460
rect 83320 241448 83326 241460
rect 64846 241420 83326 241448
rect 57698 241340 57704 241392
rect 57756 241380 57762 241392
rect 64846 241380 64874 241420
rect 83320 241408 83326 241420
rect 83378 241408 83384 241460
rect 57756 241352 64874 241380
rect 57756 241340 57762 241352
rect 156368 241340 156374 241392
rect 156426 241380 156432 241392
rect 160186 241380 160192 241392
rect 156426 241352 160192 241380
rect 156426 241340 156432 241352
rect 160186 241340 160192 241352
rect 160244 241340 160250 241392
rect 3510 241068 3516 241120
rect 3568 241108 3574 241120
rect 7558 241108 7564 241120
rect 3568 241080 7564 241108
rect 3568 241068 3574 241080
rect 7558 241068 7564 241080
rect 7616 241068 7622 241120
rect 166258 240796 166264 240848
rect 166316 240836 166322 240848
rect 200114 240836 200120 240848
rect 166316 240808 200120 240836
rect 166316 240796 166322 240808
rect 200114 240796 200120 240808
rect 200172 240796 200178 240848
rect 300118 240796 300124 240848
rect 300176 240836 300182 240848
rect 309870 240836 309876 240848
rect 300176 240808 309876 240836
rect 300176 240796 300182 240808
rect 309870 240796 309876 240808
rect 309928 240796 309934 240848
rect 18598 240728 18604 240780
rect 18656 240768 18662 240780
rect 57790 240768 57796 240780
rect 18656 240740 57796 240768
rect 18656 240728 18662 240740
rect 57790 240728 57796 240740
rect 57848 240728 57854 240780
rect 66070 240728 66076 240780
rect 66128 240768 66134 240780
rect 86218 240768 86224 240780
rect 66128 240740 86224 240768
rect 66128 240728 66134 240740
rect 86218 240728 86224 240740
rect 86276 240728 86282 240780
rect 128814 240728 128820 240780
rect 128872 240768 128878 240780
rect 167822 240768 167828 240780
rect 128872 240740 167828 240768
rect 128872 240728 128878 240740
rect 167822 240728 167828 240740
rect 167880 240728 167886 240780
rect 260190 240728 260196 240780
rect 260248 240768 260254 240780
rect 420178 240768 420184 240780
rect 260248 240740 420184 240768
rect 260248 240728 260254 240740
rect 420178 240728 420184 240740
rect 420236 240728 420242 240780
rect 155494 240388 155500 240440
rect 155552 240428 155558 240440
rect 156690 240428 156696 240440
rect 155552 240400 156696 240428
rect 155552 240388 155558 240400
rect 156690 240388 156696 240400
rect 156748 240388 156754 240440
rect 199654 240388 199660 240440
rect 199712 240428 199718 240440
rect 199712 240400 202828 240428
rect 199712 240388 199718 240400
rect 199562 240320 199568 240372
rect 199620 240360 199626 240372
rect 199620 240332 202368 240360
rect 199620 240320 199626 240332
rect 103606 240184 103612 240236
rect 103664 240224 103670 240236
rect 104802 240224 104808 240236
rect 103664 240196 104808 240224
rect 103664 240184 103670 240196
rect 104802 240184 104808 240196
rect 104860 240224 104866 240236
rect 104860 240196 113174 240224
rect 104860 240184 104866 240196
rect 67726 240116 67732 240168
rect 67784 240156 67790 240168
rect 68462 240156 68468 240168
rect 67784 240128 68468 240156
rect 67784 240116 67790 240128
rect 68462 240116 68468 240128
rect 68520 240116 68526 240168
rect 77294 240116 77300 240168
rect 77352 240156 77358 240168
rect 77846 240156 77852 240168
rect 77352 240128 77852 240156
rect 77352 240116 77358 240128
rect 77846 240116 77852 240128
rect 77904 240116 77910 240168
rect 82906 240116 82912 240168
rect 82964 240156 82970 240168
rect 83734 240156 83740 240168
rect 82964 240128 83740 240156
rect 82964 240116 82970 240128
rect 83734 240116 83740 240128
rect 83792 240116 83798 240168
rect 91094 240116 91100 240168
rect 91152 240156 91158 240168
rect 91830 240156 91836 240168
rect 91152 240128 91836 240156
rect 91152 240116 91158 240128
rect 91830 240116 91836 240128
rect 91888 240116 91894 240168
rect 107654 240116 107660 240168
rect 107712 240156 107718 240168
rect 108574 240156 108580 240168
rect 107712 240128 108580 240156
rect 107712 240116 107718 240128
rect 108574 240116 108580 240128
rect 108632 240116 108638 240168
rect 113146 240156 113174 240196
rect 202340 240168 202368 240332
rect 115198 240156 115204 240168
rect 113146 240128 115204 240156
rect 115198 240116 115204 240128
rect 115256 240116 115262 240168
rect 170582 240116 170588 240168
rect 170640 240156 170646 240168
rect 201218 240156 201224 240168
rect 170640 240128 201224 240156
rect 170640 240116 170646 240128
rect 201218 240116 201224 240128
rect 201276 240116 201282 240168
rect 202322 240116 202328 240168
rect 202380 240116 202386 240168
rect 202800 240156 202828 240400
rect 244090 240292 244096 240304
rect 229066 240264 244096 240292
rect 229066 240224 229094 240264
rect 244090 240252 244096 240264
rect 244148 240252 244154 240304
rect 226812 240196 229094 240224
rect 226812 240168 226840 240196
rect 243906 240184 243912 240236
rect 243964 240224 243970 240236
rect 289906 240224 289912 240236
rect 243964 240196 289912 240224
rect 243964 240184 243970 240196
rect 289906 240184 289912 240196
rect 289964 240224 289970 240236
rect 298830 240224 298836 240236
rect 289964 240196 298836 240224
rect 289964 240184 289970 240196
rect 298830 240184 298836 240196
rect 298888 240184 298894 240236
rect 203978 240156 203984 240168
rect 202800 240128 203984 240156
rect 203978 240116 203984 240128
rect 204036 240116 204042 240168
rect 208394 240116 208400 240168
rect 208452 240156 208458 240168
rect 225046 240156 225052 240168
rect 208452 240128 225052 240156
rect 208452 240116 208458 240128
rect 225046 240116 225052 240128
rect 225104 240116 225110 240168
rect 226794 240116 226800 240168
rect 226852 240116 226858 240168
rect 228358 240116 228364 240168
rect 228416 240156 228422 240168
rect 231026 240156 231032 240168
rect 228416 240128 231032 240156
rect 228416 240116 228422 240128
rect 231026 240116 231032 240128
rect 231084 240116 231090 240168
rect 241882 240116 241888 240168
rect 241940 240156 241946 240168
rect 247126 240156 247132 240168
rect 241940 240128 247132 240156
rect 241940 240116 241946 240128
rect 247126 240116 247132 240128
rect 247184 240116 247190 240168
rect 69566 240048 69572 240100
rect 69624 240088 69630 240100
rect 72510 240088 72516 240100
rect 69624 240060 72516 240088
rect 69624 240048 69630 240060
rect 72510 240048 72516 240060
rect 72568 240048 72574 240100
rect 75178 240048 75184 240100
rect 75236 240088 75242 240100
rect 75914 240088 75920 240100
rect 75236 240060 75920 240088
rect 75236 240048 75242 240060
rect 75914 240048 75920 240060
rect 75972 240048 75978 240100
rect 82722 240048 82728 240100
rect 82780 240088 82786 240100
rect 83550 240088 83556 240100
rect 82780 240060 83556 240088
rect 82780 240048 82786 240060
rect 83550 240048 83556 240060
rect 83608 240048 83614 240100
rect 85114 240048 85120 240100
rect 85172 240088 85178 240100
rect 92566 240088 92572 240100
rect 85172 240060 92572 240088
rect 85172 240048 85178 240060
rect 92566 240048 92572 240060
rect 92624 240048 92630 240100
rect 117866 240048 117872 240100
rect 117924 240088 117930 240100
rect 118602 240088 118608 240100
rect 117924 240060 118608 240088
rect 117924 240048 117930 240060
rect 118602 240048 118608 240060
rect 118660 240048 118666 240100
rect 119338 240048 119344 240100
rect 119396 240088 119402 240100
rect 119982 240088 119988 240100
rect 119396 240060 119988 240088
rect 119396 240048 119402 240060
rect 119982 240048 119988 240060
rect 120040 240048 120046 240100
rect 128630 240048 128636 240100
rect 128688 240088 128694 240100
rect 129642 240088 129648 240100
rect 128688 240060 129648 240088
rect 128688 240048 128694 240060
rect 129642 240048 129648 240060
rect 129700 240048 129706 240100
rect 131850 240048 131856 240100
rect 131908 240088 131914 240100
rect 132402 240088 132408 240100
rect 131908 240060 132408 240088
rect 131908 240048 131914 240060
rect 132402 240048 132408 240060
rect 132460 240048 132466 240100
rect 133322 240048 133328 240100
rect 133380 240088 133386 240100
rect 133782 240088 133788 240100
rect 133380 240060 133788 240088
rect 133380 240048 133386 240060
rect 133782 240048 133788 240060
rect 133840 240048 133846 240100
rect 135346 240048 135352 240100
rect 135404 240088 135410 240100
rect 136542 240088 136548 240100
rect 135404 240060 136548 240088
rect 135404 240048 135410 240060
rect 136542 240048 136548 240060
rect 136600 240048 136606 240100
rect 138474 240048 138480 240100
rect 138532 240088 138538 240100
rect 139302 240088 139308 240100
rect 138532 240060 139308 240088
rect 138532 240048 138538 240060
rect 139302 240048 139308 240060
rect 139360 240048 139366 240100
rect 142890 240048 142896 240100
rect 142948 240088 142954 240100
rect 143350 240088 143356 240100
rect 142948 240060 143356 240088
rect 142948 240048 142954 240060
rect 143350 240048 143356 240060
rect 143408 240048 143414 240100
rect 145650 240048 145656 240100
rect 145708 240088 145714 240100
rect 146110 240088 146116 240100
rect 145708 240060 146116 240088
rect 145708 240048 145714 240060
rect 146110 240048 146116 240060
rect 146168 240048 146174 240100
rect 153470 240048 153476 240100
rect 153528 240088 153534 240100
rect 154482 240088 154488 240100
rect 153528 240060 154488 240088
rect 153528 240048 153534 240060
rect 154482 240048 154488 240060
rect 154540 240048 154546 240100
rect 228726 240048 228732 240100
rect 228784 240088 228790 240100
rect 243906 240088 243912 240100
rect 228784 240060 243912 240088
rect 228784 240048 228790 240060
rect 243906 240048 243912 240060
rect 243964 240048 243970 240100
rect 67450 239980 67456 240032
rect 67508 240020 67514 240032
rect 69750 240020 69756 240032
rect 67508 239992 69756 240020
rect 67508 239980 67514 239992
rect 69750 239980 69756 239992
rect 69808 239980 69814 240032
rect 113634 239980 113640 240032
rect 113692 240020 113698 240032
rect 118510 240020 118516 240032
rect 113692 239992 118516 240020
rect 113692 239980 113698 239992
rect 118510 239980 118516 239992
rect 118568 239980 118574 240032
rect 142246 239980 142252 240032
rect 142304 240020 142310 240032
rect 142982 240020 142988 240032
rect 142304 239992 142988 240020
rect 142304 239980 142310 239992
rect 142982 239980 142988 239992
rect 143040 239980 143046 240032
rect 237374 239980 237380 240032
rect 237432 240020 237438 240032
rect 238110 240020 238116 240032
rect 237432 239992 238116 240020
rect 237432 239980 237438 239992
rect 238110 239980 238116 239992
rect 238168 240020 238174 240032
rect 244550 240020 244556 240032
rect 238168 239992 244556 240020
rect 238168 239980 238174 239992
rect 244550 239980 244556 239992
rect 244608 239980 244614 240032
rect 82170 239776 82176 239828
rect 82228 239816 82234 239828
rect 82722 239816 82728 239828
rect 82228 239788 82728 239816
rect 82228 239776 82234 239788
rect 82722 239776 82728 239788
rect 82780 239776 82786 239828
rect 70302 239436 70308 239488
rect 70360 239476 70366 239488
rect 97258 239476 97264 239488
rect 70360 239448 97264 239476
rect 70360 239436 70366 239448
rect 97258 239436 97264 239448
rect 97316 239436 97322 239488
rect 97442 239436 97448 239488
rect 97500 239476 97506 239488
rect 97500 239448 103514 239476
rect 97500 239436 97506 239448
rect 88794 239368 88800 239420
rect 88852 239408 88858 239420
rect 89530 239408 89536 239420
rect 88852 239380 89536 239408
rect 88852 239368 88858 239380
rect 89530 239368 89536 239380
rect 89588 239368 89594 239420
rect 101950 239368 101956 239420
rect 102008 239408 102014 239420
rect 102686 239408 102692 239420
rect 102008 239380 102692 239408
rect 102008 239368 102014 239380
rect 102686 239368 102692 239380
rect 102744 239368 102750 239420
rect 103486 239408 103514 239448
rect 122282 239436 122288 239488
rect 122340 239476 122346 239488
rect 220814 239476 220820 239488
rect 122340 239448 220820 239476
rect 122340 239436 122346 239448
rect 220814 239436 220820 239448
rect 220872 239436 220878 239488
rect 305086 239436 305092 239488
rect 305144 239476 305150 239488
rect 322934 239476 322940 239488
rect 305144 239448 322940 239476
rect 305144 239436 305150 239448
rect 322934 239436 322940 239448
rect 322992 239436 322998 239488
rect 214190 239408 214196 239420
rect 103486 239380 214196 239408
rect 214190 239368 214196 239380
rect 214248 239368 214254 239420
rect 260742 239368 260748 239420
rect 260800 239408 260806 239420
rect 273898 239408 273904 239420
rect 260800 239380 273904 239408
rect 260800 239368 260806 239380
rect 273898 239368 273904 239380
rect 273956 239368 273962 239420
rect 313918 239368 313924 239420
rect 313976 239408 313982 239420
rect 345658 239408 345664 239420
rect 313976 239380 345664 239408
rect 313976 239368 313982 239380
rect 345658 239368 345664 239380
rect 345716 239368 345722 239420
rect 116578 239300 116584 239352
rect 116636 239340 116642 239352
rect 117130 239340 117136 239352
rect 116636 239312 117136 239340
rect 116636 239300 116642 239312
rect 117130 239300 117136 239312
rect 117188 239300 117194 239352
rect 120810 239300 120816 239352
rect 120868 239340 120874 239352
rect 121362 239340 121368 239352
rect 120868 239312 121368 239340
rect 120868 239300 120874 239312
rect 121362 239300 121368 239312
rect 121420 239300 121426 239352
rect 143534 239300 143540 239352
rect 143592 239340 143598 239352
rect 144270 239340 144276 239352
rect 143592 239312 144276 239340
rect 143592 239300 143598 239312
rect 144270 239300 144276 239312
rect 144328 239300 144334 239352
rect 80698 239232 80704 239284
rect 80756 239272 80762 239284
rect 81342 239272 81348 239284
rect 80756 239244 81348 239272
rect 80756 239232 80762 239244
rect 81342 239232 81348 239244
rect 81400 239232 81406 239284
rect 105538 239232 105544 239284
rect 105596 239272 105602 239284
rect 106182 239272 106188 239284
rect 105596 239244 106188 239272
rect 105596 239232 105602 239244
rect 106182 239232 106188 239244
rect 106240 239232 106246 239284
rect 131206 239232 131212 239284
rect 131264 239272 131270 239284
rect 131942 239272 131948 239284
rect 131264 239244 131948 239272
rect 131264 239232 131270 239244
rect 131942 239232 131948 239244
rect 132000 239232 132006 239284
rect 138014 239232 138020 239284
rect 138072 239272 138078 239284
rect 138566 239272 138572 239284
rect 138072 239244 138572 239272
rect 138072 239232 138078 239244
rect 138566 239232 138572 239244
rect 138624 239232 138630 239284
rect 104066 239164 104072 239216
rect 104124 239204 104130 239216
rect 104802 239204 104808 239216
rect 104124 239176 104808 239204
rect 104124 239164 104130 239176
rect 104802 239164 104808 239176
rect 104860 239164 104866 239216
rect 219434 238756 219440 238808
rect 219492 238796 219498 238808
rect 238018 238796 238024 238808
rect 219492 238768 238024 238796
rect 219492 238756 219498 238768
rect 238018 238756 238024 238768
rect 238076 238756 238082 238808
rect 73154 238688 73160 238740
rect 73212 238728 73218 238740
rect 202598 238728 202604 238740
rect 73212 238700 202604 238728
rect 73212 238688 73218 238700
rect 202598 238688 202604 238700
rect 202656 238688 202662 238740
rect 240318 238688 240324 238740
rect 240376 238728 240382 238740
rect 252462 238728 252468 238740
rect 240376 238700 252468 238728
rect 240376 238688 240382 238700
rect 252462 238688 252468 238700
rect 252520 238688 252526 238740
rect 55030 238620 55036 238672
rect 55088 238660 55094 238672
rect 75178 238660 75184 238672
rect 55088 238632 75184 238660
rect 55088 238620 55094 238632
rect 75178 238620 75184 238632
rect 75236 238620 75242 238672
rect 118510 238620 118516 238672
rect 118568 238660 118574 238672
rect 222286 238660 222292 238672
rect 118568 238632 222292 238660
rect 118568 238620 118574 238632
rect 222286 238620 222292 238632
rect 222344 238620 222350 238672
rect 242066 238620 242072 238672
rect 242124 238660 242130 238672
rect 252646 238660 252652 238672
rect 242124 238632 252652 238660
rect 242124 238620 242130 238632
rect 252646 238620 252652 238632
rect 252704 238620 252710 238672
rect 224862 238076 224868 238128
rect 224920 238116 224926 238128
rect 227530 238116 227536 238128
rect 224920 238088 227536 238116
rect 224920 238076 224926 238088
rect 227530 238076 227536 238088
rect 227588 238076 227594 238128
rect 252462 238076 252468 238128
rect 252520 238116 252526 238128
rect 262858 238116 262864 238128
rect 252520 238088 262864 238116
rect 252520 238076 252526 238088
rect 262858 238076 262864 238088
rect 262916 238076 262922 238128
rect 260098 238008 260104 238060
rect 260156 238048 260162 238060
rect 280798 238048 280804 238060
rect 260156 238020 280804 238048
rect 260156 238008 260162 238020
rect 280798 238008 280804 238020
rect 280856 238008 280862 238060
rect 295242 238008 295248 238060
rect 295300 238048 295306 238060
rect 384298 238048 384304 238060
rect 295300 238020 384304 238048
rect 295300 238008 295306 238020
rect 384298 238008 384304 238020
rect 384356 238008 384362 238060
rect 223390 237804 223396 237856
rect 223448 237844 223454 237856
rect 229370 237844 229376 237856
rect 223448 237816 229376 237844
rect 223448 237804 223454 237816
rect 229370 237804 229376 237816
rect 229428 237804 229434 237856
rect 229830 237668 229836 237720
rect 229888 237708 229894 237720
rect 236822 237708 236828 237720
rect 229888 237680 236828 237708
rect 229888 237668 229894 237680
rect 236822 237668 236828 237680
rect 236880 237668 236886 237720
rect 240042 237464 240048 237516
rect 240100 237504 240106 237516
rect 242710 237504 242716 237516
rect 240100 237476 242716 237504
rect 240100 237464 240106 237476
rect 242710 237464 242716 237476
rect 242768 237464 242774 237516
rect 202138 237396 202144 237448
rect 202196 237436 202202 237448
rect 202598 237436 202604 237448
rect 202196 237408 202604 237436
rect 202196 237396 202202 237408
rect 202598 237396 202604 237408
rect 202656 237396 202662 237448
rect 202874 237396 202880 237448
rect 202932 237436 202938 237448
rect 204990 237436 204996 237448
rect 202932 237408 204996 237436
rect 202932 237396 202938 237408
rect 204990 237396 204996 237408
rect 205048 237396 205054 237448
rect 207106 237396 207112 237448
rect 207164 237436 207170 237448
rect 207934 237436 207940 237448
rect 207164 237408 207940 237436
rect 207164 237396 207170 237408
rect 207934 237396 207940 237408
rect 207992 237396 207998 237448
rect 209682 237396 209688 237448
rect 209740 237436 209746 237448
rect 210326 237436 210332 237448
rect 209740 237408 210332 237436
rect 209740 237396 209746 237408
rect 210326 237396 210332 237408
rect 210384 237396 210390 237448
rect 230198 237396 230204 237448
rect 230256 237436 230262 237448
rect 232498 237436 232504 237448
rect 230256 237408 232504 237436
rect 230256 237396 230262 237408
rect 232498 237396 232504 237408
rect 232556 237396 232562 237448
rect 239214 237396 239220 237448
rect 239272 237436 239278 237448
rect 240962 237436 240968 237448
rect 239272 237408 240968 237436
rect 239272 237396 239278 237408
rect 240962 237396 240968 237408
rect 241020 237396 241026 237448
rect 125594 237328 125600 237380
rect 125652 237368 125658 237380
rect 181530 237368 181536 237380
rect 125652 237340 181536 237368
rect 125652 237328 125658 237340
rect 181530 237328 181536 237340
rect 181588 237368 181594 237380
rect 182082 237368 182088 237380
rect 181588 237340 182088 237368
rect 181588 237328 181594 237340
rect 182082 237328 182088 237340
rect 182140 237328 182146 237380
rect 200114 237328 200120 237380
rect 200172 237368 200178 237380
rect 223758 237368 223764 237380
rect 200172 237340 223764 237368
rect 200172 237328 200178 237340
rect 223758 237328 223764 237340
rect 223816 237328 223822 237380
rect 241238 237328 241244 237380
rect 241296 237368 241302 237380
rect 287698 237368 287704 237380
rect 241296 237340 287704 237368
rect 241296 237328 241302 237340
rect 287698 237328 287704 237340
rect 287756 237328 287762 237380
rect 149054 237260 149060 237312
rect 149112 237300 149118 237312
rect 162210 237300 162216 237312
rect 149112 237272 162216 237300
rect 149112 237260 149118 237272
rect 162210 237260 162216 237272
rect 162268 237260 162274 237312
rect 196802 237260 196808 237312
rect 196860 237300 196866 237312
rect 202782 237300 202788 237312
rect 196860 237272 202788 237300
rect 196860 237260 196866 237272
rect 202782 237260 202788 237272
rect 202840 237260 202846 237312
rect 194318 236716 194324 236768
rect 194376 236756 194382 236768
rect 199378 236756 199384 236768
rect 194376 236728 199384 236756
rect 194376 236716 194382 236728
rect 199378 236716 199384 236728
rect 199436 236716 199442 236768
rect 229094 236716 229100 236768
rect 229152 236756 229158 236768
rect 242250 236756 242256 236768
rect 229152 236728 242256 236756
rect 229152 236716 229158 236728
rect 242250 236716 242256 236728
rect 242308 236716 242314 236768
rect 187418 236648 187424 236700
rect 187476 236688 187482 236700
rect 195238 236688 195244 236700
rect 187476 236660 195244 236688
rect 187476 236648 187482 236660
rect 195238 236648 195244 236660
rect 195296 236648 195302 236700
rect 199930 236648 199936 236700
rect 199988 236688 199994 236700
rect 200758 236688 200764 236700
rect 199988 236660 200764 236688
rect 199988 236648 199994 236660
rect 200758 236648 200764 236660
rect 200816 236648 200822 236700
rect 208302 236648 208308 236700
rect 208360 236688 208366 236700
rect 239490 236688 239496 236700
rect 208360 236660 239496 236688
rect 208360 236648 208366 236660
rect 239490 236648 239496 236660
rect 239548 236648 239554 236700
rect 260926 236648 260932 236700
rect 260984 236688 260990 236700
rect 410518 236688 410524 236700
rect 260984 236660 410524 236688
rect 260984 236648 260990 236660
rect 410518 236648 410524 236660
rect 410576 236648 410582 236700
rect 4798 235968 4804 236020
rect 4856 236008 4862 236020
rect 93854 236008 93860 236020
rect 4856 235980 93860 236008
rect 4856 235968 4862 235980
rect 93854 235968 93860 235980
rect 93912 236008 93918 236020
rect 94498 236008 94504 236020
rect 93912 235980 94504 236008
rect 93912 235968 93918 235980
rect 94498 235968 94504 235980
rect 94556 235968 94562 236020
rect 240778 235968 240784 236020
rect 240836 236008 240842 236020
rect 241238 236008 241244 236020
rect 240836 235980 241244 236008
rect 240836 235968 240842 235980
rect 241238 235968 241244 235980
rect 241296 235968 241302 236020
rect 61746 235900 61752 235952
rect 61804 235940 61810 235952
rect 130102 235940 130108 235952
rect 61804 235912 130108 235940
rect 61804 235900 61810 235912
rect 130102 235900 130108 235912
rect 130160 235900 130166 235952
rect 196710 235900 196716 235952
rect 196768 235940 196774 235952
rect 220262 235940 220268 235952
rect 196768 235912 220268 235940
rect 196768 235900 196774 235912
rect 220262 235900 220268 235912
rect 220320 235900 220326 235952
rect 232038 235900 232044 235952
rect 232096 235940 232102 235952
rect 268378 235940 268384 235952
rect 232096 235912 268384 235940
rect 232096 235900 232102 235912
rect 268378 235900 268384 235912
rect 268436 235900 268442 235952
rect 50890 235832 50896 235884
rect 50948 235872 50954 235884
rect 77386 235872 77392 235884
rect 50948 235844 77392 235872
rect 50948 235832 50954 235844
rect 77386 235832 77392 235844
rect 77444 235832 77450 235884
rect 114646 235832 114652 235884
rect 114704 235872 114710 235884
rect 152458 235872 152464 235884
rect 114704 235844 152464 235872
rect 114704 235832 114710 235844
rect 152458 235832 152464 235844
rect 152516 235872 152522 235884
rect 152734 235872 152740 235884
rect 152516 235844 152740 235872
rect 152516 235832 152522 235844
rect 152734 235832 152740 235844
rect 152792 235832 152798 235884
rect 185670 235832 185676 235884
rect 185728 235872 185734 235884
rect 206830 235872 206836 235884
rect 185728 235844 206836 235872
rect 185728 235832 185734 235844
rect 206830 235832 206836 235844
rect 206888 235832 206894 235884
rect 152366 235696 152372 235748
rect 152424 235736 152430 235748
rect 155954 235736 155960 235748
rect 152424 235708 155960 235736
rect 152424 235696 152430 235708
rect 155954 235696 155960 235708
rect 156012 235696 156018 235748
rect 222930 235288 222936 235340
rect 222988 235328 222994 235340
rect 232038 235328 232044 235340
rect 222988 235300 232044 235328
rect 222988 235288 222994 235300
rect 232038 235288 232044 235300
rect 232096 235288 232102 235340
rect 131206 235220 131212 235272
rect 131264 235260 131270 235272
rect 184750 235260 184756 235272
rect 131264 235232 184756 235260
rect 131264 235220 131270 235232
rect 184750 235220 184756 235232
rect 184808 235260 184814 235272
rect 185578 235260 185584 235272
rect 184808 235232 185584 235260
rect 184808 235220 184814 235232
rect 185578 235220 185584 235232
rect 185636 235220 185642 235272
rect 205634 235220 205640 235272
rect 205692 235260 205698 235272
rect 224218 235260 224224 235272
rect 205692 235232 224224 235260
rect 205692 235220 205698 235232
rect 224218 235220 224224 235232
rect 224276 235220 224282 235272
rect 168190 234648 168196 234660
rect 167012 234620 168196 234648
rect 57606 234540 57612 234592
rect 57664 234580 57670 234592
rect 128722 234580 128728 234592
rect 57664 234552 128728 234580
rect 57664 234540 57670 234552
rect 128722 234540 128728 234552
rect 128780 234540 128786 234592
rect 150434 234540 150440 234592
rect 150492 234580 150498 234592
rect 167012 234580 167040 234620
rect 168190 234608 168196 234620
rect 168248 234648 168254 234660
rect 174538 234648 174544 234660
rect 168248 234620 174544 234648
rect 168248 234608 168254 234620
rect 174538 234608 174544 234620
rect 174596 234608 174602 234660
rect 186958 234608 186964 234660
rect 187016 234648 187022 234660
rect 188430 234648 188436 234660
rect 187016 234620 188436 234648
rect 187016 234608 187022 234620
rect 188430 234608 188436 234620
rect 188488 234608 188494 234660
rect 206370 234608 206376 234660
rect 206428 234648 206434 234660
rect 206830 234648 206836 234660
rect 206428 234620 206836 234648
rect 206428 234608 206434 234620
rect 206830 234608 206836 234620
rect 206888 234608 206894 234660
rect 231578 234608 231584 234660
rect 231636 234648 231642 234660
rect 234062 234648 234068 234660
rect 231636 234620 234068 234648
rect 231636 234608 231642 234620
rect 234062 234608 234068 234620
rect 234120 234608 234126 234660
rect 240870 234608 240876 234660
rect 240928 234648 240934 234660
rect 243262 234648 243268 234660
rect 240928 234620 243268 234648
rect 240928 234608 240934 234620
rect 243262 234608 243268 234620
rect 243320 234608 243326 234660
rect 150492 234552 167040 234580
rect 150492 234540 150498 234552
rect 152090 234472 152096 234524
rect 152148 234512 152154 234524
rect 155678 234512 155684 234524
rect 152148 234484 155684 234512
rect 152148 234472 152154 234484
rect 155678 234472 155684 234484
rect 155736 234472 155742 234524
rect 191466 234132 191472 234184
rect 191524 234172 191530 234184
rect 192570 234172 192576 234184
rect 191524 234144 192576 234172
rect 191524 234132 191530 234144
rect 192570 234132 192576 234144
rect 192628 234132 192634 234184
rect 242250 233996 242256 234048
rect 242308 234036 242314 234048
rect 265618 234036 265624 234048
rect 242308 234008 265624 234036
rect 242308 233996 242314 234008
rect 265618 233996 265624 234008
rect 265676 233996 265682 234048
rect 133138 233928 133144 233980
rect 133196 233968 133202 233980
rect 152918 233968 152924 233980
rect 133196 233940 152924 233968
rect 133196 233928 133202 233940
rect 152918 233928 152924 233940
rect 152976 233928 152982 233980
rect 176194 233928 176200 233980
rect 176252 233968 176258 233980
rect 187050 233968 187056 233980
rect 176252 233940 187056 233968
rect 176252 233928 176258 233940
rect 187050 233928 187056 233940
rect 187108 233928 187114 233980
rect 195238 233928 195244 233980
rect 195296 233968 195302 233980
rect 210602 233968 210608 233980
rect 195296 233940 210608 233968
rect 195296 233928 195302 233940
rect 210602 233928 210608 233940
rect 210660 233928 210666 233980
rect 215294 233928 215300 233980
rect 215352 233968 215358 233980
rect 247218 233968 247224 233980
rect 215352 233940 247224 233968
rect 215352 233928 215358 233940
rect 247218 233928 247224 233940
rect 247276 233928 247282 233980
rect 111886 233860 111892 233912
rect 111944 233900 111950 233912
rect 139578 233900 139584 233912
rect 111944 233872 139584 233900
rect 111944 233860 111950 233872
rect 139578 233860 139584 233872
rect 139636 233860 139642 233912
rect 155218 233860 155224 233912
rect 155276 233900 155282 233912
rect 176654 233900 176660 233912
rect 155276 233872 176660 233900
rect 155276 233860 155282 233872
rect 176654 233860 176660 233872
rect 176712 233860 176718 233912
rect 184290 233860 184296 233912
rect 184348 233900 184354 233912
rect 235994 233900 236000 233912
rect 184348 233872 236000 233900
rect 184348 233860 184354 233872
rect 235994 233860 236000 233872
rect 236052 233860 236058 233912
rect 256694 233860 256700 233912
rect 256752 233900 256758 233912
rect 322290 233900 322296 233912
rect 256752 233872 322296 233900
rect 256752 233860 256758 233872
rect 322290 233860 322296 233872
rect 322348 233860 322354 233912
rect 280798 233288 280804 233300
rect 271616 233260 280804 233288
rect 14458 233180 14464 233232
rect 14516 233220 14522 233232
rect 92658 233220 92664 233232
rect 14516 233192 92664 233220
rect 14516 233180 14522 233192
rect 92658 233180 92664 233192
rect 92716 233180 92722 233232
rect 143626 233180 143632 233232
rect 143684 233220 143690 233232
rect 156874 233220 156880 233232
rect 143684 233192 156880 233220
rect 143684 233180 143690 233192
rect 156874 233180 156880 233192
rect 156932 233180 156938 233232
rect 192938 233180 192944 233232
rect 192996 233220 193002 233232
rect 270494 233220 270500 233232
rect 192996 233192 270500 233220
rect 192996 233180 193002 233192
rect 270494 233180 270500 233192
rect 270552 233220 270558 233232
rect 271616 233220 271644 233260
rect 280798 233248 280804 233260
rect 280856 233248 280862 233300
rect 270552 233192 271644 233220
rect 270552 233180 270558 233192
rect 155862 233112 155868 233164
rect 155920 233152 155926 233164
rect 158254 233152 158260 233164
rect 155920 233124 158260 233152
rect 155920 233112 155926 233124
rect 158254 233112 158260 233124
rect 158312 233112 158318 233164
rect 190454 233112 190460 233164
rect 190512 233152 190518 233164
rect 205358 233152 205364 233164
rect 190512 233124 205364 233152
rect 190512 233112 190518 233124
rect 205358 233112 205364 233124
rect 205416 233112 205422 233164
rect 211798 233112 211804 233164
rect 211856 233152 211862 233164
rect 212810 233152 212816 233164
rect 211856 233124 212816 233152
rect 211856 233112 211862 233124
rect 212810 233112 212816 233124
rect 212868 233112 212874 233164
rect 235994 233112 236000 233164
rect 236052 233152 236058 233164
rect 236638 233152 236644 233164
rect 236052 233124 236644 233152
rect 236052 233112 236058 233124
rect 236638 233112 236644 233124
rect 236696 233152 236702 233164
rect 244458 233152 244464 233164
rect 236696 233124 244464 233152
rect 236696 233112 236702 233124
rect 244458 233112 244464 233124
rect 244516 233112 244522 233164
rect 92658 232704 92664 232756
rect 92716 232744 92722 232756
rect 93118 232744 93124 232756
rect 92716 232716 93124 232744
rect 92716 232704 92722 232716
rect 93118 232704 93124 232716
rect 93176 232704 93182 232756
rect 156598 232704 156604 232756
rect 156656 232744 156662 232756
rect 159174 232744 159180 232756
rect 156656 232716 159180 232744
rect 156656 232704 156662 232716
rect 159174 232704 159180 232716
rect 159232 232704 159238 232756
rect 140866 232568 140872 232620
rect 140924 232608 140930 232620
rect 155862 232608 155868 232620
rect 140924 232580 155868 232608
rect 140924 232568 140930 232580
rect 155862 232568 155868 232580
rect 155920 232568 155926 232620
rect 44082 232500 44088 232552
rect 44140 232540 44146 232552
rect 143534 232540 143540 232552
rect 44140 232512 143540 232540
rect 44140 232500 44146 232512
rect 143534 232500 143540 232512
rect 143592 232500 143598 232552
rect 157334 232500 157340 232552
rect 157392 232540 157398 232552
rect 187418 232540 187424 232552
rect 157392 232512 187424 232540
rect 157392 232500 157398 232512
rect 187418 232500 187424 232512
rect 187476 232540 187482 232552
rect 191098 232540 191104 232552
rect 187476 232512 191104 232540
rect 187476 232500 187482 232512
rect 191098 232500 191104 232512
rect 191156 232500 191162 232552
rect 216030 232500 216036 232552
rect 216088 232540 216094 232552
rect 227714 232540 227720 232552
rect 216088 232512 227720 232540
rect 216088 232500 216094 232512
rect 227714 232500 227720 232512
rect 227772 232500 227778 232552
rect 282178 232500 282184 232552
rect 282236 232540 282242 232552
rect 465074 232540 465080 232552
rect 282236 232512 465080 232540
rect 282236 232500 282242 232512
rect 465074 232500 465080 232512
rect 465132 232500 465138 232552
rect 158714 231820 158720 231872
rect 158772 231860 158778 231872
rect 184290 231860 184296 231872
rect 158772 231832 184296 231860
rect 158772 231820 158778 231832
rect 184290 231820 184296 231832
rect 184348 231820 184354 231872
rect 69750 231752 69756 231804
rect 69808 231792 69814 231804
rect 156966 231792 156972 231804
rect 69808 231764 156972 231792
rect 69808 231752 69814 231764
rect 156966 231752 156972 231764
rect 157024 231752 157030 231804
rect 124306 231684 124312 231736
rect 124364 231724 124370 231736
rect 198734 231724 198740 231736
rect 124364 231696 198740 231724
rect 124364 231684 124370 231696
rect 198734 231684 198740 231696
rect 198792 231684 198798 231736
rect 205634 231548 205640 231600
rect 205692 231588 205698 231600
rect 206462 231588 206468 231600
rect 205692 231560 206468 231588
rect 205692 231548 205698 231560
rect 206462 231548 206468 231560
rect 206520 231548 206526 231600
rect 198734 231140 198740 231192
rect 198792 231180 198798 231192
rect 199838 231180 199844 231192
rect 198792 231152 199844 231180
rect 198792 231140 198798 231152
rect 199838 231140 199844 231152
rect 199896 231180 199902 231192
rect 230474 231180 230480 231192
rect 199896 231152 230480 231180
rect 199896 231140 199902 231152
rect 230474 231140 230480 231152
rect 230532 231140 230538 231192
rect 204070 231072 204076 231124
rect 204128 231112 204134 231124
rect 224218 231112 224224 231124
rect 204128 231084 224224 231112
rect 204128 231072 204134 231084
rect 224218 231072 224224 231084
rect 224276 231072 224282 231124
rect 228174 231072 228180 231124
rect 228232 231112 228238 231124
rect 398926 231112 398932 231124
rect 228232 231084 398932 231112
rect 228232 231072 228238 231084
rect 398926 231072 398932 231084
rect 398984 231072 398990 231124
rect 208394 230936 208400 230988
rect 208452 230976 208458 230988
rect 209222 230976 209228 230988
rect 208452 230948 209228 230976
rect 208452 230936 208458 230948
rect 209222 230936 209228 230948
rect 209280 230936 209286 230988
rect 270402 230500 270408 230512
rect 270315 230472 270408 230500
rect 270402 230460 270408 230472
rect 270460 230500 270466 230512
rect 282178 230500 282184 230512
rect 270460 230472 282184 230500
rect 270460 230460 270466 230472
rect 282178 230460 282184 230472
rect 282236 230460 282242 230512
rect 143350 230392 143356 230444
rect 143408 230432 143414 230444
rect 231578 230432 231584 230444
rect 143408 230404 231584 230432
rect 143408 230392 143414 230404
rect 231578 230392 231584 230404
rect 231636 230392 231642 230444
rect 139302 230324 139308 230376
rect 139360 230364 139366 230376
rect 165430 230364 165436 230376
rect 139360 230336 165436 230364
rect 139360 230324 139366 230336
rect 165430 230324 165436 230336
rect 165488 230324 165494 230376
rect 166350 230324 166356 230376
rect 166408 230364 166414 230376
rect 195238 230364 195244 230376
rect 166408 230336 195244 230364
rect 166408 230324 166414 230336
rect 195238 230324 195244 230336
rect 195296 230324 195302 230376
rect 202322 230324 202328 230376
rect 202380 230364 202386 230376
rect 207566 230364 207572 230376
rect 202380 230336 207572 230364
rect 202380 230324 202386 230336
rect 207566 230324 207572 230336
rect 207624 230324 207630 230376
rect 222286 230324 222292 230376
rect 222344 230364 222350 230376
rect 270420 230364 270448 230460
rect 222344 230336 270448 230364
rect 222344 230324 222350 230336
rect 83642 229780 83648 229832
rect 83700 229820 83706 229832
rect 141418 229820 141424 229832
rect 83700 229792 141424 229820
rect 83700 229780 83706 229792
rect 141418 229780 141424 229792
rect 141476 229780 141482 229832
rect 64690 229712 64696 229764
rect 64748 229752 64754 229764
rect 137922 229752 137928 229764
rect 64748 229724 137928 229752
rect 64748 229712 64754 229724
rect 137922 229712 137928 229724
rect 137980 229712 137986 229764
rect 165430 229576 165436 229628
rect 165488 229616 165494 229628
rect 166258 229616 166264 229628
rect 165488 229588 166264 229616
rect 165488 229576 165494 229588
rect 166258 229576 166264 229588
rect 166316 229576 166322 229628
rect 243538 229100 243544 229152
rect 243596 229140 243602 229152
rect 248506 229140 248512 229152
rect 243596 229112 248512 229140
rect 243596 229100 243602 229112
rect 248506 229100 248512 229112
rect 248564 229100 248570 229152
rect 117314 229032 117320 229084
rect 117372 229072 117378 229084
rect 224310 229072 224316 229084
rect 117372 229044 224316 229072
rect 117372 229032 117378 229044
rect 224310 229032 224316 229044
rect 224368 229032 224374 229084
rect 94498 228964 94504 229016
rect 94556 229004 94562 229016
rect 174630 229004 174636 229016
rect 94556 228976 174636 229004
rect 94556 228964 94562 228976
rect 174630 228964 174636 228976
rect 174688 228964 174694 229016
rect 175918 228964 175924 229016
rect 175976 229004 175982 229016
rect 242894 229004 242900 229016
rect 175976 228976 242900 229004
rect 175976 228964 175982 228976
rect 242894 228964 242900 228976
rect 242952 228964 242958 229016
rect 242894 228556 242900 228608
rect 242952 228596 242958 228608
rect 243906 228596 243912 228608
rect 242952 228568 243912 228596
rect 242952 228556 242958 228568
rect 243906 228556 243912 228568
rect 243964 228556 243970 228608
rect 327074 228352 327080 228404
rect 327132 228392 327138 228404
rect 403066 228392 403072 228404
rect 327132 228364 403072 228392
rect 327132 228352 327138 228364
rect 403066 228352 403072 228364
rect 403124 228352 403130 228404
rect 242802 227740 242808 227792
rect 242860 227780 242866 227792
rect 258258 227780 258264 227792
rect 242860 227752 258264 227780
rect 242860 227740 242866 227752
rect 258258 227740 258264 227752
rect 258316 227780 258322 227792
rect 258718 227780 258724 227792
rect 258316 227752 258724 227780
rect 258316 227740 258322 227752
rect 258718 227740 258724 227752
rect 258776 227740 258782 227792
rect 137922 227672 137928 227724
rect 137980 227712 137986 227724
rect 173158 227712 173164 227724
rect 137980 227684 173164 227712
rect 137980 227672 137986 227684
rect 173158 227672 173164 227684
rect 173216 227672 173222 227724
rect 181714 227672 181720 227724
rect 181772 227712 181778 227724
rect 222838 227712 222844 227724
rect 181772 227684 222844 227712
rect 181772 227672 181778 227684
rect 222838 227672 222844 227684
rect 222896 227672 222902 227724
rect 224310 227060 224316 227112
rect 224368 227100 224374 227112
rect 240686 227100 240692 227112
rect 224368 227072 240692 227100
rect 224368 227060 224374 227072
rect 240686 227060 240692 227072
rect 240744 227060 240750 227112
rect 54938 226992 54944 227044
rect 54996 227032 55002 227044
rect 194318 227032 194324 227044
rect 54996 227004 194324 227032
rect 54996 226992 55002 227004
rect 194318 226992 194324 227004
rect 194376 226992 194382 227044
rect 217134 226992 217140 227044
rect 217192 227032 217198 227044
rect 226334 227032 226340 227044
rect 217192 227004 226340 227032
rect 217192 226992 217198 227004
rect 226334 226992 226340 227004
rect 226392 226992 226398 227044
rect 239490 226992 239496 227044
rect 239548 227032 239554 227044
rect 298278 227032 298284 227044
rect 239548 227004 298284 227032
rect 239548 226992 239554 227004
rect 298278 226992 298284 227004
rect 298336 226992 298342 227044
rect 204898 226312 204904 226364
rect 204956 226352 204962 226364
rect 209682 226352 209688 226364
rect 204956 226324 209688 226352
rect 204956 226312 204962 226324
rect 209682 226312 209688 226324
rect 209740 226312 209746 226364
rect 71774 226244 71780 226296
rect 71832 226284 71838 226296
rect 158070 226284 158076 226296
rect 71832 226256 158076 226284
rect 71832 226244 71838 226256
rect 158070 226244 158076 226256
rect 158128 226244 158134 226296
rect 187050 226244 187056 226296
rect 187108 226284 187114 226296
rect 213638 226284 213644 226296
rect 187108 226256 213644 226284
rect 187108 226244 187114 226256
rect 213638 226244 213644 226256
rect 213696 226244 213702 226296
rect 139394 226176 139400 226228
rect 139452 226216 139458 226228
rect 222930 226216 222936 226228
rect 139452 226188 222936 226216
rect 139452 226176 139458 226188
rect 222930 226176 222936 226188
rect 222988 226176 222994 226228
rect 240686 225632 240692 225684
rect 240744 225672 240750 225684
rect 284478 225672 284484 225684
rect 240744 225644 284484 225672
rect 240744 225632 240750 225644
rect 284478 225632 284484 225644
rect 284536 225632 284542 225684
rect 68278 225564 68284 225616
rect 68336 225604 68342 225616
rect 104158 225604 104164 225616
rect 68336 225576 104164 225604
rect 68336 225564 68342 225576
rect 104158 225564 104164 225576
rect 104216 225564 104222 225616
rect 219894 225564 219900 225616
rect 219952 225604 219958 225616
rect 220354 225604 220360 225616
rect 219952 225576 220360 225604
rect 219952 225564 219958 225576
rect 220354 225564 220360 225576
rect 220412 225604 220418 225616
rect 266998 225604 267004 225616
rect 220412 225576 267004 225604
rect 220412 225564 220418 225576
rect 266998 225564 267004 225576
rect 267056 225564 267062 225616
rect 292482 225564 292488 225616
rect 292540 225604 292546 225616
rect 307110 225604 307116 225616
rect 292540 225576 307116 225604
rect 292540 225564 292546 225576
rect 307110 225564 307116 225576
rect 307168 225564 307174 225616
rect 213178 225428 213184 225480
rect 213236 225468 213242 225480
rect 213638 225468 213644 225480
rect 213236 225440 213644 225468
rect 213236 225428 213242 225440
rect 213638 225428 213644 225440
rect 213696 225428 213702 225480
rect 284478 224952 284484 225004
rect 284536 224992 284542 225004
rect 285674 224992 285680 225004
rect 284536 224964 285680 224992
rect 284536 224952 284542 224964
rect 285674 224952 285680 224964
rect 285732 224952 285738 225004
rect 111702 224884 111708 224936
rect 111760 224924 111766 224936
rect 192938 224924 192944 224936
rect 111760 224896 192944 224924
rect 111760 224884 111766 224896
rect 192938 224884 192944 224896
rect 192996 224884 193002 224936
rect 221458 224884 221464 224936
rect 221516 224924 221522 224936
rect 276014 224924 276020 224936
rect 221516 224896 276020 224924
rect 221516 224884 221522 224896
rect 276014 224884 276020 224896
rect 276072 224884 276078 224936
rect 246298 224612 246304 224664
rect 246356 224652 246362 224664
rect 247218 224652 247224 224664
rect 246356 224624 247224 224652
rect 246356 224612 246362 224624
rect 247218 224612 247224 224624
rect 247276 224612 247282 224664
rect 95326 224204 95332 224256
rect 95384 224244 95390 224256
rect 95384 224216 142154 224244
rect 95384 224204 95390 224216
rect 142126 224176 142154 224216
rect 157334 224204 157340 224256
rect 157392 224244 157398 224256
rect 178034 224244 178040 224256
rect 157392 224216 178040 224244
rect 157392 224204 157398 224216
rect 178034 224204 178040 224216
rect 178092 224204 178098 224256
rect 193950 224204 193956 224256
rect 194008 224244 194014 224256
rect 223482 224244 223488 224256
rect 194008 224216 223488 224244
rect 194008 224204 194014 224216
rect 223482 224204 223488 224216
rect 223540 224204 223546 224256
rect 276014 224204 276020 224256
rect 276072 224244 276078 224256
rect 285674 224244 285680 224256
rect 276072 224216 285680 224244
rect 276072 224204 276078 224216
rect 285674 224204 285680 224216
rect 285732 224204 285738 224256
rect 158162 224176 158168 224188
rect 142126 224148 158168 224176
rect 158162 224136 158168 224148
rect 158220 224136 158226 224188
rect 79962 223524 79968 223576
rect 80020 223564 80026 223576
rect 211890 223564 211896 223576
rect 80020 223536 211896 223564
rect 80020 223524 80026 223536
rect 211890 223524 211896 223536
rect 211948 223524 211954 223576
rect 124214 222844 124220 222896
rect 124272 222884 124278 222896
rect 186314 222884 186320 222896
rect 124272 222856 186320 222884
rect 124272 222844 124278 222856
rect 186314 222844 186320 222856
rect 186372 222844 186378 222896
rect 201494 222844 201500 222896
rect 201552 222884 201558 222896
rect 302326 222884 302332 222896
rect 201552 222856 302332 222884
rect 201552 222844 201558 222856
rect 302326 222844 302332 222856
rect 302384 222884 302390 222896
rect 338758 222884 338764 222896
rect 302384 222856 338764 222884
rect 302384 222844 302390 222856
rect 338758 222844 338764 222856
rect 338816 222844 338822 222896
rect 65978 222096 65984 222148
rect 66036 222136 66042 222148
rect 159634 222136 159640 222148
rect 66036 222108 159640 222136
rect 66036 222096 66042 222108
rect 159634 222096 159640 222108
rect 159692 222096 159698 222148
rect 194318 222096 194324 222148
rect 194376 222136 194382 222148
rect 213270 222136 213276 222148
rect 194376 222108 213276 222136
rect 194376 222096 194382 222108
rect 213270 222096 213276 222108
rect 213328 222096 213334 222148
rect 223482 222096 223488 222148
rect 223540 222136 223546 222148
rect 248598 222136 248604 222148
rect 223540 222108 248604 222136
rect 223540 222096 223546 222108
rect 248598 222096 248604 222108
rect 248656 222096 248662 222148
rect 106274 222028 106280 222080
rect 106332 222068 106338 222080
rect 171778 222068 171784 222080
rect 106332 222040 171784 222068
rect 106332 222028 106338 222040
rect 171778 222028 171784 222040
rect 171836 222028 171842 222080
rect 203058 221824 203064 221876
rect 203116 221864 203122 221876
rect 203610 221864 203616 221876
rect 203116 221836 203616 221864
rect 203116 221824 203122 221836
rect 203610 221824 203616 221836
rect 203668 221824 203674 221876
rect 166994 221416 167000 221468
rect 167052 221456 167058 221468
rect 167730 221456 167736 221468
rect 167052 221428 167736 221456
rect 167052 221416 167058 221428
rect 167730 221416 167736 221428
rect 167788 221456 167794 221468
rect 203058 221456 203064 221468
rect 167788 221428 203064 221456
rect 167788 221416 167794 221428
rect 203058 221416 203064 221428
rect 203116 221416 203122 221468
rect 208394 221416 208400 221468
rect 208452 221456 208458 221468
rect 228726 221456 228732 221468
rect 208452 221428 228732 221456
rect 208452 221416 208458 221428
rect 228726 221416 228732 221428
rect 228784 221416 228790 221468
rect 260742 221416 260748 221468
rect 260800 221456 260806 221468
rect 387058 221456 387064 221468
rect 260800 221428 387064 221456
rect 260800 221416 260806 221428
rect 387058 221416 387064 221428
rect 387116 221416 387122 221468
rect 104894 220736 104900 220788
rect 104952 220776 104958 220788
rect 180242 220776 180248 220788
rect 104952 220748 180248 220776
rect 104952 220736 104958 220748
rect 180242 220736 180248 220748
rect 180300 220736 180306 220788
rect 186314 220736 186320 220788
rect 186372 220776 186378 220788
rect 220078 220776 220084 220788
rect 186372 220748 220084 220776
rect 186372 220736 186378 220748
rect 220078 220736 220084 220748
rect 220136 220736 220142 220788
rect 227254 220736 227260 220788
rect 227312 220776 227318 220788
rect 260742 220776 260748 220788
rect 227312 220748 260748 220776
rect 227312 220736 227318 220748
rect 260742 220736 260748 220748
rect 260800 220736 260806 220788
rect 195698 220668 195704 220720
rect 195756 220708 195762 220720
rect 199470 220708 199476 220720
rect 195756 220680 199476 220708
rect 195756 220668 195762 220680
rect 199470 220668 199476 220680
rect 199528 220668 199534 220720
rect 127250 220056 127256 220108
rect 127308 220096 127314 220108
rect 194410 220096 194416 220108
rect 127308 220068 194416 220096
rect 127308 220056 127314 220068
rect 194410 220056 194416 220068
rect 194468 220056 194474 220108
rect 260742 220056 260748 220108
rect 260800 220096 260806 220108
rect 276934 220096 276940 220108
rect 260800 220068 276940 220096
rect 260800 220056 260806 220068
rect 276934 220056 276940 220068
rect 276992 220056 276998 220108
rect 278130 220056 278136 220108
rect 278188 220096 278194 220108
rect 294046 220096 294052 220108
rect 278188 220068 294052 220096
rect 278188 220056 278194 220068
rect 294046 220056 294052 220068
rect 294104 220056 294110 220108
rect 200022 219444 200028 219496
rect 200080 219484 200086 219496
rect 201494 219484 201500 219496
rect 200080 219456 201500 219484
rect 200080 219444 200086 219456
rect 201494 219444 201500 219456
rect 201552 219484 201558 219496
rect 217318 219484 217324 219496
rect 201552 219456 217324 219484
rect 201552 219444 201558 219456
rect 217318 219444 217324 219456
rect 217376 219444 217382 219496
rect 221366 219376 221372 219428
rect 221424 219416 221430 219428
rect 258074 219416 258080 219428
rect 221424 219388 258080 219416
rect 221424 219376 221430 219388
rect 258074 219376 258080 219388
rect 258132 219416 258138 219428
rect 259270 219416 259276 219428
rect 258132 219388 259276 219416
rect 258132 219376 258138 219388
rect 259270 219376 259276 219388
rect 259328 219376 259334 219428
rect 194410 219308 194416 219360
rect 194468 219348 194474 219360
rect 227254 219348 227260 219360
rect 194468 219320 227260 219348
rect 194468 219308 194474 219320
rect 227254 219308 227260 219320
rect 227312 219308 227318 219360
rect 236454 219308 236460 219360
rect 236512 219348 236518 219360
rect 269758 219348 269764 219360
rect 236512 219320 269764 219348
rect 236512 219308 236518 219320
rect 269758 219308 269764 219320
rect 269816 219308 269822 219360
rect 106182 218764 106188 218816
rect 106240 218804 106246 218816
rect 133138 218804 133144 218816
rect 106240 218776 133144 218804
rect 106240 218764 106246 218776
rect 133138 218764 133144 218776
rect 133196 218764 133202 218816
rect 136634 218764 136640 218816
rect 136692 218804 136698 218816
rect 182266 218804 182272 218816
rect 136692 218776 182272 218804
rect 136692 218764 136698 218776
rect 182266 218764 182272 218776
rect 182324 218764 182330 218816
rect 269758 218764 269764 218816
rect 269816 218804 269822 218816
rect 304258 218804 304264 218816
rect 269816 218776 304264 218804
rect 269816 218764 269822 218776
rect 304258 218764 304264 218776
rect 304316 218764 304322 218816
rect 82722 218696 82728 218748
rect 82780 218736 82786 218748
rect 142798 218736 142804 218748
rect 82780 218708 142804 218736
rect 82780 218696 82786 218708
rect 142798 218696 142804 218708
rect 142856 218696 142862 218748
rect 207658 218696 207664 218748
rect 207716 218736 207722 218748
rect 222102 218736 222108 218748
rect 207716 218708 222108 218736
rect 207716 218696 207722 218708
rect 222102 218696 222108 218708
rect 222160 218696 222166 218748
rect 259270 218696 259276 218748
rect 259328 218736 259334 218748
rect 414014 218736 414020 218748
rect 259328 218708 414020 218736
rect 259328 218696 259334 218708
rect 414014 218696 414020 218708
rect 414072 218696 414078 218748
rect 143442 218016 143448 218068
rect 143500 218056 143506 218068
rect 195238 218056 195244 218068
rect 143500 218028 195244 218056
rect 143500 218016 143506 218028
rect 195238 218016 195244 218028
rect 195296 218016 195302 218068
rect 126974 217948 126980 218000
rect 127032 217988 127038 218000
rect 208394 217988 208400 218000
rect 127032 217960 208400 217988
rect 127032 217948 127038 217960
rect 208394 217948 208400 217960
rect 208452 217948 208458 218000
rect 184474 217880 184480 217932
rect 184532 217920 184538 217932
rect 225230 217920 225236 217932
rect 184532 217892 225236 217920
rect 184532 217880 184538 217892
rect 225230 217880 225236 217892
rect 225288 217880 225294 217932
rect 83550 217268 83556 217320
rect 83608 217308 83614 217320
rect 83608 217280 161474 217308
rect 83608 217268 83614 217280
rect 161446 217172 161474 217280
rect 177850 217172 177856 217184
rect 161446 217144 177856 217172
rect 177850 217132 177856 217144
rect 177908 217172 177914 217184
rect 178770 217172 178776 217184
rect 177908 217144 178776 217172
rect 177908 217132 177914 217144
rect 178770 217132 178776 217144
rect 178828 217132 178834 217184
rect 234982 216656 234988 216708
rect 235040 216696 235046 216708
rect 394050 216696 394056 216708
rect 235040 216668 394056 216696
rect 235040 216656 235046 216668
rect 394050 216656 394056 216668
rect 394108 216656 394114 216708
rect 107654 216588 107660 216640
rect 107712 216628 107718 216640
rect 220354 216628 220360 216640
rect 107712 216600 220360 216628
rect 107712 216588 107718 216600
rect 220354 216588 220360 216600
rect 220412 216588 220418 216640
rect 132402 216520 132408 216572
rect 132460 216560 132466 216572
rect 181438 216560 181444 216572
rect 132460 216532 181444 216560
rect 132460 216520 132466 216532
rect 181438 216520 181444 216532
rect 181496 216520 181502 216572
rect 220262 215976 220268 216028
rect 220320 216016 220326 216028
rect 233326 216016 233332 216028
rect 220320 215988 233332 216016
rect 220320 215976 220326 215988
rect 233326 215976 233332 215988
rect 233384 215976 233390 216028
rect 232590 215908 232596 215960
rect 232648 215948 232654 215960
rect 321554 215948 321560 215960
rect 232648 215920 321560 215948
rect 232648 215908 232654 215920
rect 321554 215908 321560 215920
rect 321612 215908 321618 215960
rect 3326 215228 3332 215280
rect 3384 215268 3390 215280
rect 35158 215268 35164 215280
rect 3384 215240 35164 215268
rect 3384 215228 3390 215240
rect 35158 215228 35164 215240
rect 35216 215228 35222 215280
rect 87138 215228 87144 215280
rect 87196 215268 87202 215280
rect 186958 215268 186964 215280
rect 87196 215240 186964 215268
rect 87196 215228 87202 215240
rect 186958 215228 186964 215240
rect 187016 215228 187022 215280
rect 219342 215228 219348 215280
rect 219400 215268 219406 215280
rect 267734 215268 267740 215280
rect 219400 215240 267740 215268
rect 219400 215228 219406 215240
rect 267734 215228 267740 215240
rect 267792 215268 267798 215280
rect 269022 215268 269028 215280
rect 267792 215240 269028 215268
rect 267792 215228 267798 215240
rect 269022 215228 269028 215240
rect 269080 215228 269086 215280
rect 201126 214616 201132 214668
rect 201184 214656 201190 214668
rect 206462 214656 206468 214668
rect 201184 214628 206468 214656
rect 201184 214616 201190 214628
rect 206462 214616 206468 214628
rect 206520 214616 206526 214668
rect 182266 214548 182272 214600
rect 182324 214588 182330 214600
rect 223482 214588 223488 214600
rect 182324 214560 223488 214588
rect 182324 214548 182330 214560
rect 223482 214548 223488 214560
rect 223540 214548 223546 214600
rect 269022 214548 269028 214600
rect 269080 214588 269086 214600
rect 287238 214588 287244 214600
rect 269080 214560 287244 214588
rect 269080 214548 269086 214560
rect 287238 214548 287244 214560
rect 287296 214548 287302 214600
rect 317322 214548 317328 214600
rect 317380 214588 317386 214600
rect 447226 214588 447232 214600
rect 317380 214560 447232 214588
rect 317380 214548 317386 214560
rect 447226 214548 447232 214560
rect 447284 214548 447290 214600
rect 97258 213868 97264 213920
rect 97316 213908 97322 213920
rect 202230 213908 202236 213920
rect 97316 213880 202236 213908
rect 97316 213868 97322 213880
rect 202230 213868 202236 213880
rect 202288 213868 202294 213920
rect 223482 213868 223488 213920
rect 223540 213908 223546 213920
rect 245654 213908 245660 213920
rect 223540 213880 245660 213908
rect 223540 213868 223546 213880
rect 245654 213868 245660 213880
rect 245712 213868 245718 213920
rect 118694 213800 118700 213852
rect 118752 213840 118758 213852
rect 169018 213840 169024 213852
rect 118752 213812 169024 213840
rect 118752 213800 118758 213812
rect 169018 213800 169024 213812
rect 169076 213800 169082 213852
rect 205634 213256 205640 213308
rect 205692 213296 205698 213308
rect 215294 213296 215300 213308
rect 205692 213268 215300 213296
rect 205692 213256 205698 213268
rect 215294 213256 215300 213268
rect 215352 213256 215358 213308
rect 202414 213188 202420 213240
rect 202472 213228 202478 213240
rect 229738 213228 229744 213240
rect 202472 213200 229744 213228
rect 202472 213188 202478 213200
rect 229738 213188 229744 213200
rect 229796 213188 229802 213240
rect 249702 212508 249708 212560
rect 249760 212548 249766 212560
rect 456794 212548 456800 212560
rect 249760 212520 456800 212548
rect 249760 212508 249766 212520
rect 456794 212508 456800 212520
rect 456852 212508 456858 212560
rect 124122 212440 124128 212492
rect 124180 212480 124186 212492
rect 225138 212480 225144 212492
rect 124180 212452 225144 212480
rect 124180 212440 124186 212452
rect 225138 212440 225144 212452
rect 225196 212480 225202 212492
rect 225598 212480 225604 212492
rect 225196 212452 225604 212480
rect 225196 212440 225202 212452
rect 225598 212440 225604 212452
rect 225656 212440 225662 212492
rect 215110 212372 215116 212424
rect 215168 212412 215174 212424
rect 215662 212412 215668 212424
rect 215168 212384 215668 212412
rect 215168 212372 215174 212384
rect 215662 212372 215668 212384
rect 215720 212372 215726 212424
rect 263594 211828 263600 211880
rect 263652 211868 263658 211880
rect 283558 211868 283564 211880
rect 263652 211840 283564 211868
rect 263652 211828 263658 211840
rect 283558 211828 283564 211840
rect 283616 211828 283622 211880
rect 70394 211760 70400 211812
rect 70452 211800 70458 211812
rect 215110 211800 215116 211812
rect 70452 211772 215116 211800
rect 70452 211760 70458 211772
rect 215110 211760 215116 211772
rect 215168 211760 215174 211812
rect 233510 211760 233516 211812
rect 233568 211800 233574 211812
rect 380158 211800 380164 211812
rect 233568 211772 380164 211800
rect 233568 211760 233574 211772
rect 380158 211760 380164 211772
rect 380216 211760 380222 211812
rect 77294 211080 77300 211132
rect 77352 211120 77358 211132
rect 215294 211120 215300 211132
rect 77352 211092 215300 211120
rect 77352 211080 77358 211092
rect 215294 211080 215300 211092
rect 215352 211080 215358 211132
rect 158162 211012 158168 211064
rect 158220 211052 158226 211064
rect 248690 211052 248696 211064
rect 158220 211024 248696 211052
rect 158220 211012 158226 211024
rect 248690 211012 248696 211024
rect 248748 211012 248754 211064
rect 238846 209788 238852 209840
rect 238904 209828 238910 209840
rect 239766 209828 239772 209840
rect 238904 209800 239772 209828
rect 238904 209788 238910 209800
rect 239766 209788 239772 209800
rect 239824 209828 239830 209840
rect 309962 209828 309968 209840
rect 239824 209800 309968 209828
rect 239824 209788 239830 209800
rect 309962 209788 309968 209800
rect 310020 209788 310026 209840
rect 104158 209720 104164 209772
rect 104216 209760 104222 209772
rect 226334 209760 226340 209772
rect 104216 209732 226340 209760
rect 104216 209720 104222 209732
rect 226334 209720 226340 209732
rect 226392 209720 226398 209772
rect 90910 209652 90916 209704
rect 90968 209692 90974 209704
rect 189718 209692 189724 209704
rect 90968 209664 189724 209692
rect 90968 209652 90974 209664
rect 189718 209652 189724 209664
rect 189776 209652 189782 209704
rect 204714 209040 204720 209092
rect 204772 209080 204778 209092
rect 234430 209080 234436 209092
rect 204772 209052 234436 209080
rect 204772 209040 204778 209052
rect 234430 209040 234436 209052
rect 234488 209040 234494 209092
rect 267826 209040 267832 209092
rect 267884 209080 267890 209092
rect 445846 209080 445852 209092
rect 267884 209052 445852 209080
rect 267884 209040 267890 209052
rect 445846 209040 445852 209052
rect 445904 209040 445910 209092
rect 89714 208972 89720 209024
rect 89772 209012 89778 209024
rect 90910 209012 90916 209024
rect 89772 208984 90916 209012
rect 89772 208972 89778 208984
rect 90910 208972 90916 208984
rect 90968 208972 90974 209024
rect 226334 208360 226340 208412
rect 226392 208400 226398 208412
rect 227070 208400 227076 208412
rect 226392 208372 227076 208400
rect 226392 208360 226398 208372
rect 227070 208360 227076 208372
rect 227128 208360 227134 208412
rect 48130 208292 48136 208344
rect 48188 208332 48194 208344
rect 240226 208332 240232 208344
rect 48188 208304 240232 208332
rect 48188 208292 48194 208304
rect 240226 208292 240232 208304
rect 240284 208332 240290 208344
rect 240870 208332 240876 208344
rect 240284 208304 240876 208332
rect 240284 208292 240290 208304
rect 240870 208292 240876 208304
rect 240928 208292 240934 208344
rect 100662 208224 100668 208276
rect 100720 208264 100726 208276
rect 181622 208264 181628 208276
rect 100720 208236 181628 208264
rect 100720 208224 100726 208236
rect 181622 208224 181628 208236
rect 181680 208224 181686 208276
rect 99374 207748 99380 207800
rect 99432 207788 99438 207800
rect 100662 207788 100668 207800
rect 99432 207760 100668 207788
rect 99432 207748 99438 207760
rect 100662 207748 100668 207760
rect 100720 207748 100726 207800
rect 262858 207680 262864 207732
rect 262916 207720 262922 207732
rect 278130 207720 278136 207732
rect 262916 207692 278136 207720
rect 262916 207680 262922 207692
rect 278130 207680 278136 207692
rect 278188 207680 278194 207732
rect 229738 207612 229744 207664
rect 229796 207652 229802 207664
rect 272610 207652 272616 207664
rect 229796 207624 272616 207652
rect 229796 207612 229802 207624
rect 272610 207612 272616 207624
rect 272668 207612 272674 207664
rect 181622 207000 181628 207052
rect 181680 207040 181686 207052
rect 228358 207040 228364 207052
rect 181680 207012 228364 207040
rect 181680 207000 181686 207012
rect 228358 207000 228364 207012
rect 228416 207000 228422 207052
rect 114462 206932 114468 206984
rect 114520 206972 114526 206984
rect 247218 206972 247224 206984
rect 114520 206944 247224 206972
rect 114520 206932 114526 206944
rect 247218 206932 247224 206944
rect 247276 206932 247282 206984
rect 133782 206864 133788 206916
rect 133840 206904 133846 206916
rect 227714 206904 227720 206916
rect 133840 206876 227720 206904
rect 133840 206864 133846 206876
rect 227714 206864 227720 206876
rect 227772 206904 227778 206916
rect 247126 206904 247132 206916
rect 227772 206876 247132 206904
rect 227772 206864 227778 206876
rect 247126 206864 247132 206876
rect 247184 206864 247190 206916
rect 86954 205572 86960 205624
rect 87012 205612 87018 205624
rect 214466 205612 214472 205624
rect 87012 205584 214472 205612
rect 87012 205572 87018 205584
rect 214466 205572 214472 205584
rect 214524 205572 214530 205624
rect 142798 205504 142804 205556
rect 142856 205544 142862 205556
rect 249886 205544 249892 205556
rect 142856 205516 249892 205544
rect 142856 205504 142862 205516
rect 249886 205504 249892 205516
rect 249944 205504 249950 205556
rect 51074 204892 51080 204944
rect 51132 204932 51138 204944
rect 137278 204932 137284 204944
rect 51132 204904 137284 204932
rect 51132 204892 51138 204904
rect 137278 204892 137284 204904
rect 137336 204892 137342 204944
rect 225690 204892 225696 204944
rect 225748 204932 225754 204944
rect 284386 204932 284392 204944
rect 225748 204904 284392 204932
rect 225748 204892 225754 204904
rect 284386 204892 284392 204904
rect 284444 204892 284450 204944
rect 214466 204280 214472 204332
rect 214524 204320 214530 204332
rect 224310 204320 224316 204332
rect 214524 204292 224316 204320
rect 214524 204280 214530 204292
rect 224310 204280 224316 204292
rect 224368 204280 224374 204332
rect 91094 204212 91100 204264
rect 91152 204252 91158 204264
rect 212442 204252 212448 204264
rect 91152 204224 212448 204252
rect 91152 204212 91158 204224
rect 212442 204212 212448 204224
rect 212500 204212 212506 204264
rect 100754 204144 100760 204196
rect 100812 204184 100818 204196
rect 212810 204184 212816 204196
rect 100812 204156 212816 204184
rect 100812 204144 100818 204156
rect 212810 204144 212816 204156
rect 212868 204184 212874 204196
rect 213822 204184 213828 204196
rect 212868 204156 213828 204184
rect 212868 204144 212874 204156
rect 213822 204144 213828 204156
rect 213880 204144 213886 204196
rect 213822 203600 213828 203652
rect 213880 203640 213886 203652
rect 238754 203640 238760 203652
rect 213880 203612 238760 203640
rect 213880 203600 213886 203612
rect 238754 203600 238760 203612
rect 238812 203600 238818 203652
rect 212442 203532 212448 203584
rect 212500 203572 212506 203584
rect 272518 203572 272524 203584
rect 212500 203544 272524 203572
rect 212500 203532 212506 203544
rect 272518 203532 272524 203544
rect 272576 203532 272582 203584
rect 3050 202784 3056 202836
rect 3108 202824 3114 202836
rect 51074 202824 51080 202836
rect 3108 202796 51080 202824
rect 3108 202784 3114 202796
rect 51074 202784 51080 202796
rect 51132 202784 51138 202836
rect 59262 202784 59268 202836
rect 59320 202824 59326 202836
rect 211798 202824 211804 202836
rect 59320 202796 211804 202824
rect 59320 202784 59326 202796
rect 211798 202784 211804 202796
rect 211856 202824 211862 202836
rect 212166 202824 212172 202836
rect 211856 202796 212172 202824
rect 211856 202784 211862 202796
rect 212166 202784 212172 202796
rect 212224 202784 212230 202836
rect 72510 202716 72516 202768
rect 72568 202756 72574 202768
rect 181622 202756 181628 202768
rect 72568 202728 181628 202756
rect 72568 202716 72574 202728
rect 181622 202716 181628 202728
rect 181680 202716 181686 202768
rect 213178 202172 213184 202224
rect 213236 202212 213242 202224
rect 237374 202212 237380 202224
rect 213236 202184 237380 202212
rect 213236 202172 213242 202184
rect 237374 202172 237380 202184
rect 237432 202172 237438 202224
rect 197170 202104 197176 202156
rect 197228 202144 197234 202156
rect 370590 202144 370596 202156
rect 197228 202116 370596 202144
rect 197228 202104 197234 202116
rect 370590 202104 370596 202116
rect 370648 202104 370654 202156
rect 288710 201492 288716 201544
rect 288768 201532 288774 201544
rect 437474 201532 437480 201544
rect 288768 201504 437480 201532
rect 288768 201492 288774 201504
rect 437474 201492 437480 201504
rect 437532 201492 437538 201544
rect 67634 200812 67640 200864
rect 67692 200852 67698 200864
rect 169754 200852 169760 200864
rect 67692 200824 169760 200852
rect 67692 200812 67698 200824
rect 169754 200812 169760 200824
rect 169812 200812 169818 200864
rect 193122 200812 193128 200864
rect 193180 200852 193186 200864
rect 203610 200852 203616 200864
rect 193180 200824 203616 200852
rect 193180 200812 193186 200824
rect 203610 200812 203616 200824
rect 203668 200812 203674 200864
rect 126882 200744 126888 200796
rect 126940 200784 126946 200796
rect 234614 200784 234620 200796
rect 126940 200756 234620 200784
rect 126940 200744 126946 200756
rect 234614 200744 234620 200756
rect 234672 200784 234678 200796
rect 255314 200784 255320 200796
rect 234672 200756 255320 200784
rect 234672 200744 234678 200756
rect 255314 200744 255320 200756
rect 255372 200744 255378 200796
rect 205542 200132 205548 200184
rect 205600 200172 205606 200184
rect 215846 200172 215852 200184
rect 205600 200144 215852 200172
rect 205600 200132 205606 200144
rect 215846 200132 215852 200144
rect 215904 200132 215910 200184
rect 232590 200172 232596 200184
rect 217336 200144 232596 200172
rect 169754 200064 169760 200116
rect 169812 200104 169818 200116
rect 205560 200104 205588 200132
rect 169812 200076 205588 200104
rect 169812 200064 169818 200076
rect 206462 200064 206468 200116
rect 206520 200104 206526 200116
rect 217336 200104 217364 200144
rect 232590 200132 232596 200144
rect 232648 200132 232654 200184
rect 206520 200076 217364 200104
rect 206520 200064 206526 200076
rect 147582 199452 147588 199504
rect 147640 199492 147646 199504
rect 194318 199492 194324 199504
rect 147640 199464 194324 199492
rect 147640 199452 147646 199464
rect 194318 199452 194324 199464
rect 194376 199452 194382 199504
rect 63402 199384 63408 199436
rect 63460 199424 63466 199436
rect 168374 199424 168380 199436
rect 63460 199396 168380 199424
rect 63460 199384 63466 199396
rect 168374 199384 168380 199396
rect 168432 199384 168438 199436
rect 217318 199384 217324 199436
rect 217376 199424 217382 199436
rect 307846 199424 307852 199436
rect 217376 199396 307852 199424
rect 217376 199384 217382 199396
rect 307846 199384 307852 199396
rect 307904 199384 307910 199436
rect 53466 198636 53472 198688
rect 53524 198676 53530 198688
rect 160738 198676 160744 198688
rect 53524 198648 160744 198676
rect 53524 198636 53530 198648
rect 160738 198636 160744 198648
rect 160796 198636 160802 198688
rect 168374 198636 168380 198688
rect 168432 198676 168438 198688
rect 201494 198676 201500 198688
rect 168432 198648 201500 198676
rect 168432 198636 168438 198648
rect 201494 198636 201500 198648
rect 201552 198636 201558 198688
rect 120074 198568 120080 198620
rect 120132 198608 120138 198620
rect 156782 198608 156788 198620
rect 120132 198580 156788 198608
rect 120132 198568 120138 198580
rect 156782 198568 156788 198580
rect 156840 198568 156846 198620
rect 166994 198024 167000 198076
rect 167052 198064 167058 198076
rect 213270 198064 213276 198076
rect 167052 198036 213276 198064
rect 167052 198024 167058 198036
rect 213270 198024 213276 198036
rect 213328 198024 213334 198076
rect 215110 198024 215116 198076
rect 215168 198064 215174 198076
rect 241606 198064 241612 198076
rect 215168 198036 241612 198064
rect 215168 198024 215174 198036
rect 241606 198024 241612 198036
rect 241664 198024 241670 198076
rect 202138 197956 202144 198008
rect 202196 197996 202202 198008
rect 295518 197996 295524 198008
rect 202196 197968 295524 197996
rect 202196 197956 202202 197968
rect 295518 197956 295524 197968
rect 295576 197956 295582 198008
rect 118602 197276 118608 197328
rect 118660 197316 118666 197328
rect 170490 197316 170496 197328
rect 118660 197288 170496 197316
rect 118660 197276 118666 197288
rect 170490 197276 170496 197288
rect 170548 197276 170554 197328
rect 188522 196664 188528 196716
rect 188580 196704 188586 196716
rect 196802 196704 196808 196716
rect 188580 196676 196808 196704
rect 188580 196664 188586 196676
rect 196802 196664 196808 196676
rect 196860 196664 196866 196716
rect 201310 196664 201316 196716
rect 201368 196704 201374 196716
rect 240134 196704 240140 196716
rect 201368 196676 240140 196704
rect 201368 196664 201374 196676
rect 240134 196664 240140 196676
rect 240192 196664 240198 196716
rect 255958 196664 255964 196716
rect 256016 196704 256022 196716
rect 285858 196704 285864 196716
rect 256016 196676 285864 196704
rect 256016 196664 256022 196676
rect 285858 196664 285864 196676
rect 285916 196664 285922 196716
rect 112990 196596 112996 196648
rect 113048 196636 113054 196648
rect 185578 196636 185584 196648
rect 113048 196608 185584 196636
rect 113048 196596 113054 196608
rect 185578 196596 185584 196608
rect 185636 196596 185642 196648
rect 195790 196596 195796 196648
rect 195848 196636 195854 196648
rect 279602 196636 279608 196648
rect 195848 196608 279608 196636
rect 195848 196596 195854 196608
rect 279602 196596 279608 196608
rect 279660 196596 279666 196648
rect 191926 195916 191932 195968
rect 191984 195956 191990 195968
rect 255406 195956 255412 195968
rect 191984 195928 255412 195956
rect 191984 195916 191990 195928
rect 255406 195916 255412 195928
rect 255464 195916 255470 195968
rect 158714 195848 158720 195900
rect 158772 195888 158778 195900
rect 159358 195888 159364 195900
rect 158772 195860 159364 195888
rect 158772 195848 158778 195860
rect 159358 195848 159364 195860
rect 159416 195888 159422 195900
rect 193122 195888 193128 195900
rect 159416 195860 193128 195888
rect 159416 195848 159422 195860
rect 193122 195848 193128 195860
rect 193180 195848 193186 195900
rect 194318 195848 194324 195900
rect 194376 195888 194382 195900
rect 252738 195888 252744 195900
rect 194376 195860 252744 195888
rect 194376 195848 194382 195860
rect 252738 195848 252744 195860
rect 252796 195848 252802 195900
rect 318150 195304 318156 195356
rect 318208 195344 318214 195356
rect 326338 195344 326344 195356
rect 318208 195316 326344 195344
rect 318208 195304 318214 195316
rect 326338 195304 326344 195316
rect 326396 195304 326402 195356
rect 133138 195236 133144 195288
rect 133196 195276 133202 195288
rect 158714 195276 158720 195288
rect 133196 195248 158720 195276
rect 133196 195236 133202 195248
rect 158714 195236 158720 195248
rect 158772 195236 158778 195288
rect 272610 195236 272616 195288
rect 272668 195276 272674 195288
rect 292666 195276 292672 195288
rect 272668 195248 292672 195276
rect 272668 195236 272674 195248
rect 292666 195236 292672 195248
rect 292724 195236 292730 195288
rect 325602 195236 325608 195288
rect 325660 195276 325666 195288
rect 349890 195276 349896 195288
rect 325660 195248 349896 195276
rect 325660 195236 325666 195248
rect 349890 195236 349896 195248
rect 349948 195236 349954 195288
rect 17218 195032 17224 195084
rect 17276 195072 17282 195084
rect 17862 195072 17868 195084
rect 17276 195044 17868 195072
rect 17276 195032 17282 195044
rect 17862 195032 17868 195044
rect 17920 195032 17926 195084
rect 17862 194556 17868 194608
rect 17920 194596 17926 194608
rect 181530 194596 181536 194608
rect 17920 194568 181536 194596
rect 17920 194556 17926 194568
rect 181530 194556 181536 194568
rect 181588 194556 181594 194608
rect 200758 194488 200764 194540
rect 200816 194528 200822 194540
rect 204254 194528 204260 194540
rect 200816 194500 204260 194528
rect 200816 194488 200822 194500
rect 204254 194488 204260 194500
rect 204312 194488 204318 194540
rect 50798 193876 50804 193928
rect 50856 193916 50862 193928
rect 139394 193916 139400 193928
rect 50856 193888 139400 193916
rect 50856 193876 50862 193888
rect 139394 193876 139400 193888
rect 139452 193876 139458 193928
rect 206278 193876 206284 193928
rect 206336 193916 206342 193928
rect 281626 193916 281632 193928
rect 206336 193888 281632 193916
rect 206336 193876 206342 193888
rect 281626 193876 281632 193888
rect 281684 193876 281690 193928
rect 89622 193808 89628 193860
rect 89680 193848 89686 193860
rect 209222 193848 209228 193860
rect 89680 193820 209228 193848
rect 89680 193808 89686 193820
rect 209222 193808 209228 193820
rect 209280 193808 209286 193860
rect 266998 193808 267004 193860
rect 267056 193848 267062 193860
rect 276750 193848 276756 193860
rect 267056 193820 276756 193848
rect 267056 193808 267062 193820
rect 276750 193808 276756 193820
rect 276808 193808 276814 193860
rect 286962 193808 286968 193860
rect 287020 193848 287026 193860
rect 294138 193848 294144 193860
rect 287020 193820 294144 193848
rect 287020 193808 287026 193820
rect 294138 193808 294144 193820
rect 294196 193808 294202 193860
rect 93118 193128 93124 193180
rect 93176 193168 93182 193180
rect 166994 193168 167000 193180
rect 93176 193140 167000 193168
rect 93176 193128 93182 193140
rect 166994 193128 167000 193140
rect 167052 193128 167058 193180
rect 139394 193060 139400 193112
rect 139452 193100 139458 193112
rect 198734 193100 198740 193112
rect 139452 193072 198740 193100
rect 139452 193060 139458 193072
rect 198734 193060 198740 193072
rect 198792 193060 198798 193112
rect 198734 192516 198740 192568
rect 198792 192556 198798 192568
rect 223482 192556 223488 192568
rect 198792 192528 223488 192556
rect 198792 192516 198798 192528
rect 223482 192516 223488 192528
rect 223540 192516 223546 192568
rect 224310 192516 224316 192568
rect 224368 192556 224374 192568
rect 245746 192556 245752 192568
rect 224368 192528 245752 192556
rect 224368 192516 224374 192528
rect 245746 192516 245752 192528
rect 245804 192516 245810 192568
rect 276934 192516 276940 192568
rect 276992 192556 276998 192568
rect 298186 192556 298192 192568
rect 276992 192528 298192 192556
rect 276992 192516 276998 192528
rect 298186 192516 298192 192528
rect 298244 192516 298250 192568
rect 204254 192448 204260 192500
rect 204312 192488 204318 192500
rect 238110 192488 238116 192500
rect 204312 192460 238116 192488
rect 204312 192448 204318 192460
rect 238110 192448 238116 192460
rect 238168 192448 238174 192500
rect 253198 192448 253204 192500
rect 253256 192488 253262 192500
rect 443086 192488 443092 192500
rect 253256 192460 443092 192488
rect 253256 192448 253262 192460
rect 443086 192448 443092 192460
rect 443144 192448 443150 192500
rect 33778 191768 33784 191820
rect 33836 191808 33842 191820
rect 34330 191808 34336 191820
rect 33836 191780 34336 191808
rect 33836 191768 33842 191780
rect 34330 191768 34336 191780
rect 34388 191808 34394 191820
rect 165522 191808 165528 191820
rect 34388 191780 165528 191808
rect 34388 191768 34394 191780
rect 165522 191768 165528 191780
rect 165580 191808 165586 191820
rect 196710 191808 196716 191820
rect 165580 191780 196716 191808
rect 165580 191768 165586 191780
rect 196710 191768 196716 191780
rect 196768 191768 196774 191820
rect 199470 191156 199476 191208
rect 199528 191196 199534 191208
rect 235994 191196 236000 191208
rect 199528 191168 236000 191196
rect 199528 191156 199534 191168
rect 235994 191156 236000 191168
rect 236052 191156 236058 191208
rect 197998 191088 198004 191140
rect 198056 191128 198062 191140
rect 290090 191128 290096 191140
rect 198056 191100 290096 191128
rect 198056 191088 198062 191100
rect 290090 191088 290096 191100
rect 290148 191088 290154 191140
rect 177298 189796 177304 189848
rect 177356 189836 177362 189848
rect 202138 189836 202144 189848
rect 177356 189808 202144 189836
rect 177356 189796 177362 189808
rect 202138 189796 202144 189808
rect 202196 189796 202202 189848
rect 224218 189796 224224 189848
rect 224276 189836 224282 189848
rect 242986 189836 242992 189848
rect 224276 189808 242992 189836
rect 224276 189796 224282 189808
rect 242986 189796 242992 189808
rect 243044 189796 243050 189848
rect 155862 189728 155868 189780
rect 155920 189768 155926 189780
rect 164878 189768 164884 189780
rect 155920 189740 164884 189768
rect 155920 189728 155926 189740
rect 164878 189728 164884 189740
rect 164936 189728 164942 189780
rect 193858 189728 193864 189780
rect 193916 189768 193922 189780
rect 231118 189768 231124 189780
rect 193916 189740 231124 189768
rect 193916 189728 193922 189740
rect 231118 189728 231124 189740
rect 231176 189728 231182 189780
rect 110322 189048 110328 189100
rect 110380 189088 110386 189100
rect 175918 189088 175924 189100
rect 110380 189060 175924 189088
rect 110380 189048 110386 189060
rect 175918 189048 175924 189060
rect 175976 189048 175982 189100
rect 3510 188980 3516 189032
rect 3568 189020 3574 189032
rect 29638 189020 29644 189032
rect 3568 188992 29644 189020
rect 3568 188980 3574 188992
rect 29638 188980 29644 188992
rect 29696 188980 29702 189032
rect 180702 188300 180708 188352
rect 180760 188340 180766 188352
rect 204898 188340 204904 188352
rect 180760 188312 204904 188340
rect 180760 188300 180766 188312
rect 204898 188300 204904 188312
rect 204956 188300 204962 188352
rect 268378 188300 268384 188352
rect 268436 188340 268442 188352
rect 285766 188340 285772 188352
rect 268436 188312 285772 188340
rect 268436 188300 268442 188312
rect 285766 188300 285772 188312
rect 285824 188300 285830 188352
rect 129090 187688 129096 187740
rect 129148 187728 129154 187740
rect 177298 187728 177304 187740
rect 129148 187700 177304 187728
rect 129148 187688 129154 187700
rect 177298 187688 177304 187700
rect 177356 187688 177362 187740
rect 205634 187688 205640 187740
rect 205692 187728 205698 187740
rect 244458 187728 244464 187740
rect 205692 187700 244464 187728
rect 205692 187688 205698 187700
rect 244458 187688 244464 187700
rect 244516 187688 244522 187740
rect 222838 187620 222844 187672
rect 222896 187660 222902 187672
rect 229738 187660 229744 187672
rect 222896 187632 229744 187660
rect 222896 187620 222902 187632
rect 229738 187620 229744 187632
rect 229796 187620 229802 187672
rect 177942 187008 177948 187060
rect 178000 187048 178006 187060
rect 206278 187048 206284 187060
rect 178000 187020 206284 187048
rect 178000 187008 178006 187020
rect 206278 187008 206284 187020
rect 206336 187008 206342 187060
rect 56502 186940 56508 186992
rect 56560 186980 56566 186992
rect 217226 186980 217232 186992
rect 56560 186952 217232 186980
rect 56560 186940 56566 186952
rect 217226 186940 217232 186952
rect 217284 186940 217290 186992
rect 275278 186940 275284 186992
rect 275336 186980 275342 186992
rect 296806 186980 296812 186992
rect 275336 186952 296812 186980
rect 275336 186940 275342 186952
rect 296806 186940 296812 186952
rect 296864 186940 296870 186992
rect 217226 186396 217232 186448
rect 217284 186436 217290 186448
rect 218146 186436 218152 186448
rect 217284 186408 218152 186436
rect 217284 186396 217290 186408
rect 218146 186396 218152 186408
rect 218204 186396 218210 186448
rect 133782 186328 133788 186380
rect 133840 186368 133846 186380
rect 176010 186368 176016 186380
rect 133840 186340 176016 186368
rect 133840 186328 133846 186340
rect 176010 186328 176016 186340
rect 176068 186328 176074 186380
rect 218054 186328 218060 186380
rect 218112 186368 218118 186380
rect 238938 186368 238944 186380
rect 218112 186340 238944 186368
rect 218112 186328 218118 186340
rect 238938 186328 238944 186340
rect 238996 186328 239002 186380
rect 186222 185648 186228 185700
rect 186280 185688 186286 185700
rect 236086 185688 236092 185700
rect 186280 185660 236092 185688
rect 186280 185648 186286 185660
rect 236086 185648 236092 185660
rect 236144 185648 236150 185700
rect 258718 185648 258724 185700
rect 258776 185688 258782 185700
rect 281718 185688 281724 185700
rect 258776 185660 281724 185688
rect 258776 185648 258782 185660
rect 281718 185648 281724 185660
rect 281776 185648 281782 185700
rect 207658 185580 207664 185632
rect 207716 185620 207722 185632
rect 279418 185620 279424 185632
rect 207716 185592 279424 185620
rect 207716 185580 207722 185592
rect 279418 185580 279424 185592
rect 279476 185580 279482 185632
rect 114462 184968 114468 185020
rect 114520 185008 114526 185020
rect 185762 185008 185768 185020
rect 114520 184980 185768 185008
rect 114520 184968 114526 184980
rect 185762 184968 185768 184980
rect 185820 184968 185826 185020
rect 100662 184900 100668 184952
rect 100720 184940 100726 184952
rect 178678 184940 178684 184952
rect 100720 184912 178684 184940
rect 100720 184900 100726 184912
rect 178678 184900 178684 184912
rect 178736 184900 178742 184952
rect 177850 184220 177856 184272
rect 177908 184260 177914 184272
rect 204162 184260 204168 184272
rect 177908 184232 204168 184260
rect 177908 184220 177914 184232
rect 204162 184220 204168 184232
rect 204220 184220 204226 184272
rect 204898 184220 204904 184272
rect 204956 184260 204962 184272
rect 232038 184260 232044 184272
rect 204956 184232 232044 184260
rect 204956 184220 204962 184232
rect 232038 184220 232044 184232
rect 232096 184220 232102 184272
rect 184750 184152 184756 184204
rect 184808 184192 184814 184204
rect 232498 184192 232504 184204
rect 184808 184164 232504 184192
rect 184808 184152 184814 184164
rect 232498 184152 232504 184164
rect 232556 184152 232562 184204
rect 232590 184152 232596 184204
rect 232648 184192 232654 184204
rect 254026 184192 254032 184204
rect 232648 184164 254032 184192
rect 232648 184152 232654 184164
rect 254026 184152 254032 184164
rect 254084 184152 254090 184204
rect 280798 184152 280804 184204
rect 280856 184192 280862 184204
rect 301130 184192 301136 184204
rect 280856 184164 301136 184192
rect 280856 184152 280862 184164
rect 301130 184152 301136 184164
rect 301188 184152 301194 184204
rect 117222 183608 117228 183660
rect 117280 183648 117286 183660
rect 169386 183648 169392 183660
rect 117280 183620 169392 183648
rect 117280 183608 117286 183620
rect 169386 183608 169392 183620
rect 169444 183608 169450 183660
rect 108942 183540 108948 183592
rect 109000 183580 109006 183592
rect 171962 183580 171968 183592
rect 109000 183552 171968 183580
rect 109000 183540 109006 183552
rect 171962 183540 171968 183552
rect 172020 183540 172026 183592
rect 204162 183472 204168 183524
rect 204220 183512 204226 183524
rect 218054 183512 218060 183524
rect 204220 183484 218060 183512
rect 204220 183472 204226 183484
rect 218054 183472 218060 183484
rect 218112 183472 218118 183524
rect 224954 182928 224960 182980
rect 225012 182968 225018 182980
rect 227714 182968 227720 182980
rect 225012 182940 227720 182968
rect 225012 182928 225018 182940
rect 227714 182928 227720 182940
rect 227772 182928 227778 182980
rect 184842 182860 184848 182912
rect 184900 182900 184906 182912
rect 193858 182900 193864 182912
rect 184900 182872 193864 182900
rect 184900 182860 184906 182872
rect 193858 182860 193864 182872
rect 193916 182860 193922 182912
rect 199378 182860 199384 182912
rect 199436 182900 199442 182912
rect 225690 182900 225696 182912
rect 199436 182872 225696 182900
rect 199436 182860 199442 182872
rect 225690 182860 225696 182872
rect 225748 182860 225754 182912
rect 240778 182860 240784 182912
rect 240836 182900 240842 182912
rect 280430 182900 280436 182912
rect 240836 182872 280436 182900
rect 240836 182860 240842 182872
rect 280430 182860 280436 182872
rect 280488 182860 280494 182912
rect 170490 182792 170496 182844
rect 170548 182832 170554 182844
rect 200758 182832 200764 182844
rect 170548 182804 200764 182832
rect 170548 182792 170554 182804
rect 200758 182792 200764 182804
rect 200816 182792 200822 182844
rect 220078 182792 220084 182844
rect 220136 182832 220142 182844
rect 233510 182832 233516 182844
rect 220136 182804 233516 182832
rect 220136 182792 220142 182804
rect 233510 182792 233516 182804
rect 233568 182792 233574 182844
rect 246298 182792 246304 182844
rect 246356 182832 246362 182844
rect 432046 182832 432052 182844
rect 246356 182804 432052 182832
rect 246356 182792 246362 182804
rect 432046 182792 432052 182804
rect 432104 182792 432110 182844
rect 134794 182248 134800 182300
rect 134852 182288 134858 182300
rect 162854 182288 162860 182300
rect 134852 182260 162860 182288
rect 134852 182248 134858 182260
rect 162854 182248 162860 182260
rect 162912 182248 162918 182300
rect 123478 182180 123484 182232
rect 123536 182220 123542 182232
rect 170490 182220 170496 182232
rect 123536 182192 170496 182220
rect 123536 182180 123542 182192
rect 170490 182180 170496 182192
rect 170548 182180 170554 182232
rect 178770 181500 178776 181552
rect 178828 181540 178834 181552
rect 204898 181540 204904 181552
rect 178828 181512 204904 181540
rect 178828 181500 178834 181512
rect 204898 181500 204904 181512
rect 204956 181500 204962 181552
rect 206370 181500 206376 181552
rect 206428 181540 206434 181552
rect 238846 181540 238852 181552
rect 206428 181512 238852 181540
rect 206428 181500 206434 181512
rect 238846 181500 238852 181512
rect 238904 181500 238910 181552
rect 181438 181432 181444 181484
rect 181496 181472 181502 181484
rect 227806 181472 227812 181484
rect 181496 181444 227812 181472
rect 181496 181432 181502 181444
rect 227806 181432 227812 181444
rect 227864 181432 227870 181484
rect 260742 181432 260748 181484
rect 260800 181472 260806 181484
rect 269206 181472 269212 181484
rect 260800 181444 269212 181472
rect 260800 181432 260806 181444
rect 269206 181432 269212 181444
rect 269264 181432 269270 181484
rect 279510 181432 279516 181484
rect 279568 181472 279574 181484
rect 287330 181472 287336 181484
rect 279568 181444 287336 181472
rect 279568 181432 279574 181444
rect 287330 181432 287336 181444
rect 287388 181432 287394 181484
rect 148226 180888 148232 180940
rect 148284 180928 148290 180940
rect 174538 180928 174544 180940
rect 148284 180900 174544 180928
rect 148284 180888 148290 180900
rect 174538 180888 174544 180900
rect 174596 180888 174602 180940
rect 115842 180820 115848 180872
rect 115900 180860 115906 180872
rect 166442 180860 166448 180872
rect 115900 180832 166448 180860
rect 115900 180820 115906 180832
rect 166442 180820 166448 180832
rect 166500 180820 166506 180872
rect 275278 180820 275284 180872
rect 275336 180860 275342 180872
rect 303798 180860 303804 180872
rect 275336 180832 303804 180860
rect 275336 180820 275342 180832
rect 303798 180820 303804 180832
rect 303856 180820 303862 180872
rect 182910 180752 182916 180804
rect 182968 180792 182974 180804
rect 225874 180792 225880 180804
rect 182968 180764 225880 180792
rect 182968 180752 182974 180764
rect 225874 180752 225880 180764
rect 225932 180752 225938 180804
rect 228634 180752 228640 180804
rect 228692 180792 228698 180804
rect 278682 180792 278688 180804
rect 228692 180764 278688 180792
rect 228692 180752 228698 180764
rect 278682 180752 278688 180764
rect 278740 180752 278746 180804
rect 278130 180616 278136 180668
rect 278188 180656 278194 180668
rect 280338 180656 280344 180668
rect 278188 180628 280344 180656
rect 278188 180616 278194 180628
rect 280338 180616 280344 180628
rect 280396 180616 280402 180668
rect 214558 180072 214564 180124
rect 214616 180112 214622 180124
rect 230382 180112 230388 180124
rect 214616 180084 230388 180112
rect 214616 180072 214622 180084
rect 230382 180072 230388 180084
rect 230440 180072 230446 180124
rect 254578 180072 254584 180124
rect 254636 180112 254642 180124
rect 262214 180112 262220 180124
rect 254636 180084 262220 180112
rect 254636 180072 254642 180084
rect 262214 180072 262220 180084
rect 262272 180072 262278 180124
rect 272518 180072 272524 180124
rect 272576 180112 272582 180124
rect 292758 180112 292764 180124
rect 272576 180084 292764 180112
rect 272576 180072 272582 180084
rect 292758 180072 292764 180084
rect 292816 180072 292822 180124
rect 282178 179732 282184 179784
rect 282236 179772 282242 179784
rect 285950 179772 285956 179784
rect 282236 179744 285956 179772
rect 282236 179732 282242 179744
rect 285950 179732 285956 179744
rect 286008 179732 286014 179784
rect 119798 179460 119804 179512
rect 119856 179500 119862 179512
rect 167730 179500 167736 179512
rect 119856 179472 167736 179500
rect 119856 179460 119862 179472
rect 167730 179460 167736 179472
rect 167788 179460 167794 179512
rect 128170 179392 128176 179444
rect 128228 179432 128234 179444
rect 214098 179432 214104 179444
rect 128228 179404 214104 179432
rect 128228 179392 128234 179404
rect 214098 179392 214104 179404
rect 214156 179392 214162 179444
rect 231118 179324 231124 179376
rect 231176 179364 231182 179376
rect 275278 179364 275284 179376
rect 231176 179336 275284 179364
rect 231176 179324 231182 179336
rect 275278 179324 275284 179336
rect 275336 179324 275342 179376
rect 215110 178712 215116 178764
rect 215168 178752 215174 178764
rect 229278 178752 229284 178764
rect 215168 178724 229284 178752
rect 215168 178712 215174 178724
rect 229278 178712 229284 178724
rect 229336 178712 229342 178764
rect 276750 178712 276756 178764
rect 276808 178752 276814 178764
rect 279234 178752 279240 178764
rect 276808 178724 279240 178752
rect 276808 178712 276814 178724
rect 279234 178712 279240 178724
rect 279292 178712 279298 178764
rect 196802 178644 196808 178696
rect 196860 178684 196866 178696
rect 237466 178684 237472 178696
rect 196860 178656 237472 178684
rect 196860 178644 196866 178656
rect 237466 178644 237472 178656
rect 237524 178644 237530 178696
rect 265618 178644 265624 178696
rect 265676 178684 265682 178696
rect 283006 178684 283012 178696
rect 265676 178656 283012 178684
rect 265676 178644 265682 178656
rect 283006 178644 283012 178656
rect 283064 178644 283070 178696
rect 285030 178644 285036 178696
rect 285088 178684 285094 178696
rect 299658 178684 299664 178696
rect 285088 178656 299664 178684
rect 285088 178644 285094 178656
rect 299658 178644 299664 178656
rect 299716 178644 299722 178696
rect 300210 178644 300216 178696
rect 300268 178684 300274 178696
rect 414106 178684 414112 178696
rect 300268 178656 414112 178684
rect 300268 178644 300274 178656
rect 414106 178644 414112 178656
rect 414164 178644 414170 178696
rect 132402 178100 132408 178152
rect 132460 178140 132466 178152
rect 165522 178140 165528 178152
rect 132460 178112 165528 178140
rect 132460 178100 132466 178112
rect 165522 178100 165528 178112
rect 165580 178100 165586 178152
rect 125042 178032 125048 178084
rect 125100 178072 125106 178084
rect 198090 178072 198096 178084
rect 125100 178044 198096 178072
rect 125100 178032 125106 178044
rect 198090 178032 198096 178044
rect 198148 178032 198154 178084
rect 102042 177964 102048 178016
rect 102100 178004 102106 178016
rect 129090 178004 129096 178016
rect 102100 177976 129096 178004
rect 102100 177964 102106 177976
rect 129090 177964 129096 177976
rect 129148 177964 129154 178016
rect 225690 177964 225696 178016
rect 225748 178004 225754 178016
rect 229094 178004 229100 178016
rect 225748 177976 229100 178004
rect 225748 177964 225754 177976
rect 229094 177964 229100 177976
rect 229152 177964 229158 178016
rect 276658 177964 276664 178016
rect 276716 178004 276722 178016
rect 279326 178004 279332 178016
rect 276716 177976 279332 178004
rect 276716 177964 276722 177976
rect 279326 177964 279332 177976
rect 279384 177964 279390 178016
rect 284938 177964 284944 178016
rect 284996 178004 285002 178016
rect 288434 178004 288440 178016
rect 284996 177976 288440 178004
rect 284996 177964 285002 177976
rect 288434 177964 288440 177976
rect 288492 177964 288498 178016
rect 215386 177352 215392 177404
rect 215444 177392 215450 177404
rect 226242 177392 226248 177404
rect 215444 177364 226248 177392
rect 215444 177352 215450 177364
rect 226242 177352 226248 177364
rect 226300 177352 226306 177404
rect 238110 177352 238116 177404
rect 238168 177392 238174 177404
rect 241514 177392 241520 177404
rect 238168 177364 241520 177392
rect 238168 177352 238174 177364
rect 241514 177352 241520 177364
rect 241572 177352 241578 177404
rect 198642 177284 198648 177336
rect 198700 177324 198706 177336
rect 279510 177324 279516 177336
rect 198700 177296 279516 177324
rect 198700 177284 198706 177296
rect 279510 177284 279516 177296
rect 279568 177284 279574 177336
rect 136082 176740 136088 176792
rect 136140 176780 136146 176792
rect 140774 176780 140780 176792
rect 136140 176752 140780 176780
rect 136140 176740 136146 176752
rect 140774 176740 140780 176752
rect 140832 176740 140838 176792
rect 158990 176740 158996 176792
rect 159048 176780 159054 176792
rect 170398 176780 170404 176792
rect 159048 176752 170404 176780
rect 159048 176740 159054 176752
rect 170398 176740 170404 176752
rect 170456 176740 170462 176792
rect 130746 176672 130752 176724
rect 130804 176712 130810 176724
rect 212442 176712 212448 176724
rect 130804 176684 212448 176712
rect 130804 176672 130810 176684
rect 212442 176672 212448 176684
rect 212500 176672 212506 176724
rect 140774 176604 140780 176656
rect 140832 176644 140838 176656
rect 213914 176644 213920 176656
rect 140832 176616 213920 176644
rect 140832 176604 140838 176616
rect 213914 176604 213920 176616
rect 213972 176604 213978 176656
rect 269850 176604 269856 176656
rect 269908 176644 269914 176656
rect 279878 176644 279884 176656
rect 269908 176616 279884 176644
rect 269908 176604 269914 176616
rect 279878 176604 279884 176616
rect 279936 176604 279942 176656
rect 276842 176536 276848 176588
rect 276900 176576 276906 176588
rect 280062 176576 280068 176588
rect 276900 176548 280068 176576
rect 276900 176536 276906 176548
rect 280062 176536 280068 176548
rect 280120 176536 280126 176588
rect 227530 175992 227536 176044
rect 227588 176032 227594 176044
rect 234706 176032 234712 176044
rect 227588 176004 234712 176032
rect 227588 175992 227594 176004
rect 234706 175992 234712 176004
rect 234764 175992 234770 176044
rect 47578 175924 47584 175976
rect 47636 175964 47642 175976
rect 128998 175964 129004 175976
rect 47636 175936 129004 175964
rect 47636 175924 47642 175936
rect 128998 175924 129004 175936
rect 129056 175924 129062 175976
rect 129458 175924 129464 175976
rect 129516 175964 129522 175976
rect 169754 175964 169760 175976
rect 129516 175936 169760 175964
rect 129516 175924 129522 175936
rect 169754 175924 169760 175936
rect 169812 175924 169818 175976
rect 185762 175924 185768 175976
rect 185820 175964 185826 175976
rect 214466 175964 214472 175976
rect 185820 175936 214472 175964
rect 185820 175924 185826 175936
rect 214466 175924 214472 175936
rect 214524 175924 214530 175976
rect 227714 175924 227720 175976
rect 227772 175964 227778 175976
rect 247218 175964 247224 175976
rect 227772 175936 247224 175964
rect 227772 175924 227778 175936
rect 247218 175924 247224 175936
rect 247276 175924 247282 175976
rect 279602 175924 279608 175976
rect 279660 175964 279666 175976
rect 280154 175964 280160 175976
rect 279660 175936 280160 175964
rect 279660 175924 279666 175936
rect 280154 175924 280160 175936
rect 280212 175924 280218 175976
rect 314010 175924 314016 175976
rect 314068 175964 314074 175976
rect 335998 175964 336004 175976
rect 314068 175936 336004 175964
rect 314068 175924 314074 175936
rect 335998 175924 336004 175936
rect 336056 175924 336062 175976
rect 227806 175896 227812 175908
rect 219406 175868 227812 175896
rect 215294 175244 215300 175296
rect 215352 175284 215358 175296
rect 219406 175284 219434 175868
rect 227806 175856 227812 175868
rect 227864 175856 227870 175908
rect 221182 175788 221188 175840
rect 221240 175788 221246 175840
rect 224218 175788 224224 175840
rect 224276 175788 224282 175840
rect 215352 175256 219434 175284
rect 215352 175244 215358 175256
rect 162854 175176 162860 175228
rect 162912 175216 162918 175228
rect 213914 175216 213920 175228
rect 162912 175188 213920 175216
rect 162912 175176 162918 175188
rect 213914 175176 213920 175188
rect 213972 175176 213978 175228
rect 214558 175176 214564 175228
rect 214616 175216 214622 175228
rect 221200 175216 221228 175788
rect 214616 175188 221228 175216
rect 224236 175216 224264 175788
rect 235350 175244 235356 175296
rect 235408 175284 235414 175296
rect 264974 175284 264980 175296
rect 235408 175256 264980 175284
rect 235408 175244 235414 175256
rect 264974 175244 264980 175256
rect 265032 175244 265038 175296
rect 281810 175244 281816 175296
rect 281868 175284 281874 175296
rect 314010 175284 314016 175296
rect 281868 175256 314016 175284
rect 281868 175244 281874 175256
rect 314010 175244 314016 175256
rect 314068 175244 314074 175296
rect 224236 175188 229048 175216
rect 214616 175176 214622 175188
rect 229020 175160 229048 175188
rect 231118 175176 231124 175228
rect 231176 175216 231182 175228
rect 232038 175216 232044 175228
rect 231176 175188 232044 175216
rect 231176 175176 231182 175188
rect 232038 175176 232044 175188
rect 232096 175176 232102 175228
rect 176010 175108 176016 175160
rect 176068 175148 176074 175160
rect 214006 175148 214012 175160
rect 176068 175120 214012 175148
rect 176068 175108 176074 175120
rect 214006 175108 214012 175120
rect 214064 175108 214070 175160
rect 229002 175108 229008 175160
rect 229060 175108 229066 175160
rect 282822 175108 282828 175160
rect 282880 175148 282886 175160
rect 300946 175148 300952 175160
rect 282880 175120 300952 175148
rect 282880 175108 282886 175120
rect 300946 175108 300952 175120
rect 301004 175108 301010 175160
rect 244918 174496 244924 174548
rect 244976 174536 244982 174548
rect 258166 174536 258172 174548
rect 244976 174508 258172 174536
rect 244976 174496 244982 174508
rect 258166 174496 258172 174508
rect 258224 174496 258230 174548
rect 229002 174020 229008 174072
rect 229060 174060 229066 174072
rect 229186 174060 229192 174072
rect 229060 174032 229192 174060
rect 229060 174020 229066 174032
rect 229186 174020 229192 174032
rect 229244 174020 229250 174072
rect 258718 173952 258724 174004
rect 258776 173992 258782 174004
rect 265066 173992 265072 174004
rect 258776 173964 265072 173992
rect 258776 173952 258782 173964
rect 265066 173952 265072 173964
rect 265124 173952 265130 174004
rect 214558 173884 214564 173936
rect 214616 173924 214622 173936
rect 233418 173924 233424 173936
rect 214616 173896 233424 173924
rect 214616 173884 214622 173896
rect 233418 173884 233424 173896
rect 233476 173884 233482 173936
rect 240870 173884 240876 173936
rect 240928 173924 240934 173936
rect 264974 173924 264980 173936
rect 240928 173896 264980 173924
rect 240928 173884 240934 173896
rect 264974 173884 264980 173896
rect 265032 173884 265038 173936
rect 165522 173816 165528 173868
rect 165580 173856 165586 173868
rect 213914 173856 213920 173868
rect 165580 173828 213920 173856
rect 165580 173816 165586 173828
rect 213914 173816 213920 173828
rect 213972 173816 213978 173868
rect 212442 173748 212448 173800
rect 212500 173788 212506 173800
rect 214006 173788 214012 173800
rect 212500 173760 214012 173788
rect 212500 173748 212506 173760
rect 214006 173748 214012 173760
rect 214064 173748 214070 173800
rect 167822 173408 167828 173460
rect 167880 173448 167886 173460
rect 173434 173448 173440 173460
rect 167880 173420 173440 173448
rect 167880 173408 167886 173420
rect 173434 173408 173440 173420
rect 173492 173408 173498 173460
rect 230750 173340 230756 173392
rect 230808 173380 230814 173392
rect 233234 173380 233240 173392
rect 230808 173352 233240 173380
rect 230808 173340 230814 173352
rect 233234 173340 233240 173352
rect 233292 173340 233298 173392
rect 177298 173136 177304 173188
rect 177356 173176 177362 173188
rect 197998 173176 198004 173188
rect 177356 173148 198004 173176
rect 177356 173136 177362 173148
rect 197998 173136 198004 173148
rect 198056 173136 198062 173188
rect 238110 173136 238116 173188
rect 238168 173176 238174 173188
rect 252554 173176 252560 173188
rect 238168 173148 252560 173176
rect 238168 173136 238174 173148
rect 252554 173136 252560 173148
rect 252612 173136 252618 173188
rect 258994 172592 259000 172644
rect 259052 172632 259058 172644
rect 265066 172632 265072 172644
rect 259052 172604 265072 172632
rect 259052 172592 259058 172604
rect 265066 172592 265072 172604
rect 265124 172592 265130 172644
rect 254670 172524 254676 172576
rect 254728 172564 254734 172576
rect 264974 172564 264980 172576
rect 254728 172536 264980 172564
rect 254728 172524 254734 172536
rect 264974 172524 264980 172536
rect 265032 172524 265038 172576
rect 169754 172456 169760 172508
rect 169812 172496 169818 172508
rect 213914 172496 213920 172508
rect 169812 172468 213920 172496
rect 169812 172456 169818 172468
rect 213914 172456 213920 172468
rect 213972 172456 213978 172508
rect 231578 172456 231584 172508
rect 231636 172496 231642 172508
rect 240226 172496 240232 172508
rect 231636 172468 240232 172496
rect 231636 172456 231642 172468
rect 240226 172456 240232 172468
rect 240284 172456 240290 172508
rect 173158 172388 173164 172440
rect 173216 172428 173222 172440
rect 215294 172428 215300 172440
rect 173216 172400 215300 172428
rect 173216 172388 173222 172400
rect 215294 172388 215300 172400
rect 215352 172388 215358 172440
rect 231762 172116 231768 172168
rect 231820 172156 231826 172168
rect 234614 172156 234620 172168
rect 231820 172128 234620 172156
rect 231820 172116 231826 172128
rect 234614 172116 234620 172128
rect 234672 172116 234678 172168
rect 247954 171164 247960 171216
rect 248012 171204 248018 171216
rect 264974 171204 264980 171216
rect 248012 171176 264980 171204
rect 248012 171164 248018 171176
rect 264974 171164 264980 171176
rect 265032 171164 265038 171216
rect 240962 171096 240968 171148
rect 241020 171136 241026 171148
rect 265066 171136 265072 171148
rect 241020 171108 265072 171136
rect 241020 171096 241026 171108
rect 265066 171096 265072 171108
rect 265124 171096 265130 171148
rect 165154 171028 165160 171080
rect 165212 171068 165218 171080
rect 214006 171068 214012 171080
rect 165212 171040 214012 171068
rect 165212 171028 165218 171040
rect 214006 171028 214012 171040
rect 214064 171028 214070 171080
rect 231762 171028 231768 171080
rect 231820 171068 231826 171080
rect 241514 171068 241520 171080
rect 231820 171040 241520 171068
rect 231820 171028 231826 171040
rect 241514 171028 241520 171040
rect 241572 171028 241578 171080
rect 164970 170960 164976 171012
rect 165028 171000 165034 171012
rect 213914 171000 213920 171012
rect 165028 170972 213920 171000
rect 165028 170960 165034 170972
rect 213914 170960 213920 170972
rect 213972 170960 213978 171012
rect 230750 170960 230756 171012
rect 230808 171000 230814 171012
rect 232498 171000 232504 171012
rect 230808 170972 232504 171000
rect 230808 170960 230814 170972
rect 232498 170960 232504 170972
rect 232556 170960 232562 171012
rect 281810 170960 281816 171012
rect 281868 171000 281874 171012
rect 283190 171000 283196 171012
rect 281868 170972 283196 171000
rect 281868 170960 281874 170972
rect 283190 170960 283196 170972
rect 283248 170960 283254 171012
rect 371970 170348 371976 170400
rect 372028 170388 372034 170400
rect 433978 170388 433984 170400
rect 372028 170360 433984 170388
rect 372028 170348 372034 170360
rect 433978 170348 433984 170360
rect 434036 170348 434042 170400
rect 243814 169736 243820 169788
rect 243872 169776 243878 169788
rect 264974 169776 264980 169788
rect 243872 169748 264980 169776
rect 243872 169736 243878 169748
rect 264974 169736 264980 169748
rect 265032 169736 265038 169788
rect 170490 169668 170496 169720
rect 170548 169708 170554 169720
rect 214006 169708 214012 169720
rect 170548 169680 214012 169708
rect 170548 169668 170554 169680
rect 214006 169668 214012 169680
rect 214064 169668 214070 169720
rect 231762 169668 231768 169720
rect 231820 169708 231826 169720
rect 243538 169708 243544 169720
rect 231820 169680 243544 169708
rect 231820 169668 231826 169680
rect 243538 169668 243544 169680
rect 243596 169668 243602 169720
rect 282822 169668 282828 169720
rect 282880 169708 282886 169720
rect 295518 169708 295524 169720
rect 282880 169680 295524 169708
rect 282880 169668 282886 169680
rect 295518 169668 295524 169680
rect 295576 169668 295582 169720
rect 198090 169600 198096 169652
rect 198148 169640 198154 169652
rect 213914 169640 213920 169652
rect 198148 169612 213920 169640
rect 198148 169600 198154 169612
rect 213914 169600 213920 169612
rect 213972 169600 213978 169652
rect 231210 169192 231216 169244
rect 231268 169232 231274 169244
rect 233326 169232 233332 169244
rect 231268 169204 233332 169232
rect 231268 169192 231274 169204
rect 233326 169192 233332 169204
rect 233384 169192 233390 169244
rect 250714 168444 250720 168496
rect 250772 168484 250778 168496
rect 264974 168484 264980 168496
rect 250772 168456 264980 168484
rect 250772 168444 250778 168456
rect 264974 168444 264980 168456
rect 265032 168444 265038 168496
rect 240778 168376 240784 168428
rect 240836 168416 240842 168428
rect 265066 168416 265072 168428
rect 240836 168388 265072 168416
rect 240836 168376 240842 168388
rect 265066 168376 265072 168388
rect 265124 168376 265130 168428
rect 167914 168308 167920 168360
rect 167972 168348 167978 168360
rect 213914 168348 213920 168360
rect 167972 168320 213920 168348
rect 167972 168308 167978 168320
rect 213914 168308 213920 168320
rect 213972 168308 213978 168360
rect 282730 168308 282736 168360
rect 282788 168348 282794 168360
rect 290090 168348 290096 168360
rect 282788 168320 290096 168348
rect 282788 168308 282794 168320
rect 290090 168308 290096 168320
rect 290148 168308 290154 168360
rect 169202 168240 169208 168292
rect 169260 168280 169266 168292
rect 214006 168280 214012 168292
rect 169260 168252 214012 168280
rect 169260 168240 169266 168252
rect 214006 168240 214012 168252
rect 214064 168240 214070 168292
rect 230566 168240 230572 168292
rect 230624 168280 230630 168292
rect 230842 168280 230848 168292
rect 230624 168252 230848 168280
rect 230624 168240 230630 168252
rect 230842 168240 230848 168252
rect 230900 168240 230906 168292
rect 231394 168172 231400 168224
rect 231452 168212 231458 168224
rect 237466 168212 237472 168224
rect 231452 168184 237472 168212
rect 231452 168172 231458 168184
rect 237466 168172 237472 168184
rect 237524 168172 237530 168224
rect 282822 167968 282828 168020
rect 282880 168008 282886 168020
rect 288434 168008 288440 168020
rect 282880 167980 288440 168008
rect 282880 167968 282886 167980
rect 288434 167968 288440 167980
rect 288492 167968 288498 168020
rect 391198 167628 391204 167680
rect 391256 167668 391262 167680
rect 430666 167668 430672 167680
rect 391256 167640 430672 167668
rect 391256 167628 391262 167640
rect 430666 167628 430672 167640
rect 430724 167628 430730 167680
rect 256050 167084 256056 167136
rect 256108 167124 256114 167136
rect 264974 167124 264980 167136
rect 256108 167096 264980 167124
rect 256108 167084 256114 167096
rect 264974 167084 264980 167096
rect 265032 167084 265038 167136
rect 252094 167016 252100 167068
rect 252152 167056 252158 167068
rect 265066 167056 265072 167068
rect 252152 167028 265072 167056
rect 252152 167016 252158 167028
rect 265066 167016 265072 167028
rect 265124 167016 265130 167068
rect 167730 166948 167736 167000
rect 167788 166988 167794 167000
rect 213914 166988 213920 167000
rect 167788 166960 213920 166988
rect 167788 166948 167794 166960
rect 213914 166948 213920 166960
rect 213972 166948 213978 167000
rect 177390 166880 177396 166932
rect 177448 166920 177454 166932
rect 214006 166920 214012 166932
rect 177448 166892 214012 166920
rect 177448 166880 177454 166892
rect 214006 166880 214012 166892
rect 214064 166880 214070 166932
rect 231762 166676 231768 166728
rect 231820 166716 231826 166728
rect 235258 166716 235264 166728
rect 231820 166688 235264 166716
rect 231820 166676 231826 166688
rect 235258 166676 235264 166688
rect 235316 166676 235322 166728
rect 230474 166268 230480 166320
rect 230532 166308 230538 166320
rect 230750 166308 230756 166320
rect 230532 166280 230756 166308
rect 230532 166268 230538 166280
rect 230750 166268 230756 166280
rect 230808 166268 230814 166320
rect 236730 166268 236736 166320
rect 236788 166308 236794 166320
rect 265710 166308 265716 166320
rect 236788 166280 265716 166308
rect 236788 166268 236794 166280
rect 265710 166268 265716 166280
rect 265768 166268 265774 166320
rect 370498 166268 370504 166320
rect 370556 166308 370562 166320
rect 439866 166308 439872 166320
rect 370556 166280 439872 166308
rect 370556 166268 370562 166280
rect 439866 166268 439872 166280
rect 439924 166268 439930 166320
rect 232774 165588 232780 165640
rect 232832 165628 232838 165640
rect 264974 165628 264980 165640
rect 232832 165600 264980 165628
rect 232832 165588 232838 165600
rect 264974 165588 264980 165600
rect 265032 165588 265038 165640
rect 166442 165520 166448 165572
rect 166500 165560 166506 165572
rect 213914 165560 213920 165572
rect 166500 165532 213920 165560
rect 166500 165520 166506 165532
rect 213914 165520 213920 165532
rect 213972 165520 213978 165572
rect 166534 165452 166540 165504
rect 166592 165492 166598 165504
rect 214006 165492 214012 165504
rect 166592 165464 214012 165492
rect 166592 165452 166598 165464
rect 214006 165452 214012 165464
rect 214064 165452 214070 165504
rect 231486 165452 231492 165504
rect 231544 165492 231550 165504
rect 235994 165492 236000 165504
rect 231544 165464 236000 165492
rect 231544 165452 231550 165464
rect 235994 165452 236000 165464
rect 236052 165452 236058 165504
rect 282822 165180 282828 165232
rect 282880 165220 282886 165232
rect 287054 165220 287060 165232
rect 282880 165192 287060 165220
rect 282880 165180 282886 165192
rect 287054 165180 287060 165192
rect 287112 165180 287118 165232
rect 3510 164840 3516 164892
rect 3568 164880 3574 164892
rect 17218 164880 17224 164892
rect 3568 164852 17224 164880
rect 3568 164840 3574 164852
rect 17218 164840 17224 164852
rect 17276 164840 17282 164892
rect 406378 164840 406384 164892
rect 406436 164880 406442 164892
rect 420270 164880 420276 164892
rect 406436 164852 420276 164880
rect 406436 164840 406442 164852
rect 420270 164840 420276 164852
rect 420328 164840 420334 164892
rect 238294 164296 238300 164348
rect 238352 164336 238358 164348
rect 264974 164336 264980 164348
rect 238352 164308 264980 164336
rect 238352 164296 238358 164308
rect 264974 164296 264980 164308
rect 265032 164296 265038 164348
rect 234062 164228 234068 164280
rect 234120 164268 234126 164280
rect 265066 164268 265072 164280
rect 234120 164240 265072 164268
rect 234120 164228 234126 164240
rect 265066 164228 265072 164240
rect 265124 164228 265130 164280
rect 184382 164160 184388 164212
rect 184440 164200 184446 164212
rect 213914 164200 213920 164212
rect 184440 164172 213920 164200
rect 184440 164160 184446 164172
rect 213914 164160 213920 164172
rect 213972 164160 213978 164212
rect 231762 164160 231768 164212
rect 231820 164200 231826 164212
rect 247402 164200 247408 164212
rect 231820 164172 247408 164200
rect 231820 164160 231826 164172
rect 247402 164160 247408 164172
rect 247460 164160 247466 164212
rect 282178 164160 282184 164212
rect 282236 164200 282242 164212
rect 309134 164200 309140 164212
rect 282236 164172 309140 164200
rect 282236 164160 282242 164172
rect 309134 164160 309140 164172
rect 309192 164160 309198 164212
rect 231670 164092 231676 164144
rect 231728 164132 231734 164144
rect 242894 164132 242900 164144
rect 231728 164104 242900 164132
rect 231728 164092 231734 164104
rect 242894 164092 242900 164104
rect 242952 164092 242958 164144
rect 281810 164092 281816 164144
rect 281868 164132 281874 164144
rect 284478 164132 284484 164144
rect 281868 164104 284484 164132
rect 281868 164092 281874 164104
rect 284478 164092 284484 164104
rect 284536 164092 284542 164144
rect 197998 163480 198004 163532
rect 198056 163520 198062 163532
rect 214834 163520 214840 163532
rect 198056 163492 214840 163520
rect 198056 163480 198062 163492
rect 214834 163480 214840 163492
rect 214892 163480 214898 163532
rect 319438 163480 319444 163532
rect 319496 163520 319502 163532
rect 371970 163520 371976 163532
rect 319496 163492 371976 163520
rect 319496 163480 319502 163492
rect 371970 163480 371976 163492
rect 372028 163480 372034 163532
rect 380158 163480 380164 163532
rect 380216 163520 380222 163532
rect 447410 163520 447416 163532
rect 380216 163492 447416 163520
rect 380216 163480 380222 163492
rect 447410 163480 447416 163492
rect 447468 163480 447474 163532
rect 255958 162936 255964 162988
rect 256016 162976 256022 162988
rect 265066 162976 265072 162988
rect 256016 162948 265072 162976
rect 256016 162936 256022 162948
rect 265066 162936 265072 162948
rect 265124 162936 265130 162988
rect 245010 162868 245016 162920
rect 245068 162908 245074 162920
rect 264974 162908 264980 162920
rect 245068 162880 264980 162908
rect 245068 162868 245074 162880
rect 264974 162868 264980 162880
rect 265032 162868 265038 162920
rect 167638 162800 167644 162852
rect 167696 162840 167702 162852
rect 213914 162840 213920 162852
rect 167696 162812 213920 162840
rect 167696 162800 167702 162812
rect 213914 162800 213920 162812
rect 213972 162800 213978 162852
rect 175918 162732 175924 162784
rect 175976 162772 175982 162784
rect 214006 162772 214012 162784
rect 175976 162744 214012 162772
rect 175976 162732 175982 162744
rect 214006 162732 214012 162744
rect 214064 162732 214070 162784
rect 282270 162732 282276 162784
rect 282328 162772 282334 162784
rect 329834 162772 329840 162784
rect 282328 162744 329840 162772
rect 282328 162732 282334 162744
rect 329834 162732 329840 162744
rect 329892 162732 329898 162784
rect 230934 162664 230940 162716
rect 230992 162704 230998 162716
rect 233418 162704 233424 162716
rect 230992 162676 233424 162704
rect 230992 162664 230998 162676
rect 233418 162664 233424 162676
rect 233476 162664 233482 162716
rect 378870 162120 378876 162172
rect 378928 162160 378934 162172
rect 418246 162160 418252 162172
rect 378928 162132 418252 162160
rect 378928 162120 378934 162132
rect 418246 162120 418252 162132
rect 418304 162120 418310 162172
rect 247770 161508 247776 161560
rect 247828 161548 247834 161560
rect 264974 161548 264980 161560
rect 247828 161520 264980 161548
rect 247828 161508 247834 161520
rect 264974 161508 264980 161520
rect 265032 161508 265038 161560
rect 235442 161440 235448 161492
rect 235500 161480 235506 161492
rect 265066 161480 265072 161492
rect 235500 161452 265072 161480
rect 235500 161440 235506 161452
rect 265066 161440 265072 161452
rect 265124 161440 265130 161492
rect 171962 161372 171968 161424
rect 172020 161412 172026 161424
rect 213914 161412 213920 161424
rect 172020 161384 213920 161412
rect 172020 161372 172026 161384
rect 213914 161372 213920 161384
rect 213972 161372 213978 161424
rect 282638 161372 282644 161424
rect 282696 161412 282702 161424
rect 325694 161412 325700 161424
rect 282696 161384 325700 161412
rect 282696 161372 282702 161384
rect 325694 161372 325700 161384
rect 325752 161372 325758 161424
rect 173342 161304 173348 161356
rect 173400 161344 173406 161356
rect 214006 161344 214012 161356
rect 173400 161316 214012 161344
rect 173400 161304 173406 161316
rect 214006 161304 214012 161316
rect 214064 161304 214070 161356
rect 231762 160692 231768 160744
rect 231820 160732 231826 160744
rect 241514 160732 241520 160744
rect 231820 160704 241520 160732
rect 231820 160692 231826 160704
rect 241514 160692 241520 160704
rect 241572 160692 241578 160744
rect 243722 160148 243728 160200
rect 243780 160188 243786 160200
rect 264974 160188 264980 160200
rect 243780 160160 264980 160188
rect 243780 160148 243786 160160
rect 264974 160148 264980 160160
rect 265032 160148 265038 160200
rect 236914 160080 236920 160132
rect 236972 160120 236978 160132
rect 265066 160120 265072 160132
rect 236972 160092 265072 160120
rect 236972 160080 236978 160092
rect 265066 160080 265072 160092
rect 265124 160080 265130 160132
rect 181530 160012 181536 160064
rect 181588 160052 181594 160064
rect 213914 160052 213920 160064
rect 181588 160024 213920 160052
rect 181588 160012 181594 160024
rect 213914 160012 213920 160024
rect 213972 160012 213978 160064
rect 282822 160012 282828 160064
rect 282880 160052 282886 160064
rect 320174 160052 320180 160064
rect 282880 160024 320180 160052
rect 282880 160012 282886 160024
rect 320174 160012 320180 160024
rect 320232 160012 320238 160064
rect 196710 159944 196716 159996
rect 196768 159984 196774 159996
rect 214006 159984 214012 159996
rect 196768 159956 214012 159984
rect 196768 159944 196774 159956
rect 214006 159944 214012 159956
rect 214064 159944 214070 159996
rect 282730 159944 282736 159996
rect 282788 159984 282794 159996
rect 296898 159984 296904 159996
rect 282788 159956 296904 159984
rect 282788 159944 282794 159956
rect 296898 159944 296904 159956
rect 296956 159944 296962 159996
rect 167822 159332 167828 159384
rect 167880 159372 167886 159384
rect 181438 159372 181444 159384
rect 167880 159344 181444 159372
rect 167880 159332 167886 159344
rect 181438 159332 181444 159344
rect 181496 159332 181502 159384
rect 230566 159332 230572 159384
rect 230624 159372 230630 159384
rect 244918 159372 244924 159384
rect 230624 159344 244924 159372
rect 230624 159332 230630 159344
rect 244918 159332 244924 159344
rect 244976 159332 244982 159384
rect 309042 159332 309048 159384
rect 309100 159372 309106 159384
rect 425054 159372 425060 159384
rect 309100 159344 425060 159372
rect 309100 159332 309106 159344
rect 425054 159332 425060 159344
rect 425112 159332 425118 159384
rect 231118 159264 231124 159316
rect 231176 159304 231182 159316
rect 238386 159304 238392 159316
rect 231176 159276 238392 159304
rect 231176 159264 231182 159276
rect 238386 159264 238392 159276
rect 238444 159264 238450 159316
rect 248046 158788 248052 158840
rect 248104 158828 248110 158840
rect 265066 158828 265072 158840
rect 248104 158800 265072 158828
rect 248104 158788 248110 158800
rect 265066 158788 265072 158800
rect 265124 158788 265130 158840
rect 238202 158720 238208 158772
rect 238260 158760 238266 158772
rect 264974 158760 264980 158772
rect 238260 158732 264980 158760
rect 238260 158720 238266 158732
rect 264974 158720 264980 158732
rect 265032 158720 265038 158772
rect 180334 158652 180340 158704
rect 180392 158692 180398 158704
rect 213914 158692 213920 158704
rect 180392 158664 213920 158692
rect 180392 158652 180398 158664
rect 213914 158652 213920 158664
rect 213972 158652 213978 158704
rect 282086 158652 282092 158704
rect 282144 158692 282150 158704
rect 288618 158692 288624 158704
rect 282144 158664 288624 158692
rect 282144 158652 282150 158664
rect 288618 158652 288624 158664
rect 288676 158652 288682 158704
rect 170398 157972 170404 158024
rect 170456 158012 170462 158024
rect 214558 158012 214564 158024
rect 170456 157984 214564 158012
rect 170456 157972 170462 157984
rect 214558 157972 214564 157984
rect 214616 157972 214622 158024
rect 231302 157972 231308 158024
rect 231360 158012 231366 158024
rect 238754 158012 238760 158024
rect 231360 157984 238760 158012
rect 231360 157972 231366 157984
rect 238754 157972 238760 157984
rect 238812 157972 238818 158024
rect 282178 157972 282184 158024
rect 282236 158012 282242 158024
rect 306466 158012 306472 158024
rect 282236 157984 306472 158012
rect 282236 157972 282242 157984
rect 306466 157972 306472 157984
rect 306524 157972 306530 158024
rect 353938 157972 353944 158024
rect 353996 158012 354002 158024
rect 414198 158012 414204 158024
rect 353996 157984 414204 158012
rect 353996 157972 354002 157984
rect 414198 157972 414204 157984
rect 414256 157972 414262 158024
rect 244918 157428 244924 157480
rect 244976 157468 244982 157480
rect 264974 157468 264980 157480
rect 244976 157440 264980 157468
rect 244976 157428 244982 157440
rect 264974 157428 264980 157440
rect 265032 157428 265038 157480
rect 233970 157360 233976 157412
rect 234028 157400 234034 157412
rect 265066 157400 265072 157412
rect 234028 157372 265072 157400
rect 234028 157360 234034 157372
rect 265066 157360 265072 157372
rect 265124 157360 265130 157412
rect 280062 157360 280068 157412
rect 280120 157400 280126 157412
rect 281534 157400 281540 157412
rect 280120 157372 281540 157400
rect 280120 157360 280126 157372
rect 281534 157360 281540 157372
rect 281592 157360 281598 157412
rect 166350 157292 166356 157344
rect 166408 157332 166414 157344
rect 213914 157332 213920 157344
rect 166408 157304 213920 157332
rect 166408 157292 166414 157304
rect 213914 157292 213920 157304
rect 213972 157292 213978 157344
rect 178678 157224 178684 157276
rect 178736 157264 178742 157276
rect 214006 157264 214012 157276
rect 178736 157236 214012 157264
rect 178736 157224 178742 157236
rect 214006 157224 214012 157236
rect 214064 157224 214070 157276
rect 283558 156680 283564 156732
rect 283616 156720 283622 156732
rect 294230 156720 294236 156732
rect 283616 156692 294236 156720
rect 283616 156680 283622 156692
rect 294230 156680 294236 156692
rect 294288 156680 294294 156732
rect 231118 156612 231124 156664
rect 231176 156652 231182 156664
rect 231946 156652 231952 156664
rect 231176 156624 231952 156652
rect 231176 156612 231182 156624
rect 231946 156612 231952 156624
rect 232004 156612 232010 156664
rect 282822 156612 282828 156664
rect 282880 156652 282886 156664
rect 303798 156652 303804 156664
rect 282880 156624 303804 156652
rect 282880 156612 282886 156624
rect 303798 156612 303804 156624
rect 303856 156612 303862 156664
rect 398742 156612 398748 156664
rect 398800 156652 398806 156664
rect 582742 156652 582748 156664
rect 398800 156624 582748 156652
rect 398800 156612 398806 156624
rect 582742 156612 582748 156624
rect 582800 156612 582806 156664
rect 231762 156544 231768 156596
rect 231820 156584 231826 156596
rect 244458 156584 244464 156596
rect 231820 156556 244464 156584
rect 231820 156544 231826 156556
rect 244458 156544 244464 156556
rect 244516 156544 244522 156596
rect 253290 156000 253296 156052
rect 253348 156040 253354 156052
rect 264974 156040 264980 156052
rect 253348 156012 264980 156040
rect 253348 156000 253354 156012
rect 264974 156000 264980 156012
rect 265032 156000 265038 156052
rect 239858 155932 239864 155984
rect 239916 155972 239922 155984
rect 265066 155972 265072 155984
rect 239916 155944 265072 155972
rect 239916 155932 239922 155944
rect 265066 155932 265072 155944
rect 265124 155932 265130 155984
rect 169110 155864 169116 155916
rect 169168 155904 169174 155916
rect 213914 155904 213920 155916
rect 169168 155876 213920 155904
rect 169168 155864 169174 155876
rect 213914 155864 213920 155876
rect 213972 155864 213978 155916
rect 185670 155796 185676 155848
rect 185728 155836 185734 155848
rect 214006 155836 214012 155848
rect 185728 155808 214012 155836
rect 185728 155796 185734 155808
rect 214006 155796 214012 155808
rect 214064 155796 214070 155848
rect 282546 155660 282552 155712
rect 282604 155700 282610 155712
rect 285950 155700 285956 155712
rect 282604 155672 285956 155700
rect 282604 155660 282610 155672
rect 285950 155660 285956 155672
rect 286008 155660 286014 155712
rect 230014 155184 230020 155236
rect 230072 155224 230078 155236
rect 265250 155224 265256 155236
rect 230072 155196 265256 155224
rect 230072 155184 230078 155196
rect 265250 155184 265256 155196
rect 265308 155184 265314 155236
rect 398650 155184 398656 155236
rect 398708 155224 398714 155236
rect 583570 155224 583576 155236
rect 398708 155196 583576 155224
rect 398708 155184 398714 155196
rect 583570 155184 583576 155196
rect 583628 155184 583634 155236
rect 235534 154572 235540 154624
rect 235592 154612 235598 154624
rect 265158 154612 265164 154624
rect 235592 154584 265164 154612
rect 235592 154572 235598 154584
rect 265158 154572 265164 154584
rect 265216 154572 265222 154624
rect 231578 154504 231584 154556
rect 231636 154544 231642 154556
rect 240134 154544 240140 154556
rect 231636 154516 240140 154544
rect 231636 154504 231642 154516
rect 240134 154504 240140 154516
rect 240192 154504 240198 154556
rect 282362 154504 282368 154556
rect 282420 154544 282426 154556
rect 313458 154544 313464 154556
rect 282420 154516 313464 154544
rect 282420 154504 282426 154516
rect 313458 154504 313464 154516
rect 313516 154504 313522 154556
rect 230658 153892 230664 153944
rect 230716 153932 230722 153944
rect 241606 153932 241612 153944
rect 230716 153904 241612 153932
rect 230716 153892 230722 153904
rect 241606 153892 241612 153904
rect 241664 153892 241670 153944
rect 241054 153824 241060 153876
rect 241112 153864 241118 153876
rect 264974 153864 264980 153876
rect 241112 153836 264980 153864
rect 241112 153824 241118 153836
rect 264974 153824 264980 153836
rect 265032 153824 265038 153876
rect 282730 153824 282736 153876
rect 282788 153864 282794 153876
rect 289906 153864 289912 153876
rect 282788 153836 289912 153864
rect 282788 153824 282794 153836
rect 289906 153824 289912 153836
rect 289964 153824 289970 153876
rect 331950 153824 331956 153876
rect 332008 153864 332014 153876
rect 385770 153864 385776 153876
rect 332008 153836 385776 153864
rect 332008 153824 332014 153836
rect 385770 153824 385776 153836
rect 385828 153824 385834 153876
rect 389910 153824 389916 153876
rect 389968 153864 389974 153876
rect 438946 153864 438952 153876
rect 389968 153836 438952 153864
rect 389968 153824 389974 153836
rect 438946 153824 438952 153836
rect 439004 153824 439010 153876
rect 211890 153280 211896 153332
rect 211948 153320 211954 153332
rect 214006 153320 214012 153332
rect 211948 153292 214012 153320
rect 211948 153280 211954 153292
rect 214006 153280 214012 153292
rect 214064 153280 214070 153332
rect 166350 153212 166356 153264
rect 166408 153252 166414 153264
rect 213914 153252 213920 153264
rect 166408 153224 213920 153252
rect 166408 153212 166414 153224
rect 213914 153212 213920 153224
rect 213972 153212 213978 153264
rect 260282 153212 260288 153264
rect 260340 153252 260346 153264
rect 264974 153252 264980 153264
rect 260340 153224 264980 153252
rect 260340 153212 260346 153224
rect 264974 153212 264980 153224
rect 265032 153212 265038 153264
rect 282822 153144 282828 153196
rect 282880 153184 282886 153196
rect 298278 153184 298284 153196
rect 282880 153156 298284 153184
rect 282880 153144 282886 153156
rect 298278 153144 298284 153156
rect 298336 153144 298342 153196
rect 230750 152464 230756 152516
rect 230808 152504 230814 152516
rect 260834 152504 260840 152516
rect 230808 152476 260840 152504
rect 230808 152464 230814 152476
rect 260834 152464 260840 152476
rect 260892 152464 260898 152516
rect 297358 152464 297364 152516
rect 297416 152504 297422 152516
rect 443178 152504 443184 152516
rect 297416 152476 443184 152504
rect 297416 152464 297422 152476
rect 443178 152464 443184 152476
rect 443236 152464 443242 152516
rect 177298 151784 177304 151836
rect 177356 151824 177362 151836
rect 213914 151824 213920 151836
rect 177356 151796 213920 151824
rect 177356 151784 177362 151796
rect 213914 151784 213920 151796
rect 213972 151784 213978 151836
rect 232590 151784 232596 151836
rect 232648 151824 232654 151836
rect 264974 151824 264980 151836
rect 232648 151796 264980 151824
rect 232648 151784 232654 151796
rect 264974 151784 264980 151796
rect 265032 151784 265038 151836
rect 246482 151104 246488 151156
rect 246540 151144 246546 151156
rect 265802 151144 265808 151156
rect 246540 151116 265808 151144
rect 246540 151104 246546 151116
rect 265802 151104 265808 151116
rect 265860 151104 265866 151156
rect 171870 151036 171876 151088
rect 171928 151076 171934 151088
rect 202230 151076 202236 151088
rect 171928 151048 202236 151076
rect 171928 151036 171934 151048
rect 202230 151036 202236 151048
rect 202288 151036 202294 151088
rect 230382 151036 230388 151088
rect 230440 151076 230446 151088
rect 249794 151076 249800 151088
rect 230440 151048 249800 151076
rect 230440 151036 230446 151048
rect 249794 151036 249800 151048
rect 249852 151036 249858 151088
rect 282730 151036 282736 151088
rect 282788 151076 282794 151088
rect 311986 151076 311992 151088
rect 282788 151048 311992 151076
rect 282788 151036 282794 151048
rect 311986 151036 311992 151048
rect 312044 151036 312050 151088
rect 374730 151036 374736 151088
rect 374788 151076 374794 151088
rect 395430 151076 395436 151088
rect 374788 151048 395436 151076
rect 374788 151036 374794 151048
rect 395430 151036 395436 151048
rect 395488 151036 395494 151088
rect 198090 150424 198096 150476
rect 198148 150464 198154 150476
rect 213914 150464 213920 150476
rect 198148 150436 213920 150464
rect 198148 150424 198154 150436
rect 213914 150424 213920 150436
rect 213972 150424 213978 150476
rect 245654 150464 245660 150476
rect 242176 150436 245660 150464
rect 174538 150356 174544 150408
rect 174596 150396 174602 150408
rect 214006 150396 214012 150408
rect 174596 150368 214012 150396
rect 174596 150356 174602 150368
rect 214006 150356 214012 150368
rect 214064 150356 214070 150408
rect 230566 150356 230572 150408
rect 230624 150396 230630 150408
rect 242176 150396 242204 150436
rect 245654 150424 245660 150436
rect 245712 150424 245718 150476
rect 252002 150424 252008 150476
rect 252060 150464 252066 150476
rect 264974 150464 264980 150476
rect 252060 150436 264980 150464
rect 252060 150424 252066 150436
rect 264974 150424 264980 150436
rect 265032 150424 265038 150476
rect 334710 150424 334716 150476
rect 334768 150464 334774 150476
rect 407206 150464 407212 150476
rect 334768 150436 407212 150464
rect 334768 150424 334774 150436
rect 407206 150424 407212 150436
rect 407264 150424 407270 150476
rect 230624 150368 242204 150396
rect 230624 150356 230630 150368
rect 281902 150356 281908 150408
rect 281960 150396 281966 150408
rect 317414 150396 317420 150408
rect 281960 150368 317420 150396
rect 281960 150356 281966 150368
rect 317414 150356 317420 150368
rect 317472 150356 317478 150408
rect 421098 150356 421104 150408
rect 421156 150396 421162 150408
rect 421558 150396 421564 150408
rect 421156 150368 421564 150396
rect 421156 150356 421162 150368
rect 421558 150356 421564 150368
rect 421616 150396 421622 150408
rect 583386 150396 583392 150408
rect 421616 150368 583392 150396
rect 421616 150356 421622 150368
rect 583386 150356 583392 150368
rect 583444 150356 583450 150408
rect 2774 150288 2780 150340
rect 2832 150328 2838 150340
rect 4798 150328 4804 150340
rect 2832 150300 4804 150328
rect 2832 150288 2838 150300
rect 4798 150288 4804 150300
rect 4856 150288 4862 150340
rect 181438 150288 181444 150340
rect 181496 150328 181502 150340
rect 213914 150328 213920 150340
rect 181496 150300 213920 150328
rect 181496 150288 181502 150300
rect 213914 150288 213920 150300
rect 213972 150288 213978 150340
rect 282822 150288 282828 150340
rect 282880 150328 282886 150340
rect 299750 150328 299756 150340
rect 282880 150300 299756 150328
rect 282880 150288 282886 150300
rect 299750 150288 299756 150300
rect 299808 150288 299814 150340
rect 231210 149676 231216 149728
rect 231268 149716 231274 149728
rect 258718 149716 258724 149728
rect 231268 149688 258724 149716
rect 231268 149676 231274 149688
rect 258718 149676 258724 149688
rect 258776 149676 258782 149728
rect 309778 149676 309784 149728
rect 309836 149716 309842 149728
rect 425790 149716 425796 149728
rect 309836 149688 425796 149716
rect 309836 149676 309842 149688
rect 425790 149676 425796 149688
rect 425848 149676 425854 149728
rect 253382 149064 253388 149116
rect 253440 149104 253446 149116
rect 264974 149104 264980 149116
rect 253440 149076 264980 149104
rect 253440 149064 253446 149076
rect 264974 149064 264980 149076
rect 265032 149064 265038 149116
rect 230566 148996 230572 149048
rect 230624 149036 230630 149048
rect 252646 149036 252652 149048
rect 230624 149008 252652 149036
rect 230624 148996 230630 149008
rect 252646 148996 252652 149008
rect 252704 148996 252710 149048
rect 282822 148996 282828 149048
rect 282880 149036 282886 149048
rect 292574 149036 292580 149048
rect 282880 149008 292580 149036
rect 282880 148996 282886 149008
rect 292574 148996 292580 149008
rect 292632 148996 292638 149048
rect 449986 148996 449992 149048
rect 450044 149036 450050 149048
rect 450538 149036 450544 149048
rect 450044 149008 450544 149036
rect 450044 148996 450050 149008
rect 450538 148996 450544 149008
rect 450596 149036 450602 149048
rect 583018 149036 583024 149048
rect 450596 149008 583024 149036
rect 450596 148996 450602 149008
rect 583018 148996 583024 149008
rect 583076 148996 583082 149048
rect 411898 148384 411904 148436
rect 411956 148424 411962 148436
rect 434070 148424 434076 148436
rect 411956 148396 434076 148424
rect 411956 148384 411962 148396
rect 434070 148384 434076 148396
rect 434128 148384 434134 148436
rect 173250 148316 173256 148368
rect 173308 148356 173314 148368
rect 186958 148356 186964 148368
rect 173308 148328 186964 148356
rect 173308 148316 173314 148328
rect 186958 148316 186964 148328
rect 187016 148316 187022 148368
rect 356698 148316 356704 148368
rect 356756 148356 356762 148368
rect 442258 148356 442264 148368
rect 356756 148328 442264 148356
rect 356756 148316 356762 148328
rect 442258 148316 442264 148328
rect 442316 148316 442322 148368
rect 256234 147704 256240 147756
rect 256292 147744 256298 147756
rect 264974 147744 264980 147756
rect 256292 147716 264980 147744
rect 256292 147704 256298 147716
rect 264974 147704 264980 147716
rect 265032 147704 265038 147756
rect 184382 147636 184388 147688
rect 184440 147676 184446 147688
rect 213914 147676 213920 147688
rect 184440 147648 213920 147676
rect 184440 147636 184446 147648
rect 213914 147636 213920 147648
rect 213972 147636 213978 147688
rect 238110 147636 238116 147688
rect 238168 147676 238174 147688
rect 265066 147676 265072 147688
rect 238168 147648 265072 147676
rect 238168 147636 238174 147648
rect 265066 147636 265072 147648
rect 265124 147636 265130 147688
rect 299382 147636 299388 147688
rect 299440 147676 299446 147688
rect 407666 147676 407672 147688
rect 299440 147648 407672 147676
rect 299440 147636 299446 147648
rect 407666 147636 407672 147648
rect 407724 147636 407730 147688
rect 580902 147636 580908 147688
rect 580960 147676 580966 147688
rect 582374 147676 582380 147688
rect 580960 147648 582380 147676
rect 580960 147636 580966 147648
rect 582374 147636 582380 147648
rect 582432 147636 582438 147688
rect 230750 147568 230756 147620
rect 230808 147608 230814 147620
rect 233510 147608 233516 147620
rect 230808 147580 233516 147608
rect 230808 147568 230814 147580
rect 233510 147568 233516 147580
rect 233568 147568 233574 147620
rect 282730 147568 282736 147620
rect 282788 147608 282794 147620
rect 323026 147608 323032 147620
rect 282788 147580 323032 147608
rect 282788 147568 282794 147580
rect 323026 147568 323032 147580
rect 323084 147568 323090 147620
rect 282822 147500 282828 147552
rect 282880 147540 282886 147552
rect 292758 147540 292764 147552
rect 282880 147512 292764 147540
rect 282880 147500 282886 147512
rect 292758 147500 292764 147512
rect 292816 147500 292822 147552
rect 233786 146956 233792 147008
rect 233844 146996 233850 147008
rect 247218 146996 247224 147008
rect 233844 146968 247224 146996
rect 233844 146956 233850 146968
rect 247218 146956 247224 146968
rect 247276 146956 247282 147008
rect 231118 146888 231124 146940
rect 231176 146928 231182 146940
rect 250714 146928 250720 146940
rect 231176 146900 250720 146928
rect 231176 146888 231182 146900
rect 250714 146888 250720 146900
rect 250772 146888 250778 146940
rect 398466 146888 398472 146940
rect 398524 146928 398530 146940
rect 583294 146928 583300 146940
rect 398524 146900 583300 146928
rect 398524 146888 398530 146900
rect 583294 146888 583300 146900
rect 583352 146888 583358 146940
rect 250622 146344 250628 146396
rect 250680 146384 250686 146396
rect 264974 146384 264980 146396
rect 250680 146356 264980 146384
rect 250680 146344 250686 146356
rect 264974 146344 264980 146356
rect 265032 146344 265038 146396
rect 178678 146276 178684 146328
rect 178736 146316 178742 146328
rect 213914 146316 213920 146328
rect 178736 146288 213920 146316
rect 178736 146276 178742 146288
rect 213914 146276 213920 146288
rect 213972 146276 213978 146328
rect 249150 146276 249156 146328
rect 249208 146316 249214 146328
rect 265066 146316 265072 146328
rect 249208 146288 265072 146316
rect 249208 146276 249214 146288
rect 265066 146276 265072 146288
rect 265124 146276 265130 146328
rect 387150 146276 387156 146328
rect 387208 146316 387214 146328
rect 436646 146316 436652 146328
rect 387208 146288 436652 146316
rect 387208 146276 387214 146288
rect 436646 146276 436652 146288
rect 436704 146276 436710 146328
rect 230658 146208 230664 146260
rect 230716 146248 230722 146260
rect 238846 146248 238852 146260
rect 230716 146220 238852 146248
rect 230716 146208 230722 146220
rect 238846 146208 238852 146220
rect 238904 146208 238910 146260
rect 282546 146208 282552 146260
rect 282604 146248 282610 146260
rect 299658 146248 299664 146260
rect 282604 146220 299664 146248
rect 282604 146208 282610 146220
rect 299658 146208 299664 146220
rect 299716 146208 299722 146260
rect 420178 146208 420184 146260
rect 420236 146248 420242 146260
rect 422938 146248 422944 146260
rect 420236 146220 422944 146248
rect 420236 146208 420242 146220
rect 422938 146208 422944 146220
rect 422996 146208 423002 146260
rect 282822 146140 282828 146192
rect 282880 146180 282886 146192
rect 294138 146180 294144 146192
rect 282880 146152 294144 146180
rect 282880 146140 282886 146152
rect 294138 146140 294144 146152
rect 294196 146140 294202 146192
rect 382918 145596 382924 145648
rect 382976 145636 382982 145648
rect 412726 145636 412732 145648
rect 382976 145608 412732 145636
rect 382976 145596 382982 145608
rect 412726 145596 412732 145608
rect 412784 145596 412790 145648
rect 231394 145528 231400 145580
rect 231452 145568 231458 145580
rect 240962 145568 240968 145580
rect 231452 145540 240968 145568
rect 231452 145528 231458 145540
rect 240962 145528 240968 145540
rect 241020 145528 241026 145580
rect 322198 145528 322204 145580
rect 322256 145568 322262 145580
rect 409966 145568 409972 145580
rect 322256 145540 409972 145568
rect 322256 145528 322262 145540
rect 409966 145528 409972 145540
rect 410024 145528 410030 145580
rect 411990 145528 411996 145580
rect 412048 145568 412054 145580
rect 422386 145568 422392 145580
rect 412048 145540 422392 145568
rect 412048 145528 412054 145540
rect 422386 145528 422392 145540
rect 422444 145528 422450 145580
rect 177390 144984 177396 145036
rect 177448 145024 177454 145036
rect 214006 145024 214012 145036
rect 177448 144996 214012 145024
rect 177448 144984 177454 144996
rect 214006 144984 214012 144996
rect 214064 144984 214070 145036
rect 243630 144984 243636 145036
rect 243688 145024 243694 145036
rect 265066 145024 265072 145036
rect 243688 144996 265072 145024
rect 243688 144984 243694 144996
rect 265066 144984 265072 144996
rect 265124 144984 265130 145036
rect 167638 144916 167644 144968
rect 167696 144956 167702 144968
rect 213914 144956 213920 144968
rect 167696 144928 213920 144956
rect 167696 144916 167702 144928
rect 213914 144916 213920 144928
rect 213972 144916 213978 144968
rect 239582 144916 239588 144968
rect 239640 144956 239646 144968
rect 264974 144956 264980 144968
rect 239640 144928 264980 144956
rect 239640 144916 239646 144928
rect 264974 144916 264980 144928
rect 265032 144916 265038 144968
rect 231762 144848 231768 144900
rect 231820 144888 231826 144900
rect 242158 144888 242164 144900
rect 231820 144860 242164 144888
rect 231820 144848 231826 144860
rect 242158 144848 242164 144860
rect 242216 144848 242222 144900
rect 282454 144848 282460 144900
rect 282512 144888 282518 144900
rect 303614 144888 303620 144900
rect 282512 144860 303620 144888
rect 282512 144848 282518 144860
rect 303614 144848 303620 144860
rect 303672 144848 303678 144900
rect 302970 144236 302976 144288
rect 303028 144276 303034 144288
rect 441982 144276 441988 144288
rect 303028 144248 441988 144276
rect 303028 144236 303034 144248
rect 441982 144236 441988 144248
rect 442040 144236 442046 144288
rect 403618 144168 403624 144220
rect 403676 144208 403682 144220
rect 419718 144208 419724 144220
rect 403676 144180 419724 144208
rect 403676 144168 403682 144180
rect 419718 144168 419724 144180
rect 419776 144168 419782 144220
rect 424686 144168 424692 144220
rect 424744 144208 424750 144220
rect 582558 144208 582564 144220
rect 424744 144180 582564 144208
rect 424744 144168 424750 144180
rect 582558 144168 582564 144180
rect 582616 144168 582622 144220
rect 246390 143624 246396 143676
rect 246448 143664 246454 143676
rect 264974 143664 264980 143676
rect 246448 143636 264980 143664
rect 246448 143624 246454 143636
rect 264974 143624 264980 143636
rect 265032 143624 265038 143676
rect 180242 143556 180248 143608
rect 180300 143596 180306 143608
rect 213914 143596 213920 143608
rect 180300 143568 213920 143596
rect 180300 143556 180306 143568
rect 213914 143556 213920 143568
rect 213972 143556 213978 143608
rect 240962 143556 240968 143608
rect 241020 143596 241026 143608
rect 265066 143596 265072 143608
rect 241020 143568 265072 143596
rect 241020 143556 241026 143568
rect 265066 143556 265072 143568
rect 265124 143556 265130 143608
rect 329098 143488 329104 143540
rect 329156 143528 329162 143540
rect 330478 143528 330484 143540
rect 329156 143500 330484 143528
rect 329156 143488 329162 143500
rect 330478 143488 330484 143500
rect 330536 143488 330542 143540
rect 407206 143488 407212 143540
rect 407264 143528 407270 143540
rect 408862 143528 408868 143540
rect 407264 143500 408868 143528
rect 407264 143488 407270 143500
rect 408862 143488 408868 143500
rect 408920 143488 408926 143540
rect 410518 143488 410524 143540
rect 410576 143528 410582 143540
rect 411990 143528 411996 143540
rect 410576 143500 411996 143528
rect 410576 143488 410582 143500
rect 411990 143488 411996 143500
rect 412048 143488 412054 143540
rect 414750 143488 414756 143540
rect 414808 143528 414814 143540
rect 416406 143528 416412 143540
rect 414808 143500 416412 143528
rect 414808 143488 414814 143500
rect 416406 143488 416412 143500
rect 416464 143488 416470 143540
rect 430574 143488 430580 143540
rect 430632 143528 430638 143540
rect 431310 143528 431316 143540
rect 430632 143500 431316 143528
rect 430632 143488 430638 143500
rect 431310 143488 431316 143500
rect 431368 143488 431374 143540
rect 231762 143420 231768 143472
rect 231820 143460 231826 143472
rect 236638 143460 236644 143472
rect 231820 143432 236644 143460
rect 231820 143420 231826 143432
rect 236638 143420 236644 143432
rect 236696 143420 236702 143472
rect 413278 143420 413284 143472
rect 413336 143460 413342 143472
rect 418430 143460 418436 143472
rect 413336 143432 418436 143460
rect 413336 143420 413342 143432
rect 418430 143420 418436 143432
rect 418488 143420 418494 143472
rect 237006 142808 237012 142860
rect 237064 142848 237070 142860
rect 265618 142848 265624 142860
rect 237064 142820 265624 142848
rect 237064 142808 237070 142820
rect 265618 142808 265624 142820
rect 265676 142808 265682 142860
rect 415854 142808 415860 142860
rect 415912 142848 415918 142860
rect 416774 142848 416780 142860
rect 415912 142820 416780 142848
rect 415912 142808 415918 142820
rect 416774 142808 416780 142820
rect 416832 142808 416838 142860
rect 438670 142808 438676 142860
rect 438728 142848 438734 142860
rect 449986 142848 449992 142860
rect 438728 142820 449992 142848
rect 438728 142808 438734 142820
rect 449986 142808 449992 142820
rect 450044 142808 450050 142860
rect 282822 142400 282828 142452
rect 282880 142440 282886 142452
rect 287330 142440 287336 142452
rect 282880 142412 287336 142440
rect 282880 142400 282886 142412
rect 287330 142400 287336 142412
rect 287388 142400 287394 142452
rect 209222 142196 209228 142248
rect 209280 142236 209286 142248
rect 213914 142236 213920 142248
rect 209280 142208 213920 142236
rect 209280 142196 209286 142208
rect 213914 142196 213920 142208
rect 213972 142196 213978 142248
rect 171778 142128 171784 142180
rect 171836 142168 171842 142180
rect 214006 142168 214012 142180
rect 171836 142140 214012 142168
rect 171836 142128 171842 142140
rect 214006 142128 214012 142140
rect 214064 142128 214070 142180
rect 232498 142128 232504 142180
rect 232556 142168 232562 142180
rect 264974 142168 264980 142180
rect 232556 142140 264980 142168
rect 232556 142128 232562 142140
rect 264974 142128 264980 142140
rect 265032 142128 265038 142180
rect 381538 142128 381544 142180
rect 381596 142168 381602 142180
rect 405182 142168 405188 142180
rect 381596 142140 405188 142168
rect 381596 142128 381602 142140
rect 405182 142128 405188 142140
rect 405240 142128 405246 142180
rect 418798 142128 418804 142180
rect 418856 142168 418862 142180
rect 424134 142168 424140 142180
rect 418856 142140 424140 142168
rect 418856 142128 418862 142140
rect 424134 142128 424140 142140
rect 424192 142128 424198 142180
rect 425698 142128 425704 142180
rect 425756 142168 425762 142180
rect 433518 142168 433524 142180
rect 425756 142140 433524 142168
rect 425756 142128 425762 142140
rect 433518 142128 433524 142140
rect 433576 142128 433582 142180
rect 434070 142128 434076 142180
rect 434128 142168 434134 142180
rect 583018 142168 583024 142180
rect 434128 142140 583024 142168
rect 434128 142128 434134 142140
rect 583018 142128 583024 142140
rect 583076 142128 583082 142180
rect 282822 142060 282828 142112
rect 282880 142100 282886 142112
rect 313274 142100 313280 142112
rect 282880 142072 313280 142100
rect 282880 142060 282886 142072
rect 313274 142060 313280 142072
rect 313332 142060 313338 142112
rect 374638 142060 374644 142112
rect 374696 142100 374702 142112
rect 376754 142100 376760 142112
rect 374696 142072 376760 142100
rect 374696 142060 374702 142072
rect 376754 142060 376760 142072
rect 376812 142060 376818 142112
rect 282730 141992 282736 142044
rect 282788 142032 282794 142044
rect 295426 142032 295432 142044
rect 282788 142004 295432 142032
rect 282788 141992 282794 142004
rect 295426 141992 295432 142004
rect 295484 141992 295490 142044
rect 249334 141448 249340 141500
rect 249392 141488 249398 141500
rect 265986 141488 265992 141500
rect 249392 141460 265992 141488
rect 249392 141448 249398 141460
rect 265986 141448 265992 141460
rect 266044 141448 266050 141500
rect 181530 141380 181536 141432
rect 181588 141420 181594 141432
rect 214650 141420 214656 141432
rect 181588 141392 214656 141420
rect 181588 141380 181594 141392
rect 214650 141380 214656 141392
rect 214708 141380 214714 141432
rect 231578 141380 231584 141432
rect 231636 141420 231642 141432
rect 251818 141420 251824 141432
rect 231636 141392 251824 141420
rect 231636 141380 231642 141392
rect 251818 141380 251824 141392
rect 251876 141380 251882 141432
rect 383102 140836 383108 140888
rect 383160 140876 383166 140888
rect 417142 140876 417148 140888
rect 383160 140848 417148 140876
rect 383160 140836 383166 140848
rect 417142 140836 417148 140848
rect 417200 140836 417206 140888
rect 425422 140836 425428 140888
rect 425480 140876 425486 140888
rect 425790 140876 425796 140888
rect 425480 140848 425796 140876
rect 425480 140836 425486 140848
rect 425790 140836 425796 140848
rect 425848 140876 425854 140888
rect 464338 140876 464344 140888
rect 425848 140848 464344 140876
rect 425848 140836 425854 140848
rect 464338 140836 464344 140848
rect 464396 140836 464402 140888
rect 205266 140768 205272 140820
rect 205324 140808 205330 140820
rect 213914 140808 213920 140820
rect 205324 140780 213920 140808
rect 205324 140768 205330 140780
rect 213914 140768 213920 140780
rect 213972 140768 213978 140820
rect 261662 140768 261668 140820
rect 261720 140808 261726 140820
rect 264974 140808 264980 140820
rect 261720 140780 264980 140808
rect 261720 140768 261726 140780
rect 264974 140768 264980 140780
rect 265032 140768 265038 140820
rect 303614 140768 303620 140820
rect 303672 140808 303678 140820
rect 409598 140808 409604 140820
rect 303672 140780 409604 140808
rect 303672 140768 303678 140780
rect 409598 140768 409604 140780
rect 409656 140768 409662 140820
rect 428550 140768 428556 140820
rect 428608 140808 428614 140820
rect 582650 140808 582656 140820
rect 428608 140780 582656 140808
rect 428608 140768 428614 140780
rect 582650 140768 582656 140780
rect 582708 140768 582714 140820
rect 282822 140700 282828 140752
rect 282880 140740 282886 140752
rect 289814 140740 289820 140752
rect 282880 140712 289820 140740
rect 282880 140700 282886 140712
rect 289814 140700 289820 140712
rect 289872 140700 289878 140752
rect 405734 140700 405740 140752
rect 405792 140740 405798 140752
rect 406654 140740 406660 140752
rect 405792 140712 406660 140740
rect 405792 140700 405798 140712
rect 406654 140700 406660 140712
rect 406712 140700 406718 140752
rect 412634 140700 412640 140752
rect 412692 140740 412698 140752
rect 412910 140740 412916 140752
rect 412692 140712 412916 140740
rect 412692 140700 412698 140712
rect 412910 140700 412916 140712
rect 412968 140700 412974 140752
rect 400214 140292 400220 140344
rect 400272 140332 400278 140344
rect 401318 140332 401324 140344
rect 400272 140304 401324 140332
rect 400272 140292 400278 140304
rect 401318 140292 401324 140304
rect 401376 140292 401382 140344
rect 234154 140088 234160 140140
rect 234212 140128 234218 140140
rect 243814 140128 243820 140140
rect 234212 140100 243820 140128
rect 234212 140088 234218 140100
rect 243814 140088 243820 140100
rect 243872 140088 243878 140140
rect 242526 140020 242532 140072
rect 242584 140060 242590 140072
rect 264330 140060 264336 140072
rect 242584 140032 264336 140060
rect 242584 140020 242590 140032
rect 264330 140020 264336 140032
rect 264388 140020 264394 140072
rect 417418 140020 417424 140072
rect 417476 140060 417482 140072
rect 441706 140060 441712 140072
rect 417476 140032 441712 140060
rect 417476 140020 417482 140032
rect 441706 140020 441712 140032
rect 441764 140020 441770 140072
rect 417326 139652 417332 139664
rect 393286 139624 417332 139652
rect 342898 139476 342904 139528
rect 342956 139516 342962 139528
rect 393286 139516 393314 139624
rect 417326 139612 417332 139624
rect 417384 139612 417390 139664
rect 401502 139544 401508 139596
rect 401560 139584 401566 139596
rect 401560 139556 407712 139584
rect 401560 139544 401566 139556
rect 342956 139488 393314 139516
rect 342956 139476 342962 139488
rect 170398 139408 170404 139460
rect 170456 139448 170462 139460
rect 213914 139448 213920 139460
rect 170456 139420 213920 139448
rect 170456 139408 170462 139420
rect 213914 139408 213920 139420
rect 213972 139408 213978 139460
rect 254578 139408 254584 139460
rect 254636 139448 254642 139460
rect 264974 139448 264980 139460
rect 254636 139420 264980 139448
rect 254636 139408 254642 139420
rect 264974 139408 264980 139420
rect 265032 139408 265038 139460
rect 399478 139408 399484 139460
rect 399536 139448 399542 139460
rect 402974 139448 402980 139460
rect 399536 139420 402980 139448
rect 399536 139408 399542 139420
rect 402974 139408 402980 139420
rect 403032 139408 403038 139460
rect 407684 139448 407712 139556
rect 580166 139448 580172 139460
rect 407684 139420 580172 139448
rect 580166 139408 580172 139420
rect 580224 139408 580230 139460
rect 231762 139340 231768 139392
rect 231820 139380 231826 139392
rect 254026 139380 254032 139392
rect 231820 139352 254032 139380
rect 231820 139340 231826 139352
rect 254026 139340 254032 139352
rect 254084 139340 254090 139392
rect 282638 139340 282644 139392
rect 282696 139380 282702 139392
rect 301130 139380 301136 139392
rect 282696 139352 301136 139380
rect 282696 139340 282702 139352
rect 301130 139340 301136 139352
rect 301188 139340 301194 139392
rect 395430 139340 395436 139392
rect 395488 139380 395494 139392
rect 397546 139380 397552 139392
rect 395488 139352 397552 139380
rect 395488 139340 395494 139352
rect 397546 139340 397552 139352
rect 397604 139340 397610 139392
rect 399846 139340 399852 139392
rect 399904 139380 399910 139392
rect 404078 139380 404084 139392
rect 399904 139352 404084 139380
rect 399904 139340 399910 139352
rect 404078 139340 404084 139352
rect 404136 139340 404142 139392
rect 442166 139340 442172 139392
rect 442224 139380 442230 139392
rect 460934 139380 460940 139392
rect 442224 139352 460940 139380
rect 442224 139340 442230 139352
rect 460934 139340 460940 139352
rect 460992 139380 460998 139392
rect 583478 139380 583484 139392
rect 460992 139352 583484 139380
rect 460992 139340 460998 139352
rect 583478 139340 583484 139352
rect 583536 139340 583542 139392
rect 281718 138932 281724 138984
rect 281776 138972 281782 138984
rect 284570 138972 284576 138984
rect 281776 138944 284576 138972
rect 281776 138932 281782 138944
rect 284570 138932 284576 138944
rect 284628 138932 284634 138984
rect 169110 138660 169116 138712
rect 169168 138700 169174 138712
rect 214374 138700 214380 138712
rect 169168 138672 214380 138700
rect 169168 138660 169174 138672
rect 214374 138660 214380 138672
rect 214432 138660 214438 138712
rect 195422 137980 195428 138032
rect 195480 138020 195486 138032
rect 213914 138020 213920 138032
rect 195480 137992 213920 138020
rect 195480 137980 195486 137992
rect 213914 137980 213920 137992
rect 213972 137980 213978 138032
rect 229830 137980 229836 138032
rect 229888 138020 229894 138032
rect 264974 138020 264980 138032
rect 229888 137992 264980 138020
rect 229888 137980 229894 137992
rect 264974 137980 264980 137992
rect 265032 137980 265038 138032
rect 3510 137912 3516 137964
rect 3568 137952 3574 137964
rect 22738 137952 22744 137964
rect 3568 137924 22744 137952
rect 3568 137912 3574 137924
rect 22738 137912 22744 137924
rect 22796 137912 22802 137964
rect 231762 137912 231768 137964
rect 231820 137952 231826 137964
rect 244366 137952 244372 137964
rect 231820 137924 244372 137952
rect 231820 137912 231826 137924
rect 244366 137912 244372 137924
rect 244424 137912 244430 137964
rect 282822 137912 282828 137964
rect 282880 137952 282886 137964
rect 306374 137952 306380 137964
rect 282880 137924 306380 137952
rect 282880 137912 282886 137924
rect 306374 137912 306380 137924
rect 306432 137912 306438 137964
rect 442902 137232 442908 137284
rect 442960 137272 442966 137284
rect 447134 137272 447140 137284
rect 442960 137244 447140 137272
rect 442960 137232 442966 137244
rect 447134 137232 447140 137244
rect 447192 137272 447198 137284
rect 582558 137272 582564 137284
rect 447192 137244 582564 137272
rect 447192 137232 447198 137244
rect 582558 137232 582564 137244
rect 582616 137232 582622 137284
rect 187142 136620 187148 136672
rect 187200 136660 187206 136672
rect 213914 136660 213920 136672
rect 187200 136632 213920 136660
rect 187200 136620 187206 136632
rect 213914 136620 213920 136632
rect 213972 136620 213978 136672
rect 258718 136620 258724 136672
rect 258776 136660 258782 136672
rect 264974 136660 264980 136672
rect 258776 136632 264980 136660
rect 258776 136620 258782 136632
rect 264974 136620 264980 136632
rect 265032 136620 265038 136672
rect 395614 136620 395620 136672
rect 395672 136660 395678 136672
rect 397914 136660 397920 136672
rect 395672 136632 397920 136660
rect 395672 136620 395678 136632
rect 397914 136620 397920 136632
rect 397972 136620 397978 136672
rect 230566 136552 230572 136604
rect 230624 136592 230630 136604
rect 245838 136592 245844 136604
rect 230624 136564 245844 136592
rect 230624 136552 230630 136564
rect 245838 136552 245844 136564
rect 245896 136552 245902 136604
rect 282822 136552 282828 136604
rect 282880 136592 282886 136604
rect 292666 136592 292672 136604
rect 282880 136564 292672 136592
rect 282880 136552 282886 136564
rect 292666 136552 292672 136564
rect 292724 136552 292730 136604
rect 231302 136144 231308 136196
rect 231360 136184 231366 136196
rect 236730 136184 236736 136196
rect 231360 136156 236736 136184
rect 231360 136144 231366 136156
rect 236730 136144 236736 136156
rect 236788 136144 236794 136196
rect 196710 135940 196716 135992
rect 196768 135980 196774 135992
rect 214006 135980 214012 135992
rect 196768 135952 214012 135980
rect 196768 135940 196774 135952
rect 214006 135940 214012 135952
rect 214064 135940 214070 135992
rect 167730 135872 167736 135924
rect 167788 135912 167794 135924
rect 213362 135912 213368 135924
rect 167788 135884 213368 135912
rect 167788 135872 167794 135884
rect 213362 135872 213368 135884
rect 213420 135872 213426 135924
rect 282270 135872 282276 135924
rect 282328 135912 282334 135924
rect 327166 135912 327172 135924
rect 282328 135884 327172 135912
rect 282328 135872 282334 135884
rect 327166 135872 327172 135884
rect 327224 135872 327230 135924
rect 331950 135872 331956 135924
rect 332008 135912 332014 135924
rect 387150 135912 387156 135924
rect 332008 135884 387156 135912
rect 332008 135872 332014 135884
rect 387150 135872 387156 135884
rect 387208 135872 387214 135924
rect 442902 135464 442908 135516
rect 442960 135504 442966 135516
rect 448698 135504 448704 135516
rect 442960 135476 448704 135504
rect 442960 135464 442966 135476
rect 448698 135464 448704 135476
rect 448756 135464 448762 135516
rect 258810 135328 258816 135380
rect 258868 135368 258874 135380
rect 265066 135368 265072 135380
rect 258868 135340 265072 135368
rect 258868 135328 258874 135340
rect 265066 135328 265072 135340
rect 265124 135328 265130 135380
rect 388530 135328 388536 135380
rect 388588 135368 388594 135380
rect 397638 135368 397644 135380
rect 388588 135340 397644 135368
rect 388588 135328 388594 135340
rect 397638 135328 397644 135340
rect 397696 135328 397702 135380
rect 231302 135260 231308 135312
rect 231360 135300 231366 135312
rect 231578 135300 231584 135312
rect 231360 135272 231584 135300
rect 231360 135260 231366 135272
rect 231578 135260 231584 135272
rect 231636 135260 231642 135312
rect 260190 135260 260196 135312
rect 260248 135300 260254 135312
rect 264974 135300 264980 135312
rect 260248 135272 264980 135300
rect 260248 135260 260254 135272
rect 264974 135260 264980 135272
rect 265032 135260 265038 135312
rect 374730 135260 374736 135312
rect 374788 135300 374794 135312
rect 397546 135300 397552 135312
rect 374788 135272 397552 135300
rect 374788 135260 374794 135272
rect 397546 135260 397552 135272
rect 397604 135260 397610 135312
rect 231486 135192 231492 135244
rect 231544 135232 231550 135244
rect 258994 135232 259000 135244
rect 231544 135204 259000 135232
rect 231544 135192 231550 135204
rect 258994 135192 259000 135204
rect 259052 135192 259058 135244
rect 282822 135192 282828 135244
rect 282880 135232 282886 135244
rect 318794 135232 318800 135244
rect 282880 135204 318800 135232
rect 282880 135192 282886 135204
rect 318794 135192 318800 135204
rect 318852 135192 318858 135244
rect 231762 135124 231768 135176
rect 231820 135164 231826 135176
rect 249242 135164 249248 135176
rect 231820 135136 249248 135164
rect 231820 135124 231826 135136
rect 249242 135124 249248 135136
rect 249300 135124 249306 135176
rect 282454 134920 282460 134972
rect 282512 134960 282518 134972
rect 285858 134960 285864 134972
rect 282512 134932 285864 134960
rect 282512 134920 282518 134932
rect 285858 134920 285864 134932
rect 285916 134920 285922 134972
rect 169202 134512 169208 134564
rect 169260 134552 169266 134564
rect 214098 134552 214104 134564
rect 169260 134524 214104 134552
rect 169260 134512 169266 134524
rect 214098 134512 214104 134524
rect 214156 134512 214162 134564
rect 363598 134512 363604 134564
rect 363656 134552 363662 134564
rect 381630 134552 381636 134564
rect 363656 134524 381636 134552
rect 363656 134512 363662 134524
rect 381630 134512 381636 134524
rect 381688 134512 381694 134564
rect 210418 133900 210424 133952
rect 210476 133940 210482 133952
rect 213914 133940 213920 133952
rect 210476 133912 213920 133940
rect 210476 133900 210482 133912
rect 213914 133900 213920 133912
rect 213972 133900 213978 133952
rect 378870 133900 378876 133952
rect 378928 133940 378934 133952
rect 397638 133940 397644 133952
rect 378928 133912 397644 133940
rect 378928 133900 378934 133912
rect 397638 133900 397644 133912
rect 397696 133900 397702 133952
rect 231486 133832 231492 133884
rect 231544 133872 231550 133884
rect 254670 133872 254676 133884
rect 231544 133844 254676 133872
rect 231544 133832 231550 133844
rect 254670 133832 254676 133844
rect 254728 133832 254734 133884
rect 444374 133832 444380 133884
rect 444432 133872 444438 133884
rect 448606 133872 448612 133884
rect 444432 133844 448612 133872
rect 444432 133832 444438 133844
rect 448606 133832 448612 133844
rect 448664 133832 448670 133884
rect 442902 133220 442908 133272
rect 442960 133260 442966 133272
rect 444374 133260 444380 133272
rect 442960 133232 444380 133260
rect 442960 133220 442966 133232
rect 444374 133220 444380 133232
rect 444432 133220 444438 133272
rect 230658 133152 230664 133204
rect 230716 133192 230722 133204
rect 256050 133192 256056 133204
rect 230716 133164 256056 133192
rect 230716 133152 230722 133164
rect 256050 133152 256056 133164
rect 256108 133152 256114 133204
rect 358170 133152 358176 133204
rect 358228 133192 358234 133204
rect 391198 133192 391204 133204
rect 358228 133164 391204 133192
rect 358228 133152 358234 133164
rect 391198 133152 391204 133164
rect 391256 133152 391262 133204
rect 209130 132540 209136 132592
rect 209188 132580 209194 132592
rect 213914 132580 213920 132592
rect 209188 132552 213920 132580
rect 209188 132540 209194 132552
rect 213914 132540 213920 132552
rect 213972 132540 213978 132592
rect 192662 132472 192668 132524
rect 192720 132512 192726 132524
rect 214006 132512 214012 132524
rect 192720 132484 214012 132512
rect 192720 132472 192726 132484
rect 214006 132472 214012 132484
rect 214064 132472 214070 132524
rect 255958 132472 255964 132524
rect 256016 132512 256022 132524
rect 264974 132512 264980 132524
rect 256016 132484 264980 132512
rect 256016 132472 256022 132484
rect 264974 132472 264980 132484
rect 265032 132472 265038 132524
rect 392762 132472 392768 132524
rect 392820 132512 392826 132524
rect 397546 132512 397552 132524
rect 392820 132484 397552 132512
rect 392820 132472 392826 132484
rect 397546 132472 397552 132484
rect 397604 132472 397610 132524
rect 231762 132404 231768 132456
rect 231820 132444 231826 132456
rect 247954 132444 247960 132456
rect 231820 132416 247960 132444
rect 231820 132404 231826 132416
rect 247954 132404 247960 132416
rect 248012 132404 248018 132456
rect 282822 132404 282828 132456
rect 282880 132444 282886 132456
rect 324314 132444 324320 132456
rect 282880 132416 324320 132444
rect 282880 132404 282886 132416
rect 324314 132404 324320 132416
rect 324372 132404 324378 132456
rect 371878 132404 371884 132456
rect 371936 132444 371942 132456
rect 398466 132444 398472 132456
rect 371936 132416 398472 132444
rect 371936 132404 371942 132416
rect 398466 132404 398472 132416
rect 398524 132404 398530 132456
rect 442902 132404 442908 132456
rect 442960 132444 442966 132456
rect 583754 132444 583760 132456
rect 442960 132416 583760 132444
rect 442960 132404 442966 132416
rect 583754 132404 583760 132416
rect 583812 132404 583818 132456
rect 181438 131724 181444 131776
rect 181496 131764 181502 131776
rect 211890 131764 211896 131776
rect 181496 131736 211896 131764
rect 181496 131724 181502 131736
rect 211890 131724 211896 131736
rect 211948 131724 211954 131776
rect 305730 131724 305736 131776
rect 305788 131764 305794 131776
rect 327074 131764 327080 131776
rect 305788 131736 327080 131764
rect 305788 131724 305794 131736
rect 327074 131724 327080 131736
rect 327132 131764 327138 131776
rect 395614 131764 395620 131776
rect 327132 131736 395620 131764
rect 327132 131724 327138 131736
rect 395614 131724 395620 131736
rect 395672 131724 395678 131776
rect 231394 131656 231400 131708
rect 231452 131696 231458 131708
rect 234154 131696 234160 131708
rect 231452 131668 234160 131696
rect 231452 131656 231458 131668
rect 234154 131656 234160 131668
rect 234212 131656 234218 131708
rect 251818 131180 251824 131232
rect 251876 131220 251882 131232
rect 264974 131220 264980 131232
rect 251876 131192 264980 131220
rect 251876 131180 251882 131192
rect 264974 131180 264980 131192
rect 265032 131180 265038 131232
rect 185670 131112 185676 131164
rect 185728 131152 185734 131164
rect 213914 131152 213920 131164
rect 185728 131124 213920 131152
rect 185728 131112 185734 131124
rect 213914 131112 213920 131124
rect 213972 131112 213978 131164
rect 247678 131112 247684 131164
rect 247736 131152 247742 131164
rect 265066 131152 265072 131164
rect 247736 131124 265072 131152
rect 247736 131112 247742 131124
rect 265066 131112 265072 131124
rect 265124 131112 265130 131164
rect 231762 131044 231768 131096
rect 231820 131084 231826 131096
rect 264238 131084 264244 131096
rect 231820 131056 264244 131084
rect 231820 131044 231826 131056
rect 264238 131044 264244 131056
rect 264296 131044 264302 131096
rect 282270 131044 282276 131096
rect 282328 131084 282334 131096
rect 310606 131084 310612 131096
rect 282328 131056 310612 131084
rect 282328 131044 282334 131056
rect 310606 131044 310612 131056
rect 310664 131044 310670 131096
rect 231118 130976 231124 131028
rect 231176 131016 231182 131028
rect 260098 131016 260104 131028
rect 231176 130988 260104 131016
rect 231176 130976 231182 130988
rect 260098 130976 260104 130988
rect 260156 130976 260162 131028
rect 282638 130976 282644 131028
rect 282696 131016 282702 131028
rect 307846 131016 307852 131028
rect 282696 130988 307852 131016
rect 282696 130976 282702 130988
rect 307846 130976 307852 130988
rect 307904 130976 307910 131028
rect 192570 130364 192576 130416
rect 192628 130404 192634 130416
rect 206462 130404 206468 130416
rect 192628 130376 206468 130404
rect 192628 130364 192634 130376
rect 206462 130364 206468 130376
rect 206520 130364 206526 130416
rect 210510 129820 210516 129872
rect 210568 129860 210574 129872
rect 214006 129860 214012 129872
rect 210568 129832 214012 129860
rect 210568 129820 210574 129832
rect 214006 129820 214012 129832
rect 214064 129820 214070 129872
rect 200850 129752 200856 129804
rect 200908 129792 200914 129804
rect 213914 129792 213920 129804
rect 200908 129764 213920 129792
rect 200908 129752 200914 129764
rect 213914 129752 213920 129764
rect 213972 129752 213978 129804
rect 389910 129752 389916 129804
rect 389968 129792 389974 129804
rect 398834 129792 398840 129804
rect 389968 129764 398840 129792
rect 389968 129752 389974 129764
rect 398834 129752 398840 129764
rect 398892 129752 398898 129804
rect 230750 129684 230756 129736
rect 230808 129724 230814 129736
rect 240778 129724 240784 129736
rect 230808 129696 240784 129724
rect 230808 129684 230814 129696
rect 240778 129684 240784 129696
rect 240836 129684 240842 129736
rect 370498 129684 370504 129736
rect 370556 129724 370562 129736
rect 372614 129724 372620 129736
rect 370556 129696 372620 129724
rect 370556 129684 370562 129696
rect 372614 129684 372620 129696
rect 372672 129724 372678 129736
rect 397546 129724 397552 129736
rect 372672 129696 397552 129724
rect 372672 129684 372678 129696
rect 397546 129684 397552 129696
rect 397604 129684 397610 129736
rect 318242 129004 318248 129056
rect 318300 129044 318306 129056
rect 398190 129044 398196 129056
rect 318300 129016 398196 129044
rect 318300 129004 318306 129016
rect 398190 129004 398196 129016
rect 398248 129004 398254 129056
rect 205174 128392 205180 128444
rect 205232 128432 205238 128444
rect 213914 128432 213920 128444
rect 205232 128404 213920 128432
rect 205232 128392 205238 128404
rect 213914 128392 213920 128404
rect 213972 128392 213978 128444
rect 264974 128432 264980 128444
rect 258046 128404 264980 128432
rect 202414 128324 202420 128376
rect 202472 128364 202478 128376
rect 214006 128364 214012 128376
rect 202472 128336 214012 128364
rect 202472 128324 202478 128336
rect 214006 128324 214012 128336
rect 214064 128324 214070 128376
rect 254854 128324 254860 128376
rect 254912 128364 254918 128376
rect 258046 128364 258074 128404
rect 264974 128392 264980 128404
rect 265032 128392 265038 128444
rect 254912 128336 258074 128364
rect 254912 128324 254918 128336
rect 264606 128324 264612 128376
rect 264664 128364 264670 128376
rect 265710 128364 265716 128376
rect 264664 128336 265716 128364
rect 264664 128324 264670 128336
rect 265710 128324 265716 128336
rect 265768 128324 265774 128376
rect 231762 128256 231768 128308
rect 231820 128296 231826 128308
rect 252094 128296 252100 128308
rect 231820 128268 252100 128296
rect 231820 128256 231826 128268
rect 252094 128256 252100 128268
rect 252152 128256 252158 128308
rect 340230 128256 340236 128308
rect 340288 128296 340294 128308
rect 397546 128296 397552 128308
rect 340288 128268 397552 128296
rect 340288 128256 340294 128268
rect 397546 128256 397552 128268
rect 397604 128256 397610 128308
rect 231670 128188 231676 128240
rect 231728 128228 231734 128240
rect 236822 128228 236828 128240
rect 231728 128200 236828 128228
rect 231728 128188 231734 128200
rect 236822 128188 236828 128200
rect 236880 128188 236886 128240
rect 282822 128188 282828 128240
rect 282880 128228 282886 128240
rect 316034 128228 316040 128240
rect 282880 128200 316040 128228
rect 282880 128188 282886 128200
rect 316034 128188 316040 128200
rect 316092 128188 316098 128240
rect 182910 127576 182916 127628
rect 182968 127616 182974 127628
rect 214834 127616 214840 127628
rect 182968 127588 214840 127616
rect 182968 127576 182974 127588
rect 214834 127576 214840 127588
rect 214892 127576 214898 127628
rect 442902 127576 442908 127628
rect 442960 127616 442966 127628
rect 449986 127616 449992 127628
rect 442960 127588 449992 127616
rect 442960 127576 442966 127588
rect 449986 127576 449992 127588
rect 450044 127576 450050 127628
rect 261570 127032 261576 127084
rect 261628 127072 261634 127084
rect 265066 127072 265072 127084
rect 261628 127044 265072 127072
rect 261628 127032 261634 127044
rect 265066 127032 265072 127044
rect 265124 127032 265130 127084
rect 62022 126964 62028 127016
rect 62080 127004 62086 127016
rect 65518 127004 65524 127016
rect 62080 126976 65524 127004
rect 62080 126964 62086 126976
rect 65518 126964 65524 126976
rect 65576 126964 65582 127016
rect 197998 126964 198004 127016
rect 198056 127004 198062 127016
rect 213914 127004 213920 127016
rect 198056 126976 213920 127004
rect 198056 126964 198062 126976
rect 213914 126964 213920 126976
rect 213972 126964 213978 127016
rect 236730 126964 236736 127016
rect 236788 127004 236794 127016
rect 264974 127004 264980 127016
rect 236788 126976 264980 127004
rect 236788 126964 236794 126976
rect 264974 126964 264980 126976
rect 265032 126964 265038 127016
rect 363598 126964 363604 127016
rect 363656 127004 363662 127016
rect 397546 127004 397552 127016
rect 363656 126976 397552 127004
rect 363656 126964 363662 126976
rect 397546 126964 397552 126976
rect 397604 126964 397610 127016
rect 231302 126896 231308 126948
rect 231360 126936 231366 126948
rect 250438 126936 250444 126948
rect 231360 126908 250444 126936
rect 231360 126896 231366 126908
rect 250438 126896 250444 126908
rect 250496 126896 250502 126948
rect 263042 126896 263048 126948
rect 263100 126936 263106 126948
rect 266078 126936 266084 126948
rect 263100 126908 266084 126936
rect 263100 126896 263106 126908
rect 266078 126896 266084 126908
rect 266136 126896 266142 126948
rect 282822 126896 282828 126948
rect 282880 126936 282886 126948
rect 291194 126936 291200 126948
rect 282880 126908 291200 126936
rect 282880 126896 282886 126908
rect 291194 126896 291200 126908
rect 291252 126896 291258 126948
rect 464338 126896 464344 126948
rect 464396 126936 464402 126948
rect 580166 126936 580172 126948
rect 464396 126908 580172 126936
rect 464396 126896 464402 126908
rect 580166 126896 580172 126908
rect 580224 126896 580230 126948
rect 230566 126692 230572 126744
rect 230624 126732 230630 126744
rect 232774 126732 232780 126744
rect 230624 126704 232780 126732
rect 230624 126692 230630 126704
rect 232774 126692 232780 126704
rect 232832 126692 232838 126744
rect 166442 126216 166448 126268
rect 166500 126256 166506 126268
rect 213270 126256 213276 126268
rect 166500 126228 213276 126256
rect 166500 126216 166506 126228
rect 213270 126216 213276 126228
rect 213328 126216 213334 126268
rect 238386 126216 238392 126268
rect 238444 126256 238450 126268
rect 245286 126256 245292 126268
rect 238444 126228 245292 126256
rect 238444 126216 238450 126228
rect 245286 126216 245292 126228
rect 245344 126216 245350 126268
rect 282086 126216 282092 126268
rect 282144 126256 282150 126268
rect 313366 126256 313372 126268
rect 282144 126228 313372 126256
rect 282144 126216 282150 126228
rect 313366 126216 313372 126228
rect 313424 126216 313430 126268
rect 353938 126216 353944 126268
rect 353996 126256 354002 126268
rect 354582 126256 354588 126268
rect 353996 126228 354588 126256
rect 353996 126216 354002 126228
rect 354582 126216 354588 126228
rect 354640 126256 354646 126268
rect 397546 126256 397552 126268
rect 354640 126228 397552 126256
rect 354640 126216 354646 126228
rect 397546 126216 397552 126228
rect 397604 126216 397610 126268
rect 195514 125604 195520 125656
rect 195572 125644 195578 125656
rect 213914 125644 213920 125656
rect 195572 125616 213920 125644
rect 195572 125604 195578 125616
rect 213914 125604 213920 125616
rect 213972 125604 213978 125656
rect 245102 125604 245108 125656
rect 245160 125644 245166 125656
rect 264974 125644 264980 125656
rect 245160 125616 264980 125644
rect 245160 125604 245166 125616
rect 264974 125604 264980 125616
rect 265032 125604 265038 125656
rect 442902 125604 442908 125656
rect 442960 125644 442966 125656
rect 454034 125644 454040 125656
rect 442960 125616 454040 125644
rect 442960 125604 442966 125616
rect 454034 125604 454040 125616
rect 454092 125604 454098 125656
rect 230750 125536 230756 125588
rect 230808 125576 230814 125588
rect 238294 125576 238300 125588
rect 230808 125548 238300 125576
rect 230808 125536 230814 125548
rect 238294 125536 238300 125548
rect 238352 125536 238358 125588
rect 281626 125536 281632 125588
rect 281684 125576 281690 125588
rect 303706 125576 303712 125588
rect 281684 125548 303712 125576
rect 281684 125536 281690 125548
rect 303706 125536 303712 125548
rect 303764 125536 303770 125588
rect 315298 125536 315304 125588
rect 315356 125576 315362 125588
rect 397638 125576 397644 125588
rect 315356 125548 397644 125576
rect 315356 125536 315362 125548
rect 397638 125536 397644 125548
rect 397696 125536 397702 125588
rect 392670 125468 392676 125520
rect 392728 125508 392734 125520
rect 397546 125508 397552 125520
rect 392728 125480 397552 125508
rect 392728 125468 392734 125480
rect 397546 125468 397552 125480
rect 397604 125468 397610 125520
rect 231486 125128 231492 125180
rect 231544 125168 231550 125180
rect 234062 125168 234068 125180
rect 231544 125140 234068 125168
rect 231544 125128 231550 125140
rect 234062 125128 234068 125140
rect 234120 125128 234126 125180
rect 207750 124244 207756 124296
rect 207808 124284 207814 124296
rect 214006 124284 214012 124296
rect 207808 124256 214012 124284
rect 207808 124244 207814 124256
rect 214006 124244 214012 124256
rect 214064 124244 214070 124296
rect 238018 124244 238024 124296
rect 238076 124284 238082 124296
rect 264974 124284 264980 124296
rect 238076 124256 264980 124284
rect 238076 124244 238082 124256
rect 264974 124244 264980 124256
rect 265032 124244 265038 124296
rect 171962 124176 171968 124228
rect 172020 124216 172026 124228
rect 213914 124216 213920 124228
rect 172020 124188 213920 124216
rect 172020 124176 172026 124188
rect 213914 124176 213920 124188
rect 213972 124176 213978 124228
rect 236638 124176 236644 124228
rect 236696 124216 236702 124228
rect 265066 124216 265072 124228
rect 236696 124188 265072 124216
rect 236696 124176 236702 124188
rect 265066 124176 265072 124188
rect 265124 124176 265130 124228
rect 282638 124108 282644 124160
rect 282696 124148 282702 124160
rect 307754 124148 307760 124160
rect 282696 124120 307760 124148
rect 282696 124108 282702 124120
rect 307754 124108 307760 124120
rect 307812 124108 307818 124160
rect 309962 124108 309968 124160
rect 310020 124148 310026 124160
rect 397546 124148 397552 124160
rect 310020 124120 397552 124148
rect 310020 124108 310026 124120
rect 397546 124108 397552 124120
rect 397604 124108 397610 124160
rect 442902 124108 442908 124160
rect 442960 124148 442966 124160
rect 582926 124148 582932 124160
rect 442960 124120 582932 124148
rect 442960 124108 442966 124120
rect 582926 124108 582932 124120
rect 582984 124108 582990 124160
rect 442810 124040 442816 124092
rect 442868 124080 442874 124092
rect 447226 124080 447232 124092
rect 442868 124052 447232 124080
rect 442868 124040 442874 124052
rect 447226 124040 447232 124052
rect 447284 124040 447290 124092
rect 231118 123904 231124 123956
rect 231176 123944 231182 123956
rect 235534 123944 235540 123956
rect 231176 123916 235540 123944
rect 231176 123904 231182 123916
rect 235534 123904 235540 123916
rect 235592 123904 235598 123956
rect 230658 123428 230664 123480
rect 230716 123468 230722 123480
rect 248046 123468 248052 123480
rect 230716 123440 248052 123468
rect 230716 123428 230722 123440
rect 248046 123428 248052 123440
rect 248104 123428 248110 123480
rect 171870 122816 171876 122868
rect 171928 122856 171934 122868
rect 213914 122856 213920 122868
rect 171928 122828 213920 122856
rect 171928 122816 171934 122828
rect 213914 122816 213920 122828
rect 213972 122816 213978 122868
rect 235442 122816 235448 122868
rect 235500 122856 235506 122868
rect 264974 122856 264980 122868
rect 235500 122828 264980 122856
rect 235500 122816 235506 122828
rect 264974 122816 264980 122828
rect 265032 122816 265038 122868
rect 231762 122748 231768 122800
rect 231820 122788 231826 122800
rect 257430 122788 257436 122800
rect 231820 122760 257436 122788
rect 231820 122748 231826 122760
rect 257430 122748 257436 122760
rect 257488 122748 257494 122800
rect 309870 122748 309876 122800
rect 309928 122788 309934 122800
rect 374730 122788 374736 122800
rect 309928 122760 374736 122788
rect 309928 122748 309934 122760
rect 374730 122748 374736 122760
rect 374788 122748 374794 122800
rect 442258 122748 442264 122800
rect 442316 122788 442322 122800
rect 442902 122788 442908 122800
rect 442316 122760 442908 122788
rect 442316 122748 442322 122760
rect 442902 122748 442908 122760
rect 442960 122788 442966 122800
rect 582466 122788 582472 122800
rect 442960 122760 582472 122788
rect 442960 122748 442966 122760
rect 582466 122748 582472 122760
rect 582524 122748 582530 122800
rect 231026 122680 231032 122732
rect 231084 122720 231090 122732
rect 245010 122720 245016 122732
rect 231084 122692 245016 122720
rect 231084 122680 231090 122692
rect 245010 122680 245016 122692
rect 245068 122680 245074 122732
rect 252094 122068 252100 122120
rect 252152 122108 252158 122120
rect 265066 122108 265072 122120
rect 252152 122080 265072 122108
rect 252152 122068 252158 122080
rect 265066 122068 265072 122080
rect 265124 122068 265130 122120
rect 282822 121592 282828 121644
rect 282880 121632 282886 121644
rect 288710 121632 288716 121644
rect 282880 121604 288716 121632
rect 282880 121592 282886 121604
rect 288710 121592 288716 121604
rect 288768 121592 288774 121644
rect 196802 121524 196808 121576
rect 196860 121564 196866 121576
rect 213914 121564 213920 121576
rect 196860 121536 213920 121564
rect 196860 121524 196866 121536
rect 213914 121524 213920 121536
rect 213972 121524 213978 121576
rect 63402 121456 63408 121508
rect 63460 121496 63466 121508
rect 65978 121496 65984 121508
rect 63460 121468 65984 121496
rect 63460 121456 63466 121468
rect 65978 121456 65984 121468
rect 66036 121456 66042 121508
rect 175918 121456 175924 121508
rect 175976 121496 175982 121508
rect 214006 121496 214012 121508
rect 175976 121468 214012 121496
rect 175976 121456 175982 121468
rect 214006 121456 214012 121468
rect 214064 121456 214070 121508
rect 309134 121456 309140 121508
rect 309192 121496 309198 121508
rect 309870 121496 309876 121508
rect 309192 121468 309876 121496
rect 309192 121456 309198 121468
rect 309870 121456 309876 121468
rect 309928 121456 309934 121508
rect 374638 121456 374644 121508
rect 374696 121496 374702 121508
rect 397546 121496 397552 121508
rect 374696 121468 397552 121496
rect 374696 121456 374702 121468
rect 397546 121456 397552 121468
rect 397604 121456 397610 121508
rect 231762 121388 231768 121440
rect 231820 121428 231826 121440
rect 247770 121428 247776 121440
rect 231820 121400 247776 121428
rect 231820 121388 231826 121400
rect 247770 121388 247776 121400
rect 247828 121388 247834 121440
rect 342990 121388 342996 121440
rect 343048 121428 343054 121440
rect 398742 121428 398748 121440
rect 343048 121400 398748 121428
rect 343048 121388 343054 121400
rect 398742 121388 398748 121400
rect 398800 121388 398806 121440
rect 441614 121388 441620 121440
rect 441672 121428 441678 121440
rect 442626 121428 442632 121440
rect 441672 121400 442632 121428
rect 441672 121388 441678 121400
rect 442626 121388 442632 121400
rect 442684 121428 442690 121440
rect 582374 121428 582380 121440
rect 442684 121400 582380 121428
rect 442684 121388 442690 121400
rect 582374 121388 582380 121400
rect 582432 121388 582438 121440
rect 249242 120708 249248 120760
rect 249300 120748 249306 120760
rect 264974 120748 264980 120760
rect 249300 120720 264980 120748
rect 249300 120708 249306 120720
rect 264974 120708 264980 120720
rect 265032 120708 265038 120760
rect 231486 120640 231492 120692
rect 231544 120680 231550 120692
rect 236914 120680 236920 120692
rect 231544 120652 236920 120680
rect 231544 120640 231550 120652
rect 236914 120640 236920 120652
rect 236972 120640 236978 120692
rect 193950 120164 193956 120216
rect 194008 120204 194014 120216
rect 213914 120204 213920 120216
rect 194008 120176 213920 120204
rect 194008 120164 194014 120176
rect 213914 120164 213920 120176
rect 213972 120164 213978 120216
rect 170490 120096 170496 120148
rect 170548 120136 170554 120148
rect 214006 120136 214012 120148
rect 170548 120108 214012 120136
rect 170548 120096 170554 120108
rect 214006 120096 214012 120108
rect 214064 120096 214070 120148
rect 258994 120096 259000 120148
rect 259052 120136 259058 120148
rect 265066 120136 265072 120148
rect 259052 120108 265072 120136
rect 259052 120096 259058 120108
rect 265066 120096 265072 120108
rect 265124 120096 265130 120148
rect 231762 120028 231768 120080
rect 231820 120068 231826 120080
rect 243722 120068 243728 120080
rect 231820 120040 243728 120068
rect 231820 120028 231826 120040
rect 243722 120028 243728 120040
rect 243780 120028 243786 120080
rect 282822 120028 282828 120080
rect 282880 120068 282886 120080
rect 288526 120068 288532 120080
rect 282880 120040 288532 120068
rect 282880 120028 282886 120040
rect 288526 120028 288532 120040
rect 288584 120028 288590 120080
rect 378778 120028 378784 120080
rect 378836 120068 378842 120080
rect 397546 120068 397552 120080
rect 378836 120040 397552 120068
rect 378836 120028 378842 120040
rect 397546 120028 397552 120040
rect 397604 120028 397610 120080
rect 442902 119688 442908 119740
rect 442960 119728 442966 119740
rect 447410 119728 447416 119740
rect 442960 119700 447416 119728
rect 442960 119688 442966 119700
rect 447410 119688 447416 119700
rect 447468 119688 447474 119740
rect 247954 119348 247960 119400
rect 248012 119388 248018 119400
rect 262858 119388 262864 119400
rect 248012 119360 262864 119388
rect 248012 119348 248018 119360
rect 262858 119348 262864 119360
rect 262916 119348 262922 119400
rect 282178 119348 282184 119400
rect 282236 119388 282242 119400
rect 299566 119388 299572 119400
rect 282236 119360 299572 119388
rect 282236 119348 282242 119360
rect 299566 119348 299572 119360
rect 299624 119348 299630 119400
rect 338206 119348 338212 119400
rect 338264 119388 338270 119400
rect 395430 119388 395436 119400
rect 338264 119360 395436 119388
rect 338264 119348 338270 119360
rect 395430 119348 395436 119360
rect 395488 119348 395494 119400
rect 203702 118736 203708 118788
rect 203760 118776 203766 118788
rect 213914 118776 213920 118788
rect 203760 118748 213920 118776
rect 203760 118736 203766 118748
rect 213914 118736 213920 118748
rect 213972 118736 213978 118788
rect 195330 118668 195336 118720
rect 195388 118708 195394 118720
rect 214006 118708 214012 118720
rect 195388 118680 214012 118708
rect 195388 118668 195394 118680
rect 214006 118668 214012 118680
rect 214064 118668 214070 118720
rect 259270 118668 259276 118720
rect 259328 118708 259334 118720
rect 264974 118708 264980 118720
rect 259328 118680 264980 118708
rect 259328 118668 259334 118680
rect 264974 118668 264980 118680
rect 265032 118668 265038 118720
rect 230566 118600 230572 118652
rect 230624 118640 230630 118652
rect 233970 118640 233976 118652
rect 230624 118612 233976 118640
rect 230624 118600 230630 118612
rect 233970 118600 233976 118612
rect 234028 118600 234034 118652
rect 282822 118600 282828 118652
rect 282880 118640 282886 118652
rect 298186 118640 298192 118652
rect 282880 118612 298192 118640
rect 282880 118600 282886 118612
rect 298186 118600 298192 118612
rect 298244 118600 298250 118652
rect 352558 118600 352564 118652
rect 352616 118640 352622 118652
rect 397638 118640 397644 118652
rect 352616 118612 397644 118640
rect 352616 118600 352622 118612
rect 397638 118600 397644 118612
rect 397696 118600 397702 118652
rect 360838 118532 360844 118584
rect 360896 118572 360902 118584
rect 397546 118572 397552 118584
rect 360896 118544 397552 118572
rect 360896 118532 360902 118544
rect 397546 118532 397552 118544
rect 397604 118532 397610 118584
rect 282822 118056 282828 118108
rect 282880 118096 282886 118108
rect 287238 118096 287244 118108
rect 282880 118068 287244 118096
rect 282880 118056 282886 118068
rect 287238 118056 287244 118068
rect 287296 118056 287302 118108
rect 231670 117988 231676 118040
rect 231728 118028 231734 118040
rect 246482 118028 246488 118040
rect 231728 118000 246488 118028
rect 231728 117988 231734 118000
rect 246482 117988 246488 118000
rect 246540 117988 246546 118040
rect 238294 117920 238300 117972
rect 238352 117960 238358 117972
rect 265802 117960 265808 117972
rect 238352 117932 265808 117960
rect 238352 117920 238358 117932
rect 265802 117920 265808 117932
rect 265860 117920 265866 117972
rect 198274 117376 198280 117428
rect 198332 117416 198338 117428
rect 214006 117416 214012 117428
rect 198332 117388 214012 117416
rect 198332 117376 198338 117388
rect 214006 117376 214012 117388
rect 214064 117376 214070 117428
rect 169294 117308 169300 117360
rect 169352 117348 169358 117360
rect 213914 117348 213920 117360
rect 169352 117320 213920 117348
rect 169352 117308 169358 117320
rect 213914 117308 213920 117320
rect 213972 117308 213978 117360
rect 250438 117308 250444 117360
rect 250496 117348 250502 117360
rect 264974 117348 264980 117360
rect 250496 117320 264980 117348
rect 250496 117308 250502 117320
rect 264974 117308 264980 117320
rect 265032 117308 265038 117360
rect 282822 117240 282828 117292
rect 282880 117280 282886 117292
rect 289998 117280 290004 117292
rect 282880 117252 290004 117280
rect 282880 117240 282886 117252
rect 289998 117240 290004 117252
rect 290056 117280 290062 117292
rect 291102 117280 291108 117292
rect 290056 117252 291108 117280
rect 290056 117240 290062 117252
rect 291102 117240 291108 117252
rect 291160 117240 291166 117292
rect 391198 117240 391204 117292
rect 391256 117280 391262 117292
rect 397546 117280 397552 117292
rect 391256 117252 397552 117280
rect 391256 117240 391262 117252
rect 397546 117240 397552 117252
rect 397604 117240 397610 117292
rect 231762 117172 231768 117224
rect 231820 117212 231826 117224
rect 244918 117212 244924 117224
rect 231820 117184 244924 117212
rect 231820 117172 231826 117184
rect 244918 117172 244924 117184
rect 244976 117172 244982 117224
rect 230842 117104 230848 117156
rect 230900 117144 230906 117156
rect 232682 117144 232688 117156
rect 230900 117116 232688 117144
rect 230900 117104 230906 117116
rect 232682 117104 232688 117116
rect 232740 117104 232746 117156
rect 282270 116696 282276 116748
rect 282328 116736 282334 116748
rect 285766 116736 285772 116748
rect 282328 116708 285772 116736
rect 282328 116696 282334 116708
rect 285766 116696 285772 116708
rect 285824 116696 285830 116748
rect 167822 116560 167828 116612
rect 167880 116600 167886 116612
rect 198090 116600 198096 116612
rect 167880 116572 198096 116600
rect 167880 116560 167886 116572
rect 198090 116560 198096 116572
rect 198148 116560 198154 116612
rect 200942 116016 200948 116068
rect 201000 116056 201006 116068
rect 214006 116056 214012 116068
rect 201000 116028 214012 116056
rect 201000 116016 201006 116028
rect 214006 116016 214012 116028
rect 214064 116016 214070 116068
rect 257430 116016 257436 116068
rect 257488 116056 257494 116068
rect 264974 116056 264980 116068
rect 257488 116028 264980 116056
rect 257488 116016 257494 116028
rect 264974 116016 264980 116028
rect 265032 116016 265038 116068
rect 189902 115948 189908 116000
rect 189960 115988 189966 116000
rect 213914 115988 213920 116000
rect 189960 115960 213920 115988
rect 189960 115948 189966 115960
rect 213914 115948 213920 115960
rect 213972 115948 213978 116000
rect 240778 115948 240784 116000
rect 240836 115988 240842 116000
rect 265066 115988 265072 116000
rect 240836 115960 265072 115988
rect 240836 115948 240842 115960
rect 265066 115948 265072 115960
rect 265124 115948 265130 116000
rect 231486 115880 231492 115932
rect 231544 115920 231550 115932
rect 253290 115920 253296 115932
rect 231544 115892 253296 115920
rect 231544 115880 231550 115892
rect 253290 115880 253296 115892
rect 253348 115880 253354 115932
rect 281718 115880 281724 115932
rect 281776 115920 281782 115932
rect 302326 115920 302332 115932
rect 281776 115892 302332 115920
rect 281776 115880 281782 115892
rect 302326 115880 302332 115892
rect 302384 115880 302390 115932
rect 356790 115880 356796 115932
rect 356848 115920 356854 115932
rect 397546 115920 397552 115932
rect 356848 115892 397552 115920
rect 356848 115880 356854 115892
rect 397546 115880 397552 115892
rect 397604 115880 397610 115932
rect 282454 115812 282460 115864
rect 282512 115852 282518 115864
rect 295334 115852 295340 115864
rect 282512 115824 295340 115852
rect 282512 115812 282518 115824
rect 295334 115812 295340 115824
rect 295392 115812 295398 115864
rect 184290 115200 184296 115252
rect 184348 115240 184354 115252
rect 200850 115240 200856 115252
rect 184348 115212 200856 115240
rect 184348 115200 184354 115212
rect 200850 115200 200856 115212
rect 200908 115200 200914 115252
rect 230658 115200 230664 115252
rect 230716 115240 230722 115252
rect 251910 115240 251916 115252
rect 230716 115212 251916 115240
rect 230716 115200 230722 115212
rect 251910 115200 251916 115212
rect 251968 115200 251974 115252
rect 363690 115200 363696 115252
rect 363748 115240 363754 115252
rect 397362 115240 397368 115252
rect 363748 115212 397368 115240
rect 363748 115200 363754 115212
rect 397362 115200 397368 115212
rect 397420 115200 397426 115252
rect 203610 114588 203616 114640
rect 203668 114628 203674 114640
rect 214006 114628 214012 114640
rect 203668 114600 214012 114628
rect 203668 114588 203674 114600
rect 214006 114588 214012 114600
rect 214064 114588 214070 114640
rect 258902 114588 258908 114640
rect 258960 114628 258966 114640
rect 265066 114628 265072 114640
rect 258960 114600 265072 114628
rect 258960 114588 258966 114600
rect 265066 114588 265072 114600
rect 265124 114588 265130 114640
rect 198090 114520 198096 114572
rect 198148 114560 198154 114572
rect 213914 114560 213920 114572
rect 198148 114532 213920 114560
rect 198148 114520 198154 114532
rect 213914 114520 213920 114532
rect 213972 114520 213978 114572
rect 256234 114520 256240 114572
rect 256292 114560 256298 114572
rect 264974 114560 264980 114572
rect 256292 114532 264980 114560
rect 256292 114520 256298 114532
rect 264974 114520 264980 114532
rect 265032 114520 265038 114572
rect 442902 114520 442908 114572
rect 442960 114560 442966 114572
rect 445938 114560 445944 114572
rect 442960 114532 445944 114560
rect 442960 114520 442966 114532
rect 445938 114520 445944 114532
rect 445996 114560 446002 114572
rect 452654 114560 452660 114572
rect 445996 114532 452660 114560
rect 445996 114520 446002 114532
rect 452654 114520 452660 114532
rect 452712 114520 452718 114572
rect 231670 114452 231676 114504
rect 231728 114492 231734 114504
rect 241054 114492 241060 114504
rect 231728 114464 241060 114492
rect 231728 114452 231734 114464
rect 241054 114452 241060 114464
rect 241112 114452 241118 114504
rect 323578 114452 323584 114504
rect 323636 114492 323642 114504
rect 397546 114492 397552 114504
rect 323636 114464 397552 114492
rect 323636 114452 323642 114464
rect 397546 114452 397552 114464
rect 397604 114452 397610 114504
rect 231486 114180 231492 114232
rect 231544 114220 231550 114232
rect 233878 114220 233884 114232
rect 231544 114192 233884 114220
rect 231544 114180 231550 114192
rect 233878 114180 233884 114192
rect 233936 114180 233942 114232
rect 282270 114112 282276 114164
rect 282328 114152 282334 114164
rect 285674 114152 285680 114164
rect 282328 114124 285680 114152
rect 282328 114112 282334 114124
rect 285674 114112 285680 114124
rect 285732 114112 285738 114164
rect 442350 113908 442356 113960
rect 442408 113948 442414 113960
rect 449894 113948 449900 113960
rect 442408 113920 449900 113948
rect 442408 113908 442414 113920
rect 449894 113908 449900 113920
rect 449952 113908 449958 113960
rect 241146 113772 241152 113824
rect 241204 113812 241210 113824
rect 254854 113812 254860 113824
rect 241204 113784 254860 113812
rect 241204 113772 241210 113784
rect 254854 113772 254860 113784
rect 254912 113772 254918 113824
rect 385770 113772 385776 113824
rect 385828 113812 385834 113824
rect 397914 113812 397920 113824
rect 385828 113784 397920 113812
rect 385828 113772 385834 113784
rect 397914 113772 397920 113784
rect 397972 113772 397978 113824
rect 188522 113228 188528 113280
rect 188580 113268 188586 113280
rect 213914 113268 213920 113280
rect 188580 113240 213920 113268
rect 188580 113228 188586 113240
rect 213914 113228 213920 113240
rect 213972 113228 213978 113280
rect 181622 113160 181628 113212
rect 181680 113200 181686 113212
rect 214006 113200 214012 113212
rect 181680 113172 214012 113200
rect 181680 113160 181686 113172
rect 214006 113160 214012 113172
rect 214064 113160 214070 113212
rect 253474 113160 253480 113212
rect 253532 113200 253538 113212
rect 264974 113200 264980 113212
rect 253532 113172 264980 113200
rect 253532 113160 253538 113172
rect 264974 113160 264980 113172
rect 265032 113160 265038 113212
rect 231762 113092 231768 113144
rect 231820 113132 231826 113144
rect 260282 113132 260288 113144
rect 231820 113104 260288 113132
rect 231820 113092 231826 113104
rect 260282 113092 260288 113104
rect 260340 113092 260346 113144
rect 282822 113092 282828 113144
rect 282880 113132 282886 113144
rect 321554 113132 321560 113144
rect 282880 113104 321560 113132
rect 282880 113092 282886 113104
rect 321554 113092 321560 113104
rect 321612 113132 321618 113144
rect 367094 113132 367100 113144
rect 321612 113104 367100 113132
rect 321612 113092 321618 113104
rect 367094 113092 367100 113104
rect 367152 113092 367158 113144
rect 231026 113024 231032 113076
rect 231084 113064 231090 113076
rect 249334 113064 249340 113076
rect 231084 113036 249340 113064
rect 231084 113024 231090 113036
rect 249334 113024 249340 113036
rect 249392 113024 249398 113076
rect 282822 112616 282828 112668
rect 282880 112656 282886 112668
rect 287146 112656 287152 112668
rect 282880 112628 287152 112656
rect 282880 112616 282886 112628
rect 287146 112616 287152 112628
rect 287204 112616 287210 112668
rect 178770 111868 178776 111920
rect 178828 111908 178834 111920
rect 214006 111908 214012 111920
rect 178828 111880 214012 111908
rect 178828 111868 178834 111880
rect 214006 111868 214012 111880
rect 214064 111868 214070 111920
rect 263134 111868 263140 111920
rect 263192 111908 263198 111920
rect 265250 111908 265256 111920
rect 263192 111880 265256 111908
rect 263192 111868 263198 111880
rect 265250 111868 265256 111880
rect 265308 111868 265314 111920
rect 377490 111868 377496 111920
rect 377548 111908 377554 111920
rect 397638 111908 397644 111920
rect 377548 111880 397644 111908
rect 377548 111868 377554 111880
rect 397638 111868 397644 111880
rect 397696 111868 397702 111920
rect 173342 111800 173348 111852
rect 173400 111840 173406 111852
rect 213914 111840 213920 111852
rect 173400 111812 213920 111840
rect 173400 111800 173406 111812
rect 213914 111800 213920 111812
rect 213972 111800 213978 111852
rect 251910 111800 251916 111852
rect 251968 111840 251974 111852
rect 264974 111840 264980 111852
rect 251968 111812 264980 111840
rect 251968 111800 251974 111812
rect 264974 111800 264980 111812
rect 265032 111800 265038 111852
rect 359550 111800 359556 111852
rect 359608 111840 359614 111852
rect 397730 111840 397736 111852
rect 359608 111812 397736 111840
rect 359608 111800 359614 111812
rect 397730 111800 397736 111812
rect 397788 111800 397794 111852
rect 3142 111732 3148 111784
rect 3200 111772 3206 111784
rect 35158 111772 35164 111784
rect 3200 111744 35164 111772
rect 3200 111732 3206 111744
rect 35158 111732 35164 111744
rect 35216 111732 35222 111784
rect 230566 111732 230572 111784
rect 230624 111772 230630 111784
rect 232590 111772 232596 111784
rect 230624 111744 232596 111772
rect 230624 111732 230630 111744
rect 232590 111732 232596 111744
rect 232648 111732 232654 111784
rect 282270 111732 282276 111784
rect 282328 111772 282334 111784
rect 293954 111772 293960 111784
rect 282328 111744 293960 111772
rect 282328 111732 282334 111744
rect 293954 111732 293960 111744
rect 294012 111732 294018 111784
rect 336090 111732 336096 111784
rect 336148 111772 336154 111784
rect 397454 111772 397460 111784
rect 336148 111744 397460 111772
rect 336148 111732 336154 111744
rect 397454 111732 397460 111744
rect 397512 111732 397518 111784
rect 231762 111664 231768 111716
rect 231820 111704 231826 111716
rect 242526 111704 242532 111716
rect 231820 111676 242532 111704
rect 231820 111664 231826 111676
rect 242526 111664 242532 111676
rect 242584 111664 242590 111716
rect 442350 111528 442356 111580
rect 442408 111568 442414 111580
rect 445846 111568 445852 111580
rect 442408 111540 445852 111568
rect 442408 111528 442414 111540
rect 445846 111528 445852 111540
rect 445904 111528 445910 111580
rect 359458 111052 359464 111104
rect 359516 111092 359522 111104
rect 397638 111092 397644 111104
rect 359516 111064 397644 111092
rect 359516 111052 359522 111064
rect 397638 111052 397644 111064
rect 397696 111052 397702 111104
rect 442166 111052 442172 111104
rect 442224 111092 442230 111104
rect 447134 111092 447140 111104
rect 442224 111064 447140 111092
rect 442224 111052 442230 111064
rect 447134 111052 447140 111064
rect 447192 111052 447198 111104
rect 193858 110508 193864 110560
rect 193916 110548 193922 110560
rect 214006 110548 214012 110560
rect 193916 110520 214012 110548
rect 193916 110508 193922 110520
rect 214006 110508 214012 110520
rect 214064 110508 214070 110560
rect 249058 110508 249064 110560
rect 249116 110548 249122 110560
rect 265066 110548 265072 110560
rect 249116 110520 265072 110548
rect 249116 110508 249122 110520
rect 265066 110508 265072 110520
rect 265124 110508 265130 110560
rect 166534 110440 166540 110492
rect 166592 110480 166598 110492
rect 213914 110480 213920 110492
rect 166592 110452 213920 110480
rect 166592 110440 166598 110452
rect 213914 110440 213920 110452
rect 213972 110440 213978 110492
rect 243722 110440 243728 110492
rect 243780 110480 243786 110492
rect 264974 110480 264980 110492
rect 243780 110452 264980 110480
rect 243780 110440 243786 110452
rect 264974 110440 264980 110452
rect 265032 110440 265038 110492
rect 167822 110372 167828 110424
rect 167880 110412 167886 110424
rect 181530 110412 181536 110424
rect 167880 110384 181536 110412
rect 167880 110372 167886 110384
rect 181530 110372 181536 110384
rect 181588 110372 181594 110424
rect 231762 110372 231768 110424
rect 231820 110412 231826 110424
rect 252002 110412 252008 110424
rect 231820 110384 252008 110412
rect 231820 110372 231826 110384
rect 252002 110372 252008 110384
rect 252060 110372 252066 110424
rect 282822 110372 282828 110424
rect 282880 110412 282886 110424
rect 298094 110412 298100 110424
rect 282880 110384 298100 110412
rect 282880 110372 282886 110384
rect 298094 110372 298100 110384
rect 298152 110372 298158 110424
rect 231670 109692 231676 109744
rect 231728 109732 231734 109744
rect 246390 109732 246396 109744
rect 231728 109704 246396 109732
rect 231728 109692 231734 109704
rect 246390 109692 246396 109704
rect 246448 109692 246454 109744
rect 360838 109692 360844 109744
rect 360896 109732 360902 109744
rect 397546 109732 397552 109744
rect 360896 109704 397552 109732
rect 360896 109692 360902 109704
rect 397546 109692 397552 109704
rect 397604 109692 397610 109744
rect 192478 109080 192484 109132
rect 192536 109120 192542 109132
rect 214006 109120 214012 109132
rect 192536 109092 214012 109120
rect 192536 109080 192542 109092
rect 214006 109080 214012 109092
rect 214064 109080 214070 109132
rect 256050 109080 256056 109132
rect 256108 109120 256114 109132
rect 264974 109120 264980 109132
rect 256108 109092 264980 109120
rect 256108 109080 256114 109092
rect 264974 109080 264980 109092
rect 265032 109080 265038 109132
rect 180334 109012 180340 109064
rect 180392 109052 180398 109064
rect 213914 109052 213920 109064
rect 180392 109024 213920 109052
rect 180392 109012 180398 109024
rect 213914 109012 213920 109024
rect 213972 109012 213978 109064
rect 250530 109012 250536 109064
rect 250588 109052 250594 109064
rect 265066 109052 265072 109064
rect 250588 109024 265072 109052
rect 250588 109012 250594 109024
rect 265066 109012 265072 109024
rect 265124 109012 265130 109064
rect 385770 109012 385776 109064
rect 385828 109052 385834 109064
rect 397454 109052 397460 109064
rect 385828 109024 397460 109052
rect 385828 109012 385834 109024
rect 397454 109012 397460 109024
rect 397512 109012 397518 109064
rect 231486 108944 231492 108996
rect 231544 108984 231550 108996
rect 253382 108984 253388 108996
rect 231544 108956 253388 108984
rect 231544 108944 231550 108956
rect 253382 108944 253388 108956
rect 253440 108944 253446 108996
rect 282362 108944 282368 108996
rect 282420 108984 282426 108996
rect 305086 108984 305092 108996
rect 282420 108956 305092 108984
rect 282420 108944 282426 108956
rect 305086 108944 305092 108956
rect 305144 108944 305150 108996
rect 231762 108876 231768 108928
rect 231820 108916 231826 108928
rect 242434 108916 242440 108928
rect 231820 108888 242440 108916
rect 231820 108876 231826 108888
rect 242434 108876 242440 108888
rect 242492 108876 242498 108928
rect 257614 108264 257620 108316
rect 257672 108304 257678 108316
rect 264330 108304 264336 108316
rect 257672 108276 264336 108304
rect 257672 108264 257678 108276
rect 264330 108264 264336 108276
rect 264388 108264 264394 108316
rect 302878 108264 302884 108316
rect 302936 108304 302942 108316
rect 398190 108304 398196 108316
rect 302936 108276 398196 108304
rect 302936 108264 302942 108276
rect 398190 108264 398196 108276
rect 398248 108264 398254 108316
rect 207658 107720 207664 107772
rect 207716 107760 207722 107772
rect 214006 107760 214012 107772
rect 207716 107732 214012 107760
rect 207716 107720 207722 107732
rect 214006 107720 214012 107732
rect 214064 107720 214070 107772
rect 173250 107652 173256 107704
rect 173308 107692 173314 107704
rect 213914 107692 213920 107704
rect 173308 107664 213920 107692
rect 173308 107652 173314 107664
rect 213914 107652 213920 107664
rect 213972 107652 213978 107704
rect 367830 107652 367836 107704
rect 367888 107692 367894 107704
rect 397454 107692 397460 107704
rect 367888 107664 397460 107692
rect 367888 107652 367894 107664
rect 397454 107652 397460 107664
rect 397512 107652 397518 107704
rect 442902 107652 442908 107704
rect 442960 107692 442966 107704
rect 452654 107692 452660 107704
rect 442960 107664 452660 107692
rect 442960 107652 442966 107664
rect 452654 107652 452660 107664
rect 452712 107652 452718 107704
rect 231578 107584 231584 107636
rect 231636 107624 231642 107636
rect 264606 107624 264612 107636
rect 231636 107596 264612 107624
rect 231636 107584 231642 107596
rect 264606 107584 264612 107596
rect 264664 107584 264670 107636
rect 304258 107584 304264 107636
rect 304316 107624 304322 107636
rect 397546 107624 397552 107636
rect 304316 107596 397552 107624
rect 304316 107584 304322 107596
rect 397546 107584 397552 107596
rect 397604 107584 397610 107636
rect 442534 107584 442540 107636
rect 442592 107624 442598 107636
rect 456794 107624 456800 107636
rect 442592 107596 456800 107624
rect 442592 107584 442598 107596
rect 456794 107584 456800 107596
rect 456852 107584 456858 107636
rect 230934 107516 230940 107568
rect 230992 107556 230998 107568
rect 238110 107556 238116 107568
rect 230992 107528 238116 107556
rect 230992 107516 230998 107528
rect 238110 107516 238116 107528
rect 238168 107516 238174 107568
rect 381630 107516 381636 107568
rect 381688 107556 381694 107568
rect 397454 107556 397460 107568
rect 381688 107528 397460 107556
rect 381688 107516 381694 107528
rect 397454 107516 397460 107528
rect 397512 107516 397518 107568
rect 178862 106904 178868 106956
rect 178920 106944 178926 106956
rect 205266 106944 205272 106956
rect 178920 106916 205272 106944
rect 178920 106904 178926 106916
rect 205266 106904 205272 106916
rect 205324 106904 205330 106956
rect 205082 106360 205088 106412
rect 205140 106400 205146 106412
rect 214006 106400 214012 106412
rect 205140 106372 214012 106400
rect 205140 106360 205146 106372
rect 214006 106360 214012 106372
rect 214064 106360 214070 106412
rect 167822 106292 167828 106344
rect 167880 106332 167886 106344
rect 213914 106332 213920 106344
rect 167880 106304 213920 106332
rect 167880 106292 167886 106304
rect 213914 106292 213920 106304
rect 213972 106292 213978 106344
rect 246482 106292 246488 106344
rect 246540 106332 246546 106344
rect 264974 106332 264980 106344
rect 246540 106304 264980 106332
rect 246540 106292 246546 106304
rect 264974 106292 264980 106304
rect 265032 106292 265038 106344
rect 231578 106224 231584 106276
rect 231636 106264 231642 106276
rect 249150 106264 249156 106276
rect 231636 106236 249156 106264
rect 231636 106224 231642 106236
rect 249150 106224 249156 106236
rect 249208 106224 249214 106276
rect 320910 106224 320916 106276
rect 320968 106264 320974 106276
rect 397454 106264 397460 106276
rect 320968 106236 397460 106264
rect 320968 106224 320974 106236
rect 397454 106224 397460 106236
rect 397512 106224 397518 106276
rect 167730 105544 167736 105596
rect 167788 105584 167794 105596
rect 195514 105584 195520 105596
rect 167788 105556 195520 105584
rect 167788 105544 167794 105556
rect 195514 105544 195520 105556
rect 195572 105544 195578 105596
rect 371970 105544 371976 105596
rect 372028 105584 372034 105596
rect 399754 105584 399760 105596
rect 372028 105556 399760 105584
rect 372028 105544 372034 105556
rect 399754 105544 399760 105556
rect 399812 105544 399818 105596
rect 260282 104932 260288 104984
rect 260340 104972 260346 104984
rect 265066 104972 265072 104984
rect 260340 104944 265072 104972
rect 260340 104932 260346 104944
rect 265066 104932 265072 104944
rect 265124 104932 265130 104984
rect 198182 104864 198188 104916
rect 198240 104904 198246 104916
rect 213914 104904 213920 104916
rect 198240 104876 213920 104904
rect 198240 104864 198246 104876
rect 213914 104864 213920 104876
rect 213972 104864 213978 104916
rect 245010 104864 245016 104916
rect 245068 104904 245074 104916
rect 264974 104904 264980 104916
rect 245068 104876 264980 104904
rect 245068 104864 245074 104876
rect 264974 104864 264980 104876
rect 265032 104864 265038 104916
rect 231762 104796 231768 104848
rect 231820 104836 231826 104848
rect 250622 104836 250628 104848
rect 231820 104808 250628 104836
rect 231820 104796 231826 104808
rect 250622 104796 250628 104808
rect 250680 104796 250686 104848
rect 281902 104796 281908 104848
rect 281960 104836 281966 104848
rect 284386 104836 284392 104848
rect 281960 104808 284392 104836
rect 281960 104796 281966 104808
rect 284386 104796 284392 104808
rect 284444 104796 284450 104848
rect 327718 104796 327724 104848
rect 327776 104836 327782 104848
rect 397454 104836 397460 104848
rect 327776 104808 397460 104836
rect 327776 104796 327782 104808
rect 397454 104796 397460 104808
rect 397512 104796 397518 104848
rect 231486 104728 231492 104780
rect 231544 104768 231550 104780
rect 243630 104768 243636 104780
rect 231544 104740 243636 104768
rect 231544 104728 231550 104740
rect 243630 104728 243636 104740
rect 243688 104728 243694 104780
rect 172054 104184 172060 104236
rect 172112 104224 172118 104236
rect 198274 104224 198280 104236
rect 172112 104196 198280 104224
rect 172112 104184 172118 104196
rect 198274 104184 198280 104196
rect 198332 104184 198338 104236
rect 166258 104116 166264 104168
rect 166316 104156 166322 104168
rect 214558 104156 214564 104168
rect 166316 104128 214564 104156
rect 166316 104116 166322 104128
rect 214558 104116 214564 104128
rect 214616 104116 214622 104168
rect 383010 104116 383016 104168
rect 383068 104156 383074 104168
rect 399846 104156 399852 104168
rect 383068 104128 399852 104156
rect 383068 104116 383074 104128
rect 399846 104116 399852 104128
rect 399904 104116 399910 104168
rect 441982 104116 441988 104168
rect 442040 104156 442046 104168
rect 451274 104156 451280 104168
rect 442040 104128 451280 104156
rect 442040 104116 442046 104128
rect 451274 104116 451280 104128
rect 451332 104116 451338 104168
rect 211890 103504 211896 103556
rect 211948 103544 211954 103556
rect 213914 103544 213920 103556
rect 211948 103516 213920 103544
rect 211948 103504 211954 103516
rect 213914 103504 213920 103516
rect 213972 103504 213978 103556
rect 254762 103504 254768 103556
rect 254820 103544 254826 103556
rect 264974 103544 264980 103556
rect 254820 103516 264980 103544
rect 254820 103504 254826 103516
rect 264974 103504 264980 103516
rect 265032 103504 265038 103556
rect 231762 103436 231768 103488
rect 231820 103476 231826 103488
rect 240962 103476 240968 103488
rect 231820 103448 240968 103476
rect 231820 103436 231826 103448
rect 240962 103436 240968 103448
rect 241020 103436 241026 103488
rect 282822 103436 282828 103488
rect 282880 103476 282886 103488
rect 314654 103476 314660 103488
rect 282880 103448 314660 103476
rect 282880 103436 282886 103448
rect 314654 103436 314660 103448
rect 314712 103436 314718 103488
rect 322290 103436 322296 103488
rect 322348 103476 322354 103488
rect 397454 103476 397460 103488
rect 322348 103448 397460 103476
rect 322348 103436 322354 103448
rect 397454 103436 397460 103448
rect 397512 103436 397518 103488
rect 231394 103368 231400 103420
rect 231452 103408 231458 103420
rect 239582 103408 239588 103420
rect 231452 103380 239588 103408
rect 231452 103368 231458 103380
rect 239582 103368 239588 103380
rect 239640 103368 239646 103420
rect 281718 103164 281724 103216
rect 281776 103204 281782 103216
rect 283558 103204 283564 103216
rect 281776 103176 283564 103204
rect 281776 103164 281782 103176
rect 283558 103164 283564 103176
rect 283616 103164 283622 103216
rect 442718 102756 442724 102808
rect 442776 102796 442782 102808
rect 444466 102796 444472 102808
rect 442776 102768 444472 102796
rect 442776 102756 442782 102768
rect 444466 102756 444472 102768
rect 444524 102756 444530 102808
rect 187050 102212 187056 102264
rect 187108 102252 187114 102264
rect 214006 102252 214012 102264
rect 187108 102224 214012 102252
rect 187108 102212 187114 102224
rect 214006 102212 214012 102224
rect 214064 102212 214070 102264
rect 169018 102144 169024 102196
rect 169076 102184 169082 102196
rect 213914 102184 213920 102196
rect 169076 102156 213920 102184
rect 169076 102144 169082 102156
rect 213914 102144 213920 102156
rect 213972 102144 213978 102196
rect 249150 102144 249156 102196
rect 249208 102184 249214 102196
rect 264974 102184 264980 102196
rect 249208 102156 264980 102184
rect 249208 102144 249214 102156
rect 264974 102144 264980 102156
rect 265032 102144 265038 102196
rect 231762 102076 231768 102128
rect 231820 102116 231826 102128
rect 247862 102116 247868 102128
rect 231820 102088 247868 102116
rect 231820 102076 231826 102088
rect 247862 102076 247868 102088
rect 247920 102076 247926 102128
rect 170674 101464 170680 101516
rect 170732 101504 170738 101516
rect 196710 101504 196716 101516
rect 170732 101476 196716 101504
rect 170732 101464 170738 101476
rect 196710 101464 196716 101476
rect 196768 101464 196774 101516
rect 230474 101464 230480 101516
rect 230532 101504 230538 101516
rect 238294 101504 238300 101516
rect 230532 101476 238300 101504
rect 230532 101464 230538 101476
rect 238294 101464 238300 101476
rect 238352 101464 238358 101516
rect 177482 101396 177488 101448
rect 177540 101436 177546 101448
rect 213454 101436 213460 101448
rect 177540 101408 213460 101436
rect 177540 101396 177546 101408
rect 213454 101396 213460 101408
rect 213512 101396 213518 101448
rect 439958 101396 439964 101448
rect 440016 101436 440022 101448
rect 463694 101436 463700 101448
rect 440016 101408 463700 101436
rect 440016 101396 440022 101408
rect 463694 101396 463700 101408
rect 463752 101396 463758 101448
rect 261754 100784 261760 100836
rect 261812 100824 261818 100836
rect 265066 100824 265072 100836
rect 261812 100796 265072 100824
rect 261812 100784 261818 100796
rect 265066 100784 265072 100796
rect 265124 100784 265130 100836
rect 176010 100716 176016 100768
rect 176068 100756 176074 100768
rect 177390 100756 177396 100768
rect 176068 100728 177396 100756
rect 176068 100716 176074 100728
rect 177390 100716 177396 100728
rect 177448 100716 177454 100768
rect 196894 100716 196900 100768
rect 196952 100756 196958 100768
rect 213914 100756 213920 100768
rect 196952 100728 213920 100756
rect 196952 100716 196958 100728
rect 213914 100716 213920 100728
rect 213972 100716 213978 100768
rect 241054 100716 241060 100768
rect 241112 100756 241118 100768
rect 264974 100756 264980 100768
rect 241112 100728 264980 100756
rect 241112 100716 241118 100728
rect 264974 100716 264980 100728
rect 265032 100716 265038 100768
rect 395430 100716 395436 100768
rect 395488 100756 395494 100768
rect 397546 100756 397552 100768
rect 395488 100728 397552 100756
rect 395488 100716 395494 100728
rect 397546 100716 397552 100728
rect 397604 100716 397610 100768
rect 398190 100716 398196 100768
rect 398248 100756 398254 100768
rect 439958 100756 439964 100768
rect 398248 100728 404676 100756
rect 398248 100716 398254 100728
rect 404648 100700 404676 100728
rect 439332 100728 439964 100756
rect 439332 100700 439360 100728
rect 439958 100716 439964 100728
rect 440016 100716 440022 100768
rect 399846 100648 399852 100700
rect 399904 100688 399910 100700
rect 403342 100688 403348 100700
rect 399904 100660 403348 100688
rect 399904 100648 399910 100660
rect 403342 100648 403348 100660
rect 403400 100648 403406 100700
rect 404630 100648 404636 100700
rect 404688 100648 404694 100700
rect 439314 100648 439320 100700
rect 439372 100648 439378 100700
rect 231762 100580 231768 100632
rect 231820 100620 231826 100632
rect 256142 100620 256148 100632
rect 231820 100592 256148 100620
rect 231820 100580 231826 100592
rect 256142 100580 256148 100592
rect 256200 100580 256206 100632
rect 399754 100580 399760 100632
rect 399812 100620 399818 100632
rect 402974 100620 402980 100632
rect 399812 100592 402980 100620
rect 399812 100580 399818 100592
rect 402974 100580 402980 100592
rect 403032 100580 403038 100632
rect 405274 99968 405280 100020
rect 405332 100008 405338 100020
rect 580166 100008 580172 100020
rect 405332 99980 580172 100008
rect 405332 99968 405338 99980
rect 580166 99968 580172 99980
rect 580224 99968 580230 100020
rect 230566 99696 230572 99748
rect 230624 99736 230630 99748
rect 232498 99736 232504 99748
rect 230624 99708 232504 99736
rect 230624 99696 230630 99708
rect 232498 99696 232504 99708
rect 232556 99696 232562 99748
rect 211982 99424 211988 99476
rect 212040 99464 212046 99476
rect 214466 99464 214472 99476
rect 212040 99436 214472 99464
rect 212040 99424 212046 99436
rect 214466 99424 214472 99436
rect 214524 99424 214530 99476
rect 257522 99424 257528 99476
rect 257580 99464 257586 99476
rect 265066 99464 265072 99476
rect 257580 99436 265072 99464
rect 257580 99424 257586 99436
rect 265066 99424 265072 99436
rect 265124 99424 265130 99476
rect 181714 99356 181720 99408
rect 181772 99396 181778 99408
rect 213914 99396 213920 99408
rect 181772 99368 213920 99396
rect 181772 99356 181778 99368
rect 213914 99356 213920 99368
rect 213972 99356 213978 99408
rect 233970 99356 233976 99408
rect 234028 99396 234034 99408
rect 264974 99396 264980 99408
rect 234028 99368 264980 99396
rect 234028 99356 234034 99368
rect 264974 99356 264980 99368
rect 265032 99356 265038 99408
rect 395338 99356 395344 99408
rect 395396 99396 395402 99408
rect 432782 99396 432788 99408
rect 395396 99368 432788 99396
rect 395396 99356 395402 99368
rect 432782 99356 432788 99368
rect 432840 99356 432846 99408
rect 435542 99356 435548 99408
rect 435600 99396 435606 99408
rect 440510 99396 440516 99408
rect 435600 99368 440516 99396
rect 435600 99356 435606 99368
rect 440510 99356 440516 99368
rect 440568 99356 440574 99408
rect 231026 99288 231032 99340
rect 231084 99328 231090 99340
rect 263042 99328 263048 99340
rect 231084 99300 263048 99328
rect 231084 99288 231090 99300
rect 263042 99288 263048 99300
rect 263100 99288 263106 99340
rect 281994 99288 282000 99340
rect 282052 99328 282058 99340
rect 296806 99328 296812 99340
rect 282052 99300 296812 99328
rect 282052 99288 282058 99300
rect 296806 99288 296812 99300
rect 296864 99288 296870 99340
rect 376018 99288 376024 99340
rect 376076 99328 376082 99340
rect 417694 99328 417700 99340
rect 376076 99300 417700 99328
rect 376076 99288 376082 99300
rect 417694 99288 417700 99300
rect 417752 99328 417758 99340
rect 582742 99328 582748 99340
rect 417752 99300 582748 99328
rect 417752 99288 417758 99300
rect 582742 99288 582748 99300
rect 582800 99288 582806 99340
rect 282822 99220 282828 99272
rect 282880 99260 282886 99272
rect 294046 99260 294052 99272
rect 282880 99232 294052 99260
rect 282880 99220 282886 99232
rect 294046 99220 294052 99232
rect 294104 99220 294110 99272
rect 384298 99220 384304 99272
rect 384356 99260 384362 99272
rect 411990 99260 411996 99272
rect 384356 99232 411996 99260
rect 384356 99220 384362 99232
rect 411990 99220 411996 99232
rect 412048 99220 412054 99272
rect 433518 99220 433524 99272
rect 433576 99260 433582 99272
rect 445754 99260 445760 99272
rect 433576 99232 445760 99260
rect 433576 99220 433582 99232
rect 445754 99220 445760 99232
rect 445812 99220 445818 99272
rect 230750 98812 230756 98864
rect 230808 98852 230814 98864
rect 234154 98852 234160 98864
rect 230808 98824 234160 98852
rect 230808 98812 230814 98824
rect 234154 98812 234160 98824
rect 234212 98812 234218 98864
rect 358078 98608 358084 98660
rect 358136 98648 358142 98660
rect 381630 98648 381636 98660
rect 358136 98620 381636 98648
rect 358136 98608 358142 98620
rect 381630 98608 381636 98620
rect 381688 98608 381694 98660
rect 173434 98064 173440 98116
rect 173492 98104 173498 98116
rect 214006 98104 214012 98116
rect 173492 98076 214012 98104
rect 173492 98064 173498 98076
rect 214006 98064 214012 98076
rect 214064 98064 214070 98116
rect 164878 97996 164884 98048
rect 164936 98036 164942 98048
rect 213914 98036 213920 98048
rect 164936 98008 213920 98036
rect 164936 97996 164942 98008
rect 213914 97996 213920 98008
rect 213972 97996 213978 98048
rect 261846 97996 261852 98048
rect 261904 98036 261910 98048
rect 264974 98036 264980 98048
rect 261904 98008 264980 98036
rect 261904 97996 261910 98008
rect 264974 97996 264980 98008
rect 265032 97996 265038 98048
rect 3510 97928 3516 97980
rect 3568 97968 3574 97980
rect 15838 97968 15844 97980
rect 3568 97940 15844 97968
rect 3568 97928 3574 97940
rect 15838 97928 15844 97940
rect 15896 97928 15902 97980
rect 215294 97928 215300 97980
rect 215352 97968 215358 97980
rect 215352 97940 224954 97968
rect 215352 97928 215358 97940
rect 182818 97248 182824 97300
rect 182876 97288 182882 97300
rect 213270 97288 213276 97300
rect 182876 97260 213276 97288
rect 182876 97248 182882 97260
rect 213270 97248 213276 97260
rect 213328 97248 213334 97300
rect 165522 96636 165528 96688
rect 165580 96676 165586 96688
rect 213914 96676 213920 96688
rect 165580 96648 213920 96676
rect 165580 96636 165586 96648
rect 213914 96636 213920 96648
rect 213972 96636 213978 96688
rect 224926 96064 224954 97940
rect 282822 97928 282828 97980
rect 282880 97968 282886 97980
rect 302234 97968 302240 97980
rect 282880 97940 302240 97968
rect 282880 97928 282886 97940
rect 302234 97928 302240 97940
rect 302292 97928 302298 97980
rect 434622 97928 434628 97980
rect 434680 97968 434686 97980
rect 465074 97968 465080 97980
rect 434680 97940 465080 97968
rect 434680 97928 434686 97940
rect 465074 97928 465080 97940
rect 465132 97968 465138 97980
rect 583110 97968 583116 97980
rect 465132 97940 583116 97968
rect 465132 97928 465138 97940
rect 583110 97928 583116 97940
rect 583168 97928 583174 97980
rect 282730 97860 282736 97912
rect 282788 97900 282794 97912
rect 291378 97900 291384 97912
rect 282788 97872 291384 97900
rect 282788 97860 282794 97872
rect 291378 97860 291384 97872
rect 291436 97860 291442 97912
rect 401410 97860 401416 97912
rect 401468 97900 401474 97912
rect 432230 97900 432236 97912
rect 401468 97872 432236 97900
rect 401468 97860 401474 97872
rect 432230 97860 432236 97872
rect 432288 97860 432294 97912
rect 435358 97860 435364 97912
rect 435416 97900 435422 97912
rect 448514 97900 448520 97912
rect 435416 97872 448520 97900
rect 435416 97860 435422 97872
rect 448514 97860 448520 97872
rect 448572 97860 448578 97912
rect 403618 97792 403624 97844
rect 403676 97832 403682 97844
rect 404446 97832 404452 97844
rect 403676 97804 404452 97832
rect 403676 97792 403682 97804
rect 404446 97792 404452 97804
rect 404504 97792 404510 97844
rect 264974 97288 264980 97300
rect 234586 97260 264980 97288
rect 234586 96676 234614 97260
rect 264974 97248 264980 97260
rect 265032 97248 265038 97300
rect 300118 97248 300124 97300
rect 300176 97288 300182 97300
rect 391934 97288 391940 97300
rect 300176 97260 391940 97288
rect 300176 97248 300182 97260
rect 391934 97248 391940 97260
rect 391992 97248 391998 97300
rect 394142 96908 394148 96960
rect 394200 96948 394206 96960
rect 401134 96948 401140 96960
rect 394200 96920 401140 96948
rect 394200 96908 394206 96920
rect 401134 96908 401140 96920
rect 401192 96908 401198 96960
rect 414014 96908 414020 96960
rect 414072 96948 414078 96960
rect 414750 96948 414756 96960
rect 414072 96920 414756 96948
rect 414072 96908 414078 96920
rect 414750 96908 414756 96920
rect 414808 96908 414814 96960
rect 430574 96908 430580 96960
rect 430632 96948 430638 96960
rect 431126 96948 431132 96960
rect 430632 96920 431132 96948
rect 430632 96908 430638 96920
rect 431126 96908 431132 96920
rect 431184 96908 431190 96960
rect 421558 96840 421564 96892
rect 421616 96880 421622 96892
rect 423398 96880 423404 96892
rect 421616 96852 423404 96880
rect 421616 96840 421622 96852
rect 423398 96840 423404 96852
rect 423456 96840 423462 96892
rect 418798 96704 418804 96756
rect 418856 96744 418862 96756
rect 420086 96744 420092 96756
rect 418856 96716 420092 96744
rect 418856 96704 418862 96716
rect 420086 96704 420092 96716
rect 420144 96704 420150 96756
rect 226444 96648 234614 96676
rect 226444 96076 226472 96648
rect 235350 96636 235356 96688
rect 235408 96676 235414 96688
rect 265066 96676 265072 96688
rect 235408 96648 265072 96676
rect 235408 96636 235414 96648
rect 265066 96636 265072 96648
rect 265124 96636 265130 96688
rect 282822 96568 282828 96620
rect 282880 96608 282886 96620
rect 301038 96608 301044 96620
rect 282880 96580 301044 96608
rect 282880 96568 282886 96580
rect 301038 96568 301044 96580
rect 301096 96568 301102 96620
rect 334618 96568 334624 96620
rect 334676 96608 334682 96620
rect 422662 96608 422668 96620
rect 334676 96580 422668 96608
rect 334676 96568 334682 96580
rect 422662 96568 422668 96580
rect 422720 96568 422726 96620
rect 389818 96500 389824 96552
rect 389876 96540 389882 96552
rect 418982 96540 418988 96552
rect 389876 96512 418988 96540
rect 389876 96500 389882 96512
rect 418982 96500 418988 96512
rect 419040 96500 419046 96552
rect 225046 96064 225052 96076
rect 224926 96036 225052 96064
rect 225046 96024 225052 96036
rect 225104 96024 225110 96076
rect 226426 96024 226432 96076
rect 226484 96024 226490 96076
rect 168282 95956 168288 96008
rect 168340 95996 168346 96008
rect 184382 95996 184388 96008
rect 168340 95968 184388 95996
rect 168340 95956 168346 95968
rect 184382 95956 184388 95968
rect 184440 95956 184446 96008
rect 198642 95956 198648 96008
rect 198700 95996 198706 96008
rect 222470 95996 222476 96008
rect 198700 95968 222476 95996
rect 198700 95956 198706 95968
rect 222470 95956 222476 95968
rect 222528 95956 222534 96008
rect 173158 95888 173164 95940
rect 173216 95928 173222 95940
rect 213178 95928 213184 95940
rect 173216 95900 213184 95928
rect 173216 95888 173222 95900
rect 213178 95888 213184 95900
rect 213236 95888 213242 95940
rect 211798 95820 211804 95872
rect 211856 95860 211862 95872
rect 229002 95860 229008 95872
rect 211856 95832 229008 95860
rect 211856 95820 211862 95832
rect 229002 95820 229008 95832
rect 229060 95820 229066 95872
rect 230474 95480 230480 95532
rect 230532 95520 230538 95532
rect 232498 95520 232504 95532
rect 230532 95492 232504 95520
rect 230532 95480 230538 95492
rect 232498 95480 232504 95492
rect 232556 95480 232562 95532
rect 267642 95412 267648 95464
rect 267700 95452 267706 95464
rect 269206 95452 269212 95464
rect 267700 95424 269212 95452
rect 267700 95412 267706 95424
rect 269206 95412 269212 95424
rect 269264 95412 269270 95464
rect 226426 95208 226432 95260
rect 226484 95248 226490 95260
rect 241514 95248 241520 95260
rect 226484 95220 241520 95248
rect 226484 95208 226490 95220
rect 241514 95208 241520 95220
rect 241572 95208 241578 95260
rect 222470 95140 222476 95192
rect 222528 95180 222534 95192
rect 281718 95180 281724 95192
rect 222528 95152 281724 95180
rect 222528 95140 222534 95152
rect 281718 95140 281724 95152
rect 281776 95140 281782 95192
rect 370590 95140 370596 95192
rect 370648 95180 370654 95192
rect 413278 95180 413284 95192
rect 370648 95152 413284 95180
rect 370648 95140 370654 95152
rect 413278 95140 413284 95152
rect 413336 95140 413342 95192
rect 216122 95072 216128 95124
rect 216180 95112 216186 95124
rect 229186 95112 229192 95124
rect 216180 95084 229192 95112
rect 216180 95072 216186 95084
rect 229186 95072 229192 95084
rect 229244 95072 229250 95124
rect 391934 95072 391940 95124
rect 391992 95112 391998 95124
rect 418246 95112 418252 95124
rect 391992 95084 418252 95112
rect 391992 95072 391998 95084
rect 418246 95072 418252 95084
rect 418304 95072 418310 95124
rect 66070 94460 66076 94512
rect 66128 94500 66134 94512
rect 97258 94500 97264 94512
rect 66128 94472 97264 94500
rect 66128 94460 66134 94472
rect 97258 94460 97264 94472
rect 97316 94460 97322 94512
rect 162118 94460 162124 94512
rect 162176 94500 162182 94512
rect 173342 94500 173348 94512
rect 162176 94472 173348 94500
rect 162176 94460 162182 94472
rect 173342 94460 173348 94472
rect 173400 94460 173406 94512
rect 202322 94460 202328 94512
rect 202380 94500 202386 94512
rect 214650 94500 214656 94512
rect 202380 94472 214656 94500
rect 202380 94460 202386 94472
rect 214650 94460 214656 94472
rect 214708 94460 214714 94512
rect 275922 94460 275928 94512
rect 275980 94500 275986 94512
rect 331950 94500 331956 94512
rect 275980 94472 331956 94500
rect 275980 94460 275986 94472
rect 331950 94460 331956 94472
rect 332008 94460 332014 94512
rect 418246 94460 418252 94512
rect 418304 94500 418310 94512
rect 582742 94500 582748 94512
rect 418304 94472 582748 94500
rect 418304 94460 418310 94472
rect 582742 94460 582748 94472
rect 582800 94460 582806 94512
rect 398834 94120 398840 94172
rect 398892 94160 398898 94172
rect 399662 94160 399668 94172
rect 398892 94132 399668 94160
rect 398892 94120 398898 94132
rect 399662 94120 399668 94132
rect 399720 94120 399726 94172
rect 130746 93916 130752 93968
rect 130804 93956 130810 93968
rect 167638 93956 167644 93968
rect 130804 93928 167644 93956
rect 130804 93916 130810 93928
rect 167638 93916 167644 93928
rect 167696 93916 167702 93968
rect 405734 93916 405740 93968
rect 405792 93956 405798 93968
rect 406470 93956 406476 93968
rect 405792 93928 406476 93956
rect 405792 93916 405798 93928
rect 406470 93916 406476 93928
rect 406528 93916 406534 93968
rect 113174 93848 113180 93900
rect 113232 93888 113238 93900
rect 153194 93888 153200 93900
rect 113232 93860 153200 93888
rect 113232 93848 113238 93860
rect 153194 93848 153200 93860
rect 153252 93848 153258 93900
rect 187602 93780 187608 93832
rect 187660 93820 187666 93832
rect 220814 93820 220820 93832
rect 187660 93792 220820 93820
rect 187660 93780 187666 93792
rect 220814 93780 220820 93792
rect 220872 93780 220878 93832
rect 266262 93780 266268 93832
rect 266320 93820 266326 93832
rect 279326 93820 279332 93832
rect 266320 93792 279332 93820
rect 266320 93780 266326 93792
rect 279326 93780 279332 93792
rect 279384 93780 279390 93832
rect 398098 93780 398104 93832
rect 398156 93820 398162 93832
rect 434714 93820 434720 93832
rect 398156 93792 434720 93820
rect 398156 93780 398162 93792
rect 434714 93780 434720 93792
rect 434772 93780 434778 93832
rect 260742 93712 260748 93764
rect 260800 93752 260806 93764
rect 273990 93752 273996 93764
rect 260800 93724 273996 93752
rect 260800 93712 260806 93724
rect 273990 93712 273996 93724
rect 274048 93712 274054 93764
rect 123018 93168 123024 93220
rect 123076 93208 123082 93220
rect 171962 93208 171968 93220
rect 123076 93180 171968 93208
rect 123076 93168 123082 93180
rect 171962 93168 171968 93180
rect 172020 93168 172026 93220
rect 213178 93168 213184 93220
rect 213236 93208 213242 93220
rect 232590 93208 232596 93220
rect 213236 93180 232596 93208
rect 213236 93168 213242 93180
rect 232590 93168 232596 93180
rect 232648 93168 232654 93220
rect 376018 93168 376024 93220
rect 376076 93208 376082 93220
rect 419626 93208 419632 93220
rect 376076 93180 419632 93208
rect 376076 93168 376082 93180
rect 419626 93168 419632 93180
rect 419684 93168 419690 93220
rect 119706 93100 119712 93152
rect 119764 93140 119770 93152
rect 175918 93140 175924 93152
rect 119764 93112 175924 93140
rect 119764 93100 119770 93112
rect 175918 93100 175924 93112
rect 175976 93100 175982 93152
rect 200850 93100 200856 93152
rect 200908 93140 200914 93152
rect 210418 93140 210424 93152
rect 200908 93112 210424 93140
rect 200908 93100 200914 93112
rect 210418 93100 210424 93112
rect 210476 93100 210482 93152
rect 222838 93100 222844 93152
rect 222896 93140 222902 93152
rect 243722 93140 243728 93152
rect 222896 93112 243728 93140
rect 222896 93100 222902 93112
rect 243722 93100 243728 93112
rect 243780 93100 243786 93152
rect 273898 93100 273904 93152
rect 273956 93140 273962 93152
rect 395522 93140 395528 93152
rect 273956 93112 395528 93140
rect 273956 93100 273962 93112
rect 395522 93100 395528 93112
rect 395580 93100 395586 93152
rect 426618 92488 426624 92540
rect 426676 92528 426682 92540
rect 582926 92528 582932 92540
rect 426676 92500 582932 92528
rect 426676 92488 426682 92500
rect 582926 92488 582932 92500
rect 582984 92488 582990 92540
rect 134426 92420 134432 92472
rect 134484 92460 134490 92472
rect 166442 92460 166448 92472
rect 134484 92432 166448 92460
rect 134484 92420 134490 92432
rect 166442 92420 166448 92432
rect 166500 92420 166506 92472
rect 209682 92420 209688 92472
rect 209740 92460 209746 92472
rect 281810 92460 281816 92472
rect 209740 92432 281816 92460
rect 209740 92420 209746 92432
rect 281810 92420 281816 92432
rect 281868 92420 281874 92472
rect 67450 91740 67456 91792
rect 67508 91780 67514 91792
rect 100018 91780 100024 91792
rect 67508 91752 100024 91780
rect 67508 91740 67514 91752
rect 100018 91740 100024 91752
rect 100076 91740 100082 91792
rect 215938 91740 215944 91792
rect 215996 91780 216002 91792
rect 242526 91780 242532 91792
rect 215996 91752 242532 91780
rect 215996 91740 216002 91752
rect 242526 91740 242532 91752
rect 242584 91740 242590 91792
rect 298094 91740 298100 91792
rect 298152 91780 298158 91792
rect 424134 91780 424140 91792
rect 298152 91752 424140 91780
rect 298152 91740 298158 91752
rect 424134 91740 424140 91752
rect 424192 91740 424198 91792
rect 126698 91400 126704 91452
rect 126756 91440 126762 91452
rect 128998 91440 129004 91452
rect 126756 91412 129004 91440
rect 126756 91400 126762 91412
rect 128998 91400 129004 91412
rect 129056 91400 129062 91452
rect 162118 91332 162124 91384
rect 162176 91372 162182 91384
rect 168282 91372 168288 91384
rect 162176 91344 168288 91372
rect 162176 91332 162182 91344
rect 168282 91332 168288 91344
rect 168340 91332 168346 91384
rect 97350 91128 97356 91180
rect 97408 91168 97414 91180
rect 104158 91168 104164 91180
rect 97408 91140 104164 91168
rect 97408 91128 97414 91140
rect 104158 91128 104164 91140
rect 104216 91128 104222 91180
rect 133782 91168 133788 91180
rect 122806 91140 133788 91168
rect 74810 91060 74816 91112
rect 74868 91100 74874 91112
rect 89714 91100 89720 91112
rect 74868 91072 89720 91100
rect 74868 91060 74874 91072
rect 89714 91060 89720 91072
rect 89772 91060 89778 91112
rect 100110 91060 100116 91112
rect 100168 91100 100174 91112
rect 108298 91100 108304 91112
rect 100168 91072 108304 91100
rect 100168 91060 100174 91072
rect 108298 91060 108304 91072
rect 108356 91060 108362 91112
rect 108574 91060 108580 91112
rect 108632 91100 108638 91112
rect 116578 91100 116584 91112
rect 108632 91072 116584 91100
rect 108632 91060 108638 91072
rect 116578 91060 116584 91072
rect 116636 91060 116642 91112
rect 116762 91060 116768 91112
rect 116820 91100 116826 91112
rect 122806 91100 122834 91140
rect 133782 91128 133788 91140
rect 133840 91128 133846 91180
rect 116820 91072 122834 91100
rect 116820 91060 116826 91072
rect 151354 91060 151360 91112
rect 151412 91100 151418 91112
rect 158714 91100 158720 91112
rect 151412 91072 158720 91100
rect 151412 91060 151418 91072
rect 158714 91060 158720 91072
rect 158772 91060 158778 91112
rect 411346 91060 411352 91112
rect 411404 91100 411410 91112
rect 411898 91100 411904 91112
rect 411404 91072 411904 91100
rect 411404 91060 411410 91072
rect 411898 91060 411904 91072
rect 411956 91100 411962 91112
rect 582374 91100 582380 91112
rect 411956 91072 582380 91100
rect 411956 91060 411962 91072
rect 582374 91060 582380 91072
rect 582432 91060 582438 91112
rect 103146 90992 103152 91044
rect 103204 91032 103210 91044
rect 188522 91032 188528 91044
rect 103204 91004 188528 91032
rect 103204 90992 103210 91004
rect 188522 90992 188528 91004
rect 188580 90992 188586 91044
rect 381630 90992 381636 91044
rect 381688 91032 381694 91044
rect 426618 91032 426624 91044
rect 381688 91004 426624 91032
rect 381688 90992 381694 91004
rect 426618 90992 426624 91004
rect 426676 90992 426682 91044
rect 124122 90924 124128 90976
rect 124180 90964 124186 90976
rect 207750 90964 207756 90976
rect 124180 90936 207756 90964
rect 124180 90924 124186 90936
rect 207750 90924 207756 90936
rect 207808 90924 207814 90976
rect 220078 90380 220084 90432
rect 220136 90420 220142 90432
rect 238386 90420 238392 90432
rect 220136 90392 238392 90420
rect 220136 90380 220142 90392
rect 238386 90380 238392 90392
rect 238444 90380 238450 90432
rect 67358 90312 67364 90364
rect 67416 90352 67422 90364
rect 106918 90352 106924 90364
rect 67416 90324 106924 90352
rect 67416 90312 67422 90324
rect 106918 90312 106924 90324
rect 106976 90312 106982 90364
rect 206370 90312 206376 90364
rect 206428 90352 206434 90364
rect 263134 90352 263140 90364
rect 206428 90324 263140 90352
rect 206428 90312 206434 90324
rect 263134 90312 263140 90324
rect 263192 90312 263198 90364
rect 121178 89632 121184 89684
rect 121236 89672 121242 89684
rect 177482 89672 177488 89684
rect 121236 89644 177488 89672
rect 121236 89632 121242 89644
rect 177482 89632 177488 89644
rect 177540 89632 177546 89684
rect 217226 89632 217232 89684
rect 217284 89672 217290 89684
rect 279050 89672 279056 89684
rect 217284 89644 279056 89672
rect 217284 89632 217290 89644
rect 279050 89632 279056 89644
rect 279108 89632 279114 89684
rect 158714 89564 158720 89616
rect 158772 89604 158778 89616
rect 177298 89604 177304 89616
rect 158772 89576 177304 89604
rect 158772 89564 158778 89576
rect 177298 89564 177304 89576
rect 177356 89564 177362 89616
rect 209130 88952 209136 89004
rect 209188 88992 209194 89004
rect 234062 88992 234068 89004
rect 209188 88964 234068 88992
rect 209188 88952 209194 88964
rect 234062 88952 234068 88964
rect 234120 88952 234126 89004
rect 349890 88952 349896 89004
rect 349948 88992 349954 89004
rect 357434 88992 357440 89004
rect 349948 88964 357440 88992
rect 349948 88952 349954 88964
rect 357434 88952 357440 88964
rect 357492 88992 357498 89004
rect 426526 88992 426532 89004
rect 357492 88964 426532 88992
rect 357492 88952 357498 88964
rect 426526 88952 426532 88964
rect 426584 88952 426590 89004
rect 117130 88272 117136 88324
rect 117188 88312 117194 88324
rect 170490 88312 170496 88324
rect 117188 88284 170496 88312
rect 117188 88272 117194 88284
rect 170490 88272 170496 88284
rect 170548 88272 170554 88324
rect 267826 88272 267832 88324
rect 267884 88312 267890 88324
rect 410058 88312 410064 88324
rect 267884 88284 410064 88312
rect 267884 88272 267890 88284
rect 410058 88272 410064 88284
rect 410116 88272 410122 88324
rect 121822 88204 121828 88256
rect 121880 88244 121886 88256
rect 171870 88244 171876 88256
rect 121880 88216 171876 88244
rect 121880 88204 121886 88216
rect 171870 88204 171876 88216
rect 171928 88204 171934 88256
rect 379514 88204 379520 88256
rect 379572 88244 379578 88256
rect 429746 88244 429752 88256
rect 379572 88216 429752 88244
rect 379572 88204 379578 88216
rect 429746 88204 429752 88216
rect 429804 88204 429810 88256
rect 170766 87660 170772 87712
rect 170824 87700 170830 87712
rect 196894 87700 196900 87712
rect 170824 87672 196900 87700
rect 170824 87660 170830 87672
rect 196894 87660 196900 87672
rect 196952 87660 196958 87712
rect 224310 87660 224316 87712
rect 224368 87700 224374 87712
rect 256234 87700 256240 87712
rect 224368 87672 256240 87700
rect 224368 87660 224374 87672
rect 256234 87660 256240 87672
rect 256292 87660 256298 87712
rect 3510 87592 3516 87644
rect 3568 87632 3574 87644
rect 33778 87632 33784 87644
rect 3568 87604 33784 87632
rect 3568 87592 3574 87604
rect 33778 87592 33784 87604
rect 33836 87592 33842 87644
rect 95050 87592 95056 87644
rect 95108 87632 95114 87644
rect 115198 87632 115204 87644
rect 95108 87604 115204 87632
rect 95108 87592 95114 87604
rect 115198 87592 115204 87604
rect 115256 87592 115262 87644
rect 196802 87592 196808 87644
rect 196860 87632 196866 87644
rect 247954 87632 247960 87644
rect 196860 87604 247960 87632
rect 196860 87592 196866 87604
rect 247954 87592 247960 87604
rect 248012 87592 248018 87644
rect 304258 87592 304264 87644
rect 304316 87632 304322 87644
rect 379514 87632 379520 87644
rect 304316 87604 379520 87632
rect 304316 87592 304322 87604
rect 379514 87592 379520 87604
rect 379572 87592 379578 87644
rect 108482 86912 108488 86964
rect 108540 86952 108546 86964
rect 189902 86952 189908 86964
rect 108540 86924 189908 86952
rect 108540 86912 108546 86924
rect 189902 86912 189908 86924
rect 189960 86912 189966 86964
rect 257338 86912 257344 86964
rect 257396 86952 257402 86964
rect 257982 86952 257988 86964
rect 257396 86924 257988 86952
rect 257396 86912 257402 86924
rect 257982 86912 257988 86924
rect 258040 86952 258046 86964
rect 402054 86952 402060 86964
rect 258040 86924 402060 86952
rect 258040 86912 258046 86924
rect 402054 86912 402060 86924
rect 402112 86912 402118 86964
rect 152458 86844 152464 86896
rect 152516 86884 152522 86896
rect 169110 86884 169116 86896
rect 152516 86856 169116 86884
rect 152516 86844 152522 86856
rect 169110 86844 169116 86856
rect 169168 86844 169174 86896
rect 214558 86300 214564 86352
rect 214616 86340 214622 86352
rect 229830 86340 229836 86352
rect 214616 86312 229836 86340
rect 214616 86300 214622 86312
rect 229830 86300 229836 86312
rect 229888 86300 229894 86352
rect 181530 86232 181536 86284
rect 181588 86272 181594 86284
rect 261754 86272 261760 86284
rect 181588 86244 261760 86272
rect 181588 86232 181594 86244
rect 261754 86232 261760 86244
rect 261812 86232 261818 86284
rect 397362 86232 397368 86284
rect 397420 86272 397426 86284
rect 583018 86272 583024 86284
rect 397420 86244 583024 86272
rect 397420 86232 397426 86244
rect 583018 86232 583024 86244
rect 583076 86232 583082 86284
rect 582374 86028 582380 86080
rect 582432 86068 582438 86080
rect 582926 86068 582932 86080
rect 582432 86040 582932 86068
rect 582432 86028 582438 86040
rect 582926 86028 582932 86040
rect 582984 86028 582990 86080
rect 115750 85484 115756 85536
rect 115808 85524 115814 85536
rect 193950 85524 193956 85536
rect 115808 85496 193956 85524
rect 115808 85484 115814 85496
rect 193950 85484 193956 85496
rect 194008 85484 194014 85536
rect 203518 85484 203524 85536
rect 203576 85524 203582 85536
rect 280154 85524 280160 85536
rect 203576 85496 280160 85524
rect 203576 85484 203582 85496
rect 280154 85484 280160 85496
rect 280212 85484 280218 85536
rect 151722 85416 151728 85468
rect 151780 85456 151786 85468
rect 166350 85456 166356 85468
rect 151780 85428 166356 85456
rect 151780 85416 151786 85428
rect 166350 85416 166356 85428
rect 166408 85416 166414 85468
rect 63402 84804 63408 84856
rect 63460 84844 63466 84856
rect 115290 84844 115296 84856
rect 63460 84816 115296 84844
rect 63460 84804 63466 84816
rect 115290 84804 115296 84816
rect 115348 84804 115354 84856
rect 210418 84804 210424 84856
rect 210476 84844 210482 84856
rect 245102 84844 245108 84856
rect 210476 84816 245108 84844
rect 210476 84804 210482 84816
rect 245102 84804 245108 84816
rect 245160 84804 245166 84856
rect 309778 84804 309784 84856
rect 309836 84844 309842 84856
rect 441706 84844 441712 84856
rect 309836 84816 441712 84844
rect 309836 84804 309842 84816
rect 441706 84804 441712 84816
rect 441764 84804 441770 84856
rect 126790 84124 126796 84176
rect 126848 84164 126854 84176
rect 167730 84164 167736 84176
rect 126848 84136 167736 84164
rect 126848 84124 126854 84136
rect 167730 84124 167736 84136
rect 167788 84124 167794 84176
rect 189810 84124 189816 84176
rect 189868 84164 189874 84176
rect 427998 84164 428004 84176
rect 189868 84136 428004 84164
rect 189868 84124 189874 84136
rect 427998 84124 428004 84136
rect 428056 84124 428062 84176
rect 114370 84056 114376 84108
rect 114428 84096 114434 84108
rect 203702 84096 203708 84108
rect 114428 84068 203708 84096
rect 114428 84056 114434 84068
rect 203702 84056 203708 84068
rect 203760 84056 203766 84108
rect 57882 83444 57888 83496
rect 57940 83484 57946 83496
rect 98638 83484 98644 83496
rect 57940 83456 98644 83484
rect 57940 83444 57946 83456
rect 98638 83444 98644 83456
rect 98696 83444 98702 83496
rect 213270 83444 213276 83496
rect 213328 83484 213334 83496
rect 252094 83484 252100 83496
rect 213328 83456 252100 83484
rect 213328 83444 213334 83456
rect 252094 83444 252100 83456
rect 252152 83444 252158 83496
rect 324958 83444 324964 83496
rect 325016 83484 325022 83496
rect 441798 83484 441804 83496
rect 325016 83456 441804 83484
rect 325016 83444 325022 83456
rect 441798 83444 441804 83456
rect 441856 83444 441862 83496
rect 86862 82764 86868 82816
rect 86920 82804 86926 82816
rect 164878 82804 164884 82816
rect 86920 82776 164884 82804
rect 86920 82764 86926 82776
rect 164878 82764 164884 82776
rect 164936 82764 164942 82816
rect 313918 82764 313924 82816
rect 313976 82804 313982 82816
rect 435450 82804 435456 82816
rect 313976 82776 435456 82804
rect 313976 82764 313982 82776
rect 435450 82764 435456 82776
rect 435508 82764 435514 82816
rect 198090 82152 198096 82204
rect 198148 82192 198154 82204
rect 232774 82192 232780 82204
rect 198148 82164 232780 82192
rect 198148 82152 198154 82164
rect 232774 82152 232780 82164
rect 232832 82152 232838 82204
rect 160830 82084 160836 82136
rect 160888 82124 160894 82136
rect 213362 82124 213368 82136
rect 160888 82096 213368 82124
rect 160888 82084 160894 82096
rect 213362 82084 213368 82096
rect 213420 82084 213426 82136
rect 216122 82084 216128 82136
rect 216180 82124 216186 82136
rect 249242 82124 249248 82136
rect 216180 82096 249248 82124
rect 216180 82084 216186 82096
rect 249242 82084 249248 82096
rect 249300 82084 249306 82136
rect 359458 82084 359464 82136
rect 359516 82124 359522 82136
rect 441890 82124 441896 82136
rect 359516 82096 441896 82124
rect 359516 82084 359522 82096
rect 441890 82084 441896 82096
rect 441948 82084 441954 82136
rect 95142 81336 95148 81388
rect 95200 81376 95206 81388
rect 173250 81376 173256 81388
rect 95200 81348 173256 81376
rect 95200 81336 95206 81348
rect 173250 81336 173256 81348
rect 173308 81336 173314 81388
rect 204990 81336 204996 81388
rect 205048 81376 205054 81388
rect 281534 81376 281540 81388
rect 205048 81348 281540 81376
rect 205048 81336 205054 81348
rect 281534 81336 281540 81348
rect 281592 81336 281598 81388
rect 347038 81336 347044 81388
rect 347096 81376 347102 81388
rect 408494 81376 408500 81388
rect 347096 81348 408500 81376
rect 347096 81336 347102 81348
rect 408494 81336 408500 81348
rect 408552 81336 408558 81388
rect 119982 81268 119988 81320
rect 120040 81308 120046 81320
rect 170674 81308 170680 81320
rect 120040 81280 170680 81308
rect 120040 81268 120046 81280
rect 170674 81268 170680 81280
rect 170732 81268 170738 81320
rect 331214 80656 331220 80708
rect 331272 80696 331278 80708
rect 340138 80696 340144 80708
rect 331272 80668 340144 80696
rect 331272 80656 331278 80668
rect 340138 80656 340144 80668
rect 340196 80696 340202 80708
rect 355318 80696 355324 80708
rect 340196 80668 355324 80696
rect 340196 80656 340202 80668
rect 355318 80656 355324 80668
rect 355376 80656 355382 80708
rect 111610 79976 111616 80028
rect 111668 80016 111674 80028
rect 172054 80016 172060 80028
rect 111668 79988 172060 80016
rect 111668 79976 111674 79988
rect 172054 79976 172060 79988
rect 172112 79976 172118 80028
rect 200758 79976 200764 80028
rect 200816 80016 200822 80028
rect 411898 80016 411904 80028
rect 200816 79988 411904 80016
rect 200816 79976 200822 79988
rect 411898 79976 411904 79988
rect 411956 79976 411962 80028
rect 125502 79908 125508 79960
rect 125560 79948 125566 79960
rect 178862 79948 178868 79960
rect 125560 79920 178868 79948
rect 125560 79908 125566 79920
rect 178862 79908 178868 79920
rect 178920 79908 178926 79960
rect 337470 79296 337476 79348
rect 337528 79336 337534 79348
rect 440418 79336 440424 79348
rect 337528 79308 440424 79336
rect 337528 79296 337534 79308
rect 440418 79296 440424 79308
rect 440476 79296 440482 79348
rect 124030 78616 124036 78668
rect 124088 78656 124094 78668
rect 166258 78656 166264 78668
rect 124088 78628 166264 78656
rect 124088 78616 124094 78628
rect 166258 78616 166264 78628
rect 166316 78616 166322 78668
rect 270494 78616 270500 78668
rect 270552 78656 270558 78668
rect 271046 78656 271052 78668
rect 270552 78628 271052 78656
rect 270552 78616 270558 78628
rect 271046 78616 271052 78628
rect 271104 78656 271110 78668
rect 438854 78656 438860 78668
rect 271104 78628 438860 78656
rect 271104 78616 271110 78628
rect 438854 78616 438860 78628
rect 438912 78616 438918 78668
rect 240962 78004 240968 78056
rect 241020 78044 241026 78056
rect 271046 78044 271052 78056
rect 241020 78016 271052 78044
rect 241020 78004 241026 78016
rect 271046 78004 271052 78016
rect 271104 78004 271110 78056
rect 34422 77936 34428 77988
rect 34480 77976 34486 77988
rect 241054 77976 241060 77988
rect 34480 77948 241060 77976
rect 34480 77936 34486 77948
rect 241054 77936 241060 77948
rect 241112 77936 241118 77988
rect 100018 77188 100024 77240
rect 100076 77228 100082 77240
rect 170766 77228 170772 77240
rect 100076 77200 170772 77228
rect 100076 77188 100082 77200
rect 170766 77188 170772 77200
rect 170824 77188 170830 77240
rect 132402 77120 132408 77172
rect 132460 77160 132466 77172
rect 176010 77160 176016 77172
rect 132460 77132 176016 77160
rect 132460 77120 132466 77132
rect 176010 77120 176016 77132
rect 176068 77120 176074 77172
rect 246390 76508 246396 76560
rect 246448 76548 246454 76560
rect 404446 76548 404452 76560
rect 246448 76520 404452 76548
rect 246448 76508 246454 76520
rect 404446 76508 404452 76520
rect 404504 76508 404510 76560
rect 97258 75828 97264 75880
rect 97316 75868 97322 75880
rect 170582 75868 170588 75880
rect 97316 75840 170588 75868
rect 97316 75828 97322 75840
rect 170582 75828 170588 75840
rect 170640 75828 170646 75880
rect 151538 75760 151544 75812
rect 151596 75800 151602 75812
rect 181438 75800 181444 75812
rect 151596 75772 181444 75800
rect 151596 75760 151602 75772
rect 181438 75760 181444 75772
rect 181496 75760 181502 75812
rect 278682 75148 278688 75200
rect 278740 75188 278746 75200
rect 448698 75188 448704 75200
rect 278740 75160 448704 75188
rect 278740 75148 278746 75160
rect 448698 75148 448704 75160
rect 448756 75148 448762 75200
rect 129642 74468 129648 74520
rect 129700 74508 129706 74520
rect 210602 74508 210608 74520
rect 129700 74480 210608 74508
rect 129700 74468 129706 74480
rect 210602 74468 210608 74480
rect 210660 74468 210666 74520
rect 91002 74400 91008 74452
rect 91060 74440 91066 74452
rect 160830 74440 160836 74452
rect 91060 74412 160836 74440
rect 91060 74400 91066 74412
rect 160830 74400 160836 74412
rect 160888 74400 160894 74452
rect 218698 73856 218704 73908
rect 218756 73896 218762 73908
rect 239674 73896 239680 73908
rect 218756 73868 239680 73896
rect 218756 73856 218762 73868
rect 239674 73856 239680 73868
rect 239732 73856 239738 73908
rect 160738 73788 160744 73840
rect 160796 73828 160802 73840
rect 218790 73828 218796 73840
rect 160796 73800 218796 73828
rect 160796 73788 160802 73800
rect 218790 73788 218796 73800
rect 218848 73788 218854 73840
rect 106918 73108 106924 73160
rect 106976 73148 106982 73160
rect 214742 73148 214748 73160
rect 106976 73120 214748 73148
rect 106976 73108 106982 73120
rect 214742 73108 214748 73120
rect 214800 73108 214806 73160
rect 114462 73040 114468 73092
rect 114520 73080 114526 73092
rect 174538 73080 174544 73092
rect 114520 73052 174544 73080
rect 114520 73040 114526 73052
rect 174538 73040 174544 73052
rect 174596 73040 174602 73092
rect 301498 72428 301504 72480
rect 301556 72468 301562 72480
rect 398834 72468 398840 72480
rect 301556 72440 398840 72468
rect 301556 72428 301562 72440
rect 398834 72428 398840 72440
rect 398892 72428 398898 72480
rect 118602 71680 118608 71732
rect 118660 71720 118666 71732
rect 195422 71720 195428 71732
rect 118660 71692 195428 71720
rect 118660 71680 118666 71692
rect 195422 71680 195428 71692
rect 195480 71680 195486 71732
rect 102042 71612 102048 71664
rect 102100 71652 102106 71664
rect 178770 71652 178776 71664
rect 102100 71624 178776 71652
rect 102100 71612 102106 71624
rect 178770 71612 178776 71624
rect 178828 71612 178834 71664
rect 128998 70320 129004 70372
rect 129056 70360 129062 70372
rect 171778 70360 171784 70372
rect 129056 70332 171784 70360
rect 129056 70320 129062 70332
rect 171778 70320 171784 70332
rect 171836 70320 171842 70372
rect 119982 69640 119988 69692
rect 120040 69680 120046 69692
rect 251910 69680 251916 69692
rect 120040 69652 251916 69680
rect 120040 69640 120046 69652
rect 251910 69640 251916 69652
rect 251968 69640 251974 69692
rect 289078 69640 289084 69692
rect 289136 69680 289142 69692
rect 383102 69680 383108 69692
rect 289136 69652 383108 69680
rect 289136 69640 289142 69652
rect 383102 69640 383108 69652
rect 383160 69640 383166 69692
rect 85482 68960 85488 69012
rect 85540 69000 85546 69012
rect 169294 69000 169300 69012
rect 85540 68972 169300 69000
rect 85540 68960 85546 68972
rect 169294 68960 169300 68972
rect 169352 68960 169358 69012
rect 322934 68960 322940 69012
rect 322992 69000 322998 69012
rect 323670 69000 323676 69012
rect 322992 68972 323676 69000
rect 322992 68960 322998 68972
rect 323670 68960 323676 68972
rect 323728 69000 323734 69012
rect 416866 69000 416872 69012
rect 323728 68972 416872 69000
rect 323728 68960 323734 68972
rect 416866 68960 416872 68972
rect 416924 68960 416930 69012
rect 126698 68892 126704 68944
rect 126756 68932 126762 68944
rect 199378 68932 199384 68944
rect 126756 68904 199384 68932
rect 126756 68892 126762 68904
rect 199378 68892 199384 68904
rect 199436 68892 199442 68944
rect 67634 67532 67640 67584
rect 67692 67572 67698 67584
rect 187050 67572 187056 67584
rect 67692 67544 187056 67572
rect 67692 67532 67698 67544
rect 187050 67532 187056 67544
rect 187108 67532 187114 67584
rect 93670 67464 93676 67516
rect 93728 67504 93734 67516
rect 205082 67504 205088 67516
rect 93728 67476 205088 67504
rect 93728 67464 93734 67476
rect 205082 67464 205088 67476
rect 205140 67464 205146 67516
rect 330478 66852 330484 66904
rect 330536 66892 330542 66904
rect 441614 66892 441620 66904
rect 330536 66864 441620 66892
rect 330536 66852 330542 66864
rect 441614 66852 441620 66864
rect 441672 66852 441678 66904
rect 115198 66172 115204 66224
rect 115256 66212 115262 66224
rect 207658 66212 207664 66224
rect 115256 66184 207664 66212
rect 115256 66172 115262 66184
rect 207658 66172 207664 66184
rect 207716 66172 207722 66224
rect 122742 66104 122748 66156
rect 122800 66144 122806 66156
rect 170398 66144 170404 66156
rect 122800 66116 170404 66144
rect 122800 66104 122806 66116
rect 170398 66104 170404 66116
rect 170456 66104 170462 66156
rect 332594 65492 332600 65544
rect 332652 65532 332658 65544
rect 352650 65532 352656 65544
rect 332652 65504 352656 65532
rect 332652 65492 332658 65504
rect 352650 65492 352656 65504
rect 352708 65492 352714 65544
rect 104158 64812 104164 64864
rect 104216 64852 104222 64864
rect 192478 64852 192484 64864
rect 104216 64824 192484 64852
rect 104216 64812 104222 64824
rect 192478 64812 192484 64824
rect 192536 64812 192542 64864
rect 331858 64812 331864 64864
rect 331916 64852 331922 64864
rect 401594 64852 401600 64864
rect 331916 64824 401600 64852
rect 331916 64812 331922 64824
rect 401594 64812 401600 64824
rect 401652 64812 401658 64864
rect 121362 64744 121368 64796
rect 121420 64784 121426 64796
rect 173158 64784 173164 64796
rect 121420 64756 173164 64784
rect 121420 64744 121426 64756
rect 173158 64744 173164 64756
rect 173216 64744 173222 64796
rect 318150 64132 318156 64184
rect 318208 64172 318214 64184
rect 331858 64172 331864 64184
rect 318208 64144 331864 64172
rect 318208 64132 318214 64144
rect 331858 64132 331864 64144
rect 331916 64132 331922 64184
rect 108298 63452 108304 63504
rect 108356 63492 108362 63504
rect 193858 63492 193864 63504
rect 108356 63464 193864 63492
rect 108356 63452 108362 63464
rect 193858 63452 193864 63464
rect 193916 63452 193922 63504
rect 355318 63452 355324 63504
rect 355376 63492 355382 63504
rect 436094 63492 436100 63504
rect 355376 63464 436100 63492
rect 355376 63452 355382 63464
rect 436094 63452 436100 63464
rect 436152 63452 436158 63504
rect 68922 62772 68928 62824
rect 68980 62812 68986 62824
rect 253198 62812 253204 62824
rect 68980 62784 253204 62812
rect 68980 62772 68986 62784
rect 253198 62772 253204 62784
rect 253256 62772 253262 62824
rect 308398 62772 308404 62824
rect 308456 62812 308462 62824
rect 353938 62812 353944 62824
rect 308456 62784 353944 62812
rect 308456 62772 308462 62784
rect 353938 62772 353944 62784
rect 353996 62772 354002 62824
rect 111702 62024 111708 62076
rect 111760 62064 111766 62076
rect 200850 62064 200856 62076
rect 111760 62036 200856 62064
rect 111760 62024 111766 62036
rect 200850 62024 200856 62036
rect 200908 62024 200914 62076
rect 73062 61344 73068 61396
rect 73120 61384 73126 61396
rect 262950 61384 262956 61396
rect 73120 61356 262956 61384
rect 73120 61344 73126 61356
rect 262950 61344 262956 61356
rect 263008 61344 263014 61396
rect 288342 61344 288348 61396
rect 288400 61384 288406 61396
rect 419718 61384 419724 61396
rect 288400 61356 419724 61384
rect 288400 61344 288406 61356
rect 419718 61344 419724 61356
rect 419776 61344 419782 61396
rect 99282 60664 99288 60716
rect 99340 60704 99346 60716
rect 197998 60704 198004 60716
rect 99340 60676 198004 60704
rect 99340 60664 99346 60676
rect 197998 60664 198004 60676
rect 198056 60664 198062 60716
rect 271874 60664 271880 60716
rect 271932 60704 271938 60716
rect 359550 60704 359556 60716
rect 271932 60676 359556 60704
rect 271932 60664 271938 60676
rect 359550 60664 359556 60676
rect 359608 60664 359614 60716
rect 269114 60256 269120 60308
rect 269172 60296 269178 60308
rect 271874 60296 271880 60308
rect 269172 60268 271880 60296
rect 269172 60256 269178 60268
rect 271874 60256 271880 60268
rect 271932 60256 271938 60308
rect 70302 59984 70308 60036
rect 70360 60024 70366 60036
rect 245010 60024 245016 60036
rect 70360 59996 245016 60024
rect 70360 59984 70366 59996
rect 245010 59984 245016 59996
rect 245068 59984 245074 60036
rect 3050 59304 3056 59356
rect 3108 59344 3114 59356
rect 11698 59344 11704 59356
rect 3108 59316 11704 59344
rect 3108 59304 3114 59316
rect 11698 59304 11704 59316
rect 11756 59304 11762 59356
rect 103422 59304 103428 59356
rect 103480 59344 103486 59356
rect 184290 59344 184296 59356
rect 103480 59316 184296 59344
rect 103480 59304 103486 59316
rect 184290 59304 184296 59316
rect 184348 59304 184354 59356
rect 66162 58624 66168 58676
rect 66220 58664 66226 58676
rect 260282 58664 260288 58676
rect 66220 58636 260288 58664
rect 66220 58624 66226 58636
rect 260282 58624 260288 58636
rect 260340 58624 260346 58676
rect 271138 58624 271144 58676
rect 271196 58664 271202 58676
rect 423674 58664 423680 58676
rect 271196 58636 423680 58664
rect 271196 58624 271202 58636
rect 423674 58624 423680 58636
rect 423732 58624 423738 58676
rect 104802 57876 104808 57928
rect 104860 57916 104866 57928
rect 202322 57916 202328 57928
rect 104860 57888 202328 57916
rect 104860 57876 104866 57888
rect 202322 57876 202328 57888
rect 202380 57876 202386 57928
rect 91002 57196 91008 57248
rect 91060 57236 91066 57248
rect 264422 57236 264428 57248
rect 91060 57208 264428 57236
rect 91060 57196 91066 57208
rect 264422 57196 264428 57208
rect 264480 57196 264486 57248
rect 112990 56516 112996 56568
rect 113048 56556 113054 56568
rect 182818 56556 182824 56568
rect 113048 56528 182824 56556
rect 113048 56516 113054 56528
rect 182818 56516 182824 56528
rect 182876 56516 182882 56568
rect 97902 55836 97908 55888
rect 97960 55876 97966 55888
rect 256050 55876 256056 55888
rect 97960 55848 256056 55876
rect 97960 55836 97966 55848
rect 256050 55836 256056 55848
rect 256108 55836 256114 55888
rect 260374 55836 260380 55888
rect 260432 55876 260438 55888
rect 381538 55876 381544 55888
rect 260432 55848 381544 55876
rect 260432 55836 260438 55848
rect 381538 55836 381544 55848
rect 381596 55836 381602 55888
rect 381630 55836 381636 55888
rect 381688 55876 381694 55888
rect 447318 55876 447324 55888
rect 381688 55848 447324 55876
rect 381688 55836 381694 55848
rect 447318 55836 447324 55848
rect 447376 55836 447382 55888
rect 107470 55156 107476 55208
rect 107528 55196 107534 55208
rect 203610 55196 203616 55208
rect 107528 55168 203616 55196
rect 107528 55156 107534 55168
rect 203610 55156 203616 55168
rect 203668 55156 203674 55208
rect 311894 55156 311900 55208
rect 311952 55196 311958 55208
rect 405826 55196 405832 55208
rect 311952 55168 405832 55196
rect 311952 55156 311958 55168
rect 405826 55156 405832 55168
rect 405884 55156 405890 55208
rect 244274 54544 244280 54596
rect 244332 54584 244338 54596
rect 311894 54584 311900 54596
rect 244332 54556 311900 54584
rect 244332 54544 244338 54556
rect 311894 54544 311900 54556
rect 311952 54544 311958 54596
rect 102042 54476 102048 54528
rect 102100 54516 102106 54528
rect 250530 54516 250536 54528
rect 102100 54488 250536 54516
rect 102100 54476 102106 54488
rect 250530 54476 250536 54488
rect 250588 54476 250594 54528
rect 125410 53728 125416 53780
rect 125468 53768 125474 53780
rect 216030 53768 216036 53780
rect 125468 53740 216036 53768
rect 125468 53728 125474 53740
rect 216030 53728 216036 53740
rect 216088 53728 216094 53780
rect 89622 53048 89628 53100
rect 89680 53088 89686 53100
rect 258810 53088 258816 53100
rect 89680 53060 258816 53088
rect 89680 53048 89686 53060
rect 258810 53048 258816 53060
rect 258868 53048 258874 53100
rect 115842 52368 115848 52420
rect 115900 52408 115906 52420
rect 195330 52408 195336 52420
rect 115900 52380 195336 52408
rect 115900 52368 115906 52380
rect 195330 52368 195336 52380
rect 195388 52368 195394 52420
rect 104802 51688 104808 51740
rect 104860 51728 104866 51740
rect 267734 51728 267740 51740
rect 104860 51700 267740 51728
rect 104860 51688 104866 51700
rect 267734 51688 267740 51700
rect 267792 51688 267798 51740
rect 339494 51688 339500 51740
rect 339552 51728 339558 51740
rect 430666 51728 430672 51740
rect 339552 51700 430672 51728
rect 339552 51688 339558 51700
rect 430666 51688 430672 51700
rect 430724 51688 430730 51740
rect 110322 51008 110328 51060
rect 110380 51048 110386 51060
rect 189718 51048 189724 51060
rect 110380 51020 189724 51048
rect 110380 51008 110386 51020
rect 189718 51008 189724 51020
rect 189776 51008 189782 51060
rect 241514 51008 241520 51060
rect 241572 51048 241578 51060
rect 249794 51048 249800 51060
rect 241572 51020 249800 51048
rect 241572 51008 241578 51020
rect 249794 51008 249800 51020
rect 249852 51048 249858 51060
rect 433334 51048 433340 51060
rect 249852 51020 433340 51048
rect 249852 51008 249858 51020
rect 433334 51008 433340 51020
rect 433392 51008 433398 51060
rect 108942 50328 108948 50380
rect 109000 50368 109006 50380
rect 242250 50368 242256 50380
rect 109000 50340 242256 50368
rect 109000 50328 109006 50340
rect 242250 50328 242256 50340
rect 242308 50328 242314 50380
rect 128262 49648 128268 49700
rect 128320 49688 128326 49700
rect 180242 49688 180248 49700
rect 128320 49660 180248 49688
rect 128320 49648 128326 49660
rect 180242 49648 180248 49660
rect 180300 49648 180306 49700
rect 111702 48968 111708 49020
rect 111760 49008 111766 49020
rect 243538 49008 243544 49020
rect 111760 48980 243544 49008
rect 111760 48968 111766 48980
rect 243538 48968 243544 48980
rect 243596 48968 243602 49020
rect 247678 48968 247684 49020
rect 247736 49008 247742 49020
rect 414106 49008 414112 49020
rect 247736 48980 414112 49008
rect 247736 48968 247742 48980
rect 414106 48968 414112 48980
rect 414164 48968 414170 49020
rect 337378 48220 337384 48272
rect 337436 48260 337442 48272
rect 437474 48260 437480 48272
rect 337436 48232 437480 48260
rect 337436 48220 337442 48232
rect 437474 48220 437480 48232
rect 437532 48220 437538 48272
rect 335998 48016 336004 48068
rect 336056 48056 336062 48068
rect 337378 48056 337384 48068
rect 336056 48028 337384 48056
rect 336056 48016 336062 48028
rect 337378 48016 337384 48028
rect 337436 48016 337442 48068
rect 33042 47608 33048 47660
rect 33100 47648 33106 47660
rect 240870 47648 240876 47660
rect 33100 47620 240876 47648
rect 33100 47608 33106 47620
rect 240870 47608 240876 47620
rect 240928 47608 240934 47660
rect 67174 47540 67180 47592
rect 67232 47580 67238 47592
rect 280798 47580 280804 47592
rect 67232 47552 280804 47580
rect 67232 47540 67238 47552
rect 280798 47540 280804 47552
rect 280856 47540 280862 47592
rect 285674 47540 285680 47592
rect 285732 47580 285738 47592
rect 334710 47580 334716 47592
rect 285732 47552 334716 47580
rect 285732 47540 285738 47552
rect 334710 47540 334716 47552
rect 334768 47540 334774 47592
rect 74442 46180 74448 46232
rect 74500 46220 74506 46232
rect 262858 46220 262864 46232
rect 74500 46192 262864 46220
rect 74500 46180 74506 46192
rect 262858 46180 262864 46192
rect 262916 46180 262922 46232
rect 321554 46180 321560 46232
rect 321612 46220 321618 46232
rect 408494 46220 408500 46232
rect 321612 46192 408500 46220
rect 321612 46180 321618 46192
rect 408494 46180 408500 46192
rect 408552 46180 408558 46232
rect 44082 44888 44088 44940
rect 44140 44928 44146 44940
rect 211798 44928 211804 44940
rect 44140 44900 211804 44928
rect 44140 44888 44146 44900
rect 211798 44888 211804 44900
rect 211856 44888 211862 44940
rect 41322 44820 41328 44872
rect 41380 44860 41386 44872
rect 225598 44860 225604 44872
rect 41380 44832 225604 44860
rect 41380 44820 41386 44832
rect 225598 44820 225604 44832
rect 225656 44820 225662 44872
rect 314654 44820 314660 44872
rect 314712 44860 314718 44872
rect 444374 44860 444380 44872
rect 314712 44832 444380 44860
rect 314712 44820 314718 44832
rect 444374 44820 444380 44832
rect 444432 44820 444438 44872
rect 84102 43460 84108 43512
rect 84160 43500 84166 43512
rect 253290 43500 253296 43512
rect 84160 43472 253296 43500
rect 84160 43460 84166 43472
rect 253290 43460 253296 43472
rect 253348 43460 253354 43512
rect 29638 43392 29644 43444
rect 29696 43432 29702 43444
rect 265618 43432 265624 43444
rect 29696 43404 265624 43432
rect 29696 43392 29702 43404
rect 265618 43392 265624 43404
rect 265676 43392 265682 43444
rect 279418 43392 279424 43444
rect 279476 43432 279482 43444
rect 415394 43432 415400 43444
rect 279476 43404 415400 43432
rect 279476 43392 279482 43404
rect 415394 43392 415400 43404
rect 415452 43392 415458 43444
rect 62022 42032 62028 42084
rect 62080 42072 62086 42084
rect 264330 42072 264336 42084
rect 62080 42044 264336 42072
rect 62080 42032 62086 42044
rect 264330 42032 264336 42044
rect 264388 42032 264394 42084
rect 268378 42032 268384 42084
rect 268436 42072 268442 42084
rect 449986 42072 449992 42084
rect 268436 42044 449992 42072
rect 268436 42032 268442 42044
rect 449986 42032 449992 42044
rect 450044 42032 450050 42084
rect 115842 40740 115848 40792
rect 115900 40780 115906 40792
rect 249058 40780 249064 40792
rect 115900 40752 249064 40780
rect 115900 40740 115906 40752
rect 249058 40740 249064 40752
rect 249116 40740 249122 40792
rect 259362 40740 259368 40792
rect 259420 40780 259426 40792
rect 430574 40780 430580 40792
rect 259420 40752 430580 40780
rect 259420 40740 259426 40752
rect 430574 40740 430580 40752
rect 430632 40740 430638 40792
rect 38562 40672 38568 40724
rect 38620 40712 38626 40724
rect 269206 40712 269212 40724
rect 38620 40684 269212 40712
rect 38620 40672 38626 40684
rect 269206 40672 269212 40684
rect 269264 40672 269270 40724
rect 30282 39380 30288 39432
rect 30340 39420 30346 39432
rect 181530 39420 181536 39432
rect 30340 39392 181536 39420
rect 30340 39380 30346 39392
rect 181530 39380 181536 39392
rect 181588 39380 181594 39432
rect 13722 39312 13728 39364
rect 13780 39352 13786 39364
rect 244918 39352 244924 39364
rect 13780 39324 244924 39352
rect 13780 39312 13786 39324
rect 244918 39312 244924 39324
rect 244976 39312 244982 39364
rect 339402 38564 339408 38616
rect 339460 38604 339466 38616
rect 418798 38604 418804 38616
rect 339460 38576 418804 38604
rect 339460 38564 339466 38576
rect 418798 38564 418804 38576
rect 418856 38564 418862 38616
rect 333974 37884 333980 37936
rect 334032 37924 334038 37936
rect 338114 37924 338120 37936
rect 334032 37896 338120 37924
rect 334032 37884 334038 37896
rect 338114 37884 338120 37896
rect 338172 37924 338178 37936
rect 339402 37924 339408 37936
rect 338172 37896 339408 37924
rect 338172 37884 338178 37896
rect 339402 37884 339408 37896
rect 339460 37884 339466 37936
rect 209038 37204 209044 37256
rect 209096 37244 209102 37256
rect 258074 37244 258080 37256
rect 209096 37216 258080 37244
rect 209096 37204 209102 37216
rect 258074 37204 258080 37216
rect 258132 37244 258138 37256
rect 259362 37244 259368 37256
rect 258132 37216 259368 37244
rect 258132 37204 258138 37216
rect 259362 37204 259368 37216
rect 259420 37204 259426 37256
rect 122742 36592 122748 36644
rect 122800 36632 122806 36644
rect 206370 36632 206376 36644
rect 122800 36604 206376 36632
rect 122800 36592 122806 36604
rect 206370 36592 206376 36604
rect 206428 36592 206434 36644
rect 16482 36524 16488 36576
rect 16540 36564 16546 36576
rect 235350 36564 235356 36576
rect 16540 36536 235356 36564
rect 16540 36524 16546 36536
rect 235350 36524 235356 36536
rect 235408 36524 235414 36576
rect 276658 36524 276664 36576
rect 276716 36564 276722 36576
rect 414014 36564 414020 36576
rect 276716 36536 414020 36564
rect 276716 36524 276722 36536
rect 414014 36524 414020 36536
rect 414072 36524 414078 36576
rect 320818 35844 320824 35896
rect 320876 35884 320882 35896
rect 395430 35884 395436 35896
rect 320876 35856 395436 35884
rect 320876 35844 320882 35856
rect 395430 35844 395436 35856
rect 395488 35844 395494 35896
rect 130378 35232 130384 35284
rect 130436 35272 130442 35284
rect 213270 35272 213276 35284
rect 130436 35244 213276 35272
rect 130436 35232 130442 35244
rect 213270 35232 213276 35244
rect 213328 35232 213334 35284
rect 71038 35164 71044 35216
rect 71096 35204 71102 35216
rect 239490 35204 239496 35216
rect 71096 35176 239496 35204
rect 71096 35164 71102 35176
rect 239490 35164 239496 35176
rect 239548 35164 239554 35216
rect 320174 34484 320180 34536
rect 320232 34524 320238 34536
rect 320818 34524 320824 34536
rect 320232 34496 320824 34524
rect 320232 34484 320238 34496
rect 320818 34484 320824 34496
rect 320876 34484 320882 34536
rect 191190 33804 191196 33856
rect 191248 33844 191254 33856
rect 280890 33844 280896 33856
rect 191248 33816 280896 33844
rect 191248 33804 191254 33816
rect 280890 33804 280896 33816
rect 280948 33804 280954 33856
rect 70210 33736 70216 33788
rect 70268 33776 70274 33788
rect 218698 33776 218704 33788
rect 70268 33748 218704 33776
rect 70268 33736 70274 33748
rect 218698 33736 218704 33748
rect 218756 33736 218762 33788
rect 2866 33056 2872 33108
rect 2924 33096 2930 33108
rect 40678 33096 40684 33108
rect 2924 33068 40684 33096
rect 2924 33056 2930 33068
rect 40678 33056 40684 33068
rect 40736 33056 40742 33108
rect 85482 32444 85488 32496
rect 85540 32484 85546 32496
rect 246298 32484 246304 32496
rect 85540 32456 246304 32484
rect 85540 32444 85546 32456
rect 246298 32444 246304 32456
rect 246356 32444 246362 32496
rect 60642 32376 60648 32428
rect 60700 32416 60706 32428
rect 275278 32416 275284 32428
rect 60700 32388 275284 32416
rect 60700 32376 60706 32388
rect 275278 32376 275284 32388
rect 275336 32376 275342 32428
rect 275278 31764 275284 31816
rect 275336 31804 275342 31816
rect 276658 31804 276664 31816
rect 275336 31776 276664 31804
rect 275336 31764 275342 31776
rect 276658 31764 276664 31776
rect 276716 31764 276722 31816
rect 57238 31696 57244 31748
rect 57296 31736 57302 31748
rect 278774 31736 278780 31748
rect 57296 31708 278780 31736
rect 57296 31696 57302 31708
rect 278774 31696 278780 31708
rect 278832 31736 278838 31748
rect 279418 31736 279424 31748
rect 278832 31708 279424 31736
rect 278832 31696 278838 31708
rect 279418 31696 279424 31708
rect 279476 31696 279482 31748
rect 106 31016 112 31068
rect 164 31056 170 31068
rect 231302 31056 231308 31068
rect 164 31028 231308 31056
rect 164 31016 170 31028
rect 231302 31016 231308 31028
rect 231360 31016 231366 31068
rect 278038 31016 278044 31068
rect 278096 31056 278102 31068
rect 281534 31056 281540 31068
rect 278096 31028 281540 31056
rect 278096 31016 278102 31028
rect 281534 31016 281540 31028
rect 281592 31056 281598 31068
rect 388530 31056 388536 31068
rect 281592 31028 388536 31056
rect 281592 31016 281598 31028
rect 388530 31016 388536 31028
rect 388588 31016 388594 31068
rect 300854 30268 300860 30320
rect 300912 30308 300918 30320
rect 301314 30308 301320 30320
rect 300912 30280 301320 30308
rect 300912 30268 300918 30280
rect 301314 30268 301320 30280
rect 301372 30308 301378 30320
rect 432598 30308 432604 30320
rect 301372 30280 432604 30308
rect 301372 30268 301378 30280
rect 432598 30268 432604 30280
rect 432656 30268 432662 30320
rect 118602 29656 118608 29708
rect 118660 29696 118666 29708
rect 231210 29696 231216 29708
rect 118660 29668 231216 29696
rect 118660 29656 118666 29668
rect 231210 29656 231216 29668
rect 231268 29656 231274 29708
rect 56502 29588 56508 29640
rect 56560 29628 56566 29640
rect 260098 29628 260104 29640
rect 56560 29600 260104 29628
rect 56560 29588 56566 29600
rect 260098 29588 260104 29600
rect 260156 29588 260162 29640
rect 277394 29588 277400 29640
rect 277452 29628 277458 29640
rect 301314 29628 301320 29640
rect 277452 29600 301320 29628
rect 277452 29588 277458 29600
rect 301314 29588 301320 29600
rect 301372 29588 301378 29640
rect 99282 28296 99288 28348
rect 99340 28336 99346 28348
rect 229738 28336 229744 28348
rect 99340 28308 229744 28336
rect 99340 28296 99346 28308
rect 229738 28296 229744 28308
rect 229796 28296 229802 28348
rect 49602 28228 49608 28280
rect 49660 28268 49666 28280
rect 240778 28268 240784 28280
rect 49660 28240 240784 28268
rect 49660 28228 49666 28240
rect 240778 28228 240784 28240
rect 240836 28228 240842 28280
rect 271782 28228 271788 28280
rect 271840 28268 271846 28280
rect 392762 28268 392768 28280
rect 271840 28240 392768 28268
rect 271840 28228 271846 28240
rect 392762 28228 392768 28240
rect 392820 28228 392826 28280
rect 52362 27548 52368 27600
rect 52420 27588 52426 27600
rect 262214 27588 262220 27600
rect 52420 27560 262220 27588
rect 52420 27548 52426 27560
rect 262214 27548 262220 27560
rect 262272 27588 262278 27600
rect 262950 27588 262956 27600
rect 262272 27560 262956 27588
rect 262272 27548 262278 27560
rect 262950 27548 262956 27560
rect 263008 27548 263014 27600
rect 296714 27548 296720 27600
rect 296772 27588 296778 27600
rect 374638 27588 374644 27600
rect 296772 27560 374644 27588
rect 296772 27548 296778 27560
rect 374638 27548 374644 27560
rect 374696 27548 374702 27600
rect 344278 27480 344284 27532
rect 344336 27520 344342 27532
rect 405734 27520 405740 27532
rect 344336 27492 405740 27520
rect 344336 27480 344342 27492
rect 405734 27480 405740 27492
rect 405792 27480 405798 27532
rect 61930 26868 61936 26920
rect 61988 26908 61994 26920
rect 160738 26908 160744 26920
rect 61988 26880 160744 26908
rect 61988 26868 61994 26880
rect 160738 26868 160744 26880
rect 160796 26868 160802 26920
rect 263594 26868 263600 26920
rect 263652 26908 263658 26920
rect 296714 26908 296720 26920
rect 263652 26880 296720 26908
rect 263652 26868 263658 26880
rect 296714 26868 296720 26880
rect 296772 26868 296778 26920
rect 257338 25508 257344 25560
rect 257396 25548 257402 25560
rect 445938 25548 445944 25560
rect 257396 25520 445944 25548
rect 257396 25508 257402 25520
rect 445938 25508 445944 25520
rect 445996 25508 446002 25560
rect 55122 24760 55128 24812
rect 55180 24800 55186 24812
rect 307754 24800 307760 24812
rect 55180 24772 307760 24800
rect 55180 24760 55186 24772
rect 307754 24760 307760 24772
rect 307812 24800 307818 24812
rect 308398 24800 308404 24812
rect 307812 24772 308404 24800
rect 307812 24760 307818 24772
rect 308398 24760 308404 24772
rect 308456 24760 308462 24812
rect 92382 22788 92388 22840
rect 92440 22828 92446 22840
rect 209130 22828 209136 22840
rect 92440 22800 209136 22828
rect 92440 22788 92446 22800
rect 209130 22788 209136 22800
rect 209188 22788 209194 22840
rect 45462 22720 45468 22772
rect 45520 22760 45526 22772
rect 228358 22760 228364 22772
rect 45520 22732 228364 22760
rect 45520 22720 45526 22732
rect 228358 22720 228364 22732
rect 228416 22720 228422 22772
rect 250530 22720 250536 22772
rect 250588 22760 250594 22772
rect 389910 22760 389916 22772
rect 250588 22732 389916 22760
rect 250588 22720 250594 22732
rect 389910 22720 389916 22732
rect 389968 22720 389974 22772
rect 346394 21428 346400 21480
rect 346452 21468 346458 21480
rect 411438 21468 411444 21480
rect 346452 21440 411444 21468
rect 346452 21428 346458 21440
rect 411438 21428 411444 21440
rect 411496 21428 411502 21480
rect 95050 21360 95056 21412
rect 95108 21400 95114 21412
rect 264238 21400 264244 21412
rect 95108 21372 264244 21400
rect 95108 21360 95114 21372
rect 264238 21360 264244 21372
rect 264296 21360 264302 21412
rect 284938 21360 284944 21412
rect 284996 21400 285002 21412
rect 421558 21400 421564 21412
rect 284996 21372 421564 21400
rect 284996 21360 285002 21372
rect 421558 21360 421564 21372
rect 421616 21360 421622 21412
rect 224218 20612 224224 20664
rect 224276 20652 224282 20664
rect 270494 20652 270500 20664
rect 224276 20624 270500 20652
rect 224276 20612 224282 20624
rect 270494 20612 270500 20624
rect 270552 20652 270558 20664
rect 271782 20652 271788 20664
rect 270552 20624 271788 20652
rect 270552 20612 270558 20624
rect 271782 20612 271788 20624
rect 271840 20612 271846 20664
rect 316034 20612 316040 20664
rect 316092 20652 316098 20664
rect 316770 20652 316776 20664
rect 316092 20624 316776 20652
rect 316092 20612 316098 20624
rect 316770 20612 316776 20624
rect 316828 20652 316834 20664
rect 396718 20652 396724 20664
rect 316828 20624 396724 20652
rect 316828 20612 316834 20624
rect 396718 20612 396724 20624
rect 396776 20612 396782 20664
rect 305638 20544 305644 20596
rect 305696 20584 305702 20596
rect 336734 20584 336740 20596
rect 305696 20556 336740 20584
rect 305696 20544 305702 20556
rect 336734 20544 336740 20556
rect 336792 20584 336798 20596
rect 337470 20584 337476 20596
rect 336792 20556 337476 20584
rect 336792 20544 336798 20556
rect 337470 20544 337476 20556
rect 337528 20544 337534 20596
rect 88242 20000 88248 20052
rect 88300 20040 88306 20052
rect 216122 20040 216128 20052
rect 88300 20012 216128 20040
rect 88300 20000 88306 20012
rect 216122 20000 216128 20012
rect 216180 20000 216186 20052
rect 31662 19932 31668 19984
rect 31720 19972 31726 19984
rect 224310 19972 224316 19984
rect 31720 19944 224316 19972
rect 31720 19932 31726 19944
rect 224310 19932 224316 19944
rect 224368 19932 224374 19984
rect 341518 19320 341524 19372
rect 341576 19360 341582 19372
rect 346394 19360 346400 19372
rect 341576 19332 346400 19360
rect 341576 19320 341582 19332
rect 346394 19320 346400 19332
rect 346452 19320 346458 19372
rect 280798 19252 280804 19304
rect 280856 19292 280862 19304
rect 284938 19292 284944 19304
rect 280856 19264 284944 19292
rect 280856 19252 280862 19264
rect 284938 19252 284944 19264
rect 284996 19252 285002 19304
rect 124122 18640 124128 18692
rect 124180 18680 124186 18692
rect 210418 18680 210424 18692
rect 124180 18652 210424 18680
rect 124180 18640 124186 18652
rect 210418 18640 210424 18652
rect 210476 18640 210482 18692
rect 284938 18640 284944 18692
rect 284996 18680 285002 18692
rect 370498 18680 370504 18692
rect 284996 18652 370504 18680
rect 284996 18640 285002 18652
rect 370498 18640 370504 18652
rect 370556 18640 370562 18692
rect 45370 18572 45376 18624
rect 45428 18612 45434 18624
rect 198090 18612 198096 18624
rect 45428 18584 198096 18612
rect 45428 18572 45434 18584
rect 198090 18572 198096 18584
rect 198148 18572 198154 18624
rect 202138 18572 202144 18624
rect 202196 18612 202202 18624
rect 288434 18612 288440 18624
rect 202196 18584 288440 18612
rect 202196 18572 202202 18584
rect 288434 18572 288440 18584
rect 288492 18572 288498 18624
rect 280890 17892 280896 17944
rect 280948 17932 280954 17944
rect 363598 17932 363604 17944
rect 280948 17904 363604 17932
rect 280948 17892 280954 17904
rect 363598 17892 363604 17904
rect 363656 17892 363662 17944
rect 280154 17280 280160 17332
rect 280212 17320 280218 17332
rect 280890 17320 280896 17332
rect 280212 17292 280896 17320
rect 280212 17280 280218 17292
rect 280890 17280 280896 17292
rect 280948 17280 280954 17332
rect 53650 17212 53656 17264
rect 53708 17252 53714 17264
rect 242158 17252 242164 17264
rect 53708 17224 242164 17252
rect 53708 17212 53714 17224
rect 242158 17212 242164 17224
rect 242216 17212 242222 17264
rect 249150 16532 249156 16584
rect 249208 16572 249214 16584
rect 249702 16572 249708 16584
rect 249208 16544 249708 16572
rect 249208 16532 249214 16544
rect 249702 16532 249708 16544
rect 249760 16572 249766 16584
rect 367830 16572 367836 16584
rect 249760 16544 367836 16572
rect 249760 16532 249766 16544
rect 367830 16532 367836 16544
rect 367888 16532 367894 16584
rect 39574 15920 39580 15972
rect 39632 15960 39638 15972
rect 220170 15960 220176 15972
rect 39632 15932 220176 15960
rect 39632 15920 39638 15932
rect 220170 15920 220176 15932
rect 220228 15920 220234 15972
rect 9582 15852 9588 15904
rect 9640 15892 9646 15904
rect 231118 15892 231124 15904
rect 9640 15864 231124 15892
rect 9640 15852 9646 15864
rect 231118 15852 231124 15864
rect 231176 15852 231182 15904
rect 343358 15852 343364 15904
rect 343416 15892 343422 15904
rect 403618 15892 403624 15904
rect 343416 15864 403624 15892
rect 343416 15852 343422 15864
rect 403618 15852 403624 15864
rect 403676 15852 403682 15904
rect 255958 15104 255964 15156
rect 256016 15144 256022 15156
rect 256602 15144 256608 15156
rect 256016 15116 256608 15144
rect 256016 15104 256022 15116
rect 256602 15104 256608 15116
rect 256660 15144 256666 15156
rect 310514 15144 310520 15156
rect 256660 15116 310520 15144
rect 256660 15104 256666 15116
rect 310514 15104 310520 15116
rect 310572 15104 310578 15156
rect 311434 14492 311440 14544
rect 311492 14532 311498 14544
rect 360838 14532 360844 14544
rect 311492 14504 360844 14532
rect 311492 14492 311498 14504
rect 360838 14492 360844 14504
rect 360896 14492 360902 14544
rect 100662 14424 100668 14476
rect 100720 14464 100726 14476
rect 258718 14464 258724 14476
rect 100720 14436 258724 14464
rect 100720 14424 100726 14436
rect 258718 14424 258724 14436
rect 258776 14424 258782 14476
rect 328730 14424 328736 14476
rect 328788 14464 328794 14476
rect 382918 14464 382924 14476
rect 328788 14436 382924 14464
rect 328788 14424 328794 14436
rect 382918 14424 382924 14436
rect 382976 14424 382982 14476
rect 295334 13744 295340 13796
rect 295392 13784 295398 13796
rect 295886 13784 295892 13796
rect 295392 13756 295892 13784
rect 295392 13744 295398 13756
rect 295886 13744 295892 13756
rect 295944 13784 295950 13796
rect 400306 13784 400312 13796
rect 295944 13756 400312 13784
rect 295944 13744 295950 13756
rect 400306 13744 400312 13756
rect 400364 13744 400370 13796
rect 96246 13132 96252 13184
rect 96304 13172 96310 13184
rect 235258 13172 235264 13184
rect 96304 13144 235264 13172
rect 96304 13132 96310 13144
rect 235258 13132 235264 13144
rect 235316 13132 235322 13184
rect 54938 13064 54944 13116
rect 54996 13104 55002 13116
rect 238110 13104 238116 13116
rect 54996 13076 238116 13104
rect 54996 13064 55002 13076
rect 238110 13064 238116 13076
rect 238168 13064 238174 13116
rect 299658 13064 299664 13116
rect 299716 13104 299722 13116
rect 454034 13104 454040 13116
rect 299716 13076 454040 13104
rect 299716 13064 299722 13076
rect 454034 13064 454040 13076
rect 454092 13064 454098 13116
rect 264974 12452 264980 12504
rect 265032 12492 265038 12504
rect 295334 12492 295340 12504
rect 265032 12464 295340 12492
rect 265032 12452 265038 12464
rect 295334 12452 295340 12464
rect 295392 12452 295398 12504
rect 251818 12384 251824 12436
rect 251876 12424 251882 12436
rect 251876 12396 258074 12424
rect 251876 12384 251882 12396
rect 258046 12356 258074 12396
rect 276106 12384 276112 12436
rect 276164 12424 276170 12436
rect 277486 12424 277492 12436
rect 276164 12396 277492 12424
rect 276164 12384 276170 12396
rect 277486 12384 277492 12396
rect 277544 12424 277550 12436
rect 442994 12424 443000 12436
rect 277544 12396 443000 12424
rect 277544 12384 277550 12396
rect 442994 12384 443000 12396
rect 443052 12384 443058 12436
rect 385770 12356 385776 12368
rect 258046 12328 385776 12356
rect 385770 12316 385776 12328
rect 385828 12316 385834 12368
rect 251174 11908 251180 11960
rect 251232 11948 251238 11960
rect 251818 11948 251824 11960
rect 251232 11920 251824 11948
rect 251232 11908 251238 11920
rect 251818 11908 251824 11920
rect 251876 11908 251882 11960
rect 126882 11772 126888 11824
rect 126940 11812 126946 11824
rect 217318 11812 217324 11824
rect 126940 11784 217324 11812
rect 126940 11772 126946 11784
rect 217318 11772 217324 11784
rect 217376 11772 217382 11824
rect 12158 11704 12164 11756
rect 12216 11744 12222 11756
rect 233970 11744 233976 11756
rect 12216 11716 233976 11744
rect 12216 11704 12222 11716
rect 233970 11704 233976 11716
rect 234028 11704 234034 11756
rect 242894 11704 242900 11756
rect 242952 11744 242958 11756
rect 244090 11744 244096 11756
rect 242952 11716 244096 11744
rect 242952 11704 242958 11716
rect 244090 11704 244096 11716
rect 244148 11704 244154 11756
rect 135254 11636 135260 11688
rect 135312 11676 135318 11688
rect 136450 11676 136456 11688
rect 135312 11648 136456 11676
rect 135312 11636 135318 11648
rect 136450 11636 136456 11648
rect 136508 11636 136514 11688
rect 288434 10956 288440 11008
rect 288492 10996 288498 11008
rect 288986 10996 288992 11008
rect 288492 10968 288992 10996
rect 288492 10956 288498 10968
rect 288986 10956 288992 10968
rect 289044 10996 289050 11008
rect 377490 10996 377496 11008
rect 289044 10968 377496 10996
rect 289044 10956 289050 10968
rect 377490 10956 377496 10968
rect 377548 10956 377554 11008
rect 81342 10344 81348 10396
rect 81400 10384 81406 10396
rect 213178 10384 213184 10396
rect 81400 10356 213184 10384
rect 81400 10344 81406 10356
rect 213178 10344 213184 10356
rect 213236 10344 213242 10396
rect 24762 10276 24768 10328
rect 24820 10316 24826 10328
rect 222930 10316 222936 10328
rect 24820 10288 222936 10316
rect 24820 10276 24826 10288
rect 222930 10276 222936 10288
rect 222988 10276 222994 10328
rect 261754 9596 261760 9648
rect 261812 9636 261818 9648
rect 447134 9636 447140 9648
rect 261812 9608 447140 9636
rect 261812 9596 261818 9608
rect 447134 9596 447140 9608
rect 447192 9596 447198 9648
rect 85666 8984 85672 9036
rect 85724 9024 85730 9036
rect 220078 9024 220084 9036
rect 85724 8996 220084 9024
rect 85724 8984 85730 8996
rect 220078 8984 220084 8996
rect 220136 8984 220142 9036
rect 59630 8916 59636 8968
rect 59688 8956 59694 8968
rect 250438 8956 250444 8968
rect 59688 8928 250444 8956
rect 59688 8916 59694 8928
rect 250438 8916 250444 8928
rect 250496 8916 250502 8968
rect 345658 8236 345664 8288
rect 345716 8276 345722 8288
rect 394142 8276 394148 8288
rect 345716 8248 394148 8276
rect 345716 8236 345722 8248
rect 394142 8236 394148 8248
rect 394200 8236 394206 8288
rect 114002 7624 114008 7676
rect 114060 7664 114066 7676
rect 214558 7664 214564 7676
rect 114060 7636 214564 7664
rect 114060 7624 114066 7636
rect 214558 7624 214564 7636
rect 214616 7624 214622 7676
rect 66714 7556 66720 7608
rect 66772 7596 66778 7608
rect 261478 7596 261484 7608
rect 66772 7568 261484 7596
rect 66772 7556 66778 7568
rect 261478 7556 261484 7568
rect 261536 7556 261542 7608
rect 342162 7556 342168 7608
rect 342220 7596 342226 7608
rect 356698 7596 356704 7608
rect 342220 7568 356704 7596
rect 342220 7556 342226 7568
rect 356698 7556 356704 7568
rect 356756 7556 356762 7608
rect 325050 6808 325056 6860
rect 325108 6848 325114 6860
rect 409874 6848 409880 6860
rect 325108 6820 409880 6848
rect 325108 6808 325114 6820
rect 409874 6808 409880 6820
rect 409932 6808 409938 6860
rect 318058 6740 318064 6792
rect 318116 6780 318122 6792
rect 319438 6780 319444 6792
rect 318116 6752 319444 6780
rect 318116 6740 318122 6752
rect 319438 6740 319444 6752
rect 319496 6740 319502 6792
rect 121086 6196 121092 6248
rect 121144 6236 121150 6248
rect 239398 6236 239404 6248
rect 121144 6208 239404 6236
rect 121144 6196 121150 6208
rect 239398 6196 239404 6208
rect 239456 6196 239462 6248
rect 58434 6128 58440 6180
rect 58492 6168 58498 6180
rect 215938 6168 215944 6180
rect 58492 6140 215944 6168
rect 58492 6128 58498 6140
rect 215938 6128 215944 6140
rect 215996 6128 216002 6180
rect 298462 6128 298468 6180
rect 298520 6168 298526 6180
rect 378870 6168 378876 6180
rect 298520 6140 378876 6168
rect 298520 6128 298526 6140
rect 378870 6128 378876 6140
rect 378928 6128 378934 6180
rect 324406 5516 324412 5568
rect 324464 5556 324470 5568
rect 325050 5556 325056 5568
rect 324464 5528 325056 5556
rect 324464 5516 324470 5528
rect 325050 5516 325056 5528
rect 325108 5516 325114 5568
rect 316678 5448 316684 5500
rect 316736 5488 316742 5500
rect 317322 5488 317328 5500
rect 316736 5460 317328 5488
rect 316736 5448 316742 5460
rect 317322 5448 317328 5460
rect 317380 5488 317386 5500
rect 425882 5488 425888 5500
rect 317380 5460 425888 5488
rect 317380 5448 317386 5460
rect 425882 5448 425888 5460
rect 425940 5448 425946 5500
rect 109310 4768 109316 4820
rect 109368 4808 109374 4820
rect 238018 4808 238024 4820
rect 109368 4780 238024 4808
rect 109368 4768 109374 4780
rect 238018 4768 238024 4780
rect 238076 4768 238082 4820
rect 246206 4768 246212 4820
rect 246264 4808 246270 4820
rect 407114 4808 407120 4820
rect 246264 4780 407120 4808
rect 246264 4768 246270 4780
rect 407114 4768 407120 4780
rect 407172 4768 407178 4820
rect 232498 4156 232504 4208
rect 232556 4196 232562 4208
rect 235810 4196 235816 4208
rect 232556 4168 235816 4196
rect 232556 4156 232562 4168
rect 235810 4156 235816 4168
rect 235868 4156 235874 4208
rect 278682 4156 278688 4208
rect 278740 4196 278746 4208
rect 283098 4196 283104 4208
rect 278740 4168 283104 4196
rect 278740 4156 278746 4168
rect 283098 4156 283104 4168
rect 283156 4156 283162 4208
rect 191098 4088 191104 4140
rect 191156 4128 191162 4140
rect 247586 4128 247592 4140
rect 191156 4100 247592 4128
rect 191156 4088 191162 4100
rect 247586 4088 247592 4100
rect 247644 4088 247650 4140
rect 254670 4088 254676 4140
rect 254728 4128 254734 4140
rect 258074 4128 258080 4140
rect 254728 4100 258080 4128
rect 254728 4088 254734 4100
rect 258074 4088 258080 4100
rect 258132 4088 258138 4140
rect 291838 4088 291844 4140
rect 291896 4128 291902 4140
rect 301498 4128 301504 4140
rect 291896 4100 301504 4128
rect 291896 4088 291902 4100
rect 301498 4088 301504 4100
rect 301556 4088 301562 4140
rect 307110 4088 307116 4140
rect 307168 4128 307174 4140
rect 307938 4128 307944 4140
rect 307168 4100 307944 4128
rect 307168 4088 307174 4100
rect 307938 4088 307944 4100
rect 307996 4128 308002 4140
rect 309870 4128 309876 4140
rect 307996 4100 309876 4128
rect 307996 4088 308002 4100
rect 309870 4088 309876 4100
rect 309928 4088 309934 4140
rect 342898 4128 342904 4140
rect 316006 4100 342904 4128
rect 289078 4020 289084 4072
rect 289136 4060 289142 4072
rect 292574 4060 292580 4072
rect 289136 4032 292580 4060
rect 289136 4020 289142 4032
rect 292574 4020 292580 4032
rect 292632 4020 292638 4072
rect 306742 4020 306748 4072
rect 306800 4060 306806 4072
rect 316006 4060 316034 4100
rect 342898 4088 342904 4100
rect 342956 4088 342962 4140
rect 348418 4088 348424 4140
rect 348476 4128 348482 4140
rect 429838 4128 429844 4140
rect 348476 4100 429844 4128
rect 348476 4088 348482 4100
rect 429838 4088 429844 4100
rect 429896 4088 429902 4140
rect 306800 4032 316034 4060
rect 306800 4020 306806 4032
rect 332686 4020 332692 4072
rect 332744 4060 332750 4072
rect 335998 4060 336004 4072
rect 332744 4032 336004 4060
rect 332744 4020 332750 4032
rect 335998 4020 336004 4032
rect 336056 4020 336062 4072
rect 312630 3952 312636 4004
rect 312688 3992 312694 4004
rect 318150 3992 318156 4004
rect 312688 3964 318156 3992
rect 312688 3952 312694 3964
rect 318150 3952 318156 3964
rect 318208 3952 318214 4004
rect 291378 3680 291384 3732
rect 291436 3720 291442 3732
rect 291838 3720 291844 3732
rect 291436 3692 291844 3720
rect 291436 3680 291442 3692
rect 291838 3680 291844 3692
rect 291896 3680 291902 3732
rect 71038 3652 71044 3664
rect 65444 3624 71044 3652
rect 11146 3544 11152 3596
rect 11204 3584 11210 3596
rect 12250 3584 12256 3596
rect 11204 3556 12256 3584
rect 11204 3544 11210 3556
rect 12250 3544 12256 3556
rect 12308 3544 12314 3596
rect 27706 3544 27712 3596
rect 27764 3584 27770 3596
rect 28902 3584 28908 3596
rect 27764 3556 28908 3584
rect 27764 3544 27770 3556
rect 28902 3544 28908 3556
rect 28960 3544 28966 3596
rect 44266 3544 44272 3596
rect 44324 3584 44330 3596
rect 45370 3584 45376 3596
rect 44324 3556 45376 3584
rect 44324 3544 44330 3556
rect 45370 3544 45376 3556
rect 45428 3544 45434 3596
rect 64322 3544 64328 3596
rect 64380 3584 64386 3596
rect 64782 3584 64788 3596
rect 64380 3556 64788 3584
rect 64380 3544 64386 3556
rect 64782 3544 64788 3556
rect 64840 3544 64846 3596
rect 8754 3476 8760 3528
rect 8812 3516 8818 3528
rect 9582 3516 9588 3528
rect 8812 3488 9588 3516
rect 8812 3476 8818 3488
rect 9582 3476 9588 3488
rect 9640 3476 9646 3528
rect 9950 3476 9956 3528
rect 10008 3516 10014 3528
rect 10962 3516 10968 3528
rect 10008 3488 10968 3516
rect 10008 3476 10014 3488
rect 10962 3476 10968 3488
rect 11020 3476 11026 3528
rect 15930 3476 15936 3528
rect 15988 3516 15994 3528
rect 16482 3516 16488 3528
rect 15988 3488 16488 3516
rect 15988 3476 15994 3488
rect 16482 3476 16488 3488
rect 16540 3476 16546 3528
rect 17034 3476 17040 3528
rect 17092 3516 17098 3528
rect 17862 3516 17868 3528
rect 17092 3488 17868 3516
rect 17092 3476 17098 3488
rect 17862 3476 17868 3488
rect 17920 3476 17926 3528
rect 18230 3476 18236 3528
rect 18288 3516 18294 3528
rect 19242 3516 19248 3528
rect 18288 3488 19248 3516
rect 18288 3476 18294 3488
rect 19242 3476 19248 3488
rect 19300 3476 19306 3528
rect 24210 3476 24216 3528
rect 24268 3516 24274 3528
rect 24762 3516 24768 3528
rect 24268 3488 24768 3516
rect 24268 3476 24274 3488
rect 24762 3476 24768 3488
rect 24820 3476 24826 3528
rect 36538 3516 36544 3528
rect 26206 3488 36544 3516
rect 20530 3408 20536 3460
rect 20588 3448 20594 3460
rect 26206 3448 26234 3488
rect 36538 3476 36544 3488
rect 36596 3476 36602 3528
rect 40678 3476 40684 3528
rect 40736 3516 40742 3528
rect 41322 3516 41328 3528
rect 40736 3488 41328 3516
rect 40736 3476 40742 3488
rect 41322 3476 41328 3488
rect 41380 3476 41386 3528
rect 41874 3476 41880 3528
rect 41932 3516 41938 3528
rect 42702 3516 42708 3528
rect 41932 3488 42708 3516
rect 41932 3476 41938 3488
rect 42702 3476 42708 3488
rect 42760 3476 42766 3528
rect 43070 3476 43076 3528
rect 43128 3516 43134 3528
rect 44082 3516 44088 3528
rect 43128 3488 44088 3516
rect 43128 3476 43134 3488
rect 44082 3476 44088 3488
rect 44140 3476 44146 3528
rect 48958 3476 48964 3528
rect 49016 3516 49022 3528
rect 49602 3516 49608 3528
rect 49016 3488 49608 3516
rect 49016 3476 49022 3488
rect 49602 3476 49608 3488
rect 49660 3476 49666 3528
rect 50154 3476 50160 3528
rect 50212 3516 50218 3528
rect 50982 3516 50988 3528
rect 50212 3488 50988 3516
rect 50212 3476 50218 3488
rect 50982 3476 50988 3488
rect 51040 3476 51046 3528
rect 52546 3476 52552 3528
rect 52604 3516 52610 3528
rect 53650 3516 53656 3528
rect 52604 3488 53656 3516
rect 52604 3476 52610 3488
rect 53650 3476 53656 3488
rect 53708 3476 53714 3528
rect 56042 3476 56048 3528
rect 56100 3516 56106 3528
rect 56502 3516 56508 3528
rect 56100 3488 56508 3516
rect 56100 3476 56106 3488
rect 56502 3476 56508 3488
rect 56560 3476 56566 3528
rect 57238 3476 57244 3528
rect 57296 3516 57302 3528
rect 57882 3516 57888 3528
rect 57296 3488 57888 3516
rect 57296 3476 57302 3488
rect 57882 3476 57888 3488
rect 57940 3476 57946 3528
rect 63218 3476 63224 3528
rect 63276 3516 63282 3528
rect 65444 3516 65472 3624
rect 71038 3612 71044 3624
rect 71096 3612 71102 3664
rect 351178 3612 351184 3664
rect 351236 3652 351242 3664
rect 351638 3652 351644 3664
rect 351236 3624 351644 3652
rect 351236 3612 351242 3624
rect 351638 3612 351644 3624
rect 351696 3612 351702 3664
rect 69106 3544 69112 3596
rect 69164 3584 69170 3596
rect 70210 3584 70216 3596
rect 69164 3556 70216 3584
rect 69164 3544 69170 3556
rect 70210 3544 70216 3556
rect 70268 3544 70274 3596
rect 119890 3544 119896 3596
rect 119948 3584 119954 3596
rect 122098 3584 122104 3596
rect 119948 3556 122104 3584
rect 119948 3544 119954 3556
rect 122098 3544 122104 3556
rect 122156 3544 122162 3596
rect 276014 3544 276020 3596
rect 276072 3584 276078 3596
rect 277118 3584 277124 3596
rect 276072 3556 277124 3584
rect 276072 3544 276078 3556
rect 277118 3544 277124 3556
rect 277176 3544 277182 3596
rect 63276 3488 65472 3516
rect 63276 3476 63282 3488
rect 65518 3476 65524 3528
rect 65576 3516 65582 3528
rect 66162 3516 66168 3528
rect 65576 3488 66168 3516
rect 65576 3476 65582 3488
rect 66162 3476 66168 3488
rect 66220 3476 66226 3528
rect 67910 3476 67916 3528
rect 67968 3516 67974 3528
rect 68922 3516 68928 3528
rect 67968 3488 68928 3516
rect 67968 3476 67974 3488
rect 68922 3476 68928 3488
rect 68980 3476 68986 3528
rect 72602 3476 72608 3528
rect 72660 3516 72666 3528
rect 73062 3516 73068 3528
rect 72660 3488 73068 3516
rect 72660 3476 72666 3488
rect 73062 3476 73068 3488
rect 73120 3476 73126 3528
rect 73798 3476 73804 3528
rect 73856 3516 73862 3528
rect 74442 3516 74448 3528
rect 73856 3488 74448 3516
rect 73856 3476 73862 3488
rect 74442 3476 74448 3488
rect 74500 3476 74506 3528
rect 74994 3476 75000 3528
rect 75052 3516 75058 3528
rect 75822 3516 75828 3528
rect 75052 3488 75828 3516
rect 75052 3476 75058 3488
rect 75822 3476 75828 3488
rect 75880 3476 75886 3528
rect 76190 3476 76196 3528
rect 76248 3516 76254 3528
rect 77202 3516 77208 3528
rect 76248 3488 77208 3516
rect 76248 3476 76254 3488
rect 77202 3476 77208 3488
rect 77260 3476 77266 3528
rect 80882 3476 80888 3528
rect 80940 3516 80946 3528
rect 81342 3516 81348 3528
rect 80940 3488 81348 3516
rect 80940 3476 80946 3488
rect 81342 3476 81348 3488
rect 81400 3476 81406 3528
rect 90358 3476 90364 3528
rect 90416 3516 90422 3528
rect 91002 3516 91008 3528
rect 90416 3488 91008 3516
rect 90416 3476 90422 3488
rect 91002 3476 91008 3488
rect 91060 3476 91066 3528
rect 91554 3476 91560 3528
rect 91612 3516 91618 3528
rect 92382 3516 92388 3528
rect 91612 3488 92388 3516
rect 91612 3476 91618 3488
rect 92382 3476 92388 3488
rect 92440 3476 92446 3528
rect 92750 3476 92756 3528
rect 92808 3516 92814 3528
rect 93762 3516 93768 3528
rect 92808 3488 93768 3516
rect 92808 3476 92814 3488
rect 93762 3476 93768 3488
rect 93820 3476 93826 3528
rect 93946 3476 93952 3528
rect 94004 3516 94010 3528
rect 95050 3516 95056 3528
rect 94004 3488 95056 3516
rect 94004 3476 94010 3488
rect 95050 3476 95056 3488
rect 95108 3476 95114 3528
rect 97442 3476 97448 3528
rect 97500 3516 97506 3528
rect 97902 3516 97908 3528
rect 97500 3488 97908 3516
rect 97500 3476 97506 3488
rect 97902 3476 97908 3488
rect 97960 3476 97966 3528
rect 98638 3476 98644 3528
rect 98696 3516 98702 3528
rect 99282 3516 99288 3528
rect 98696 3488 99288 3516
rect 98696 3476 98702 3488
rect 99282 3476 99288 3488
rect 99340 3476 99346 3528
rect 99834 3476 99840 3528
rect 99892 3516 99898 3528
rect 100662 3516 100668 3528
rect 99892 3488 100668 3516
rect 99892 3476 99898 3488
rect 100662 3476 100668 3488
rect 100720 3476 100726 3528
rect 101030 3476 101036 3528
rect 101088 3516 101094 3528
rect 102042 3516 102048 3528
rect 101088 3488 102048 3516
rect 101088 3476 101094 3488
rect 102042 3476 102048 3488
rect 102100 3476 102106 3528
rect 105722 3476 105728 3528
rect 105780 3516 105786 3528
rect 106182 3516 106188 3528
rect 105780 3488 106188 3516
rect 105780 3476 105786 3488
rect 106182 3476 106188 3488
rect 106240 3476 106246 3528
rect 106918 3476 106924 3528
rect 106976 3516 106982 3528
rect 107562 3516 107568 3528
rect 106976 3488 107568 3516
rect 106976 3476 106982 3488
rect 107562 3476 107568 3488
rect 107620 3476 107626 3528
rect 108114 3476 108120 3528
rect 108172 3516 108178 3528
rect 108942 3516 108948 3528
rect 108172 3488 108948 3516
rect 108172 3476 108178 3488
rect 108942 3476 108948 3488
rect 109000 3476 109006 3528
rect 110506 3476 110512 3528
rect 110564 3516 110570 3528
rect 111702 3516 111708 3528
rect 110564 3488 111708 3516
rect 110564 3476 110570 3488
rect 111702 3476 111708 3488
rect 111760 3476 111766 3528
rect 115198 3476 115204 3528
rect 115256 3516 115262 3528
rect 115842 3516 115848 3528
rect 115256 3488 115848 3516
rect 115256 3476 115262 3488
rect 115842 3476 115848 3488
rect 115900 3476 115906 3528
rect 116394 3476 116400 3528
rect 116452 3516 116458 3528
rect 117222 3516 117228 3528
rect 116452 3488 117228 3516
rect 116452 3476 116458 3488
rect 117222 3476 117228 3488
rect 117280 3476 117286 3528
rect 117590 3476 117596 3528
rect 117648 3516 117654 3528
rect 118602 3516 118608 3528
rect 117648 3488 118608 3516
rect 117648 3476 117654 3488
rect 118602 3476 118608 3488
rect 118660 3476 118666 3528
rect 118786 3476 118792 3528
rect 118844 3516 118850 3528
rect 119982 3516 119988 3528
rect 118844 3488 119988 3516
rect 118844 3476 118850 3488
rect 119982 3476 119988 3488
rect 120040 3476 120046 3528
rect 122282 3476 122288 3528
rect 122340 3516 122346 3528
rect 122742 3516 122748 3528
rect 122340 3488 122748 3516
rect 122340 3476 122346 3488
rect 122742 3476 122748 3488
rect 122800 3476 122806 3528
rect 123478 3476 123484 3528
rect 123536 3516 123542 3528
rect 124122 3516 124128 3528
rect 123536 3488 124128 3516
rect 123536 3476 123542 3488
rect 124122 3476 124128 3488
rect 124180 3476 124186 3528
rect 124674 3476 124680 3528
rect 124732 3516 124738 3528
rect 125502 3516 125508 3528
rect 124732 3488 125508 3516
rect 124732 3476 124738 3488
rect 125502 3476 125508 3488
rect 125560 3476 125566 3528
rect 125870 3476 125876 3528
rect 125928 3516 125934 3528
rect 126882 3516 126888 3528
rect 125928 3488 126888 3516
rect 125928 3476 125934 3488
rect 126882 3476 126888 3488
rect 126940 3476 126946 3528
rect 140038 3476 140044 3528
rect 140096 3516 140102 3528
rect 141418 3516 141424 3528
rect 140096 3488 141424 3516
rect 140096 3476 140102 3488
rect 141418 3476 141424 3488
rect 141476 3476 141482 3528
rect 143534 3476 143540 3528
rect 143592 3516 143598 3528
rect 144822 3516 144828 3528
rect 143592 3488 144828 3516
rect 143592 3476 143598 3488
rect 144822 3476 144828 3488
rect 144880 3476 144886 3528
rect 240502 3476 240508 3528
rect 240560 3516 240566 3528
rect 246390 3516 246396 3528
rect 240560 3488 246396 3516
rect 240560 3476 240566 3488
rect 246390 3476 246396 3488
rect 246448 3476 246454 3528
rect 248782 3476 248788 3528
rect 248840 3516 248846 3528
rect 249702 3516 249708 3528
rect 248840 3488 249708 3516
rect 248840 3476 248846 3488
rect 249702 3476 249708 3488
rect 249760 3476 249766 3528
rect 252370 3476 252376 3528
rect 252428 3516 252434 3528
rect 253198 3516 253204 3528
rect 252428 3488 253204 3516
rect 252428 3476 252434 3488
rect 253198 3476 253204 3488
rect 253256 3476 253262 3528
rect 266354 3476 266360 3528
rect 266412 3516 266418 3528
rect 266538 3516 266544 3528
rect 266412 3488 266544 3516
rect 266412 3476 266418 3488
rect 266538 3476 266544 3488
rect 266596 3516 266602 3528
rect 271138 3516 271144 3528
rect 266596 3488 271144 3516
rect 266596 3476 266602 3488
rect 271138 3476 271144 3488
rect 271196 3476 271202 3528
rect 274818 3476 274824 3528
rect 274876 3516 274882 3528
rect 275278 3516 275284 3528
rect 274876 3488 275284 3516
rect 274876 3476 274882 3488
rect 275278 3476 275284 3488
rect 275336 3476 275342 3528
rect 284294 3476 284300 3528
rect 284352 3516 284358 3528
rect 285030 3516 285036 3528
rect 284352 3488 285036 3516
rect 284352 3476 284358 3488
rect 285030 3476 285036 3488
rect 285088 3476 285094 3528
rect 303522 3476 303528 3528
rect 303580 3516 303586 3528
rect 305546 3516 305552 3528
rect 303580 3488 305552 3516
rect 303580 3476 303586 3488
rect 305546 3476 305552 3488
rect 305604 3476 305610 3528
rect 332594 3476 332600 3528
rect 332652 3516 332658 3528
rect 333882 3516 333888 3528
rect 332652 3488 333888 3516
rect 332652 3476 332658 3488
rect 333882 3476 333888 3488
rect 333940 3476 333946 3528
rect 582190 3476 582196 3528
rect 582248 3516 582254 3528
rect 583202 3516 583208 3528
rect 582248 3488 583208 3516
rect 582248 3476 582254 3488
rect 583202 3476 583208 3488
rect 583260 3476 583266 3528
rect 20588 3420 26234 3448
rect 20588 3408 20594 3420
rect 26510 3408 26516 3460
rect 26568 3448 26574 3460
rect 27522 3448 27528 3460
rect 26568 3420 27528 3448
rect 26568 3408 26574 3420
rect 27522 3408 27528 3420
rect 27580 3408 27586 3460
rect 28902 3408 28908 3460
rect 28960 3448 28966 3460
rect 29638 3448 29644 3460
rect 28960 3420 29644 3448
rect 28960 3408 28966 3420
rect 29638 3408 29644 3420
rect 29696 3408 29702 3460
rect 32398 3408 32404 3460
rect 32456 3448 32462 3460
rect 33042 3448 33048 3460
rect 32456 3420 33048 3448
rect 32456 3408 32462 3420
rect 33042 3408 33048 3420
rect 33100 3408 33106 3460
rect 33594 3408 33600 3460
rect 33652 3448 33658 3460
rect 34422 3448 34428 3460
rect 33652 3420 34428 3448
rect 33652 3408 33658 3420
rect 34422 3408 34428 3420
rect 34480 3408 34486 3460
rect 34790 3408 34796 3460
rect 34848 3448 34854 3460
rect 35802 3448 35808 3460
rect 34848 3420 35808 3448
rect 34848 3408 34854 3420
rect 35802 3408 35808 3420
rect 35860 3408 35866 3460
rect 37090 3408 37096 3460
rect 37148 3448 37154 3460
rect 87598 3448 87604 3460
rect 37148 3420 87604 3448
rect 37148 3408 37154 3420
rect 87598 3408 87604 3420
rect 87656 3408 87662 3460
rect 102226 3408 102232 3460
rect 102284 3448 102290 3460
rect 130378 3448 130384 3460
rect 102284 3420 130384 3448
rect 102284 3408 102290 3420
rect 130378 3408 130384 3420
rect 130436 3408 130442 3460
rect 267734 3408 267740 3460
rect 267792 3448 267798 3460
rect 268838 3448 268844 3460
rect 267792 3420 268844 3448
rect 267792 3408 267798 3420
rect 268838 3408 268844 3420
rect 268896 3408 268902 3460
rect 349246 3408 349252 3460
rect 349304 3448 349310 3460
rect 357434 3448 357440 3460
rect 349304 3420 357440 3448
rect 349304 3408 349310 3420
rect 357434 3408 357440 3420
rect 357492 3408 357498 3460
rect 35986 3272 35992 3324
rect 36044 3312 36050 3324
rect 37182 3312 37188 3324
rect 36044 3284 37188 3312
rect 36044 3272 36050 3284
rect 37182 3272 37188 3284
rect 37240 3272 37246 3324
rect 89162 3272 89168 3324
rect 89220 3312 89226 3324
rect 89622 3312 89628 3324
rect 89220 3284 89628 3312
rect 89220 3272 89226 3284
rect 89622 3272 89628 3284
rect 89680 3272 89686 3324
rect 267734 3272 267740 3324
rect 267792 3312 267798 3324
rect 281626 3312 281632 3324
rect 267792 3284 281632 3312
rect 267792 3272 267798 3284
rect 281626 3272 281632 3284
rect 281684 3272 281690 3324
rect 84470 3204 84476 3256
rect 84528 3244 84534 3256
rect 85482 3244 85488 3256
rect 84528 3216 85488 3244
rect 84528 3204 84534 3216
rect 85482 3204 85488 3216
rect 85540 3204 85546 3256
rect 324958 3204 324964 3256
rect 325016 3244 325022 3256
rect 325602 3244 325608 3256
rect 325016 3216 325608 3244
rect 325016 3204 325022 3216
rect 325602 3204 325608 3216
rect 325660 3204 325666 3256
rect 341518 3204 341524 3256
rect 341576 3244 341582 3256
rect 344554 3244 344560 3256
rect 341576 3216 344560 3244
rect 341576 3204 341582 3216
rect 344554 3204 344560 3216
rect 344612 3204 344618 3256
rect 83274 3136 83280 3188
rect 83332 3176 83338 3188
rect 84102 3176 84108 3188
rect 83332 3148 84108 3176
rect 83332 3136 83338 3148
rect 84102 3136 84108 3148
rect 84160 3136 84166 3188
rect 299382 3136 299388 3188
rect 299440 3176 299446 3188
rect 301958 3176 301964 3188
rect 299440 3148 301964 3176
rect 299440 3136 299446 3148
rect 301958 3136 301964 3148
rect 302016 3136 302022 3188
rect 60826 3000 60832 3052
rect 60884 3040 60890 3052
rect 61930 3040 61936 3052
rect 60884 3012 61936 3040
rect 60884 3000 60890 3012
rect 61930 3000 61936 3012
rect 61988 3000 61994 3052
rect 82078 3000 82084 3052
rect 82136 3040 82142 3052
rect 82722 3040 82728 3052
rect 82136 3012 82728 3040
rect 82136 3000 82142 3012
rect 82722 3000 82728 3012
rect 82780 3000 82786 3052
rect 580994 3000 581000 3052
rect 581052 3040 581058 3052
rect 582834 3040 582840 3052
rect 581052 3012 582840 3040
rect 581052 3000 581058 3012
rect 582834 3000 582840 3012
rect 582892 3000 582898 3052
rect 19426 2932 19432 2984
rect 19484 2972 19490 2984
rect 20622 2972 20628 2984
rect 19484 2944 20628 2972
rect 19484 2932 19490 2944
rect 20622 2932 20628 2944
rect 20680 2932 20686 2984
rect 129366 2932 129372 2984
rect 129424 2972 129430 2984
rect 133138 2972 133144 2984
rect 129424 2944 133144 2972
rect 129424 2932 129430 2944
rect 133138 2932 133144 2944
rect 133196 2932 133202 2984
rect 239306 2932 239312 2984
rect 239364 2972 239370 2984
rect 240962 2972 240968 2984
rect 239364 2944 240968 2972
rect 239364 2932 239370 2944
rect 240962 2932 240968 2944
rect 241020 2932 241026 2984
rect 272426 2932 272432 2984
rect 272484 2972 272490 2984
rect 273990 2972 273996 2984
rect 272484 2944 273996 2972
rect 272484 2932 272490 2944
rect 273990 2932 273996 2944
rect 274048 2932 274054 2984
rect 242894 2728 242900 2780
rect 242952 2768 242958 2780
rect 412634 2768 412640 2780
rect 242952 2740 412640 2768
rect 242952 2728 242958 2740
rect 412634 2728 412640 2740
rect 412692 2728 412698 2780
rect 51350 2116 51356 2168
rect 51408 2156 51414 2168
rect 58618 2156 58624 2168
rect 51408 2128 58624 2156
rect 51408 2116 51414 2128
rect 58618 2116 58624 2128
rect 58676 2116 58682 2168
rect 111610 2116 111616 2168
rect 111668 2156 111674 2168
rect 222838 2156 222844 2168
rect 111668 2128 222844 2156
rect 111668 2116 111674 2128
rect 222838 2116 222844 2128
rect 222896 2116 222902 2168
rect 7650 2048 7656 2100
rect 7708 2088 7714 2100
rect 54478 2088 54484 2100
rect 7708 2060 54484 2088
rect 7708 2048 7714 2060
rect 54478 2048 54484 2060
rect 54536 2048 54542 2100
rect 71498 2048 71504 2100
rect 71556 2088 71562 2100
rect 233878 2088 233884 2100
rect 71556 2060 233884 2088
rect 71556 2048 71562 2060
rect 233878 2048 233884 2060
rect 233936 2048 233942 2100
rect 350442 2048 350448 2100
rect 350500 2088 350506 2100
rect 381630 2088 381636 2100
rect 350500 2060 381636 2088
rect 350500 2048 350506 2060
rect 381630 2048 381636 2060
rect 381688 2048 381694 2100
rect 307754 552 307760 604
rect 307812 592 307818 604
rect 309042 592 309048 604
rect 307812 564 309048 592
rect 307812 552 307818 564
rect 309042 552 309048 564
rect 309100 552 309106 604
<< via1 >>
rect 331220 702992 331272 703044
rect 332508 702992 332560 703044
rect 62028 702924 62080 702976
rect 267648 702924 267700 702976
rect 283840 702924 283892 702976
rect 351920 702924 351972 702976
rect 202788 702856 202840 702908
rect 273260 702856 273312 702908
rect 276664 702856 276716 702908
rect 478512 702856 478564 702908
rect 67640 702652 67692 702704
rect 170312 702652 170364 702704
rect 281540 702788 281592 702840
rect 349804 702788 349856 702840
rect 494796 702788 494848 702840
rect 233884 702720 233936 702772
rect 397368 702720 397420 702772
rect 191748 702652 191800 702704
rect 364984 702652 365036 702704
rect 378784 702652 378836 702704
rect 462320 702652 462372 702704
rect 24308 702584 24360 702636
rect 79324 702584 79376 702636
rect 95148 702584 95200 702636
rect 300124 702584 300176 702636
rect 300768 702584 300820 702636
rect 359464 702584 359516 702636
rect 543464 702584 543516 702636
rect 88248 702516 88300 702568
rect 235172 702516 235224 702568
rect 264244 702516 264296 702568
rect 559656 702516 559708 702568
rect 8116 702448 8168 702500
rect 88800 702448 88852 702500
rect 99288 702448 99340 702500
rect 527180 702448 527232 702500
rect 124864 700340 124916 700392
rect 137836 700340 137888 700392
rect 75184 700272 75236 700324
rect 105452 700272 105504 700324
rect 129004 700272 129056 700324
rect 218980 700272 219032 700324
rect 300768 700272 300820 700324
rect 341524 700272 341576 700324
rect 342904 700272 342956 700324
rect 348792 700272 348844 700324
rect 382924 700272 382976 700324
rect 429844 700272 429896 700324
rect 66168 699660 66220 699712
rect 72976 699660 73028 699712
rect 86224 699660 86276 699712
rect 89168 699660 89220 699712
rect 3424 683136 3476 683188
rect 21364 683136 21416 683188
rect 3516 670692 3568 670744
rect 22744 670692 22796 670744
rect 3516 632068 3568 632120
rect 11704 632068 11756 632120
rect 3516 618264 3568 618316
rect 14464 618264 14516 618316
rect 3516 605820 3568 605872
rect 90364 605820 90416 605872
rect 71780 605072 71832 605124
rect 86224 605072 86276 605124
rect 70308 596164 70360 596216
rect 349804 596164 349856 596216
rect 79324 595620 79376 595672
rect 80336 595620 80388 595672
rect 80336 594872 80388 594924
rect 106924 594872 106976 594924
rect 85948 594804 86000 594856
rect 141424 594804 141476 594856
rect 90364 594260 90416 594312
rect 91100 594260 91152 594312
rect 40040 594056 40092 594108
rect 89812 594056 89864 594108
rect 88248 593376 88300 593428
rect 113180 593376 113232 593428
rect 67364 592696 67416 592748
rect 75184 592696 75236 592748
rect 3424 592628 3476 592680
rect 69112 592628 69164 592680
rect 78588 592084 78640 592136
rect 103520 592084 103572 592136
rect 84108 592016 84160 592068
rect 112444 592016 112496 592068
rect 85028 591948 85080 592000
rect 88248 591948 88300 592000
rect 73068 590792 73120 590844
rect 79324 590792 79376 590844
rect 63316 590724 63368 590776
rect 73896 590724 73948 590776
rect 86868 590656 86920 590708
rect 115296 590656 115348 590708
rect 69112 589364 69164 589416
rect 89076 589364 89128 589416
rect 3424 589296 3476 589348
rect 74908 589296 74960 589348
rect 76748 589296 76800 589348
rect 101404 589296 101456 589348
rect 79324 588616 79376 588668
rect 94504 588616 94556 588668
rect 79784 588548 79836 588600
rect 105544 588548 105596 588600
rect 75920 588412 75972 588464
rect 52276 587868 52328 587920
rect 66812 587868 66864 587920
rect 88892 588344 88944 588396
rect 88892 588140 88944 588192
rect 88984 587800 89036 587852
rect 88984 586576 89036 586628
rect 98644 586576 98696 586628
rect 55128 586508 55180 586560
rect 66260 586508 66312 586560
rect 91744 586508 91796 586560
rect 95240 586508 95292 586560
rect 57796 585148 57848 585200
rect 66812 585148 66864 585200
rect 88892 584468 88944 584520
rect 116584 584468 116636 584520
rect 91376 584400 91428 584452
rect 95148 584400 95200 584452
rect 132500 584400 132552 584452
rect 91192 583652 91244 583704
rect 99288 583652 99340 583704
rect 99288 582972 99340 583024
rect 108304 582972 108356 583024
rect 50988 582360 51040 582412
rect 66812 582360 66864 582412
rect 59268 581000 59320 581052
rect 66720 581000 66772 581052
rect 91744 581000 91796 581052
rect 148416 581000 148468 581052
rect 64788 579640 64840 579692
rect 66812 579640 66864 579692
rect 91744 579640 91796 579692
rect 142804 579640 142856 579692
rect 91744 578212 91796 578264
rect 120724 578212 120776 578264
rect 95884 577464 95936 577516
rect 109040 577464 109092 577516
rect 11704 576104 11756 576156
rect 67456 576104 67508 576156
rect 91100 576104 91152 576156
rect 123116 576104 123168 576156
rect 142804 574744 142856 574796
rect 276020 574744 276072 574796
rect 276020 574404 276072 574456
rect 276664 574404 276716 574456
rect 61936 574064 61988 574116
rect 67364 574064 67416 574116
rect 91100 574064 91152 574116
rect 122196 574064 122248 574116
rect 91100 572704 91152 572756
rect 115204 572704 115256 572756
rect 49608 571344 49660 571396
rect 66812 571344 66864 571396
rect 91100 571344 91152 571396
rect 95148 571344 95200 571396
rect 91192 570596 91244 570648
rect 121552 570596 121604 570648
rect 91100 569916 91152 569968
rect 101496 569916 101548 569968
rect 95148 569168 95200 569220
rect 129740 569168 129792 569220
rect 60648 568556 60700 568608
rect 66812 568556 66864 568608
rect 91100 568556 91152 568608
rect 100024 568556 100076 568608
rect 129740 568556 129792 568608
rect 213920 568556 213972 568608
rect 120724 568488 120776 568540
rect 121368 568488 121420 568540
rect 53656 567196 53708 567248
rect 66812 567196 66864 567248
rect 121368 567196 121420 567248
rect 332600 567196 332652 567248
rect 101496 566448 101548 566500
rect 127440 566448 127492 566500
rect 184204 565904 184256 565956
rect 311900 565904 311952 565956
rect 59084 565836 59136 565888
rect 67640 565836 67692 565888
rect 91376 565836 91428 565888
rect 102784 565836 102836 565888
rect 126980 565836 127032 565888
rect 127440 565836 127492 565888
rect 291200 565836 291252 565888
rect 91468 565088 91520 565140
rect 134524 565088 134576 565140
rect 54484 564408 54536 564460
rect 66812 564408 66864 564460
rect 91376 564408 91428 564460
rect 101496 564408 101548 564460
rect 162768 564408 162820 564460
rect 309140 564408 309192 564460
rect 52368 563048 52420 563100
rect 66812 563048 66864 563100
rect 91376 563048 91428 563100
rect 194600 563116 194652 563168
rect 241520 563116 241572 563168
rect 196624 563048 196676 563100
rect 295984 563048 296036 563100
rect 115296 562504 115348 562556
rect 117964 562504 118016 562556
rect 67456 562300 67508 562352
rect 68284 562300 68336 562352
rect 166356 561756 166408 561808
rect 335360 561756 335412 561808
rect 37188 561688 37240 561740
rect 66812 561688 66864 561740
rect 111064 561688 111116 561740
rect 111708 561688 111760 561740
rect 357532 561688 357584 561740
rect 153108 560328 153160 560380
rect 215300 560328 215352 560380
rect 44088 560260 44140 560312
rect 66812 560260 66864 560312
rect 194508 560260 194560 560312
rect 268384 560260 268436 560312
rect 273260 559648 273312 559700
rect 273904 559648 273956 559700
rect 198464 558968 198516 559020
rect 273904 558968 273956 559020
rect 89628 558900 89680 558952
rect 122104 558900 122156 558952
rect 122196 558900 122248 558952
rect 122932 558900 122984 558952
rect 196716 558900 196768 558952
rect 343640 558900 343692 558952
rect 60740 558628 60792 558680
rect 62028 558628 62080 558680
rect 66260 558628 66312 558680
rect 39948 558152 40000 558204
rect 60740 558152 60792 558204
rect 198648 558152 198700 558204
rect 582932 558152 582984 558204
rect 91192 557540 91244 557592
rect 151820 557540 151872 557592
rect 191104 557540 191156 557592
rect 270500 557540 270552 557592
rect 91284 556248 91336 556300
rect 121460 556248 121512 556300
rect 195888 556248 195940 556300
rect 288440 556248 288492 556300
rect 112444 556180 112496 556232
rect 226984 556180 227036 556232
rect 187056 554820 187108 554872
rect 237380 554820 237432 554872
rect 56508 554752 56560 554804
rect 66812 554752 66864 554804
rect 198096 554752 198148 554804
rect 268292 554752 268344 554804
rect 188620 553460 188672 553512
rect 260104 553460 260156 553512
rect 3332 553392 3384 553444
rect 43444 553392 43496 553444
rect 64696 553392 64748 553444
rect 66444 553392 66496 553444
rect 91100 553392 91152 553444
rect 112536 553392 112588 553444
rect 134524 553392 134576 553444
rect 210424 553392 210476 553444
rect 91100 552100 91152 552152
rect 104256 552100 104308 552152
rect 156604 552100 156656 552152
rect 238760 552100 238812 552152
rect 92112 552032 92164 552084
rect 108396 552032 108448 552084
rect 124956 552032 125008 552084
rect 351920 552032 351972 552084
rect 117964 551964 118016 552016
rect 118608 551964 118660 552016
rect 91100 550672 91152 550724
rect 128360 550672 128412 550724
rect 180248 550672 180300 550724
rect 182088 550672 182140 550724
rect 240232 550672 240284 550724
rect 118608 550604 118660 550656
rect 212540 550604 212592 550656
rect 193956 549312 194008 549364
rect 223672 549312 223724 549364
rect 60556 549244 60608 549296
rect 66812 549244 66864 549296
rect 187608 549244 187660 549296
rect 220820 549244 220872 549296
rect 192484 547952 192536 548004
rect 287060 547952 287112 548004
rect 57704 547884 57756 547936
rect 66812 547884 66864 547936
rect 91376 547884 91428 547936
rect 245660 547884 245712 547936
rect 295340 547884 295392 547936
rect 372620 547884 372672 547936
rect 204904 546524 204956 546576
rect 251824 546524 251876 546576
rect 62028 546456 62080 546508
rect 66904 546456 66956 546508
rect 91560 546456 91612 546508
rect 104164 546456 104216 546508
rect 188436 546456 188488 546508
rect 305000 546456 305052 546508
rect 327080 546456 327132 546508
rect 361856 546456 361908 546508
rect 199384 545164 199436 545216
rect 298376 545164 298428 545216
rect 314936 545164 314988 545216
rect 363052 545164 363104 545216
rect 50896 545096 50948 545148
rect 66904 545096 66956 545148
rect 91100 545096 91152 545148
rect 94596 545096 94648 545148
rect 186964 545096 187016 545148
rect 324320 545096 324372 545148
rect 331680 545096 331732 545148
rect 364432 545096 364484 545148
rect 199476 543804 199528 543856
rect 229100 543804 229152 543856
rect 318248 543804 318300 543856
rect 365720 543804 365772 543856
rect 48228 543736 48280 543788
rect 66904 543736 66956 543788
rect 182824 543736 182876 543788
rect 321560 543736 321612 543788
rect 330024 543736 330076 543788
rect 376852 543736 376904 543788
rect 21364 542988 21416 543040
rect 34520 542988 34572 543040
rect 175924 542444 175976 542496
rect 280160 542444 280212 542496
rect 338304 542444 338356 542496
rect 367284 542444 367336 542496
rect 34520 542376 34572 542428
rect 35808 542376 35860 542428
rect 66904 542376 66956 542428
rect 91100 542376 91152 542428
rect 95884 542376 95936 542428
rect 133144 542376 133196 542428
rect 357440 542376 357492 542428
rect 22744 541628 22796 541680
rect 66996 541628 67048 541680
rect 67272 541628 67324 541680
rect 91100 541628 91152 541680
rect 124864 541628 124916 541680
rect 131580 541628 131632 541680
rect 131120 541016 131172 541068
rect 131580 541016 131632 541068
rect 258448 541016 258500 541068
rect 88892 540948 88944 541000
rect 266360 540948 266412 541000
rect 324320 540880 324372 540932
rect 324964 540880 325016 540932
rect 342904 540880 342956 540932
rect 3424 540200 3476 540252
rect 67548 539724 67600 539776
rect 91100 539656 91152 539708
rect 101588 539656 101640 539708
rect 144828 539656 144880 539708
rect 283932 539656 283984 539708
rect 328828 539656 328880 539708
rect 360476 539656 360528 539708
rect 63408 539588 63460 539640
rect 67548 539588 67600 539640
rect 69388 539588 69440 539640
rect 71872 539588 71924 539640
rect 81164 539588 81216 539640
rect 88800 539588 88852 539640
rect 88156 539520 88208 539572
rect 250628 539588 250680 539640
rect 349988 539588 350040 539640
rect 393964 539588 394016 539640
rect 268384 539520 268436 539572
rect 272340 539520 272392 539572
rect 273904 539520 273956 539572
rect 275652 539520 275704 539572
rect 278044 539520 278096 539572
rect 278964 539520 279016 539572
rect 17224 538840 17276 538892
rect 91192 538840 91244 538892
rect 172428 538840 172480 538892
rect 195244 538840 195296 538892
rect 195796 538296 195848 538348
rect 202788 538296 202840 538348
rect 221096 538296 221148 538348
rect 232412 538296 232464 538348
rect 295984 538296 296036 538348
rect 297180 538296 297232 538348
rect 323676 538296 323728 538348
rect 340788 538296 340840 538348
rect 347044 538296 347096 538348
rect 360200 538296 360252 538348
rect 67824 538228 67876 538280
rect 76564 538228 76616 538280
rect 166264 538228 166316 538280
rect 204168 538228 204220 538280
rect 208400 538228 208452 538280
rect 356336 538228 356388 538280
rect 86868 538160 86920 538212
rect 129004 538160 129056 538212
rect 340788 538160 340840 538212
rect 579896 538160 579948 538212
rect 8208 537480 8260 537532
rect 91284 537480 91336 537532
rect 198740 537480 198792 537532
rect 208400 537480 208452 537532
rect 129648 536800 129700 536852
rect 267188 536800 267240 536852
rect 43444 536732 43496 536784
rect 70492 536732 70544 536784
rect 72332 536732 72384 536784
rect 81164 536732 81216 536784
rect 68652 536664 68704 536716
rect 88156 536664 88208 536716
rect 353944 536052 353996 536104
rect 354588 536052 354640 536104
rect 359464 536052 359516 536104
rect 198004 535576 198056 535628
rect 201316 535576 201368 535628
rect 148324 535508 148376 535560
rect 293500 535508 293552 535560
rect 82728 535440 82780 535492
rect 86224 535440 86276 535492
rect 201408 535440 201460 535492
rect 580264 535440 580316 535492
rect 78312 534760 78364 534812
rect 124220 534760 124272 534812
rect 125048 534760 125100 534812
rect 177304 534760 177356 534812
rect 193956 534760 194008 534812
rect 199844 534760 199896 534812
rect 204904 535236 204956 535288
rect 355600 535236 355652 535288
rect 427820 534760 427872 534812
rect 18604 534692 18656 534744
rect 91192 534692 91244 534744
rect 180064 534692 180116 534744
rect 198740 534692 198792 534744
rect 125048 534080 125100 534132
rect 140780 534080 140832 534132
rect 193864 534080 193916 534132
rect 197360 534080 197412 534132
rect 67364 534012 67416 534064
rect 188620 534012 188672 534064
rect 81072 532652 81124 532704
rect 98000 532652 98052 532704
rect 140780 532652 140832 532704
rect 197360 532652 197412 532704
rect 3424 531972 3476 532024
rect 89720 531972 89772 532024
rect 358728 531972 358780 532024
rect 582932 531972 582984 532024
rect 98000 531292 98052 531344
rect 155224 531292 155276 531344
rect 44088 531224 44140 531276
rect 188528 531224 188580 531276
rect 64788 530544 64840 530596
rect 77944 530544 77996 530596
rect 176016 530544 176068 530596
rect 199476 530544 199528 530596
rect 124864 529864 124916 529916
rect 197360 529864 197412 529916
rect 64696 529796 64748 529848
rect 124956 529796 125008 529848
rect 79324 529728 79376 529780
rect 79968 529728 80020 529780
rect 59268 529184 59320 529236
rect 79324 529184 79376 529236
rect 358728 528572 358780 528624
rect 371240 528572 371292 528624
rect 180248 528504 180300 528556
rect 197360 528504 197412 528556
rect 70400 527484 70452 527536
rect 71044 527484 71096 527536
rect 71044 527144 71096 527196
rect 141516 527144 141568 527196
rect 358728 527144 358780 527196
rect 376760 527144 376812 527196
rect 50896 527076 50948 527128
rect 160836 527076 160888 527128
rect 173164 525036 173216 525088
rect 198004 525036 198056 525088
rect 170404 524424 170456 524476
rect 197360 524424 197412 524476
rect 358728 524424 358780 524476
rect 375472 524424 375524 524476
rect 59176 523676 59228 523728
rect 78772 523676 78824 523728
rect 66904 522248 66956 522300
rect 177396 522248 177448 522300
rect 147588 521636 147640 521688
rect 197360 521636 197412 521688
rect 34428 520888 34480 520940
rect 195244 520888 195296 520940
rect 358728 520888 358780 520940
rect 395988 520888 396040 520940
rect 395988 520276 396040 520328
rect 582472 520276 582524 520328
rect 55128 519528 55180 519580
rect 85580 519528 85632 519580
rect 358728 519528 358780 519580
rect 388444 519528 388496 519580
rect 62028 517420 62080 517472
rect 186964 517420 187016 517472
rect 180248 516128 180300 516180
rect 197360 516128 197412 516180
rect 358728 516128 358780 516180
rect 374736 516128 374788 516180
rect 3516 514768 3568 514820
rect 14464 514768 14516 514820
rect 175188 514768 175240 514820
rect 197360 514768 197412 514820
rect 60556 514700 60608 514752
rect 188436 514700 188488 514752
rect 41328 511232 41380 511284
rect 180156 511232 180208 511284
rect 141516 510552 141568 510604
rect 197360 510552 197412 510604
rect 358728 509668 358780 509720
rect 360292 509668 360344 509720
rect 46848 507084 46900 507136
rect 196808 507084 196860 507136
rect 358728 505112 358780 505164
rect 414664 505112 414716 505164
rect 164884 504364 164936 504416
rect 197360 504364 197412 504416
rect 358728 502324 358780 502376
rect 369860 502324 369912 502376
rect 3516 502256 3568 502308
rect 18604 502256 18656 502308
rect 155224 500896 155276 500948
rect 198280 500896 198332 500948
rect 155868 498788 155920 498840
rect 180248 498788 180300 498840
rect 180156 496816 180208 496868
rect 197360 496816 197412 496868
rect 357164 496748 357216 496800
rect 583024 496748 583076 496800
rect 178684 495456 178736 495508
rect 197360 495456 197412 495508
rect 358636 493960 358688 494012
rect 412640 493960 412692 494012
rect 138664 492668 138716 492720
rect 197360 492668 197412 492720
rect 127624 488520 127676 488572
rect 151820 488520 151872 488572
rect 197360 488452 197412 488504
rect 358728 486412 358780 486464
rect 385040 486412 385092 486464
rect 181628 483624 181680 483676
rect 197360 483624 197412 483676
rect 358728 481652 358780 481704
rect 364340 481652 364392 481704
rect 180248 480224 180300 480276
rect 197360 480224 197412 480276
rect 358728 480224 358780 480276
rect 378140 480224 378192 480276
rect 124864 477504 124916 477556
rect 171048 477504 171100 477556
rect 197360 477504 197412 477556
rect 358728 477504 358780 477556
rect 367192 477504 367244 477556
rect 68284 476076 68336 476128
rect 68928 476076 68980 476128
rect 147496 476008 147548 476060
rect 180064 476008 180116 476060
rect 3332 475328 3384 475380
rect 8208 475328 8260 475380
rect 15844 475328 15896 475380
rect 177396 474716 177448 474768
rect 197360 474716 197412 474768
rect 137284 473356 137336 473408
rect 197360 473356 197412 473408
rect 358544 471996 358596 472048
rect 389180 471996 389232 472048
rect 191196 471248 191248 471300
rect 198096 471248 198148 471300
rect 357900 470568 357952 470620
rect 368572 470568 368624 470620
rect 165528 467848 165580 467900
rect 197360 467848 197412 467900
rect 105544 467780 105596 467832
rect 182088 467780 182140 467832
rect 188436 467780 188488 467832
rect 104900 466420 104952 466472
rect 105544 466420 105596 466472
rect 93768 465672 93820 465724
rect 107660 465672 107712 465724
rect 131764 465060 131816 465112
rect 186964 465060 187016 465112
rect 197360 465060 197412 465112
rect 358728 465060 358780 465112
rect 376944 465060 376996 465112
rect 583024 465060 583076 465112
rect 106188 462952 106240 463004
rect 120816 462952 120868 463004
rect 3516 462340 3568 462392
rect 25504 462340 25556 462392
rect 50988 462340 51040 462392
rect 67732 462340 67784 462392
rect 68836 462340 68888 462392
rect 187148 462340 187200 462392
rect 197360 462340 197412 462392
rect 68836 461592 68888 461644
rect 81440 461592 81492 461644
rect 76012 461456 76064 461508
rect 76564 461456 76616 461508
rect 76564 460912 76616 460964
rect 159364 460912 159416 460964
rect 57888 460164 57940 460216
rect 95240 460164 95292 460216
rect 148968 460164 149020 460216
rect 197360 460164 197412 460216
rect 375288 460164 375340 460216
rect 582564 460164 582616 460216
rect 148416 459552 148468 459604
rect 148968 459552 149020 459604
rect 358452 459552 358504 459604
rect 374092 459552 374144 459604
rect 375288 459552 375340 459604
rect 14464 459484 14516 459536
rect 112444 459484 112496 459536
rect 127716 458192 127768 458244
rect 197360 458192 197412 458244
rect 52276 457444 52328 457496
rect 87052 457444 87104 457496
rect 60648 456696 60700 456748
rect 65616 456696 65668 456748
rect 57796 456016 57848 456068
rect 82820 456016 82872 456068
rect 65616 455404 65668 455456
rect 65892 455404 65944 455456
rect 195244 455404 195296 455456
rect 358728 455404 358780 455456
rect 363236 455404 363288 455456
rect 582472 455404 582524 455456
rect 172244 455336 172296 455388
rect 172428 455336 172480 455388
rect 173256 455336 173308 455388
rect 88340 454792 88392 454844
rect 88984 454792 89036 454844
rect 63316 454656 63368 454708
rect 95884 454656 95936 454708
rect 88340 454044 88392 454096
rect 133880 454044 133932 454096
rect 65984 453976 66036 454028
rect 71044 453976 71096 454028
rect 97264 453976 97316 454028
rect 102140 453976 102192 454028
rect 57612 453296 57664 453348
rect 73160 453296 73212 453348
rect 102784 453296 102836 453348
rect 125600 453296 125652 453348
rect 77944 452616 77996 452668
rect 128452 452616 128504 452668
rect 358728 452616 358780 452668
rect 398840 452616 398892 452668
rect 116584 451936 116636 451988
rect 124312 451936 124364 451988
rect 3424 451868 3476 451920
rect 121644 451868 121696 451920
rect 95884 451188 95936 451240
rect 124864 451188 124916 451240
rect 106924 451120 106976 451172
rect 127716 451120 127768 451172
rect 63224 450508 63276 450560
rect 75920 450508 75972 450560
rect 358728 449896 358780 449948
rect 375380 449896 375432 449948
rect 25504 449828 25556 449880
rect 71780 449828 71832 449880
rect 64696 449216 64748 449268
rect 78680 449216 78732 449268
rect 100024 449216 100076 449268
rect 123576 449216 123628 449268
rect 71780 449148 71832 449200
rect 72700 449148 72752 449200
rect 103520 449148 103572 449200
rect 103704 449148 103756 449200
rect 358728 449148 358780 449200
rect 365904 449148 365956 449200
rect 582656 449148 582708 449200
rect 3148 448536 3200 448588
rect 18604 448536 18656 448588
rect 119344 448536 119396 448588
rect 137376 448536 137428 448588
rect 184756 448536 184808 448588
rect 197360 448536 197412 448588
rect 94504 448468 94556 448520
rect 187148 448468 187200 448520
rect 61936 447788 61988 447840
rect 71780 447788 71832 447840
rect 68284 447176 68336 447228
rect 71872 447176 71924 447228
rect 71780 447108 71832 447160
rect 124864 447108 124916 447160
rect 68928 447040 68980 447092
rect 73160 447040 73212 447092
rect 109040 447040 109092 447092
rect 109776 447040 109828 447092
rect 148324 447040 148376 447092
rect 140780 446768 140832 446820
rect 142068 446768 142120 446820
rect 142988 446768 143040 446820
rect 71872 446700 71924 446752
rect 74816 446700 74868 446752
rect 49608 446360 49660 446412
rect 67824 446360 67876 446412
rect 68744 446360 68796 446412
rect 112444 445748 112496 445800
rect 112904 445748 112956 445800
rect 124956 445748 125008 445800
rect 195336 445748 195388 445800
rect 197360 445748 197412 445800
rect 358728 445748 358780 445800
rect 368480 445748 368532 445800
rect 130384 445000 130436 445052
rect 195336 445000 195388 445052
rect 59268 444456 59320 444508
rect 79416 444456 79468 444508
rect 101404 444456 101456 444508
rect 127716 444456 127768 444508
rect 4804 444388 4856 444440
rect 118700 444388 118752 444440
rect 120080 444388 120132 444440
rect 120724 444388 120776 444440
rect 130476 444388 130528 444440
rect 124128 444320 124180 444372
rect 124312 444320 124364 444372
rect 166356 444320 166408 444372
rect 147496 444252 147548 444304
rect 148324 444252 148376 444304
rect 191288 443980 191340 444032
rect 191748 443980 191800 444032
rect 197360 443980 197412 444032
rect 358728 442960 358780 443012
rect 372712 442960 372764 443012
rect 124128 441600 124180 441652
rect 163504 441600 163556 441652
rect 195244 441396 195296 441448
rect 197728 441396 197780 441448
rect 49608 440852 49660 440904
rect 68284 440852 68336 440904
rect 358728 440240 358780 440292
rect 367100 440240 367152 440292
rect 121644 440172 121696 440224
rect 131764 440172 131816 440224
rect 65892 439628 65944 439680
rect 66352 439628 66404 439680
rect 133144 439492 133196 439544
rect 169024 439492 169076 439544
rect 180064 438880 180116 438932
rect 197360 438880 197412 438932
rect 358728 438880 358780 438932
rect 392584 438880 392636 438932
rect 124128 438812 124180 438864
rect 132500 438812 132552 438864
rect 133788 438812 133840 438864
rect 53656 438132 53708 438184
rect 60740 438132 60792 438184
rect 133788 438132 133840 438184
rect 151084 438132 151136 438184
rect 60740 437452 60792 437504
rect 61936 437452 61988 437504
rect 66812 437452 66864 437504
rect 124956 436704 125008 436756
rect 157984 436704 158036 436756
rect 162216 436092 162268 436144
rect 197360 436092 197412 436144
rect 357900 436092 357952 436144
rect 360384 436092 360436 436144
rect 41236 435344 41288 435396
rect 59084 435344 59136 435396
rect 66260 435344 66312 435396
rect 147496 434664 147548 434716
rect 148416 434664 148468 434716
rect 44088 433304 44140 433356
rect 54484 433304 54536 433356
rect 124128 433304 124180 433356
rect 147496 433304 147548 433356
rect 358728 433304 358780 433356
rect 370044 433304 370096 433356
rect 66260 433236 66312 433288
rect 124036 431876 124088 431928
rect 142804 431876 142856 431928
rect 52368 431196 52420 431248
rect 65892 431196 65944 431248
rect 66536 431196 66588 431248
rect 183468 430584 183520 430636
rect 197360 430584 197412 430636
rect 358728 430584 358780 430636
rect 371332 430584 371384 430636
rect 121368 429156 121420 429208
rect 121644 429156 121696 429208
rect 36728 429088 36780 429140
rect 37188 429088 37240 429140
rect 66812 429088 66864 429140
rect 14464 428408 14516 428460
rect 36728 428408 36780 428460
rect 169024 427796 169076 427848
rect 197360 427796 197412 427848
rect 358728 427796 358780 427848
rect 382280 427796 382332 427848
rect 43996 427048 44048 427100
rect 52460 427048 52512 427100
rect 140044 426436 140096 426488
rect 197360 426436 197412 426488
rect 358728 426436 358780 426488
rect 369952 426436 370004 426488
rect 52460 425688 52512 425740
rect 53656 425688 53708 425740
rect 66812 425688 66864 425740
rect 59084 423648 59136 423700
rect 66076 423648 66128 423700
rect 167644 423648 167696 423700
rect 197360 423648 197412 423700
rect 3148 422900 3200 422952
rect 17224 422900 17276 422952
rect 39948 421540 40000 421592
rect 66076 421540 66128 421592
rect 66628 421540 66680 421592
rect 122932 421540 122984 421592
rect 143448 421540 143500 421592
rect 178776 421540 178828 421592
rect 358728 420928 358780 420980
rect 371424 420928 371476 420980
rect 124312 420860 124364 420912
rect 160744 420860 160796 420912
rect 358084 420180 358136 420232
rect 379520 420180 379572 420232
rect 181444 418140 181496 418192
rect 197360 418140 197412 418192
rect 358728 418140 358780 418192
rect 361672 418140 361724 418192
rect 195796 416780 195848 416832
rect 197360 416780 197412 416832
rect 358728 416780 358780 416832
rect 365812 416780 365864 416832
rect 122932 415148 122984 415200
rect 129740 415148 129792 415200
rect 57796 414672 57848 414724
rect 64788 414672 64840 414724
rect 66812 414672 66864 414724
rect 193956 413992 194008 414044
rect 197360 413992 197412 414044
rect 358728 413992 358780 414044
rect 365996 413992 366048 414044
rect 125692 413924 125744 413976
rect 126980 413924 127032 413976
rect 124128 412700 124180 412752
rect 125692 412700 125744 412752
rect 56416 411272 56468 411324
rect 66720 411272 66772 411324
rect 164148 411272 164200 411324
rect 197360 411272 197412 411324
rect 358728 411272 358780 411324
rect 374000 411272 374052 411324
rect 130476 409776 130528 409828
rect 197360 409776 197412 409828
rect 358728 408484 358780 408536
rect 367376 408484 367428 408536
rect 124128 407736 124180 407788
rect 134524 407736 134576 407788
rect 124128 406172 124180 406224
rect 125508 406172 125560 406224
rect 57704 405764 57756 405816
rect 64788 405764 64840 405816
rect 66352 405764 66404 405816
rect 189724 405696 189776 405748
rect 197360 405696 197412 405748
rect 358728 405696 358780 405748
rect 364524 405696 364576 405748
rect 48136 403588 48188 403640
rect 62028 403588 62080 403640
rect 66352 403588 66404 403640
rect 358728 403452 358780 403504
rect 363144 403452 363196 403504
rect 123852 403316 123904 403368
rect 124956 403316 125008 403368
rect 125508 402296 125560 402348
rect 127808 402296 127860 402348
rect 358728 401616 358780 401668
rect 406384 401616 406436 401668
rect 123944 400868 123996 400920
rect 194600 400868 194652 400920
rect 188988 400392 189040 400444
rect 191288 400392 191340 400444
rect 50896 400188 50948 400240
rect 55036 400188 55088 400240
rect 66352 400188 66404 400240
rect 194600 400188 194652 400240
rect 195244 400188 195296 400240
rect 191748 398896 191800 398948
rect 197360 398896 197412 398948
rect 48228 398828 48280 398880
rect 50896 398828 50948 398880
rect 66352 398828 66404 398880
rect 124128 398828 124180 398880
rect 125600 398828 125652 398880
rect 192576 398828 192628 398880
rect 358636 398828 358688 398880
rect 361764 398828 361816 398880
rect 2780 398692 2832 398744
rect 4804 398692 4856 398744
rect 125048 397468 125100 397520
rect 191288 397468 191340 397520
rect 191748 397468 191800 397520
rect 35808 396720 35860 396772
rect 66996 396720 67048 396772
rect 177856 396040 177908 396092
rect 197360 396040 197412 396092
rect 121552 395972 121604 396024
rect 127624 395972 127676 396024
rect 143356 394680 143408 394732
rect 197360 394680 197412 394732
rect 123760 393932 123812 393984
rect 160744 393932 160796 393984
rect 358728 393320 358780 393372
rect 368664 393320 368716 393372
rect 63316 391960 63368 392012
rect 66812 391960 66864 392012
rect 121460 391960 121512 392012
rect 153936 391960 153988 392012
rect 3424 391212 3476 391264
rect 73344 391008 73396 391060
rect 104072 391008 104124 391060
rect 131120 391212 131172 391264
rect 120448 390260 120500 390312
rect 120816 390260 120868 390312
rect 113088 389784 113140 389836
rect 120632 389784 120684 389836
rect 59176 389240 59228 389292
rect 87052 389240 87104 389292
rect 15844 389172 15896 389224
rect 111432 389172 111484 389224
rect 67640 389104 67692 389156
rect 68468 389104 68520 389156
rect 96160 389104 96212 389156
rect 125048 389104 125100 389156
rect 65984 389036 66036 389088
rect 73160 389036 73212 389088
rect 73804 389036 73856 389088
rect 101404 389036 101456 389088
rect 103796 389036 103848 389088
rect 57612 388968 57664 389020
rect 77852 388968 77904 389020
rect 88524 388628 88576 388680
rect 92480 388628 92532 388680
rect 79508 388492 79560 388544
rect 86224 388492 86276 388544
rect 93032 388424 93084 388476
rect 98644 388424 98696 388476
rect 118976 388424 119028 388476
rect 148416 388424 148468 388476
rect 167184 388424 167236 388476
rect 168288 388424 168340 388476
rect 180248 388424 180300 388476
rect 66168 387744 66220 387796
rect 82084 387744 82136 387796
rect 114468 387744 114520 387796
rect 128360 387744 128412 387796
rect 171876 387132 171928 387184
rect 181628 387132 181680 387184
rect 67824 387064 67876 387116
rect 146944 387064 146996 387116
rect 147496 387064 147548 387116
rect 178040 387064 178092 387116
rect 180340 387064 180392 387116
rect 196716 387064 196768 387116
rect 181536 386384 181588 386436
rect 197360 386384 197412 386436
rect 358728 386384 358780 386436
rect 385132 386384 385184 386436
rect 63224 386316 63276 386368
rect 80060 386316 80112 386368
rect 80888 386316 80940 386368
rect 99196 385704 99248 385756
rect 122932 385704 122984 385756
rect 111432 385636 111484 385688
rect 156696 385636 156748 385688
rect 123484 385024 123536 385076
rect 189080 385024 189132 385076
rect 45468 384956 45520 385008
rect 76564 384956 76616 385008
rect 73804 383664 73856 383716
rect 184296 383664 184348 383716
rect 358728 383664 358780 383716
rect 403624 383664 403676 383716
rect 17224 383596 17276 383648
rect 125600 383596 125652 383648
rect 118608 382916 118660 382968
rect 195980 382916 196032 382968
rect 80060 381488 80112 381540
rect 167000 381488 167052 381540
rect 167000 380944 167052 380996
rect 194508 380944 194560 380996
rect 3516 380876 3568 380928
rect 104992 380876 105044 380928
rect 105544 380876 105596 380928
rect 109684 380876 109736 380928
rect 171140 380876 171192 380928
rect 171876 380876 171928 380928
rect 39304 380128 39356 380180
rect 125692 380128 125744 380180
rect 160744 380128 160796 380180
rect 178132 380128 178184 380180
rect 178132 379584 178184 379636
rect 178776 379584 178828 379636
rect 197360 379584 197412 379636
rect 48228 379516 48280 379568
rect 188528 379516 188580 379568
rect 358636 379516 358688 379568
rect 361580 379516 361632 379568
rect 110236 378768 110288 378820
rect 160836 378768 160888 378820
rect 131304 378156 131356 378208
rect 184204 378156 184256 378208
rect 50896 378088 50948 378140
rect 187700 378088 187752 378140
rect 41236 378020 41288 378072
rect 124404 378020 124456 378072
rect 124956 378020 125008 378072
rect 130476 378020 130528 378072
rect 194416 377476 194468 377528
rect 201592 377476 201644 377528
rect 189080 377408 189132 377460
rect 194140 377408 194192 377460
rect 345664 377408 345716 377460
rect 357716 377408 357768 377460
rect 198740 377272 198792 377324
rect 199660 377272 199712 377324
rect 140688 376728 140740 376780
rect 198740 376728 198792 376780
rect 192576 376660 192628 376712
rect 215208 376660 215260 376712
rect 342904 376048 342956 376100
rect 357624 376048 357676 376100
rect 81348 375980 81400 376032
rect 95240 375980 95292 376032
rect 198832 375980 198884 376032
rect 204352 375980 204404 376032
rect 247040 375980 247092 376032
rect 248052 375980 248104 376032
rect 382924 375980 382976 376032
rect 104164 375436 104216 375488
rect 195428 375436 195480 375488
rect 67548 375368 67600 375420
rect 192668 375368 192720 375420
rect 195980 375300 196032 375352
rect 201684 375300 201736 375352
rect 202788 375300 202840 375352
rect 205640 375300 205692 375352
rect 206652 375300 206704 375352
rect 215208 375300 215260 375352
rect 218244 375300 218296 375352
rect 258724 375300 258776 375352
rect 261484 375300 261536 375352
rect 278136 375300 278188 375352
rect 279700 375300 279752 375352
rect 298836 375300 298888 375352
rect 301228 375300 301280 375352
rect 336004 375300 336056 375352
rect 337844 375300 337896 375352
rect 339500 375300 339552 375352
rect 378784 375300 378836 375352
rect 311900 375164 311952 375216
rect 312820 375164 312872 375216
rect 233884 375028 233936 375080
rect 238116 375028 238168 375080
rect 254676 374756 254728 374808
rect 255412 374756 255464 374808
rect 250444 374688 250496 374740
rect 251364 374688 251416 374740
rect 261484 374688 261536 374740
rect 274732 374688 274784 374740
rect 295248 374688 295300 374740
rect 296260 374688 296312 374740
rect 77944 374620 77996 374672
rect 138664 374620 138716 374672
rect 209688 374620 209740 374672
rect 216588 374620 216640 374672
rect 228364 374620 228416 374672
rect 233148 374620 233200 374672
rect 262864 374620 262916 374672
rect 294604 374620 294656 374672
rect 322204 374620 322256 374672
rect 334532 374620 334584 374672
rect 334716 374620 334768 374672
rect 339500 374620 339552 374672
rect 143540 374076 143592 374128
rect 164884 374076 164936 374128
rect 200028 374076 200080 374128
rect 201684 374076 201736 374128
rect 234620 374076 234672 374128
rect 238024 374076 238076 374128
rect 246396 374076 246448 374128
rect 255964 374076 256016 374128
rect 300216 374076 300268 374128
rect 311900 374076 311952 374128
rect 119988 374008 120040 374060
rect 295984 374008 296036 374060
rect 297916 374008 297968 374060
rect 307760 374008 307812 374060
rect 313924 374008 313976 374060
rect 326344 374008 326396 374060
rect 329104 374008 329156 374060
rect 354036 374008 354088 374060
rect 356060 374008 356112 374060
rect 234620 373940 234672 373992
rect 70308 373260 70360 373312
rect 158720 373260 158772 373312
rect 350540 373260 350592 373312
rect 452660 373260 452712 373312
rect 153936 372580 153988 372632
rect 208400 372580 208452 372632
rect 184296 371832 184348 371884
rect 206376 371832 206428 371884
rect 235264 371696 235316 371748
rect 238760 371696 238812 371748
rect 134524 371492 134576 371544
rect 135168 371492 135220 371544
rect 3240 371356 3292 371408
rect 4804 371356 4856 371408
rect 117964 371288 118016 371340
rect 169116 371288 169168 371340
rect 71688 371220 71740 371272
rect 73804 371220 73856 371272
rect 135168 371220 135220 371272
rect 196808 371220 196860 371272
rect 358176 371220 358228 371272
rect 360476 371220 360528 371272
rect 86316 371152 86368 371204
rect 148508 371152 148560 371204
rect 85580 370676 85632 370728
rect 86316 370676 86368 370728
rect 53472 370472 53524 370524
rect 143540 370472 143592 370524
rect 188528 370472 188580 370524
rect 199568 370472 199620 370524
rect 199660 370472 199712 370524
rect 242164 370472 242216 370524
rect 345020 370472 345072 370524
rect 420920 370472 420972 370524
rect 146208 369860 146260 369912
rect 207020 369860 207072 369912
rect 207664 369860 207716 369912
rect 343640 369792 343692 369844
rect 344284 369792 344336 369844
rect 580356 369792 580408 369844
rect 98644 369180 98696 369232
rect 151820 369180 151872 369232
rect 153844 369180 153896 369232
rect 169208 369180 169260 369232
rect 191288 369180 191340 369232
rect 267832 369180 267884 369232
rect 67732 369112 67784 369164
rect 123484 369112 123536 369164
rect 145564 369112 145616 369164
rect 202880 369112 202932 369164
rect 206284 369112 206336 369164
rect 232504 369112 232556 369164
rect 361672 369112 361724 369164
rect 66168 368976 66220 369028
rect 67640 368976 67692 369028
rect 197268 368432 197320 368484
rect 200212 368432 200264 368484
rect 113824 367888 113876 367940
rect 114468 367888 114520 367940
rect 348424 367820 348476 367872
rect 364432 367820 364484 367872
rect 79968 367752 80020 367804
rect 133144 367752 133196 367804
rect 345756 367752 345808 367804
rect 365720 367752 365772 367804
rect 113824 367072 113876 367124
rect 271880 367072 271932 367124
rect 340144 366392 340196 366444
rect 356244 366392 356296 366444
rect 64788 366324 64840 366376
rect 107752 366324 107804 366376
rect 341616 366324 341668 366376
rect 367284 366324 367336 366376
rect 126244 365780 126296 365832
rect 199384 365780 199436 365832
rect 144736 365712 144788 365764
rect 340144 365712 340196 365764
rect 66904 365644 66956 365696
rect 67364 365644 67416 365696
rect 359096 365644 359148 365696
rect 192760 364964 192812 365016
rect 213828 364964 213880 365016
rect 358728 364964 358780 365016
rect 370044 364964 370096 365016
rect 104900 364352 104952 364404
rect 191288 364352 191340 364404
rect 281448 363672 281500 363724
rect 413284 363672 413336 363724
rect 59084 363604 59136 363656
rect 130384 363604 130436 363656
rect 166908 363604 166960 363656
rect 309140 363604 309192 363656
rect 139308 362992 139360 363044
rect 143356 362992 143408 363044
rect 110328 362924 110380 362976
rect 196624 362924 196676 362976
rect 354588 362244 354640 362296
rect 363052 362244 363104 362296
rect 70308 362176 70360 362228
rect 175096 362176 175148 362228
rect 200764 362176 200816 362228
rect 338764 362176 338816 362228
rect 361580 362176 361632 362228
rect 111800 361564 111852 361616
rect 113088 361564 113140 361616
rect 232596 361564 232648 361616
rect 92204 360884 92256 360936
rect 120816 360884 120868 360936
rect 81624 360816 81676 360868
rect 82084 360816 82136 360868
rect 258172 360816 258224 360868
rect 258724 360816 258776 360868
rect 146116 360204 146168 360256
rect 187056 360204 187108 360256
rect 101128 359524 101180 359576
rect 177396 359524 177448 359576
rect 126980 359456 127032 359508
rect 127716 359456 127768 359508
rect 259460 359456 259512 359508
rect 146944 358708 146996 358760
rect 147588 358708 147640 358760
rect 3424 358572 3476 358624
rect 7564 358572 7616 358624
rect 167736 358096 167788 358148
rect 232504 358096 232556 358148
rect 56324 358028 56376 358080
rect 109684 358028 109736 358080
rect 147588 358028 147640 358080
rect 167092 358028 167144 358080
rect 167644 358028 167696 358080
rect 207664 358028 207716 358080
rect 307024 358028 307076 358080
rect 107752 357416 107804 357468
rect 206468 357416 206520 357468
rect 93768 357348 93820 357400
rect 131028 357348 131080 357400
rect 229100 357348 229152 357400
rect 238116 357348 238168 357400
rect 167092 356804 167144 356856
rect 191196 356804 191248 356856
rect 140780 356736 140832 356788
rect 141424 356736 141476 356788
rect 167736 356736 167788 356788
rect 194140 356736 194192 356788
rect 227076 356736 227128 356788
rect 76564 356668 76616 356720
rect 123024 356668 123076 356720
rect 124036 356668 124088 356720
rect 160744 356668 160796 356720
rect 252560 356736 252612 356788
rect 300124 356736 300176 356788
rect 282184 356668 282236 356720
rect 376944 356668 376996 356720
rect 96528 355376 96580 355428
rect 99196 355376 99248 355428
rect 245660 355376 245712 355428
rect 263600 355376 263652 355428
rect 84108 355308 84160 355360
rect 108764 355308 108816 355360
rect 111708 355308 111760 355360
rect 300216 355308 300268 355360
rect 309876 355308 309928 355360
rect 359004 355308 359056 355360
rect 201592 355172 201644 355224
rect 202144 355172 202196 355224
rect 102048 354696 102100 354748
rect 201592 354696 201644 354748
rect 72424 354016 72476 354068
rect 87052 354016 87104 354068
rect 273904 354016 273956 354068
rect 295984 354016 296036 354068
rect 67732 353948 67784 354000
rect 117964 353948 118016 354000
rect 195244 353948 195296 354000
rect 211160 353948 211212 354000
rect 226984 353948 227036 354000
rect 364524 353948 364576 354000
rect 121460 353336 121512 353388
rect 177304 353336 177356 353388
rect 114468 353268 114520 353320
rect 153844 353268 153896 353320
rect 154672 353268 154724 353320
rect 155316 353268 155368 353320
rect 234528 353268 234580 353320
rect 240140 353268 240192 353320
rect 77208 352588 77260 352640
rect 152464 352588 152516 352640
rect 152648 352588 152700 352640
rect 223580 352588 223632 352640
rect 86868 352520 86920 352572
rect 99380 352520 99432 352572
rect 105544 352520 105596 352572
rect 181628 352520 181680 352572
rect 152648 351908 152700 351960
rect 153108 351908 153160 351960
rect 223580 351908 223632 351960
rect 224316 351908 224368 351960
rect 74448 351228 74500 351280
rect 113824 351228 113876 351280
rect 90456 351160 90508 351212
rect 195244 351160 195296 351212
rect 195336 351160 195388 351212
rect 224224 351160 224276 351212
rect 120080 350548 120132 350600
rect 120816 350548 120868 350600
rect 156788 350548 156840 350600
rect 121552 349868 121604 349920
rect 126244 349868 126296 349920
rect 71596 349800 71648 349852
rect 121460 349800 121512 349852
rect 192668 349800 192720 349852
rect 202788 349800 202840 349852
rect 335360 349800 335412 349852
rect 126796 349188 126848 349240
rect 176200 349188 176252 349240
rect 63224 349120 63276 349172
rect 66904 349120 66956 349172
rect 67364 349120 67416 349172
rect 80152 349120 80204 349172
rect 81348 349120 81400 349172
rect 195336 349120 195388 349172
rect 356704 349120 356756 349172
rect 357348 349120 357400 349172
rect 400220 349120 400272 349172
rect 208492 349052 208544 349104
rect 209044 349052 209096 349104
rect 241428 348440 241480 348492
rect 357348 348440 357400 348492
rect 121736 348372 121788 348424
rect 246396 348372 246448 348424
rect 90364 347760 90416 347812
rect 209044 347760 209096 347812
rect 134984 347692 135036 347744
rect 244280 347692 244332 347744
rect 244924 347692 244976 347744
rect 108304 347080 108356 347132
rect 122104 347080 122156 347132
rect 81348 347012 81400 347064
rect 133880 347012 133932 347064
rect 134984 347012 135036 347064
rect 185584 347012 185636 347064
rect 204444 347012 204496 347064
rect 240876 347012 240928 347064
rect 582932 347012 582984 347064
rect 140136 346400 140188 346452
rect 162952 346400 163004 346452
rect 206468 346332 206520 346384
rect 240140 346332 240192 346384
rect 241428 346332 241480 346384
rect 249616 346332 249668 346384
rect 261484 346332 261536 346384
rect 124864 345652 124916 345704
rect 248512 345652 248564 345704
rect 249616 345652 249668 345704
rect 59084 345040 59136 345092
rect 197360 345040 197412 345092
rect 227628 344972 227680 345024
rect 332600 344972 332652 345024
rect 227076 344428 227128 344480
rect 227628 344428 227680 344480
rect 301320 344292 301372 344344
rect 355324 344292 355376 344344
rect 67272 343680 67324 343732
rect 156512 343680 156564 343732
rect 156696 343680 156748 343732
rect 161480 343680 161532 343732
rect 221556 343680 221608 343732
rect 54944 343612 54996 343664
rect 134800 343612 134852 343664
rect 137284 343612 137336 343664
rect 228364 343612 228416 343664
rect 240784 343612 240836 343664
rect 300952 343612 301004 343664
rect 301320 343612 301372 343664
rect 107568 343000 107620 343052
rect 157340 343000 157392 343052
rect 199568 342932 199620 342984
rect 215944 342932 215996 342984
rect 107476 342864 107528 342916
rect 202236 342864 202288 342916
rect 232596 342864 232648 342916
rect 260104 342864 260156 342916
rect 289728 342864 289780 342916
rect 375472 342864 375524 342916
rect 61752 342252 61804 342304
rect 66260 342252 66312 342304
rect 67364 342252 67416 342304
rect 77116 341504 77168 341556
rect 87604 341504 87656 341556
rect 206376 341504 206428 341556
rect 245108 341504 245160 341556
rect 117228 340960 117280 341012
rect 183008 340960 183060 341012
rect 85580 340892 85632 340944
rect 249892 340892 249944 340944
rect 78588 340212 78640 340264
rect 95148 340212 95200 340264
rect 93492 340144 93544 340196
rect 122196 340144 122248 340196
rect 135168 340144 135220 340196
rect 139492 340144 139544 340196
rect 162952 340144 163004 340196
rect 216680 340144 216732 340196
rect 156512 339872 156564 339924
rect 158812 339872 158864 339924
rect 139400 339532 139452 339584
rect 152464 339532 152516 339584
rect 95148 339464 95200 339516
rect 248420 339464 248472 339516
rect 216128 338716 216180 338768
rect 236000 338716 236052 338768
rect 236644 338716 236696 338768
rect 263784 338716 263836 338768
rect 280804 338716 280856 338768
rect 353944 338716 353996 338768
rect 85396 338376 85448 338428
rect 90456 338376 90508 338428
rect 112352 338172 112404 338224
rect 162308 338172 162360 338224
rect 106280 338104 106332 338156
rect 229192 338104 229244 338156
rect 58624 337356 58676 337408
rect 72424 337356 72476 337408
rect 97080 337356 97132 337408
rect 128452 337356 128504 337408
rect 149244 337356 149296 337408
rect 196808 337356 196860 337408
rect 260932 337356 260984 337408
rect 307116 337356 307168 337408
rect 358176 337356 358228 337408
rect 150348 336812 150400 336864
rect 199660 336812 199712 336864
rect 107844 336744 107896 336796
rect 176108 336744 176160 336796
rect 134800 336676 134852 336728
rect 154212 336676 154264 336728
rect 20 335996 72 336048
rect 50988 335996 51040 336048
rect 94228 335996 94280 336048
rect 118240 335996 118292 336048
rect 133972 335996 134024 336048
rect 140044 335996 140096 336048
rect 162952 336064 163004 336116
rect 153844 335996 153896 336048
rect 224316 335996 224368 336048
rect 228456 335996 228508 336048
rect 300860 335996 300912 336048
rect 154672 335724 154724 335776
rect 155868 335724 155920 335776
rect 158904 335724 158956 335776
rect 61936 335316 61988 335368
rect 132500 335316 132552 335368
rect 64512 334568 64564 334620
rect 108304 334568 108356 334620
rect 135168 334024 135220 334076
rect 158904 334024 158956 334076
rect 104440 333956 104492 334008
rect 170588 333956 170640 334008
rect 154764 333276 154816 333328
rect 217324 333276 217376 333328
rect 75644 333208 75696 333260
rect 140136 333208 140188 333260
rect 195980 333208 196032 333260
rect 582380 333208 582432 333260
rect 67824 332596 67876 332648
rect 71780 332596 71832 332648
rect 148140 332596 148192 332648
rect 158260 332596 158312 332648
rect 260104 332528 260156 332580
rect 344284 332528 344336 332580
rect 166356 332188 166408 332240
rect 168380 332188 168432 332240
rect 76656 332120 76708 332172
rect 77116 332120 77168 332172
rect 83096 332120 83148 332172
rect 84108 332120 84160 332172
rect 91928 332120 91980 332172
rect 92388 332120 92440 332172
rect 95608 332120 95660 332172
rect 96344 332120 96396 332172
rect 100024 332120 100076 332172
rect 100576 332120 100628 332172
rect 102968 332120 103020 332172
rect 103428 332120 103480 332172
rect 113824 332120 113876 332172
rect 114376 332120 114428 332172
rect 116768 332120 116820 332172
rect 117228 332120 117280 332172
rect 177396 331916 177448 331968
rect 200856 331916 200908 331968
rect 70768 331848 70820 331900
rect 71504 331848 71556 331900
rect 156604 331848 156656 331900
rect 166264 331848 166316 331900
rect 167644 331848 167696 331900
rect 195428 331848 195480 331900
rect 195520 331848 195572 331900
rect 261024 331848 261076 331900
rect 146760 331780 146812 331832
rect 150348 331780 150400 331832
rect 79968 331712 80020 331764
rect 84384 331712 84436 331764
rect 88248 331712 88300 331764
rect 90364 331712 90416 331764
rect 132776 331644 132828 331696
rect 133788 331644 133840 331696
rect 80244 331576 80296 331628
rect 81348 331576 81400 331628
rect 118884 331576 118936 331628
rect 119896 331576 119948 331628
rect 123392 331576 123444 331628
rect 124128 331576 124180 331628
rect 109408 331508 109460 331560
rect 110328 331508 110380 331560
rect 129280 331508 129332 331560
rect 135168 331508 135220 331560
rect 88984 331440 89036 331492
rect 89628 331440 89680 331492
rect 90456 331440 90508 331492
rect 93124 331440 93176 331492
rect 94136 331440 94188 331492
rect 95148 331440 95200 331492
rect 98552 331440 98604 331492
rect 99288 331440 99340 331492
rect 124128 331440 124180 331492
rect 124864 331440 124916 331492
rect 130016 331440 130068 331492
rect 131028 331440 131080 331492
rect 138664 331440 138716 331492
rect 139308 331440 139360 331492
rect 143080 331372 143132 331424
rect 144920 331372 144972 331424
rect 50988 331304 51040 331356
rect 69296 331304 69348 331356
rect 72240 331304 72292 331356
rect 75644 331304 75696 331356
rect 110880 331304 110932 331356
rect 111708 331304 111760 331356
rect 119988 331304 120040 331356
rect 120540 331304 120592 331356
rect 143816 331304 143868 331356
rect 144736 331304 144788 331356
rect 151176 331304 151228 331356
rect 152924 331304 152976 331356
rect 67364 331236 67416 331288
rect 154120 331304 154172 331356
rect 158996 331304 159048 331356
rect 49608 331168 49660 331220
rect 137008 331168 137060 331220
rect 137284 331168 137336 331220
rect 144920 331168 144972 331220
rect 153016 331168 153068 331220
rect 260104 331236 260156 331288
rect 260748 331236 260800 331288
rect 157432 331168 157484 331220
rect 298008 331168 298060 331220
rect 371240 331168 371292 331220
rect 152924 331100 152976 331152
rect 156052 331100 156104 331152
rect 167736 330964 167788 331016
rect 169116 330964 169168 331016
rect 162952 330828 163004 330880
rect 165620 330828 165672 330880
rect 150348 330556 150400 330608
rect 155868 330556 155920 330608
rect 165896 330556 165948 330608
rect 199568 330556 199620 330608
rect 245016 330556 245068 330608
rect 305736 330556 305788 330608
rect 36544 330488 36596 330540
rect 49608 330488 49660 330540
rect 195336 330488 195388 330540
rect 266452 330488 266504 330540
rect 7564 329808 7616 329860
rect 125600 329808 125652 329860
rect 155868 329808 155920 329860
rect 167644 329808 167696 329860
rect 149244 329740 149296 329792
rect 155960 329740 156012 329792
rect 156052 329740 156104 329792
rect 159456 329740 159508 329792
rect 169208 329740 169260 329792
rect 172612 329740 172664 329792
rect 173256 329740 173308 329792
rect 175280 329740 175332 329792
rect 194048 329740 194100 329792
rect 259552 329740 259604 329792
rect 374092 329740 374144 329792
rect 114652 329672 114704 329724
rect 115710 329672 115762 329724
rect 150440 329672 150492 329724
rect 156696 329672 156748 329724
rect 69388 329536 69440 329588
rect 76564 329536 76616 329588
rect 158904 329128 158956 329180
rect 166448 329128 166500 329180
rect 176200 329128 176252 329180
rect 184480 329128 184532 329180
rect 11704 328448 11756 328500
rect 115388 329060 115440 329112
rect 124312 329060 124364 329112
rect 139308 329060 139360 329112
rect 22744 327700 22796 327752
rect 152648 329060 152700 329112
rect 156328 329060 156380 329112
rect 165160 329060 165212 329112
rect 235264 329060 235316 329112
rect 374736 329060 374788 329112
rect 409880 329060 409932 329112
rect 156696 328788 156748 328840
rect 156880 328448 156932 328500
rect 165160 328448 165212 328500
rect 266452 328380 266504 328432
rect 267648 328380 267700 328432
rect 349160 328380 349212 328432
rect 156880 328312 156932 328364
rect 156788 328244 156840 328296
rect 158904 327836 158956 327888
rect 161480 327836 161532 327888
rect 189816 327768 189868 327820
rect 211896 327768 211948 327820
rect 168104 327700 168156 327752
rect 195980 327700 196032 327752
rect 239128 327700 239180 327752
rect 259368 327700 259420 327752
rect 156972 327292 157024 327344
rect 161480 327292 161532 327344
rect 216036 327088 216088 327140
rect 275284 327088 275336 327140
rect 259368 327020 259420 327072
rect 358084 327020 358136 327072
rect 199660 326408 199712 326460
rect 221464 326408 221516 326460
rect 165620 326340 165672 326392
rect 201592 326340 201644 326392
rect 207756 326340 207808 326392
rect 212632 326340 212684 326392
rect 214656 326340 214708 326392
rect 255412 326340 255464 326392
rect 326988 326340 327040 326392
rect 348424 326340 348476 326392
rect 55128 325660 55180 325712
rect 66904 325660 66956 325712
rect 158904 325660 158956 325712
rect 191380 325660 191432 325712
rect 238668 325660 238720 325712
rect 325700 325660 325752 325712
rect 326988 325660 327040 325712
rect 158260 325388 158312 325440
rect 163596 325388 163648 325440
rect 188528 325048 188580 325100
rect 206560 325048 206612 325100
rect 196624 324980 196676 325032
rect 228456 324980 228508 325032
rect 161480 324912 161532 324964
rect 195152 324912 195204 324964
rect 214564 324912 214616 324964
rect 341524 324912 341576 324964
rect 162952 324844 163004 324896
rect 165068 324844 165120 324896
rect 158904 324164 158956 324216
rect 160744 324164 160796 324216
rect 187056 323552 187108 323604
rect 220084 323552 220136 323604
rect 254584 323552 254636 323604
rect 282276 323552 282328 323604
rect 330300 323552 330352 323604
rect 351184 323552 351236 323604
rect 158720 323008 158772 323060
rect 243636 323008 243688 323060
rect 236644 322940 236696 322992
rect 237288 322940 237340 322992
rect 329840 322940 329892 322992
rect 330300 322940 330352 322992
rect 191288 322260 191340 322312
rect 220176 322260 220228 322312
rect 195152 322192 195204 322244
rect 234068 322192 234120 322244
rect 289728 322192 289780 322244
rect 313280 322192 313332 322244
rect 158720 321580 158772 321632
rect 166356 321580 166408 321632
rect 233976 321580 234028 321632
rect 259460 321580 259512 321632
rect 260104 321580 260156 321632
rect 4804 321512 4856 321564
rect 66904 321512 66956 321564
rect 184204 320900 184256 320952
rect 232596 320900 232648 320952
rect 166448 320832 166500 320884
rect 196624 320832 196676 320884
rect 214564 320832 214616 320884
rect 277400 320832 277452 320884
rect 285772 320832 285824 320884
rect 286968 320832 287020 320884
rect 360200 320832 360252 320884
rect 52368 320152 52420 320204
rect 66812 320152 66864 320204
rect 158720 320152 158772 320204
rect 164976 320152 165028 320204
rect 241980 320152 242032 320204
rect 285772 320152 285824 320204
rect 176016 319472 176068 319524
rect 209136 319472 209188 319524
rect 245108 319472 245160 319524
rect 255320 319472 255372 319524
rect 53656 319404 53708 319456
rect 66996 319404 67048 319456
rect 67272 319404 67324 319456
rect 158720 319404 158772 319456
rect 167000 319404 167052 319456
rect 170588 319404 170640 319456
rect 206284 319404 206336 319456
rect 253204 319404 253256 319456
rect 264980 319404 265032 319456
rect 4068 318724 4120 318776
rect 39304 318724 39356 318776
rect 63224 318520 63276 318572
rect 66812 318520 66864 318572
rect 252468 318044 252520 318096
rect 342260 318044 342312 318096
rect 169668 317500 169720 317552
rect 173164 317500 173216 317552
rect 205916 317500 205968 317552
rect 259460 317500 259512 317552
rect 61936 317432 61988 317484
rect 66720 317432 66772 317484
rect 158720 317432 158772 317484
rect 240968 317432 241020 317484
rect 158812 317364 158864 317416
rect 166448 317364 166500 317416
rect 166724 317364 166776 317416
rect 351920 316752 351972 316804
rect 352564 316752 352616 316804
rect 29644 316684 29696 316736
rect 64512 316684 64564 316736
rect 66812 316684 66864 316736
rect 166448 316684 166500 316736
rect 184296 316684 184348 316736
rect 211068 316684 211120 316736
rect 240876 316684 240928 316736
rect 320180 316684 320232 316736
rect 360292 316684 360344 316736
rect 245660 316072 245712 316124
rect 320180 316072 320232 316124
rect 61936 316004 61988 316056
rect 65524 316004 65576 316056
rect 188436 316004 188488 316056
rect 209964 316004 210016 316056
rect 211068 316004 211120 316056
rect 223028 316004 223080 316056
rect 352564 316004 352616 316056
rect 66628 315936 66680 315988
rect 209044 315256 209096 315308
rect 215852 315256 215904 315308
rect 63316 314916 63368 314968
rect 66168 314916 66220 314968
rect 66536 314916 66588 314968
rect 158720 314712 158772 314764
rect 175096 314712 175148 314764
rect 178684 314712 178736 314764
rect 164148 314644 164200 314696
rect 262312 314644 262364 314696
rect 60464 314576 60516 314628
rect 66904 314576 66956 314628
rect 158720 314576 158772 314628
rect 178684 313896 178736 313948
rect 188436 313896 188488 313948
rect 195428 313896 195480 313948
rect 212908 313896 212960 313948
rect 217324 313896 217376 313948
rect 236000 313896 236052 313948
rect 238024 313896 238076 313948
rect 251272 313896 251324 313948
rect 158720 313284 158772 313336
rect 180156 313284 180208 313336
rect 226248 313284 226300 313336
rect 269212 313284 269264 313336
rect 54944 313216 54996 313268
rect 66904 313216 66956 313268
rect 191104 312672 191156 312724
rect 221648 312672 221700 312724
rect 188528 312536 188580 312588
rect 205916 312536 205968 312588
rect 221556 312536 221608 312588
rect 252836 312536 252888 312588
rect 260104 312536 260156 312588
rect 460940 312536 460992 312588
rect 212908 311856 212960 311908
rect 327724 311856 327776 311908
rect 164976 311788 165028 311840
rect 245660 311788 245712 311840
rect 39948 311108 40000 311160
rect 67088 311108 67140 311160
rect 67456 311108 67508 311160
rect 246304 311108 246356 311160
rect 256700 311108 256752 311160
rect 4804 310496 4856 310548
rect 39948 310496 40000 310548
rect 206560 310496 206612 310548
rect 206836 310496 206888 310548
rect 276756 310496 276808 310548
rect 292580 310224 292632 310276
rect 293224 310224 293276 310276
rect 193036 309884 193088 309936
rect 216128 309884 216180 309936
rect 196716 309816 196768 309868
rect 239036 309816 239088 309868
rect 240048 309816 240100 309868
rect 32404 309748 32456 309800
rect 61752 309748 61804 309800
rect 66904 309748 66956 309800
rect 177304 309748 177356 309800
rect 188344 309748 188396 309800
rect 216036 309748 216088 309800
rect 292580 309748 292632 309800
rect 240048 309136 240100 309188
rect 358084 309136 358136 309188
rect 192576 309068 192628 309120
rect 226248 309068 226300 309120
rect 226892 309068 226944 309120
rect 228364 308388 228416 308440
rect 244280 308388 244332 308440
rect 63316 307776 63368 307828
rect 67824 307776 67876 307828
rect 198004 307776 198056 307828
rect 276664 307776 276716 307828
rect 64604 307708 64656 307760
rect 66904 307708 66956 307760
rect 199568 307096 199620 307148
rect 214564 307096 214616 307148
rect 170404 307028 170456 307080
rect 187608 307028 187660 307080
rect 200028 307028 200080 307080
rect 240784 307028 240836 307080
rect 298744 307028 298796 307080
rect 345756 307028 345808 307080
rect 158720 306348 158772 306400
rect 195336 306348 195388 306400
rect 215852 306348 215904 306400
rect 289820 306348 289872 306400
rect 3516 306280 3568 306332
rect 36544 306280 36596 306332
rect 208400 306212 208452 306264
rect 223028 306280 223080 306332
rect 223212 305056 223264 305108
rect 360844 305056 360896 305108
rect 53564 304988 53616 305040
rect 66904 304988 66956 305040
rect 158812 304988 158864 305040
rect 194048 304988 194100 305040
rect 198556 304988 198608 305040
rect 233148 304988 233200 305040
rect 233700 304988 233752 305040
rect 234528 304988 234580 305040
rect 447140 304988 447192 305040
rect 63132 304920 63184 304972
rect 66628 304920 66680 304972
rect 218060 304444 218112 304496
rect 219348 304444 219400 304496
rect 221188 304444 221240 304496
rect 191288 304308 191340 304360
rect 207756 304308 207808 304360
rect 222844 304308 222896 304360
rect 234620 304308 234672 304360
rect 159456 304240 159508 304292
rect 164976 304240 165028 304292
rect 183008 304240 183060 304292
rect 195428 304240 195480 304292
rect 206284 304240 206336 304292
rect 247132 304240 247184 304292
rect 234620 303628 234672 303680
rect 435364 303628 435416 303680
rect 160100 302880 160152 302932
rect 169208 302880 169260 302932
rect 247684 302880 247736 302932
rect 251180 302880 251232 302932
rect 188436 302268 188488 302320
rect 189080 302268 189132 302320
rect 159456 302200 159508 302252
rect 258264 302200 258316 302252
rect 53472 302132 53524 302184
rect 66720 302132 66772 302184
rect 158260 301452 158312 301504
rect 188528 301452 188580 301504
rect 201408 301452 201460 301504
rect 274180 301452 274232 301504
rect 60464 300840 60516 300892
rect 66904 300840 66956 300892
rect 185768 300840 185820 300892
rect 186228 300840 186280 300892
rect 214012 300840 214064 300892
rect 216036 300840 216088 300892
rect 411904 300840 411956 300892
rect 244924 300772 244976 300824
rect 247040 300772 247092 300824
rect 48136 300092 48188 300144
rect 66996 300092 67048 300144
rect 189908 299548 189960 299600
rect 244372 299548 244424 299600
rect 198648 299480 198700 299532
rect 284944 299480 284996 299532
rect 204996 299412 205048 299464
rect 223212 299412 223264 299464
rect 64696 298800 64748 298852
rect 66904 298800 66956 298852
rect 188344 298800 188396 298852
rect 201684 298800 201736 298852
rect 158720 298732 158772 298784
rect 244372 298732 244424 298784
rect 265164 298732 265216 298784
rect 324320 298732 324372 298784
rect 341616 298732 341668 298784
rect 244464 298664 244516 298716
rect 228364 298188 228416 298240
rect 279516 298188 279568 298240
rect 267096 298120 267148 298172
rect 324320 298120 324372 298172
rect 41236 298052 41288 298104
rect 66904 298052 66956 298104
rect 233148 297440 233200 297492
rect 309140 297440 309192 297492
rect 158720 297372 158772 297424
rect 175280 297372 175332 297424
rect 177948 297372 178000 297424
rect 204260 297372 204312 297424
rect 209044 297372 209096 297424
rect 215208 297372 215260 297424
rect 389916 297372 389968 297424
rect 175280 297168 175332 297220
rect 176016 297168 176068 297220
rect 160008 296692 160060 296744
rect 209044 296692 209096 296744
rect 191196 296012 191248 296064
rect 206652 296012 206704 296064
rect 216036 296012 216088 296064
rect 194048 295944 194100 295996
rect 236092 295944 236144 295996
rect 304264 295944 304316 295996
rect 358820 295944 358872 295996
rect 242256 295876 242308 295928
rect 243452 295876 243504 295928
rect 49608 295400 49660 295452
rect 66904 295400 66956 295452
rect 243452 295400 243504 295452
rect 303712 295400 303764 295452
rect 304264 295400 304316 295452
rect 17868 295332 17920 295384
rect 67180 295332 67232 295384
rect 226984 295332 227036 295384
rect 227628 295332 227680 295384
rect 308404 295332 308456 295384
rect 59084 295264 59136 295316
rect 66260 295264 66312 295316
rect 158720 295264 158772 295316
rect 187148 295264 187200 295316
rect 159548 294584 159600 294636
rect 178040 294584 178092 294636
rect 295340 294584 295392 294636
rect 382280 294584 382332 294636
rect 267004 294108 267056 294160
rect 269120 294108 269172 294160
rect 222476 294040 222528 294092
rect 222936 294040 222988 294092
rect 252560 294040 252612 294092
rect 187240 293972 187292 294024
rect 262404 293972 262456 294024
rect 19248 293904 19300 293956
rect 66904 293904 66956 293956
rect 194416 293224 194468 293276
rect 204352 293224 204404 293276
rect 270408 293224 270460 293276
rect 278136 293224 278188 293276
rect 315120 293224 315172 293276
rect 362960 293224 363012 293276
rect 158720 292612 158772 292664
rect 194048 292612 194100 292664
rect 204904 292612 204956 292664
rect 262956 292612 263008 292664
rect 3516 292544 3568 292596
rect 18604 292544 18656 292596
rect 158812 292544 158864 292596
rect 220636 292544 220688 292596
rect 234252 292544 234304 292596
rect 268384 292544 268436 292596
rect 60556 292476 60608 292528
rect 66904 292476 66956 292528
rect 283564 291796 283616 291848
rect 322204 291796 322256 291848
rect 389180 291796 389232 291848
rect 407120 291796 407172 291848
rect 158720 291252 158772 291304
rect 248696 291252 248748 291304
rect 174636 291184 174688 291236
rect 204904 291184 204956 291236
rect 241428 291184 241480 291236
rect 401600 291184 401652 291236
rect 52184 291116 52236 291168
rect 56416 291116 56468 291168
rect 220084 291116 220136 291168
rect 222108 291116 222160 291168
rect 166264 290436 166316 290488
rect 211436 290436 211488 290488
rect 159272 290164 159324 290216
rect 162216 290164 162268 290216
rect 224224 289960 224276 290012
rect 445760 289960 445812 290012
rect 211436 289892 211488 289944
rect 218060 289892 218112 289944
rect 222108 289892 222160 289944
rect 254584 289892 254636 289944
rect 56416 289824 56468 289876
rect 66904 289824 66956 289876
rect 158720 289824 158772 289876
rect 224408 289824 224460 289876
rect 56324 289756 56376 289808
rect 66628 289756 66680 289808
rect 165436 289756 165488 289808
rect 166356 289756 166408 289808
rect 191380 289076 191432 289128
rect 210976 289076 211028 289128
rect 240508 289076 240560 289128
rect 258172 289076 258224 289128
rect 280896 289076 280948 289128
rect 291292 289076 291344 289128
rect 369860 289076 369912 289128
rect 235172 288872 235224 288924
rect 236000 288872 236052 288924
rect 210516 288464 210568 288516
rect 210976 288464 211028 288516
rect 247408 288464 247460 288516
rect 158812 288396 158864 288448
rect 231308 288396 231360 288448
rect 165068 287648 165120 287700
rect 182916 287648 182968 287700
rect 247040 287648 247092 287700
rect 260104 287648 260156 287700
rect 287704 287648 287756 287700
rect 347780 287648 347832 287700
rect 190000 287104 190052 287156
rect 216772 287104 216824 287156
rect 220636 287104 220688 287156
rect 248512 287104 248564 287156
rect 158720 287036 158772 287088
rect 166264 287036 166316 287088
rect 187056 287036 187108 287088
rect 223580 287036 223632 287088
rect 224408 287036 224460 287088
rect 245476 287036 245528 287088
rect 158812 286968 158864 287020
rect 189908 286968 189960 287020
rect 158720 286288 158772 286340
rect 164884 286288 164936 286340
rect 214564 286288 214616 286340
rect 225052 286288 225104 286340
rect 255504 286288 255556 286340
rect 273260 286288 273312 286340
rect 194508 285812 194560 285864
rect 200764 285812 200816 285864
rect 191104 285744 191156 285796
rect 204628 285812 204680 285864
rect 201224 285744 201276 285796
rect 46848 285608 46900 285660
rect 62764 285676 62816 285728
rect 66812 285676 66864 285728
rect 182916 285676 182968 285728
rect 187240 285676 187292 285728
rect 203156 285676 203208 285728
rect 204168 285676 204220 285728
rect 204904 285676 204956 285728
rect 206100 285676 206152 285728
rect 213460 285744 213512 285796
rect 213920 285744 213972 285796
rect 215300 285744 215352 285796
rect 216588 285744 216640 285796
rect 230756 285812 230808 285864
rect 235448 285744 235500 285796
rect 237564 285812 237616 285864
rect 238668 285812 238720 285864
rect 225420 285676 225472 285728
rect 226984 285676 227036 285728
rect 233148 285676 233200 285728
rect 233976 285676 234028 285728
rect 236092 285676 236144 285728
rect 237288 285676 237340 285728
rect 244188 285744 244240 285796
rect 238484 285676 238536 285728
rect 251824 285676 251876 285728
rect 218060 285608 218112 285660
rect 218612 285608 218664 285660
rect 237380 285608 237432 285660
rect 238944 285608 238996 285660
rect 239588 285608 239640 285660
rect 267096 285608 267148 285660
rect 181628 284996 181680 285048
rect 190460 284996 190512 285048
rect 191748 284996 191800 285048
rect 234712 284996 234764 285048
rect 244556 284996 244608 285048
rect 164884 284928 164936 284980
rect 185676 284928 185728 284980
rect 195980 284928 196032 284980
rect 235448 284928 235500 284980
rect 245476 284928 245528 284980
rect 258172 284928 258224 284980
rect 63408 284316 63460 284368
rect 66260 284316 66312 284368
rect 158720 284316 158772 284368
rect 162768 284316 162820 284368
rect 166724 284316 166776 284368
rect 169024 284316 169076 284368
rect 199476 284316 199528 284368
rect 210884 284316 210936 284368
rect 61844 284248 61896 284300
rect 66996 284248 67048 284300
rect 181628 283908 181680 283960
rect 201132 283908 201184 283960
rect 201224 283908 201276 283960
rect 162216 283840 162268 283892
rect 244188 283568 244240 283620
rect 260840 283568 260892 283620
rect 282368 283568 282420 283620
rect 352564 283568 352616 283620
rect 246856 283160 246908 283212
rect 247224 283160 247276 283212
rect 249800 283160 249852 283212
rect 260748 282888 260800 282940
rect 319444 282888 319496 282940
rect 245936 282820 245988 282872
rect 278780 282820 278832 282872
rect 298100 282820 298152 282872
rect 298744 282820 298796 282872
rect 158720 282548 158772 282600
rect 162952 282548 163004 282600
rect 163596 282208 163648 282260
rect 189908 282208 189960 282260
rect 249708 282208 249760 282260
rect 254124 282208 254176 282260
rect 414664 282208 414716 282260
rect 431960 282208 432012 282260
rect 162768 282140 162820 282192
rect 193128 282140 193180 282192
rect 197360 282140 197412 282192
rect 254584 282140 254636 282192
rect 279424 282140 279476 282192
rect 302884 282140 302936 282192
rect 414756 282140 414808 282192
rect 64604 281528 64656 281580
rect 66812 281528 66864 281580
rect 281448 281460 281500 281512
rect 297364 281460 297416 281512
rect 245936 280780 245988 280832
rect 280344 280780 280396 280832
rect 281448 280780 281500 280832
rect 293224 280780 293276 280832
rect 421564 280780 421616 280832
rect 158720 280236 158772 280288
rect 169024 280236 169076 280288
rect 34336 280168 34388 280220
rect 67180 280168 67232 280220
rect 163688 280168 163740 280220
rect 197360 280168 197412 280220
rect 158720 280100 158772 280152
rect 171784 280100 171836 280152
rect 245936 280100 245988 280152
rect 255504 280100 255556 280152
rect 162308 279420 162360 279472
rect 176200 279420 176252 279472
rect 181720 279420 181772 279472
rect 196716 279420 196768 279472
rect 195336 279352 195388 279404
rect 197360 279352 197412 279404
rect 158720 278808 158772 278860
rect 162400 278808 162452 278860
rect 64696 278740 64748 278792
rect 66812 278740 66864 278792
rect 249708 278740 249760 278792
rect 309784 278740 309836 278792
rect 195428 278604 195480 278656
rect 197360 278604 197412 278656
rect 180156 278060 180208 278112
rect 185676 278060 185728 278112
rect 156880 277992 156932 278044
rect 195980 277992 196032 278044
rect 254032 277992 254084 278044
rect 374000 277992 374052 278044
rect 376024 277992 376076 278044
rect 245936 277380 245988 277432
rect 254032 277380 254084 277432
rect 169024 277312 169076 277364
rect 197360 277312 197412 277364
rect 158720 277244 158772 277296
rect 182916 277244 182968 277296
rect 4068 276632 4120 276684
rect 43444 276632 43496 276684
rect 183376 276632 183428 276684
rect 191288 276632 191340 276684
rect 268384 276632 268436 276684
rect 281448 276700 281500 276752
rect 322296 276700 322348 276752
rect 282276 276632 282328 276684
rect 296720 276632 296772 276684
rect 308404 276632 308456 276684
rect 395344 276632 395396 276684
rect 52184 276020 52236 276072
rect 66352 276020 66404 276072
rect 245752 275952 245804 276004
rect 263784 275952 263836 276004
rect 245936 275884 245988 275936
rect 253940 275884 253992 275936
rect 169668 275544 169720 275596
rect 172520 275544 172572 275596
rect 263784 275340 263836 275392
rect 353944 275340 353996 275392
rect 163596 275272 163648 275324
rect 185768 275272 185820 275324
rect 253940 275272 253992 275324
rect 417424 275272 417476 275324
rect 158720 274864 158772 274916
rect 161020 274864 161072 274916
rect 191564 274728 191616 274780
rect 195428 274728 195480 274780
rect 180156 274660 180208 274712
rect 197360 274660 197412 274712
rect 34428 274592 34480 274644
rect 65984 274592 66036 274644
rect 158720 274592 158772 274644
rect 170404 274592 170456 274644
rect 279516 274592 279568 274644
rect 358728 274592 358780 274644
rect 167644 273980 167696 274032
rect 182088 273980 182140 274032
rect 176108 273912 176160 273964
rect 195980 273912 196032 273964
rect 262956 273912 263008 273964
rect 370504 273912 370556 273964
rect 63224 273232 63276 273284
rect 66812 273232 66864 273284
rect 182088 273232 182140 273284
rect 197452 273232 197504 273284
rect 245844 273232 245896 273284
rect 253940 273232 253992 273284
rect 358728 273232 358780 273284
rect 363604 273232 363656 273284
rect 180708 273164 180760 273216
rect 197360 273164 197412 273216
rect 245936 273164 245988 273216
rect 254216 273164 254268 273216
rect 276848 273164 276900 273216
rect 277400 273164 277452 273216
rect 376852 273164 376904 273216
rect 251824 272552 251876 272604
rect 262220 272552 262272 272604
rect 188436 272484 188488 272536
rect 199476 272484 199528 272536
rect 245752 272484 245804 272536
rect 251180 272484 251232 272536
rect 254216 272484 254268 272536
rect 313372 272484 313424 272536
rect 358912 272484 358964 272536
rect 50804 271872 50856 271924
rect 66720 271872 66772 271924
rect 56508 271804 56560 271856
rect 66812 271804 66864 271856
rect 282276 271804 282328 271856
rect 385040 271804 385092 271856
rect 245936 271396 245988 271448
rect 248604 271396 248656 271448
rect 158812 271124 158864 271176
rect 167736 271124 167788 271176
rect 274180 271124 274232 271176
rect 293960 271124 294012 271176
rect 168196 270580 168248 270632
rect 197360 270580 197412 270632
rect 158720 270512 158772 270564
rect 196808 270512 196860 270564
rect 245844 270444 245896 270496
rect 262312 270444 262364 270496
rect 262680 270444 262732 270496
rect 244280 270172 244332 270224
rect 248420 270172 248472 270224
rect 169116 269832 169168 269884
rect 178684 269832 178736 269884
rect 159640 269764 159692 269816
rect 170404 269764 170456 269816
rect 172428 269764 172480 269816
rect 191196 269764 191248 269816
rect 262680 269764 262732 269816
rect 291200 269764 291252 269816
rect 178684 269084 178736 269136
rect 197360 269084 197412 269136
rect 158720 269016 158772 269068
rect 187056 269016 187108 269068
rect 178040 268948 178092 269000
rect 178776 268948 178828 269000
rect 197360 268948 197412 269000
rect 253204 268404 253256 268456
rect 264336 268404 264388 268456
rect 167644 268336 167696 268388
rect 178040 268336 178092 268388
rect 246304 268336 246356 268388
rect 323584 268336 323636 268388
rect 355324 268336 355376 268388
rect 580172 268336 580224 268388
rect 191748 268132 191800 268184
rect 197452 268132 197504 268184
rect 64788 267792 64840 267844
rect 66812 267792 66864 267844
rect 245752 267656 245804 267708
rect 265072 267656 265124 267708
rect 166448 267044 166500 267096
rect 175924 267044 175976 267096
rect 179328 267044 179380 267096
rect 188344 267044 188396 267096
rect 3516 266976 3568 267028
rect 14464 266976 14516 267028
rect 57612 266976 57664 267028
rect 66904 266976 66956 267028
rect 173348 266976 173400 267028
rect 184848 266976 184900 267028
rect 265072 266976 265124 267028
rect 302884 266976 302936 267028
rect 304448 266976 304500 267028
rect 367192 266976 367244 267028
rect 188712 266432 188764 266484
rect 195980 266432 196032 266484
rect 184848 266364 184900 266416
rect 197360 266364 197412 266416
rect 245660 265820 245712 265872
rect 249892 265820 249944 265872
rect 173348 265616 173400 265668
rect 181628 265616 181680 265668
rect 255320 265616 255372 265668
rect 371884 265616 371936 265668
rect 53472 264936 53524 264988
rect 66904 264936 66956 264988
rect 158720 264936 158772 264988
rect 180340 264936 180392 264988
rect 245844 264868 245896 264920
rect 266360 264868 266412 264920
rect 268384 264256 268436 264308
rect 316040 264256 316092 264308
rect 266360 264188 266412 264240
rect 267648 264188 267700 264240
rect 298744 264188 298796 264240
rect 304264 264188 304316 264240
rect 450544 264188 450596 264240
rect 188620 263644 188672 263696
rect 197452 263644 197504 263696
rect 59084 263576 59136 263628
rect 59268 263576 59320 263628
rect 66444 263576 66496 263628
rect 187056 263576 187108 263628
rect 197360 263576 197412 263628
rect 244096 263372 244148 263424
rect 245660 263372 245712 263424
rect 67548 262896 67600 262948
rect 68284 262896 68336 262948
rect 280896 262896 280948 262948
rect 308404 262896 308456 262948
rect 160928 262828 160980 262880
rect 165068 262828 165120 262880
rect 165436 262828 165488 262880
rect 180156 262828 180208 262880
rect 262772 262828 262824 262880
rect 378784 262828 378836 262880
rect 57704 262624 57756 262676
rect 59268 262624 59320 262676
rect 158720 262624 158772 262676
rect 160836 262624 160888 262676
rect 181628 262624 181680 262676
rect 184388 262624 184440 262676
rect 59268 262216 59320 262268
rect 66904 262216 66956 262268
rect 195336 262216 195388 262268
rect 198004 262216 198056 262268
rect 245936 262216 245988 262268
rect 255320 262216 255372 262268
rect 186320 262148 186372 262200
rect 186964 262148 187016 262200
rect 197360 262148 197412 262200
rect 185768 262080 185820 262132
rect 195428 262080 195480 262132
rect 158996 261536 159048 261588
rect 159456 261536 159508 261588
rect 170496 261536 170548 261588
rect 265624 261536 265676 261588
rect 302240 261536 302292 261588
rect 43444 261468 43496 261520
rect 65892 261468 65944 261520
rect 66536 261468 66588 261520
rect 161020 261468 161072 261520
rect 175924 261468 175976 261520
rect 299572 261468 299624 261520
rect 354036 261468 354088 261520
rect 245844 260924 245896 260976
rect 248420 260924 248472 260976
rect 248696 260924 248748 260976
rect 56508 260856 56560 260908
rect 66352 260856 66404 260908
rect 162768 260788 162820 260840
rect 182088 260788 182140 260840
rect 182916 260788 182968 260840
rect 182824 260720 182876 260772
rect 288348 260108 288400 260160
rect 375380 260108 375432 260160
rect 245752 259836 245804 259888
rect 249892 259836 249944 259888
rect 194508 259768 194560 259820
rect 196072 259768 196124 259820
rect 197268 259768 197320 259820
rect 170956 259428 171008 259480
rect 171140 259428 171192 259480
rect 183008 259428 183060 259480
rect 197360 259428 197412 259480
rect 246396 259428 246448 259480
rect 287152 259428 287204 259480
rect 288348 259428 288400 259480
rect 186228 259360 186280 259412
rect 187424 259360 187476 259412
rect 245752 259360 245804 259412
rect 265072 259360 265124 259412
rect 186228 259224 186280 259276
rect 190000 259224 190052 259276
rect 265072 258748 265124 258800
rect 292580 258748 292632 258800
rect 368480 258748 368532 258800
rect 164976 258680 165028 258732
rect 181720 258680 181772 258732
rect 288624 258680 288676 258732
rect 372712 258680 372764 258732
rect 187424 258136 187476 258188
rect 197360 258136 197412 258188
rect 53748 258000 53800 258052
rect 57244 258000 57296 258052
rect 66260 258068 66312 258120
rect 158812 258068 158864 258120
rect 186228 258068 186280 258120
rect 244556 258068 244608 258120
rect 288624 258068 288676 258120
rect 158720 258000 158772 258052
rect 163688 258000 163740 258052
rect 172336 258000 172388 258052
rect 173440 258000 173492 258052
rect 245752 258000 245804 258052
rect 256792 258000 256844 258052
rect 184296 257320 184348 257372
rect 199384 257320 199436 257372
rect 256792 257320 256844 257372
rect 295432 257320 295484 257372
rect 308404 257320 308456 257372
rect 383016 257320 383068 257372
rect 272524 256844 272576 256896
rect 279516 256844 279568 256896
rect 61844 256708 61896 256760
rect 66812 256708 66864 256760
rect 164148 256708 164200 256760
rect 189080 256708 189132 256760
rect 196808 256708 196860 256760
rect 197268 256708 197320 256760
rect 194416 256640 194468 256692
rect 197360 256640 197412 256692
rect 169024 255960 169076 256012
rect 194416 255960 194468 256012
rect 245660 255960 245712 256012
rect 302240 255960 302292 256012
rect 360384 255960 360436 256012
rect 245752 255348 245804 255400
rect 249984 255348 250036 255400
rect 251088 255348 251140 255400
rect 158536 255280 158588 255332
rect 177396 255280 177448 255332
rect 245844 255212 245896 255264
rect 252836 255212 252888 255264
rect 156696 254600 156748 254652
rect 170588 254600 170640 254652
rect 180340 254600 180392 254652
rect 196808 254600 196860 254652
rect 252836 254600 252888 254652
rect 334624 254600 334676 254652
rect 158260 254532 158312 254584
rect 191104 254532 191156 254584
rect 251088 254532 251140 254584
rect 358176 254532 358228 254584
rect 2780 254192 2832 254244
rect 4804 254192 4856 254244
rect 54944 253920 54996 253972
rect 66628 253920 66680 253972
rect 194416 253920 194468 253972
rect 197360 253920 197412 253972
rect 246028 253852 246080 253904
rect 262404 253852 262456 253904
rect 262680 253852 262732 253904
rect 245936 253784 245988 253836
rect 258264 253784 258316 253836
rect 259276 253784 259328 253836
rect 259276 253240 259328 253292
rect 307760 253240 307812 253292
rect 371332 253240 371384 253292
rect 52276 253172 52328 253224
rect 60188 253172 60240 253224
rect 67548 253172 67600 253224
rect 68376 253172 68428 253224
rect 158720 253172 158772 253224
rect 179420 253172 179472 253224
rect 185584 253172 185636 253224
rect 186136 253172 186188 253224
rect 197360 253172 197412 253224
rect 262680 253172 262732 253224
rect 306380 253172 306432 253224
rect 369952 253172 370004 253224
rect 60188 252560 60240 252612
rect 60556 252560 60608 252612
rect 66812 252560 66864 252612
rect 158720 252560 158772 252612
rect 166356 252560 166408 252612
rect 192944 252560 192996 252612
rect 197360 252560 197412 252612
rect 179420 252492 179472 252544
rect 195796 252492 195848 252544
rect 245936 252492 245988 252544
rect 261024 252492 261076 252544
rect 262128 252492 262180 252544
rect 156788 252424 156840 252476
rect 163780 252424 163832 252476
rect 180340 251812 180392 251864
rect 187056 251812 187108 251864
rect 245936 251812 245988 251864
rect 251364 251812 251416 251864
rect 252376 251812 252428 251864
rect 262128 251812 262180 251864
rect 322204 251812 322256 251864
rect 195796 251608 195848 251660
rect 197360 251608 197412 251660
rect 158904 251200 158956 251252
rect 180340 251200 180392 251252
rect 180708 251200 180760 251252
rect 252376 251200 252428 251252
rect 356704 251200 356756 251252
rect 245844 251132 245896 251184
rect 259460 251132 259512 251184
rect 260748 251132 260800 251184
rect 331956 251132 332008 251184
rect 334716 251132 334768 251184
rect 177304 250928 177356 250980
rect 180064 250928 180116 250980
rect 278228 250520 278280 250572
rect 301044 250520 301096 250572
rect 63408 250452 63460 250504
rect 67732 250452 67784 250504
rect 162492 250452 162544 250504
rect 173256 250452 173308 250504
rect 260748 250452 260800 250504
rect 310612 250452 310664 250504
rect 365812 250452 365864 250504
rect 180156 249908 180208 249960
rect 197360 249840 197412 249892
rect 64512 249772 64564 249824
rect 66812 249772 66864 249824
rect 158720 249772 158772 249824
rect 173440 249772 173492 249824
rect 178776 249772 178828 249824
rect 197452 249772 197504 249824
rect 186228 249704 186280 249756
rect 188528 249704 188580 249756
rect 245936 249704 245988 249756
rect 248696 249704 248748 249756
rect 264244 249092 264296 249144
rect 348424 249092 348476 249144
rect 167736 249024 167788 249076
rect 187608 249024 187660 249076
rect 299388 249024 299440 249076
rect 582840 249024 582892 249076
rect 196716 248684 196768 248736
rect 197820 248684 197872 248736
rect 158812 248412 158864 248464
rect 182824 248412 182876 248464
rect 187608 248412 187660 248464
rect 197360 248412 197412 248464
rect 299388 248344 299440 248396
rect 300216 248344 300268 248396
rect 162400 247732 162452 247784
rect 179420 247732 179472 247784
rect 168472 247664 168524 247716
rect 188712 247664 188764 247716
rect 245660 247664 245712 247716
rect 300216 247664 300268 247716
rect 195612 247120 195664 247172
rect 196716 247120 196768 247172
rect 185584 247052 185636 247104
rect 197360 247052 197412 247104
rect 245936 247052 245988 247104
rect 251272 247052 251324 247104
rect 377404 247052 377456 247104
rect 62028 246984 62080 247036
rect 66812 246984 66864 247036
rect 179420 246304 179472 246356
rect 196716 246304 196768 246356
rect 317236 246304 317288 246356
rect 331220 246304 331272 246356
rect 244556 245692 244608 245744
rect 281540 245692 281592 245744
rect 283564 245692 283616 245744
rect 181444 245624 181496 245676
rect 184296 245624 184348 245676
rect 184756 245624 184808 245676
rect 191840 245624 191892 245676
rect 198832 245624 198884 245676
rect 245844 245624 245896 245676
rect 255412 245624 255464 245676
rect 260104 245624 260156 245676
rect 316040 245624 316092 245676
rect 317236 245624 317288 245676
rect 48228 245556 48280 245608
rect 66812 245556 66864 245608
rect 328368 244944 328420 244996
rect 363144 244944 363196 244996
rect 161572 244876 161624 244928
rect 189816 244876 189868 244928
rect 189908 244876 189960 244928
rect 197728 244876 197780 244928
rect 252376 244876 252428 244928
rect 340236 244876 340288 244928
rect 356796 244876 356848 244928
rect 436284 244876 436336 244928
rect 158720 244264 158772 244316
rect 193864 244264 193916 244316
rect 245936 244264 245988 244316
rect 327172 244264 327224 244316
rect 328368 244264 328420 244316
rect 59176 244196 59228 244248
rect 66812 244196 66864 244248
rect 189816 244196 189868 244248
rect 193036 244196 193088 244248
rect 197360 244196 197412 244248
rect 157984 243516 158036 243568
rect 171324 243516 171376 243568
rect 171692 243516 171744 243568
rect 171784 243516 171836 243568
rect 173348 243516 173400 243568
rect 177488 243516 177540 243568
rect 192668 243516 192720 243568
rect 259276 243516 259328 243568
rect 342904 243516 342956 243568
rect 158720 242904 158772 242956
rect 184296 242904 184348 242956
rect 245844 242904 245896 242956
rect 258264 242904 258316 242956
rect 259276 242904 259328 242956
rect 260748 242904 260800 242956
rect 302976 242904 303028 242956
rect 155316 242020 155368 242072
rect 183100 242156 183152 242208
rect 311992 242156 312044 242208
rect 345664 242156 345716 242208
rect 246396 241544 246448 241596
rect 247224 241544 247276 241596
rect 311992 241544 312044 241596
rect 156972 241476 157024 241528
rect 186228 241476 186280 241528
rect 197360 241476 197412 241528
rect 245752 241476 245804 241528
rect 463700 241476 463752 241528
rect 57796 241408 57848 241460
rect 58624 241408 58676 241460
rect 57704 241340 57756 241392
rect 83326 241408 83378 241460
rect 156374 241340 156426 241392
rect 160192 241340 160244 241392
rect 3516 241068 3568 241120
rect 7564 241068 7616 241120
rect 166264 240796 166316 240848
rect 200120 240796 200172 240848
rect 300124 240796 300176 240848
rect 309876 240796 309928 240848
rect 18604 240728 18656 240780
rect 57796 240728 57848 240780
rect 66076 240728 66128 240780
rect 86224 240728 86276 240780
rect 128820 240728 128872 240780
rect 167828 240728 167880 240780
rect 260196 240728 260248 240780
rect 420184 240728 420236 240780
rect 155500 240388 155552 240440
rect 156696 240388 156748 240440
rect 199660 240388 199712 240440
rect 199568 240320 199620 240372
rect 103612 240184 103664 240236
rect 104808 240184 104860 240236
rect 67732 240116 67784 240168
rect 68468 240116 68520 240168
rect 77300 240116 77352 240168
rect 77852 240116 77904 240168
rect 82912 240116 82964 240168
rect 83740 240116 83792 240168
rect 91100 240116 91152 240168
rect 91836 240116 91888 240168
rect 107660 240116 107712 240168
rect 108580 240116 108632 240168
rect 115204 240116 115256 240168
rect 170588 240116 170640 240168
rect 201224 240116 201276 240168
rect 202328 240116 202380 240168
rect 244096 240252 244148 240304
rect 243912 240184 243964 240236
rect 289912 240184 289964 240236
rect 298836 240184 298888 240236
rect 203984 240116 204036 240168
rect 208400 240116 208452 240168
rect 225052 240116 225104 240168
rect 226800 240116 226852 240168
rect 228364 240116 228416 240168
rect 231032 240116 231084 240168
rect 241888 240116 241940 240168
rect 247132 240116 247184 240168
rect 69572 240048 69624 240100
rect 72516 240048 72568 240100
rect 75184 240048 75236 240100
rect 75920 240048 75972 240100
rect 82728 240048 82780 240100
rect 83556 240048 83608 240100
rect 85120 240048 85172 240100
rect 92572 240048 92624 240100
rect 117872 240048 117924 240100
rect 118608 240048 118660 240100
rect 119344 240048 119396 240100
rect 119988 240048 120040 240100
rect 128636 240048 128688 240100
rect 129648 240048 129700 240100
rect 131856 240048 131908 240100
rect 132408 240048 132460 240100
rect 133328 240048 133380 240100
rect 133788 240048 133840 240100
rect 135352 240048 135404 240100
rect 136548 240048 136600 240100
rect 138480 240048 138532 240100
rect 139308 240048 139360 240100
rect 142896 240048 142948 240100
rect 143356 240048 143408 240100
rect 145656 240048 145708 240100
rect 146116 240048 146168 240100
rect 153476 240048 153528 240100
rect 154488 240048 154540 240100
rect 228732 240048 228784 240100
rect 243912 240048 243964 240100
rect 67456 239980 67508 240032
rect 69756 239980 69808 240032
rect 113640 239980 113692 240032
rect 118516 239980 118568 240032
rect 142252 239980 142304 240032
rect 142988 239980 143040 240032
rect 237380 239980 237432 240032
rect 238116 239980 238168 240032
rect 244556 239980 244608 240032
rect 82176 239776 82228 239828
rect 82728 239776 82780 239828
rect 70308 239436 70360 239488
rect 97264 239436 97316 239488
rect 97448 239436 97500 239488
rect 88800 239368 88852 239420
rect 89536 239368 89588 239420
rect 101956 239368 102008 239420
rect 102692 239368 102744 239420
rect 122288 239436 122340 239488
rect 220820 239436 220872 239488
rect 305092 239436 305144 239488
rect 322940 239436 322992 239488
rect 214196 239368 214248 239420
rect 260748 239368 260800 239420
rect 273904 239368 273956 239420
rect 313924 239368 313976 239420
rect 345664 239368 345716 239420
rect 116584 239300 116636 239352
rect 117136 239300 117188 239352
rect 120816 239300 120868 239352
rect 121368 239300 121420 239352
rect 143540 239300 143592 239352
rect 144276 239300 144328 239352
rect 80704 239232 80756 239284
rect 81348 239232 81400 239284
rect 105544 239232 105596 239284
rect 106188 239232 106240 239284
rect 131212 239232 131264 239284
rect 131948 239232 132000 239284
rect 138020 239232 138072 239284
rect 138572 239232 138624 239284
rect 104072 239164 104124 239216
rect 104808 239164 104860 239216
rect 219440 238756 219492 238808
rect 238024 238756 238076 238808
rect 73160 238688 73212 238740
rect 202604 238688 202656 238740
rect 240324 238688 240376 238740
rect 252468 238688 252520 238740
rect 55036 238620 55088 238672
rect 75184 238620 75236 238672
rect 118516 238620 118568 238672
rect 222292 238620 222344 238672
rect 242072 238620 242124 238672
rect 252652 238620 252704 238672
rect 224868 238076 224920 238128
rect 227536 238076 227588 238128
rect 252468 238076 252520 238128
rect 262864 238076 262916 238128
rect 260104 238008 260156 238060
rect 280804 238008 280856 238060
rect 295248 238008 295300 238060
rect 384304 238008 384356 238060
rect 223396 237804 223448 237856
rect 229376 237804 229428 237856
rect 229836 237668 229888 237720
rect 236828 237668 236880 237720
rect 240048 237464 240100 237516
rect 242716 237464 242768 237516
rect 202144 237396 202196 237448
rect 202604 237396 202656 237448
rect 202880 237396 202932 237448
rect 204996 237396 205048 237448
rect 207112 237396 207164 237448
rect 207940 237396 207992 237448
rect 209688 237396 209740 237448
rect 210332 237396 210384 237448
rect 230204 237396 230256 237448
rect 232504 237396 232556 237448
rect 239220 237396 239272 237448
rect 240968 237396 241020 237448
rect 125600 237328 125652 237380
rect 181536 237328 181588 237380
rect 182088 237328 182140 237380
rect 200120 237328 200172 237380
rect 223764 237328 223816 237380
rect 241244 237328 241296 237380
rect 287704 237328 287756 237380
rect 149060 237260 149112 237312
rect 162216 237260 162268 237312
rect 196808 237260 196860 237312
rect 202788 237260 202840 237312
rect 194324 236716 194376 236768
rect 199384 236716 199436 236768
rect 229100 236716 229152 236768
rect 242256 236716 242308 236768
rect 187424 236648 187476 236700
rect 195244 236648 195296 236700
rect 199936 236648 199988 236700
rect 200764 236648 200816 236700
rect 208308 236648 208360 236700
rect 239496 236648 239548 236700
rect 260932 236648 260984 236700
rect 410524 236648 410576 236700
rect 4804 235968 4856 236020
rect 93860 235968 93912 236020
rect 94504 235968 94556 236020
rect 240784 235968 240836 236020
rect 241244 235968 241296 236020
rect 61752 235900 61804 235952
rect 130108 235900 130160 235952
rect 196716 235900 196768 235952
rect 220268 235900 220320 235952
rect 232044 235900 232096 235952
rect 268384 235900 268436 235952
rect 50896 235832 50948 235884
rect 77392 235832 77444 235884
rect 114652 235832 114704 235884
rect 152464 235832 152516 235884
rect 152740 235832 152792 235884
rect 185676 235832 185728 235884
rect 206836 235832 206888 235884
rect 152372 235696 152424 235748
rect 155960 235696 156012 235748
rect 222936 235288 222988 235340
rect 232044 235288 232096 235340
rect 131212 235220 131264 235272
rect 184756 235220 184808 235272
rect 185584 235220 185636 235272
rect 205640 235220 205692 235272
rect 224224 235220 224276 235272
rect 57612 234540 57664 234592
rect 128728 234540 128780 234592
rect 150440 234540 150492 234592
rect 168196 234608 168248 234660
rect 174544 234608 174596 234660
rect 186964 234608 187016 234660
rect 188436 234608 188488 234660
rect 206376 234608 206428 234660
rect 206836 234608 206888 234660
rect 231584 234608 231636 234660
rect 234068 234608 234120 234660
rect 240876 234608 240928 234660
rect 243268 234608 243320 234660
rect 152096 234472 152148 234524
rect 155684 234472 155736 234524
rect 191472 234132 191524 234184
rect 192576 234132 192628 234184
rect 242256 233996 242308 234048
rect 265624 233996 265676 234048
rect 133144 233928 133196 233980
rect 152924 233928 152976 233980
rect 176200 233928 176252 233980
rect 187056 233928 187108 233980
rect 195244 233928 195296 233980
rect 210608 233928 210660 233980
rect 215300 233928 215352 233980
rect 247224 233928 247276 233980
rect 111892 233860 111944 233912
rect 139584 233860 139636 233912
rect 155224 233860 155276 233912
rect 176660 233860 176712 233912
rect 184296 233860 184348 233912
rect 236000 233860 236052 233912
rect 256700 233860 256752 233912
rect 322296 233860 322348 233912
rect 14464 233180 14516 233232
rect 92664 233180 92716 233232
rect 143632 233180 143684 233232
rect 156880 233180 156932 233232
rect 192944 233180 192996 233232
rect 270500 233180 270552 233232
rect 280804 233248 280856 233300
rect 155868 233112 155920 233164
rect 158260 233112 158312 233164
rect 190460 233112 190512 233164
rect 205364 233112 205416 233164
rect 211804 233112 211856 233164
rect 212816 233112 212868 233164
rect 236000 233112 236052 233164
rect 236644 233112 236696 233164
rect 244464 233112 244516 233164
rect 92664 232704 92716 232756
rect 93124 232704 93176 232756
rect 156604 232704 156656 232756
rect 159180 232704 159232 232756
rect 140872 232568 140924 232620
rect 155868 232568 155920 232620
rect 44088 232500 44140 232552
rect 143540 232500 143592 232552
rect 157340 232500 157392 232552
rect 187424 232500 187476 232552
rect 191104 232500 191156 232552
rect 216036 232500 216088 232552
rect 227720 232500 227772 232552
rect 282184 232500 282236 232552
rect 465080 232500 465132 232552
rect 158720 231820 158772 231872
rect 184296 231820 184348 231872
rect 69756 231752 69808 231804
rect 156972 231752 157024 231804
rect 124312 231684 124364 231736
rect 198740 231684 198792 231736
rect 205640 231548 205692 231600
rect 206468 231548 206520 231600
rect 198740 231140 198792 231192
rect 199844 231140 199896 231192
rect 230480 231140 230532 231192
rect 204076 231072 204128 231124
rect 224224 231072 224276 231124
rect 228180 231072 228232 231124
rect 398932 231072 398984 231124
rect 208400 230936 208452 230988
rect 209228 230936 209280 230988
rect 270408 230460 270460 230512
rect 282184 230460 282236 230512
rect 143356 230392 143408 230444
rect 231584 230392 231636 230444
rect 139308 230324 139360 230376
rect 165436 230324 165488 230376
rect 166356 230324 166408 230376
rect 195244 230324 195296 230376
rect 202328 230324 202380 230376
rect 207572 230324 207624 230376
rect 222292 230324 222344 230376
rect 83648 229780 83700 229832
rect 141424 229780 141476 229832
rect 64696 229712 64748 229764
rect 137928 229712 137980 229764
rect 165436 229576 165488 229628
rect 166264 229576 166316 229628
rect 243544 229100 243596 229152
rect 248512 229100 248564 229152
rect 117320 229032 117372 229084
rect 224316 229032 224368 229084
rect 94504 228964 94556 229016
rect 174636 228964 174688 229016
rect 175924 228964 175976 229016
rect 242900 228964 242952 229016
rect 242900 228556 242952 228608
rect 243912 228556 243964 228608
rect 327080 228352 327132 228404
rect 403072 228352 403124 228404
rect 242808 227740 242860 227792
rect 258264 227740 258316 227792
rect 258724 227740 258776 227792
rect 137928 227672 137980 227724
rect 173164 227672 173216 227724
rect 181720 227672 181772 227724
rect 222844 227672 222896 227724
rect 224316 227060 224368 227112
rect 240692 227060 240744 227112
rect 54944 226992 54996 227044
rect 194324 226992 194376 227044
rect 217140 226992 217192 227044
rect 226340 226992 226392 227044
rect 239496 226992 239548 227044
rect 298284 226992 298336 227044
rect 204904 226312 204956 226364
rect 209688 226312 209740 226364
rect 71780 226244 71832 226296
rect 158076 226244 158128 226296
rect 187056 226244 187108 226296
rect 213644 226244 213696 226296
rect 139400 226176 139452 226228
rect 222936 226176 222988 226228
rect 240692 225632 240744 225684
rect 284484 225632 284536 225684
rect 68284 225564 68336 225616
rect 104164 225564 104216 225616
rect 219900 225564 219952 225616
rect 220360 225564 220412 225616
rect 267004 225564 267056 225616
rect 292488 225564 292540 225616
rect 307116 225564 307168 225616
rect 213184 225428 213236 225480
rect 213644 225428 213696 225480
rect 284484 224952 284536 225004
rect 285680 224952 285732 225004
rect 111708 224884 111760 224936
rect 192944 224884 192996 224936
rect 221464 224884 221516 224936
rect 276020 224884 276072 224936
rect 246304 224612 246356 224664
rect 247224 224612 247276 224664
rect 95332 224204 95384 224256
rect 157340 224204 157392 224256
rect 178040 224204 178092 224256
rect 193956 224204 194008 224256
rect 223488 224204 223540 224256
rect 276020 224204 276072 224256
rect 285680 224204 285732 224256
rect 158168 224136 158220 224188
rect 79968 223524 80020 223576
rect 211896 223524 211948 223576
rect 124220 222844 124272 222896
rect 186320 222844 186372 222896
rect 201500 222844 201552 222896
rect 302332 222844 302384 222896
rect 338764 222844 338816 222896
rect 65984 222096 66036 222148
rect 159640 222096 159692 222148
rect 194324 222096 194376 222148
rect 213276 222096 213328 222148
rect 223488 222096 223540 222148
rect 248604 222096 248656 222148
rect 106280 222028 106332 222080
rect 171784 222028 171836 222080
rect 203064 221824 203116 221876
rect 203616 221824 203668 221876
rect 167000 221416 167052 221468
rect 167736 221416 167788 221468
rect 203064 221416 203116 221468
rect 208400 221416 208452 221468
rect 228732 221416 228784 221468
rect 260748 221416 260800 221468
rect 387064 221416 387116 221468
rect 104900 220736 104952 220788
rect 180248 220736 180300 220788
rect 186320 220736 186372 220788
rect 220084 220736 220136 220788
rect 227260 220736 227312 220788
rect 260748 220736 260800 220788
rect 195704 220668 195756 220720
rect 199476 220668 199528 220720
rect 127256 220056 127308 220108
rect 194416 220056 194468 220108
rect 260748 220056 260800 220108
rect 276940 220056 276992 220108
rect 278136 220056 278188 220108
rect 294052 220056 294104 220108
rect 200028 219444 200080 219496
rect 201500 219444 201552 219496
rect 217324 219444 217376 219496
rect 221372 219376 221424 219428
rect 258080 219376 258132 219428
rect 259276 219376 259328 219428
rect 194416 219308 194468 219360
rect 227260 219308 227312 219360
rect 236460 219308 236512 219360
rect 269764 219308 269816 219360
rect 106188 218764 106240 218816
rect 133144 218764 133196 218816
rect 136640 218764 136692 218816
rect 182272 218764 182324 218816
rect 269764 218764 269816 218816
rect 304264 218764 304316 218816
rect 82728 218696 82780 218748
rect 142804 218696 142856 218748
rect 207664 218696 207716 218748
rect 222108 218696 222160 218748
rect 259276 218696 259328 218748
rect 414020 218696 414072 218748
rect 143448 218016 143500 218068
rect 195244 218016 195296 218068
rect 126980 217948 127032 218000
rect 208400 217948 208452 218000
rect 184480 217880 184532 217932
rect 225236 217880 225288 217932
rect 83556 217268 83608 217320
rect 177856 217132 177908 217184
rect 178776 217132 178828 217184
rect 234988 216656 235040 216708
rect 394056 216656 394108 216708
rect 107660 216588 107712 216640
rect 220360 216588 220412 216640
rect 132408 216520 132460 216572
rect 181444 216520 181496 216572
rect 220268 215976 220320 216028
rect 233332 215976 233384 216028
rect 232596 215908 232648 215960
rect 321560 215908 321612 215960
rect 3332 215228 3384 215280
rect 35164 215228 35216 215280
rect 87144 215228 87196 215280
rect 186964 215228 187016 215280
rect 219348 215228 219400 215280
rect 267740 215228 267792 215280
rect 269028 215228 269080 215280
rect 201132 214616 201184 214668
rect 206468 214616 206520 214668
rect 182272 214548 182324 214600
rect 223488 214548 223540 214600
rect 269028 214548 269080 214600
rect 287244 214548 287296 214600
rect 317328 214548 317380 214600
rect 447232 214548 447284 214600
rect 97264 213868 97316 213920
rect 202236 213868 202288 213920
rect 223488 213868 223540 213920
rect 245660 213868 245712 213920
rect 118700 213800 118752 213852
rect 169024 213800 169076 213852
rect 205640 213256 205692 213308
rect 215300 213256 215352 213308
rect 202420 213188 202472 213240
rect 229744 213188 229796 213240
rect 249708 212508 249760 212560
rect 456800 212508 456852 212560
rect 124128 212440 124180 212492
rect 225144 212440 225196 212492
rect 225604 212440 225656 212492
rect 215116 212372 215168 212424
rect 215668 212372 215720 212424
rect 263600 211828 263652 211880
rect 283564 211828 283616 211880
rect 70400 211760 70452 211812
rect 215116 211760 215168 211812
rect 233516 211760 233568 211812
rect 380164 211760 380216 211812
rect 77300 211080 77352 211132
rect 215300 211080 215352 211132
rect 158168 211012 158220 211064
rect 248696 211012 248748 211064
rect 238852 209788 238904 209840
rect 239772 209788 239824 209840
rect 309968 209788 310020 209840
rect 104164 209720 104216 209772
rect 226340 209720 226392 209772
rect 90916 209652 90968 209704
rect 189724 209652 189776 209704
rect 204720 209040 204772 209092
rect 234436 209040 234488 209092
rect 267832 209040 267884 209092
rect 445852 209040 445904 209092
rect 89720 208972 89772 209024
rect 90916 208972 90968 209024
rect 226340 208360 226392 208412
rect 227076 208360 227128 208412
rect 48136 208292 48188 208344
rect 240232 208292 240284 208344
rect 240876 208292 240928 208344
rect 100668 208224 100720 208276
rect 181628 208224 181680 208276
rect 99380 207748 99432 207800
rect 100668 207748 100720 207800
rect 262864 207680 262916 207732
rect 278136 207680 278188 207732
rect 229744 207612 229796 207664
rect 272616 207612 272668 207664
rect 181628 207000 181680 207052
rect 228364 207000 228416 207052
rect 114468 206932 114520 206984
rect 247224 206932 247276 206984
rect 133788 206864 133840 206916
rect 227720 206864 227772 206916
rect 247132 206864 247184 206916
rect 86960 205572 87012 205624
rect 214472 205572 214524 205624
rect 142804 205504 142856 205556
rect 249892 205504 249944 205556
rect 51080 204892 51132 204944
rect 137284 204892 137336 204944
rect 225696 204892 225748 204944
rect 284392 204892 284444 204944
rect 214472 204280 214524 204332
rect 224316 204280 224368 204332
rect 91100 204212 91152 204264
rect 212448 204212 212500 204264
rect 100760 204144 100812 204196
rect 212816 204144 212868 204196
rect 213828 204144 213880 204196
rect 213828 203600 213880 203652
rect 238760 203600 238812 203652
rect 212448 203532 212500 203584
rect 272524 203532 272576 203584
rect 3056 202784 3108 202836
rect 51080 202784 51132 202836
rect 59268 202784 59320 202836
rect 211804 202784 211856 202836
rect 212172 202784 212224 202836
rect 72516 202716 72568 202768
rect 181628 202716 181680 202768
rect 213184 202172 213236 202224
rect 237380 202172 237432 202224
rect 197176 202104 197228 202156
rect 370596 202104 370648 202156
rect 288716 201492 288768 201544
rect 437480 201492 437532 201544
rect 67640 200812 67692 200864
rect 169760 200812 169812 200864
rect 193128 200812 193180 200864
rect 203616 200812 203668 200864
rect 126888 200744 126940 200796
rect 234620 200744 234672 200796
rect 255320 200744 255372 200796
rect 205548 200132 205600 200184
rect 215852 200132 215904 200184
rect 169760 200064 169812 200116
rect 206468 200064 206520 200116
rect 232596 200132 232648 200184
rect 147588 199452 147640 199504
rect 194324 199452 194376 199504
rect 63408 199384 63460 199436
rect 168380 199384 168432 199436
rect 217324 199384 217376 199436
rect 307852 199384 307904 199436
rect 53472 198636 53524 198688
rect 160744 198636 160796 198688
rect 168380 198636 168432 198688
rect 201500 198636 201552 198688
rect 120080 198568 120132 198620
rect 156788 198568 156840 198620
rect 167000 198024 167052 198076
rect 213276 198024 213328 198076
rect 215116 198024 215168 198076
rect 241612 198024 241664 198076
rect 202144 197956 202196 198008
rect 295524 197956 295576 198008
rect 118608 197276 118660 197328
rect 170496 197276 170548 197328
rect 188528 196664 188580 196716
rect 196808 196664 196860 196716
rect 201316 196664 201368 196716
rect 240140 196664 240192 196716
rect 255964 196664 256016 196716
rect 285864 196664 285916 196716
rect 112996 196596 113048 196648
rect 185584 196596 185636 196648
rect 195796 196596 195848 196648
rect 279608 196596 279660 196648
rect 191932 195916 191984 195968
rect 255412 195916 255464 195968
rect 158720 195848 158772 195900
rect 159364 195848 159416 195900
rect 193128 195848 193180 195900
rect 194324 195848 194376 195900
rect 252744 195848 252796 195900
rect 318156 195304 318208 195356
rect 326344 195304 326396 195356
rect 133144 195236 133196 195288
rect 158720 195236 158772 195288
rect 272616 195236 272668 195288
rect 292672 195236 292724 195288
rect 325608 195236 325660 195288
rect 349896 195236 349948 195288
rect 17224 195032 17276 195084
rect 17868 195032 17920 195084
rect 17868 194556 17920 194608
rect 181536 194556 181588 194608
rect 200764 194488 200816 194540
rect 204260 194488 204312 194540
rect 50804 193876 50856 193928
rect 139400 193876 139452 193928
rect 206284 193876 206336 193928
rect 281632 193876 281684 193928
rect 89628 193808 89680 193860
rect 209228 193808 209280 193860
rect 267004 193808 267056 193860
rect 276756 193808 276808 193860
rect 286968 193808 287020 193860
rect 294144 193808 294196 193860
rect 93124 193128 93176 193180
rect 167000 193128 167052 193180
rect 139400 193060 139452 193112
rect 198740 193060 198792 193112
rect 198740 192516 198792 192568
rect 223488 192516 223540 192568
rect 224316 192516 224368 192568
rect 245752 192516 245804 192568
rect 276940 192516 276992 192568
rect 298192 192516 298244 192568
rect 204260 192448 204312 192500
rect 238116 192448 238168 192500
rect 253204 192448 253256 192500
rect 443092 192448 443144 192500
rect 33784 191768 33836 191820
rect 34336 191768 34388 191820
rect 165528 191768 165580 191820
rect 196716 191768 196768 191820
rect 199476 191156 199528 191208
rect 236000 191156 236052 191208
rect 198004 191088 198056 191140
rect 290096 191088 290148 191140
rect 177304 189796 177356 189848
rect 202144 189796 202196 189848
rect 224224 189796 224276 189848
rect 242992 189796 243044 189848
rect 155868 189728 155920 189780
rect 164884 189728 164936 189780
rect 193864 189728 193916 189780
rect 231124 189728 231176 189780
rect 110328 189048 110380 189100
rect 175924 189048 175976 189100
rect 3516 188980 3568 189032
rect 29644 188980 29696 189032
rect 180708 188300 180760 188352
rect 204904 188300 204956 188352
rect 268384 188300 268436 188352
rect 285772 188300 285824 188352
rect 129096 187688 129148 187740
rect 177304 187688 177356 187740
rect 205640 187688 205692 187740
rect 244464 187688 244516 187740
rect 222844 187620 222896 187672
rect 229744 187620 229796 187672
rect 177948 187008 178000 187060
rect 206284 187008 206336 187060
rect 56508 186940 56560 186992
rect 217232 186940 217284 186992
rect 275284 186940 275336 186992
rect 296812 186940 296864 186992
rect 217232 186396 217284 186448
rect 218152 186396 218204 186448
rect 133788 186328 133840 186380
rect 176016 186328 176068 186380
rect 218060 186328 218112 186380
rect 238944 186328 238996 186380
rect 186228 185648 186280 185700
rect 236092 185648 236144 185700
rect 258724 185648 258776 185700
rect 281724 185648 281776 185700
rect 207664 185580 207716 185632
rect 279424 185580 279476 185632
rect 114468 184968 114520 185020
rect 185768 184968 185820 185020
rect 100668 184900 100720 184952
rect 178684 184900 178736 184952
rect 177856 184220 177908 184272
rect 204168 184220 204220 184272
rect 204904 184220 204956 184272
rect 232044 184220 232096 184272
rect 184756 184152 184808 184204
rect 232504 184152 232556 184204
rect 232596 184152 232648 184204
rect 254032 184152 254084 184204
rect 280804 184152 280856 184204
rect 301136 184152 301188 184204
rect 117228 183608 117280 183660
rect 169392 183608 169444 183660
rect 108948 183540 109000 183592
rect 171968 183540 172020 183592
rect 204168 183472 204220 183524
rect 218060 183472 218112 183524
rect 224960 182928 225012 182980
rect 227720 182928 227772 182980
rect 184848 182860 184900 182912
rect 193864 182860 193916 182912
rect 199384 182860 199436 182912
rect 225696 182860 225748 182912
rect 240784 182860 240836 182912
rect 280436 182860 280488 182912
rect 170496 182792 170548 182844
rect 200764 182792 200816 182844
rect 220084 182792 220136 182844
rect 233516 182792 233568 182844
rect 246304 182792 246356 182844
rect 432052 182792 432104 182844
rect 134800 182248 134852 182300
rect 162860 182248 162912 182300
rect 123484 182180 123536 182232
rect 170496 182180 170548 182232
rect 178776 181500 178828 181552
rect 204904 181500 204956 181552
rect 206376 181500 206428 181552
rect 238852 181500 238904 181552
rect 181444 181432 181496 181484
rect 227812 181432 227864 181484
rect 260748 181432 260800 181484
rect 269212 181432 269264 181484
rect 279516 181432 279568 181484
rect 287336 181432 287388 181484
rect 148232 180888 148284 180940
rect 174544 180888 174596 180940
rect 115848 180820 115900 180872
rect 166448 180820 166500 180872
rect 275284 180820 275336 180872
rect 303804 180820 303856 180872
rect 182916 180752 182968 180804
rect 225880 180752 225932 180804
rect 228640 180752 228692 180804
rect 278688 180752 278740 180804
rect 278136 180616 278188 180668
rect 280344 180616 280396 180668
rect 214564 180072 214616 180124
rect 230388 180072 230440 180124
rect 254584 180072 254636 180124
rect 262220 180072 262272 180124
rect 272524 180072 272576 180124
rect 292764 180072 292816 180124
rect 282184 179732 282236 179784
rect 285956 179732 286008 179784
rect 119804 179460 119856 179512
rect 167736 179460 167788 179512
rect 128176 179392 128228 179444
rect 214104 179392 214156 179444
rect 231124 179324 231176 179376
rect 275284 179324 275336 179376
rect 215116 178712 215168 178764
rect 229284 178712 229336 178764
rect 276756 178712 276808 178764
rect 279240 178712 279292 178764
rect 196808 178644 196860 178696
rect 237472 178644 237524 178696
rect 265624 178644 265676 178696
rect 283012 178644 283064 178696
rect 285036 178644 285088 178696
rect 299664 178644 299716 178696
rect 300216 178644 300268 178696
rect 414112 178644 414164 178696
rect 132408 178100 132460 178152
rect 165528 178100 165580 178152
rect 125048 178032 125100 178084
rect 198096 178032 198148 178084
rect 102048 177964 102100 178016
rect 129096 177964 129148 178016
rect 225696 177964 225748 178016
rect 229100 177964 229152 178016
rect 276664 177964 276716 178016
rect 279332 177964 279384 178016
rect 284944 177964 284996 178016
rect 288440 177964 288492 178016
rect 215392 177352 215444 177404
rect 226248 177352 226300 177404
rect 238116 177352 238168 177404
rect 241520 177352 241572 177404
rect 198648 177284 198700 177336
rect 279516 177284 279568 177336
rect 136088 176740 136140 176792
rect 140780 176740 140832 176792
rect 158996 176740 159048 176792
rect 170404 176740 170456 176792
rect 130752 176672 130804 176724
rect 212448 176672 212500 176724
rect 140780 176604 140832 176656
rect 213920 176604 213972 176656
rect 269856 176604 269908 176656
rect 279884 176604 279936 176656
rect 276848 176536 276900 176588
rect 280068 176536 280120 176588
rect 227536 175992 227588 176044
rect 234712 175992 234764 176044
rect 47584 175924 47636 175976
rect 129004 175924 129056 175976
rect 129464 175924 129516 175976
rect 169760 175924 169812 175976
rect 185768 175924 185820 175976
rect 214472 175924 214524 175976
rect 227720 175924 227772 175976
rect 247224 175924 247276 175976
rect 279608 175924 279660 175976
rect 280160 175924 280212 175976
rect 314016 175924 314068 175976
rect 336004 175924 336056 175976
rect 215300 175244 215352 175296
rect 227812 175856 227864 175908
rect 221188 175788 221240 175840
rect 224224 175788 224276 175840
rect 162860 175176 162912 175228
rect 213920 175176 213972 175228
rect 214564 175176 214616 175228
rect 235356 175244 235408 175296
rect 264980 175244 265032 175296
rect 281816 175244 281868 175296
rect 314016 175244 314068 175296
rect 231124 175176 231176 175228
rect 232044 175176 232096 175228
rect 176016 175108 176068 175160
rect 214012 175108 214064 175160
rect 229008 175108 229060 175160
rect 282828 175108 282880 175160
rect 300952 175108 301004 175160
rect 244924 174496 244976 174548
rect 258172 174496 258224 174548
rect 229008 174020 229060 174072
rect 229192 174020 229244 174072
rect 258724 173952 258776 174004
rect 265072 173952 265124 174004
rect 214564 173884 214616 173936
rect 233424 173884 233476 173936
rect 240876 173884 240928 173936
rect 264980 173884 265032 173936
rect 165528 173816 165580 173868
rect 213920 173816 213972 173868
rect 212448 173748 212500 173800
rect 214012 173748 214064 173800
rect 167828 173408 167880 173460
rect 173440 173408 173492 173460
rect 230756 173340 230808 173392
rect 233240 173340 233292 173392
rect 177304 173136 177356 173188
rect 198004 173136 198056 173188
rect 238116 173136 238168 173188
rect 252560 173136 252612 173188
rect 259000 172592 259052 172644
rect 265072 172592 265124 172644
rect 254676 172524 254728 172576
rect 264980 172524 265032 172576
rect 169760 172456 169812 172508
rect 213920 172456 213972 172508
rect 231584 172456 231636 172508
rect 240232 172456 240284 172508
rect 173164 172388 173216 172440
rect 215300 172388 215352 172440
rect 231768 172116 231820 172168
rect 234620 172116 234672 172168
rect 247960 171164 248012 171216
rect 264980 171164 265032 171216
rect 240968 171096 241020 171148
rect 265072 171096 265124 171148
rect 165160 171028 165212 171080
rect 214012 171028 214064 171080
rect 231768 171028 231820 171080
rect 241520 171028 241572 171080
rect 164976 170960 165028 171012
rect 213920 170960 213972 171012
rect 230756 170960 230808 171012
rect 232504 170960 232556 171012
rect 281816 170960 281868 171012
rect 283196 170960 283248 171012
rect 371976 170348 372028 170400
rect 433984 170348 434036 170400
rect 243820 169736 243872 169788
rect 264980 169736 265032 169788
rect 170496 169668 170548 169720
rect 214012 169668 214064 169720
rect 231768 169668 231820 169720
rect 243544 169668 243596 169720
rect 282828 169668 282880 169720
rect 295524 169668 295576 169720
rect 198096 169600 198148 169652
rect 213920 169600 213972 169652
rect 231216 169192 231268 169244
rect 233332 169192 233384 169244
rect 250720 168444 250772 168496
rect 264980 168444 265032 168496
rect 240784 168376 240836 168428
rect 265072 168376 265124 168428
rect 167920 168308 167972 168360
rect 213920 168308 213972 168360
rect 282736 168308 282788 168360
rect 290096 168308 290148 168360
rect 169208 168240 169260 168292
rect 214012 168240 214064 168292
rect 230572 168240 230624 168292
rect 230848 168240 230900 168292
rect 231400 168172 231452 168224
rect 237472 168172 237524 168224
rect 282828 167968 282880 168020
rect 288440 167968 288492 168020
rect 391204 167628 391256 167680
rect 430672 167628 430724 167680
rect 256056 167084 256108 167136
rect 264980 167084 265032 167136
rect 252100 167016 252152 167068
rect 265072 167016 265124 167068
rect 167736 166948 167788 167000
rect 213920 166948 213972 167000
rect 177396 166880 177448 166932
rect 214012 166880 214064 166932
rect 231768 166676 231820 166728
rect 235264 166676 235316 166728
rect 230480 166268 230532 166320
rect 230756 166268 230808 166320
rect 236736 166268 236788 166320
rect 265716 166268 265768 166320
rect 370504 166268 370556 166320
rect 439872 166268 439924 166320
rect 232780 165588 232832 165640
rect 264980 165588 265032 165640
rect 166448 165520 166500 165572
rect 213920 165520 213972 165572
rect 166540 165452 166592 165504
rect 214012 165452 214064 165504
rect 231492 165452 231544 165504
rect 236000 165452 236052 165504
rect 282828 165180 282880 165232
rect 287060 165180 287112 165232
rect 3516 164840 3568 164892
rect 17224 164840 17276 164892
rect 406384 164840 406436 164892
rect 420276 164840 420328 164892
rect 238300 164296 238352 164348
rect 264980 164296 265032 164348
rect 234068 164228 234120 164280
rect 265072 164228 265124 164280
rect 184388 164160 184440 164212
rect 213920 164160 213972 164212
rect 231768 164160 231820 164212
rect 247408 164160 247460 164212
rect 282184 164160 282236 164212
rect 309140 164160 309192 164212
rect 231676 164092 231728 164144
rect 242900 164092 242952 164144
rect 281816 164092 281868 164144
rect 284484 164092 284536 164144
rect 198004 163480 198056 163532
rect 214840 163480 214892 163532
rect 319444 163480 319496 163532
rect 371976 163480 372028 163532
rect 380164 163480 380216 163532
rect 447416 163480 447468 163532
rect 255964 162936 256016 162988
rect 265072 162936 265124 162988
rect 245016 162868 245068 162920
rect 264980 162868 265032 162920
rect 167644 162800 167696 162852
rect 213920 162800 213972 162852
rect 175924 162732 175976 162784
rect 214012 162732 214064 162784
rect 282276 162732 282328 162784
rect 329840 162732 329892 162784
rect 230940 162664 230992 162716
rect 233424 162664 233476 162716
rect 378876 162120 378928 162172
rect 418252 162120 418304 162172
rect 247776 161508 247828 161560
rect 264980 161508 265032 161560
rect 235448 161440 235500 161492
rect 265072 161440 265124 161492
rect 171968 161372 172020 161424
rect 213920 161372 213972 161424
rect 282644 161372 282696 161424
rect 325700 161372 325752 161424
rect 173348 161304 173400 161356
rect 214012 161304 214064 161356
rect 231768 160692 231820 160744
rect 241520 160692 241572 160744
rect 243728 160148 243780 160200
rect 264980 160148 265032 160200
rect 236920 160080 236972 160132
rect 265072 160080 265124 160132
rect 181536 160012 181588 160064
rect 213920 160012 213972 160064
rect 282828 160012 282880 160064
rect 320180 160012 320232 160064
rect 196716 159944 196768 159996
rect 214012 159944 214064 159996
rect 282736 159944 282788 159996
rect 296904 159944 296956 159996
rect 167828 159332 167880 159384
rect 181444 159332 181496 159384
rect 230572 159332 230624 159384
rect 244924 159332 244976 159384
rect 309048 159332 309100 159384
rect 425060 159332 425112 159384
rect 231124 159264 231176 159316
rect 238392 159264 238444 159316
rect 248052 158788 248104 158840
rect 265072 158788 265124 158840
rect 238208 158720 238260 158772
rect 264980 158720 265032 158772
rect 180340 158652 180392 158704
rect 213920 158652 213972 158704
rect 282092 158652 282144 158704
rect 288624 158652 288676 158704
rect 170404 157972 170456 158024
rect 214564 157972 214616 158024
rect 231308 157972 231360 158024
rect 238760 157972 238812 158024
rect 282184 157972 282236 158024
rect 306472 157972 306524 158024
rect 353944 157972 353996 158024
rect 414204 157972 414256 158024
rect 244924 157428 244976 157480
rect 264980 157428 265032 157480
rect 233976 157360 234028 157412
rect 265072 157360 265124 157412
rect 280068 157360 280120 157412
rect 281540 157360 281592 157412
rect 166356 157292 166408 157344
rect 213920 157292 213972 157344
rect 178684 157224 178736 157276
rect 214012 157224 214064 157276
rect 283564 156680 283616 156732
rect 294236 156680 294288 156732
rect 231124 156612 231176 156664
rect 231952 156612 232004 156664
rect 282828 156612 282880 156664
rect 303804 156612 303856 156664
rect 398748 156612 398800 156664
rect 582748 156612 582800 156664
rect 231768 156544 231820 156596
rect 244464 156544 244516 156596
rect 253296 156000 253348 156052
rect 264980 156000 265032 156052
rect 239864 155932 239916 155984
rect 265072 155932 265124 155984
rect 169116 155864 169168 155916
rect 213920 155864 213972 155916
rect 185676 155796 185728 155848
rect 214012 155796 214064 155848
rect 282552 155660 282604 155712
rect 285956 155660 286008 155712
rect 230020 155184 230072 155236
rect 265256 155184 265308 155236
rect 398656 155184 398708 155236
rect 583576 155184 583628 155236
rect 235540 154572 235592 154624
rect 265164 154572 265216 154624
rect 231584 154504 231636 154556
rect 240140 154504 240192 154556
rect 282368 154504 282420 154556
rect 313464 154504 313516 154556
rect 230664 153892 230716 153944
rect 241612 153892 241664 153944
rect 241060 153824 241112 153876
rect 264980 153824 265032 153876
rect 282736 153824 282788 153876
rect 289912 153824 289964 153876
rect 331956 153824 332008 153876
rect 385776 153824 385828 153876
rect 389916 153824 389968 153876
rect 438952 153824 439004 153876
rect 211896 153280 211948 153332
rect 214012 153280 214064 153332
rect 166356 153212 166408 153264
rect 213920 153212 213972 153264
rect 260288 153212 260340 153264
rect 264980 153212 265032 153264
rect 282828 153144 282880 153196
rect 298284 153144 298336 153196
rect 230756 152464 230808 152516
rect 260840 152464 260892 152516
rect 297364 152464 297416 152516
rect 443184 152464 443236 152516
rect 177304 151784 177356 151836
rect 213920 151784 213972 151836
rect 232596 151784 232648 151836
rect 264980 151784 265032 151836
rect 246488 151104 246540 151156
rect 265808 151104 265860 151156
rect 171876 151036 171928 151088
rect 202236 151036 202288 151088
rect 230388 151036 230440 151088
rect 249800 151036 249852 151088
rect 282736 151036 282788 151088
rect 311992 151036 312044 151088
rect 374736 151036 374788 151088
rect 395436 151036 395488 151088
rect 198096 150424 198148 150476
rect 213920 150424 213972 150476
rect 174544 150356 174596 150408
rect 214012 150356 214064 150408
rect 230572 150356 230624 150408
rect 245660 150424 245712 150476
rect 252008 150424 252060 150476
rect 264980 150424 265032 150476
rect 334716 150424 334768 150476
rect 407212 150424 407264 150476
rect 281908 150356 281960 150408
rect 317420 150356 317472 150408
rect 421104 150356 421156 150408
rect 421564 150356 421616 150408
rect 583392 150356 583444 150408
rect 2780 150288 2832 150340
rect 4804 150288 4856 150340
rect 181444 150288 181496 150340
rect 213920 150288 213972 150340
rect 282828 150288 282880 150340
rect 299756 150288 299808 150340
rect 231216 149676 231268 149728
rect 258724 149676 258776 149728
rect 309784 149676 309836 149728
rect 425796 149676 425848 149728
rect 253388 149064 253440 149116
rect 264980 149064 265032 149116
rect 230572 148996 230624 149048
rect 252652 148996 252704 149048
rect 282828 148996 282880 149048
rect 292580 148996 292632 149048
rect 449992 148996 450044 149048
rect 450544 148996 450596 149048
rect 583024 148996 583076 149048
rect 411904 148384 411956 148436
rect 434076 148384 434128 148436
rect 173256 148316 173308 148368
rect 186964 148316 187016 148368
rect 356704 148316 356756 148368
rect 442264 148316 442316 148368
rect 256240 147704 256292 147756
rect 264980 147704 265032 147756
rect 184388 147636 184440 147688
rect 213920 147636 213972 147688
rect 238116 147636 238168 147688
rect 265072 147636 265124 147688
rect 299388 147636 299440 147688
rect 407672 147636 407724 147688
rect 580908 147636 580960 147688
rect 582380 147636 582432 147688
rect 230756 147568 230808 147620
rect 233516 147568 233568 147620
rect 282736 147568 282788 147620
rect 323032 147568 323084 147620
rect 282828 147500 282880 147552
rect 292764 147500 292816 147552
rect 233792 146956 233844 147008
rect 247224 146956 247276 147008
rect 231124 146888 231176 146940
rect 250720 146888 250772 146940
rect 398472 146888 398524 146940
rect 583300 146888 583352 146940
rect 250628 146344 250680 146396
rect 264980 146344 265032 146396
rect 178684 146276 178736 146328
rect 213920 146276 213972 146328
rect 249156 146276 249208 146328
rect 265072 146276 265124 146328
rect 387156 146276 387208 146328
rect 436652 146276 436704 146328
rect 230664 146208 230716 146260
rect 238852 146208 238904 146260
rect 282552 146208 282604 146260
rect 299664 146208 299716 146260
rect 420184 146208 420236 146260
rect 422944 146208 422996 146260
rect 282828 146140 282880 146192
rect 294144 146140 294196 146192
rect 382924 145596 382976 145648
rect 412732 145596 412784 145648
rect 231400 145528 231452 145580
rect 240968 145528 241020 145580
rect 322204 145528 322256 145580
rect 409972 145528 410024 145580
rect 411996 145528 412048 145580
rect 422392 145528 422444 145580
rect 177396 144984 177448 145036
rect 214012 144984 214064 145036
rect 243636 144984 243688 145036
rect 265072 144984 265124 145036
rect 167644 144916 167696 144968
rect 213920 144916 213972 144968
rect 239588 144916 239640 144968
rect 264980 144916 265032 144968
rect 231768 144848 231820 144900
rect 242164 144848 242216 144900
rect 282460 144848 282512 144900
rect 303620 144848 303672 144900
rect 302976 144236 303028 144288
rect 441988 144236 442040 144288
rect 403624 144168 403676 144220
rect 419724 144168 419776 144220
rect 424692 144168 424744 144220
rect 582564 144168 582616 144220
rect 246396 143624 246448 143676
rect 264980 143624 265032 143676
rect 180248 143556 180300 143608
rect 213920 143556 213972 143608
rect 240968 143556 241020 143608
rect 265072 143556 265124 143608
rect 329104 143488 329156 143540
rect 330484 143488 330536 143540
rect 407212 143488 407264 143540
rect 408868 143488 408920 143540
rect 410524 143488 410576 143540
rect 411996 143488 412048 143540
rect 414756 143488 414808 143540
rect 416412 143488 416464 143540
rect 430580 143488 430632 143540
rect 431316 143488 431368 143540
rect 231768 143420 231820 143472
rect 236644 143420 236696 143472
rect 413284 143420 413336 143472
rect 418436 143420 418488 143472
rect 237012 142808 237064 142860
rect 265624 142808 265676 142860
rect 415860 142808 415912 142860
rect 416780 142808 416832 142860
rect 438676 142808 438728 142860
rect 449992 142808 450044 142860
rect 282828 142400 282880 142452
rect 287336 142400 287388 142452
rect 209228 142196 209280 142248
rect 213920 142196 213972 142248
rect 171784 142128 171836 142180
rect 214012 142128 214064 142180
rect 232504 142128 232556 142180
rect 264980 142128 265032 142180
rect 381544 142128 381596 142180
rect 405188 142128 405240 142180
rect 418804 142128 418856 142180
rect 424140 142128 424192 142180
rect 425704 142128 425756 142180
rect 433524 142128 433576 142180
rect 434076 142128 434128 142180
rect 583024 142128 583076 142180
rect 282828 142060 282880 142112
rect 313280 142060 313332 142112
rect 374644 142060 374696 142112
rect 376760 142060 376812 142112
rect 282736 141992 282788 142044
rect 295432 141992 295484 142044
rect 249340 141448 249392 141500
rect 265992 141448 266044 141500
rect 181536 141380 181588 141432
rect 214656 141380 214708 141432
rect 231584 141380 231636 141432
rect 251824 141380 251876 141432
rect 383108 140836 383160 140888
rect 417148 140836 417200 140888
rect 425428 140836 425480 140888
rect 425796 140836 425848 140888
rect 464344 140836 464396 140888
rect 205272 140768 205324 140820
rect 213920 140768 213972 140820
rect 261668 140768 261720 140820
rect 264980 140768 265032 140820
rect 303620 140768 303672 140820
rect 409604 140768 409656 140820
rect 428556 140768 428608 140820
rect 582656 140768 582708 140820
rect 282828 140700 282880 140752
rect 289820 140700 289872 140752
rect 405740 140700 405792 140752
rect 406660 140700 406712 140752
rect 412640 140700 412692 140752
rect 412916 140700 412968 140752
rect 400220 140292 400272 140344
rect 401324 140292 401376 140344
rect 234160 140088 234212 140140
rect 243820 140088 243872 140140
rect 242532 140020 242584 140072
rect 264336 140020 264388 140072
rect 417424 140020 417476 140072
rect 441712 140020 441764 140072
rect 342904 139476 342956 139528
rect 417332 139612 417384 139664
rect 401508 139544 401560 139596
rect 170404 139408 170456 139460
rect 213920 139408 213972 139460
rect 254584 139408 254636 139460
rect 264980 139408 265032 139460
rect 399484 139408 399536 139460
rect 402980 139408 403032 139460
rect 580172 139408 580224 139460
rect 231768 139340 231820 139392
rect 254032 139340 254084 139392
rect 282644 139340 282696 139392
rect 301136 139340 301188 139392
rect 395436 139340 395488 139392
rect 397552 139340 397604 139392
rect 399852 139340 399904 139392
rect 404084 139340 404136 139392
rect 442172 139340 442224 139392
rect 460940 139340 460992 139392
rect 583484 139340 583536 139392
rect 281724 138932 281776 138984
rect 284576 138932 284628 138984
rect 169116 138660 169168 138712
rect 214380 138660 214432 138712
rect 195428 137980 195480 138032
rect 213920 137980 213972 138032
rect 229836 137980 229888 138032
rect 264980 137980 265032 138032
rect 3516 137912 3568 137964
rect 22744 137912 22796 137964
rect 231768 137912 231820 137964
rect 244372 137912 244424 137964
rect 282828 137912 282880 137964
rect 306380 137912 306432 137964
rect 442908 137232 442960 137284
rect 447140 137232 447192 137284
rect 582564 137232 582616 137284
rect 187148 136620 187200 136672
rect 213920 136620 213972 136672
rect 258724 136620 258776 136672
rect 264980 136620 265032 136672
rect 395620 136620 395672 136672
rect 397920 136620 397972 136672
rect 230572 136552 230624 136604
rect 245844 136552 245896 136604
rect 282828 136552 282880 136604
rect 292672 136552 292724 136604
rect 231308 136144 231360 136196
rect 236736 136144 236788 136196
rect 196716 135940 196768 135992
rect 214012 135940 214064 135992
rect 167736 135872 167788 135924
rect 213368 135872 213420 135924
rect 282276 135872 282328 135924
rect 327172 135872 327224 135924
rect 331956 135872 332008 135924
rect 387156 135872 387208 135924
rect 442908 135464 442960 135516
rect 448704 135464 448756 135516
rect 258816 135328 258868 135380
rect 265072 135328 265124 135380
rect 388536 135328 388588 135380
rect 397644 135328 397696 135380
rect 231308 135260 231360 135312
rect 231584 135260 231636 135312
rect 260196 135260 260248 135312
rect 264980 135260 265032 135312
rect 374736 135260 374788 135312
rect 397552 135260 397604 135312
rect 231492 135192 231544 135244
rect 259000 135192 259052 135244
rect 282828 135192 282880 135244
rect 318800 135192 318852 135244
rect 231768 135124 231820 135176
rect 249248 135124 249300 135176
rect 282460 134920 282512 134972
rect 285864 134920 285916 134972
rect 169208 134512 169260 134564
rect 214104 134512 214156 134564
rect 363604 134512 363656 134564
rect 381636 134512 381688 134564
rect 210424 133900 210476 133952
rect 213920 133900 213972 133952
rect 378876 133900 378928 133952
rect 397644 133900 397696 133952
rect 231492 133832 231544 133884
rect 254676 133832 254728 133884
rect 444380 133832 444432 133884
rect 448612 133832 448664 133884
rect 442908 133220 442960 133272
rect 444380 133220 444432 133272
rect 230664 133152 230716 133204
rect 256056 133152 256108 133204
rect 358176 133152 358228 133204
rect 391204 133152 391256 133204
rect 209136 132540 209188 132592
rect 213920 132540 213972 132592
rect 192668 132472 192720 132524
rect 214012 132472 214064 132524
rect 255964 132472 256016 132524
rect 264980 132472 265032 132524
rect 392768 132472 392820 132524
rect 397552 132472 397604 132524
rect 231768 132404 231820 132456
rect 247960 132404 248012 132456
rect 282828 132404 282880 132456
rect 324320 132404 324372 132456
rect 371884 132404 371936 132456
rect 398472 132404 398524 132456
rect 442908 132404 442960 132456
rect 583760 132404 583812 132456
rect 181444 131724 181496 131776
rect 211896 131724 211948 131776
rect 305736 131724 305788 131776
rect 327080 131724 327132 131776
rect 395620 131724 395672 131776
rect 231400 131656 231452 131708
rect 234160 131656 234212 131708
rect 251824 131180 251876 131232
rect 264980 131180 265032 131232
rect 185676 131112 185728 131164
rect 213920 131112 213972 131164
rect 247684 131112 247736 131164
rect 265072 131112 265124 131164
rect 231768 131044 231820 131096
rect 264244 131044 264296 131096
rect 282276 131044 282328 131096
rect 310612 131044 310664 131096
rect 231124 130976 231176 131028
rect 260104 130976 260156 131028
rect 282644 130976 282696 131028
rect 307852 130976 307904 131028
rect 192576 130364 192628 130416
rect 206468 130364 206520 130416
rect 210516 129820 210568 129872
rect 214012 129820 214064 129872
rect 200856 129752 200908 129804
rect 213920 129752 213972 129804
rect 389916 129752 389968 129804
rect 398840 129752 398892 129804
rect 230756 129684 230808 129736
rect 240784 129684 240836 129736
rect 370504 129684 370556 129736
rect 372620 129684 372672 129736
rect 397552 129684 397604 129736
rect 318248 129004 318300 129056
rect 398196 129004 398248 129056
rect 205180 128392 205232 128444
rect 213920 128392 213972 128444
rect 202420 128324 202472 128376
rect 214012 128324 214064 128376
rect 254860 128324 254912 128376
rect 264980 128392 265032 128444
rect 264612 128324 264664 128376
rect 265716 128324 265768 128376
rect 231768 128256 231820 128308
rect 252100 128256 252152 128308
rect 340236 128256 340288 128308
rect 397552 128256 397604 128308
rect 231676 128188 231728 128240
rect 236828 128188 236880 128240
rect 282828 128188 282880 128240
rect 316040 128188 316092 128240
rect 182916 127576 182968 127628
rect 214840 127576 214892 127628
rect 442908 127576 442960 127628
rect 449992 127576 450044 127628
rect 261576 127032 261628 127084
rect 265072 127032 265124 127084
rect 62028 126964 62080 127016
rect 65524 126964 65576 127016
rect 198004 126964 198056 127016
rect 213920 126964 213972 127016
rect 236736 126964 236788 127016
rect 264980 126964 265032 127016
rect 363604 126964 363656 127016
rect 397552 126964 397604 127016
rect 231308 126896 231360 126948
rect 250444 126896 250496 126948
rect 263048 126896 263100 126948
rect 266084 126896 266136 126948
rect 282828 126896 282880 126948
rect 291200 126896 291252 126948
rect 464344 126896 464396 126948
rect 580172 126896 580224 126948
rect 230572 126692 230624 126744
rect 232780 126692 232832 126744
rect 166448 126216 166500 126268
rect 213276 126216 213328 126268
rect 238392 126216 238444 126268
rect 245292 126216 245344 126268
rect 282092 126216 282144 126268
rect 313372 126216 313424 126268
rect 353944 126216 353996 126268
rect 354588 126216 354640 126268
rect 397552 126216 397604 126268
rect 195520 125604 195572 125656
rect 213920 125604 213972 125656
rect 245108 125604 245160 125656
rect 264980 125604 265032 125656
rect 442908 125604 442960 125656
rect 454040 125604 454092 125656
rect 230756 125536 230808 125588
rect 238300 125536 238352 125588
rect 281632 125536 281684 125588
rect 303712 125536 303764 125588
rect 315304 125536 315356 125588
rect 397644 125536 397696 125588
rect 392676 125468 392728 125520
rect 397552 125468 397604 125520
rect 231492 125128 231544 125180
rect 234068 125128 234120 125180
rect 207756 124244 207808 124296
rect 214012 124244 214064 124296
rect 238024 124244 238076 124296
rect 264980 124244 265032 124296
rect 171968 124176 172020 124228
rect 213920 124176 213972 124228
rect 236644 124176 236696 124228
rect 265072 124176 265124 124228
rect 282644 124108 282696 124160
rect 307760 124108 307812 124160
rect 309968 124108 310020 124160
rect 397552 124108 397604 124160
rect 442908 124108 442960 124160
rect 582932 124108 582984 124160
rect 442816 124040 442868 124092
rect 447232 124040 447284 124092
rect 231124 123904 231176 123956
rect 235540 123904 235592 123956
rect 230664 123428 230716 123480
rect 248052 123428 248104 123480
rect 171876 122816 171928 122868
rect 213920 122816 213972 122868
rect 235448 122816 235500 122868
rect 264980 122816 265032 122868
rect 231768 122748 231820 122800
rect 257436 122748 257488 122800
rect 309876 122748 309928 122800
rect 374736 122748 374788 122800
rect 442264 122748 442316 122800
rect 442908 122748 442960 122800
rect 582472 122748 582524 122800
rect 231032 122680 231084 122732
rect 245016 122680 245068 122732
rect 252100 122068 252152 122120
rect 265072 122068 265124 122120
rect 282828 121592 282880 121644
rect 288716 121592 288768 121644
rect 196808 121524 196860 121576
rect 213920 121524 213972 121576
rect 63408 121456 63460 121508
rect 65984 121456 66036 121508
rect 175924 121456 175976 121508
rect 214012 121456 214064 121508
rect 309140 121456 309192 121508
rect 309876 121456 309928 121508
rect 374644 121456 374696 121508
rect 397552 121456 397604 121508
rect 231768 121388 231820 121440
rect 247776 121388 247828 121440
rect 342996 121388 343048 121440
rect 398748 121388 398800 121440
rect 441620 121388 441672 121440
rect 442632 121388 442684 121440
rect 582380 121388 582432 121440
rect 249248 120708 249300 120760
rect 264980 120708 265032 120760
rect 231492 120640 231544 120692
rect 236920 120640 236972 120692
rect 193956 120164 194008 120216
rect 213920 120164 213972 120216
rect 170496 120096 170548 120148
rect 214012 120096 214064 120148
rect 259000 120096 259052 120148
rect 265072 120096 265124 120148
rect 231768 120028 231820 120080
rect 243728 120028 243780 120080
rect 282828 120028 282880 120080
rect 288532 120028 288584 120080
rect 378784 120028 378836 120080
rect 397552 120028 397604 120080
rect 442908 119688 442960 119740
rect 447416 119688 447468 119740
rect 247960 119348 248012 119400
rect 262864 119348 262916 119400
rect 282184 119348 282236 119400
rect 299572 119348 299624 119400
rect 338212 119348 338264 119400
rect 395436 119348 395488 119400
rect 203708 118736 203760 118788
rect 213920 118736 213972 118788
rect 195336 118668 195388 118720
rect 214012 118668 214064 118720
rect 259276 118668 259328 118720
rect 264980 118668 265032 118720
rect 230572 118600 230624 118652
rect 233976 118600 234028 118652
rect 282828 118600 282880 118652
rect 298192 118600 298244 118652
rect 352564 118600 352616 118652
rect 397644 118600 397696 118652
rect 360844 118532 360896 118584
rect 397552 118532 397604 118584
rect 282828 118056 282880 118108
rect 287244 118056 287296 118108
rect 231676 117988 231728 118040
rect 246488 117988 246540 118040
rect 238300 117920 238352 117972
rect 265808 117920 265860 117972
rect 198280 117376 198332 117428
rect 214012 117376 214064 117428
rect 169300 117308 169352 117360
rect 213920 117308 213972 117360
rect 250444 117308 250496 117360
rect 264980 117308 265032 117360
rect 282828 117240 282880 117292
rect 290004 117240 290056 117292
rect 291108 117240 291160 117292
rect 391204 117240 391256 117292
rect 397552 117240 397604 117292
rect 231768 117172 231820 117224
rect 244924 117172 244976 117224
rect 230848 117104 230900 117156
rect 232688 117104 232740 117156
rect 282276 116696 282328 116748
rect 285772 116696 285824 116748
rect 167828 116560 167880 116612
rect 198096 116560 198148 116612
rect 200948 116016 201000 116068
rect 214012 116016 214064 116068
rect 257436 116016 257488 116068
rect 264980 116016 265032 116068
rect 189908 115948 189960 116000
rect 213920 115948 213972 116000
rect 240784 115948 240836 116000
rect 265072 115948 265124 116000
rect 231492 115880 231544 115932
rect 253296 115880 253348 115932
rect 281724 115880 281776 115932
rect 302332 115880 302384 115932
rect 356796 115880 356848 115932
rect 397552 115880 397604 115932
rect 282460 115812 282512 115864
rect 295340 115812 295392 115864
rect 184296 115200 184348 115252
rect 200856 115200 200908 115252
rect 230664 115200 230716 115252
rect 251916 115200 251968 115252
rect 363696 115200 363748 115252
rect 397368 115200 397420 115252
rect 203616 114588 203668 114640
rect 214012 114588 214064 114640
rect 258908 114588 258960 114640
rect 265072 114588 265124 114640
rect 198096 114520 198148 114572
rect 213920 114520 213972 114572
rect 256240 114520 256292 114572
rect 264980 114520 265032 114572
rect 442908 114520 442960 114572
rect 445944 114520 445996 114572
rect 452660 114520 452712 114572
rect 231676 114452 231728 114504
rect 241060 114452 241112 114504
rect 323584 114452 323636 114504
rect 397552 114452 397604 114504
rect 231492 114180 231544 114232
rect 233884 114180 233936 114232
rect 282276 114112 282328 114164
rect 285680 114112 285732 114164
rect 442356 113908 442408 113960
rect 449900 113908 449952 113960
rect 241152 113772 241204 113824
rect 254860 113772 254912 113824
rect 385776 113772 385828 113824
rect 397920 113772 397972 113824
rect 188528 113228 188580 113280
rect 213920 113228 213972 113280
rect 181628 113160 181680 113212
rect 214012 113160 214064 113212
rect 253480 113160 253532 113212
rect 264980 113160 265032 113212
rect 231768 113092 231820 113144
rect 260288 113092 260340 113144
rect 282828 113092 282880 113144
rect 321560 113092 321612 113144
rect 367100 113092 367152 113144
rect 231032 113024 231084 113076
rect 249340 113024 249392 113076
rect 282828 112616 282880 112668
rect 287152 112616 287204 112668
rect 178776 111868 178828 111920
rect 214012 111868 214064 111920
rect 263140 111868 263192 111920
rect 265256 111868 265308 111920
rect 377496 111868 377548 111920
rect 397644 111868 397696 111920
rect 173348 111800 173400 111852
rect 213920 111800 213972 111852
rect 251916 111800 251968 111852
rect 264980 111800 265032 111852
rect 359556 111800 359608 111852
rect 397736 111800 397788 111852
rect 3148 111732 3200 111784
rect 35164 111732 35216 111784
rect 230572 111732 230624 111784
rect 232596 111732 232648 111784
rect 282276 111732 282328 111784
rect 293960 111732 294012 111784
rect 336096 111732 336148 111784
rect 397460 111732 397512 111784
rect 231768 111664 231820 111716
rect 242532 111664 242584 111716
rect 442356 111528 442408 111580
rect 445852 111528 445904 111580
rect 359464 111052 359516 111104
rect 397644 111052 397696 111104
rect 442172 111052 442224 111104
rect 447140 111052 447192 111104
rect 193864 110508 193916 110560
rect 214012 110508 214064 110560
rect 249064 110508 249116 110560
rect 265072 110508 265124 110560
rect 166540 110440 166592 110492
rect 213920 110440 213972 110492
rect 243728 110440 243780 110492
rect 264980 110440 265032 110492
rect 167828 110372 167880 110424
rect 181536 110372 181588 110424
rect 231768 110372 231820 110424
rect 252008 110372 252060 110424
rect 282828 110372 282880 110424
rect 298100 110372 298152 110424
rect 231676 109692 231728 109744
rect 246396 109692 246448 109744
rect 360844 109692 360896 109744
rect 397552 109692 397604 109744
rect 192484 109080 192536 109132
rect 214012 109080 214064 109132
rect 256056 109080 256108 109132
rect 264980 109080 265032 109132
rect 180340 109012 180392 109064
rect 213920 109012 213972 109064
rect 250536 109012 250588 109064
rect 265072 109012 265124 109064
rect 385776 109012 385828 109064
rect 397460 109012 397512 109064
rect 231492 108944 231544 108996
rect 253388 108944 253440 108996
rect 282368 108944 282420 108996
rect 305092 108944 305144 108996
rect 231768 108876 231820 108928
rect 242440 108876 242492 108928
rect 257620 108264 257672 108316
rect 264336 108264 264388 108316
rect 302884 108264 302936 108316
rect 398196 108264 398248 108316
rect 207664 107720 207716 107772
rect 214012 107720 214064 107772
rect 173256 107652 173308 107704
rect 213920 107652 213972 107704
rect 367836 107652 367888 107704
rect 397460 107652 397512 107704
rect 442908 107652 442960 107704
rect 452660 107652 452712 107704
rect 231584 107584 231636 107636
rect 264612 107584 264664 107636
rect 304264 107584 304316 107636
rect 397552 107584 397604 107636
rect 442540 107584 442592 107636
rect 456800 107584 456852 107636
rect 230940 107516 230992 107568
rect 238116 107516 238168 107568
rect 381636 107516 381688 107568
rect 397460 107516 397512 107568
rect 178868 106904 178920 106956
rect 205272 106904 205324 106956
rect 205088 106360 205140 106412
rect 214012 106360 214064 106412
rect 167828 106292 167880 106344
rect 213920 106292 213972 106344
rect 246488 106292 246540 106344
rect 264980 106292 265032 106344
rect 231584 106224 231636 106276
rect 249156 106224 249208 106276
rect 320916 106224 320968 106276
rect 397460 106224 397512 106276
rect 167736 105544 167788 105596
rect 195520 105544 195572 105596
rect 371976 105544 372028 105596
rect 399760 105544 399812 105596
rect 260288 104932 260340 104984
rect 265072 104932 265124 104984
rect 198188 104864 198240 104916
rect 213920 104864 213972 104916
rect 245016 104864 245068 104916
rect 264980 104864 265032 104916
rect 231768 104796 231820 104848
rect 250628 104796 250680 104848
rect 281908 104796 281960 104848
rect 284392 104796 284444 104848
rect 327724 104796 327776 104848
rect 397460 104796 397512 104848
rect 231492 104728 231544 104780
rect 243636 104728 243688 104780
rect 172060 104184 172112 104236
rect 198280 104184 198332 104236
rect 166264 104116 166316 104168
rect 214564 104116 214616 104168
rect 383016 104116 383068 104168
rect 399852 104116 399904 104168
rect 441988 104116 442040 104168
rect 451280 104116 451332 104168
rect 211896 103504 211948 103556
rect 213920 103504 213972 103556
rect 254768 103504 254820 103556
rect 264980 103504 265032 103556
rect 231768 103436 231820 103488
rect 240968 103436 241020 103488
rect 282828 103436 282880 103488
rect 314660 103436 314712 103488
rect 322296 103436 322348 103488
rect 397460 103436 397512 103488
rect 231400 103368 231452 103420
rect 239588 103368 239640 103420
rect 281724 103164 281776 103216
rect 283564 103164 283616 103216
rect 442724 102756 442776 102808
rect 444472 102756 444524 102808
rect 187056 102212 187108 102264
rect 214012 102212 214064 102264
rect 169024 102144 169076 102196
rect 213920 102144 213972 102196
rect 249156 102144 249208 102196
rect 264980 102144 265032 102196
rect 231768 102076 231820 102128
rect 247868 102076 247920 102128
rect 170680 101464 170732 101516
rect 196716 101464 196768 101516
rect 230480 101464 230532 101516
rect 238300 101464 238352 101516
rect 177488 101396 177540 101448
rect 213460 101396 213512 101448
rect 439964 101396 440016 101448
rect 463700 101396 463752 101448
rect 261760 100784 261812 100836
rect 265072 100784 265124 100836
rect 176016 100716 176068 100768
rect 177396 100716 177448 100768
rect 196900 100716 196952 100768
rect 213920 100716 213972 100768
rect 241060 100716 241112 100768
rect 264980 100716 265032 100768
rect 395436 100716 395488 100768
rect 397552 100716 397604 100768
rect 398196 100716 398248 100768
rect 439964 100716 440016 100768
rect 399852 100648 399904 100700
rect 403348 100648 403400 100700
rect 404636 100648 404688 100700
rect 439320 100648 439372 100700
rect 231768 100580 231820 100632
rect 256148 100580 256200 100632
rect 399760 100580 399812 100632
rect 402980 100580 403032 100632
rect 405280 99968 405332 100020
rect 580172 99968 580224 100020
rect 230572 99696 230624 99748
rect 232504 99696 232556 99748
rect 211988 99424 212040 99476
rect 214472 99424 214524 99476
rect 257528 99424 257580 99476
rect 265072 99424 265124 99476
rect 181720 99356 181772 99408
rect 213920 99356 213972 99408
rect 233976 99356 234028 99408
rect 264980 99356 265032 99408
rect 395344 99356 395396 99408
rect 432788 99356 432840 99408
rect 435548 99356 435600 99408
rect 440516 99356 440568 99408
rect 231032 99288 231084 99340
rect 263048 99288 263100 99340
rect 282000 99288 282052 99340
rect 296812 99288 296864 99340
rect 376024 99288 376076 99340
rect 417700 99288 417752 99340
rect 582748 99288 582800 99340
rect 282828 99220 282880 99272
rect 294052 99220 294104 99272
rect 384304 99220 384356 99272
rect 411996 99220 412048 99272
rect 433524 99220 433576 99272
rect 445760 99220 445812 99272
rect 230756 98812 230808 98864
rect 234160 98812 234212 98864
rect 358084 98608 358136 98660
rect 381636 98608 381688 98660
rect 173440 98064 173492 98116
rect 214012 98064 214064 98116
rect 164884 97996 164936 98048
rect 213920 97996 213972 98048
rect 261852 97996 261904 98048
rect 264980 97996 265032 98048
rect 3516 97928 3568 97980
rect 15844 97928 15896 97980
rect 215300 97928 215352 97980
rect 182824 97248 182876 97300
rect 213276 97248 213328 97300
rect 165528 96636 165580 96688
rect 213920 96636 213972 96688
rect 282828 97928 282880 97980
rect 302240 97928 302292 97980
rect 434628 97928 434680 97980
rect 465080 97928 465132 97980
rect 583116 97928 583168 97980
rect 282736 97860 282788 97912
rect 291384 97860 291436 97912
rect 401416 97860 401468 97912
rect 432236 97860 432288 97912
rect 435364 97860 435416 97912
rect 448520 97860 448572 97912
rect 403624 97792 403676 97844
rect 404452 97792 404504 97844
rect 264980 97248 265032 97300
rect 300124 97248 300176 97300
rect 391940 97248 391992 97300
rect 394148 96908 394200 96960
rect 401140 96908 401192 96960
rect 414020 96908 414072 96960
rect 414756 96908 414808 96960
rect 430580 96908 430632 96960
rect 431132 96908 431184 96960
rect 421564 96840 421616 96892
rect 423404 96840 423456 96892
rect 418804 96704 418856 96756
rect 420092 96704 420144 96756
rect 235356 96636 235408 96688
rect 265072 96636 265124 96688
rect 282828 96568 282880 96620
rect 301044 96568 301096 96620
rect 334624 96568 334676 96620
rect 422668 96568 422720 96620
rect 389824 96500 389876 96552
rect 418988 96500 419040 96552
rect 225052 96024 225104 96076
rect 226432 96024 226484 96076
rect 168288 95956 168340 96008
rect 184388 95956 184440 96008
rect 198648 95956 198700 96008
rect 222476 95956 222528 96008
rect 173164 95888 173216 95940
rect 213184 95888 213236 95940
rect 211804 95820 211856 95872
rect 229008 95820 229060 95872
rect 230480 95480 230532 95532
rect 232504 95480 232556 95532
rect 267648 95412 267700 95464
rect 269212 95412 269264 95464
rect 226432 95208 226484 95260
rect 241520 95208 241572 95260
rect 222476 95140 222528 95192
rect 281724 95140 281776 95192
rect 370596 95140 370648 95192
rect 413284 95140 413336 95192
rect 216128 95072 216180 95124
rect 229192 95072 229244 95124
rect 391940 95072 391992 95124
rect 418252 95072 418304 95124
rect 66076 94460 66128 94512
rect 97264 94460 97316 94512
rect 162124 94460 162176 94512
rect 173348 94460 173400 94512
rect 202328 94460 202380 94512
rect 214656 94460 214708 94512
rect 275928 94460 275980 94512
rect 331956 94460 332008 94512
rect 418252 94460 418304 94512
rect 582748 94460 582800 94512
rect 398840 94120 398892 94172
rect 399668 94120 399720 94172
rect 130752 93916 130804 93968
rect 167644 93916 167696 93968
rect 405740 93916 405792 93968
rect 406476 93916 406528 93968
rect 113180 93848 113232 93900
rect 153200 93848 153252 93900
rect 187608 93780 187660 93832
rect 220820 93780 220872 93832
rect 266268 93780 266320 93832
rect 279332 93780 279384 93832
rect 398104 93780 398156 93832
rect 434720 93780 434772 93832
rect 260748 93712 260800 93764
rect 273996 93712 274048 93764
rect 123024 93168 123076 93220
rect 171968 93168 172020 93220
rect 213184 93168 213236 93220
rect 232596 93168 232648 93220
rect 376024 93168 376076 93220
rect 419632 93168 419684 93220
rect 119712 93100 119764 93152
rect 175924 93100 175976 93152
rect 200856 93100 200908 93152
rect 210424 93100 210476 93152
rect 222844 93100 222896 93152
rect 243728 93100 243780 93152
rect 273904 93100 273956 93152
rect 395528 93100 395580 93152
rect 426624 92488 426676 92540
rect 582932 92488 582984 92540
rect 134432 92420 134484 92472
rect 166448 92420 166500 92472
rect 209688 92420 209740 92472
rect 281816 92420 281868 92472
rect 67456 91740 67508 91792
rect 100024 91740 100076 91792
rect 215944 91740 215996 91792
rect 242532 91740 242584 91792
rect 298100 91740 298152 91792
rect 424140 91740 424192 91792
rect 126704 91400 126756 91452
rect 129004 91400 129056 91452
rect 162124 91332 162176 91384
rect 168288 91332 168340 91384
rect 97356 91128 97408 91180
rect 104164 91128 104216 91180
rect 74816 91060 74868 91112
rect 89720 91060 89772 91112
rect 100116 91060 100168 91112
rect 108304 91060 108356 91112
rect 108580 91060 108632 91112
rect 116584 91060 116636 91112
rect 116768 91060 116820 91112
rect 133788 91128 133840 91180
rect 151360 91060 151412 91112
rect 158720 91060 158772 91112
rect 411352 91060 411404 91112
rect 411904 91060 411956 91112
rect 582380 91060 582432 91112
rect 103152 90992 103204 91044
rect 188528 90992 188580 91044
rect 381636 90992 381688 91044
rect 426624 90992 426676 91044
rect 124128 90924 124180 90976
rect 207756 90924 207808 90976
rect 220084 90380 220136 90432
rect 238392 90380 238444 90432
rect 67364 90312 67416 90364
rect 106924 90312 106976 90364
rect 206376 90312 206428 90364
rect 263140 90312 263192 90364
rect 121184 89632 121236 89684
rect 177488 89632 177540 89684
rect 217232 89632 217284 89684
rect 279056 89632 279108 89684
rect 158720 89564 158772 89616
rect 177304 89564 177356 89616
rect 209136 88952 209188 89004
rect 234068 88952 234120 89004
rect 349896 88952 349948 89004
rect 357440 88952 357492 89004
rect 426532 88952 426584 89004
rect 117136 88272 117188 88324
rect 170496 88272 170548 88324
rect 267832 88272 267884 88324
rect 410064 88272 410116 88324
rect 121828 88204 121880 88256
rect 171876 88204 171928 88256
rect 379520 88204 379572 88256
rect 429752 88204 429804 88256
rect 170772 87660 170824 87712
rect 196900 87660 196952 87712
rect 224316 87660 224368 87712
rect 256240 87660 256292 87712
rect 3516 87592 3568 87644
rect 33784 87592 33836 87644
rect 95056 87592 95108 87644
rect 115204 87592 115256 87644
rect 196808 87592 196860 87644
rect 247960 87592 248012 87644
rect 304264 87592 304316 87644
rect 379520 87592 379572 87644
rect 108488 86912 108540 86964
rect 189908 86912 189960 86964
rect 257344 86912 257396 86964
rect 257988 86912 258040 86964
rect 402060 86912 402112 86964
rect 152464 86844 152516 86896
rect 169116 86844 169168 86896
rect 214564 86300 214616 86352
rect 229836 86300 229888 86352
rect 181536 86232 181588 86284
rect 261760 86232 261812 86284
rect 397368 86232 397420 86284
rect 583024 86232 583076 86284
rect 582380 86028 582432 86080
rect 582932 86028 582984 86080
rect 115756 85484 115808 85536
rect 193956 85484 194008 85536
rect 203524 85484 203576 85536
rect 280160 85484 280212 85536
rect 151728 85416 151780 85468
rect 166356 85416 166408 85468
rect 63408 84804 63460 84856
rect 115296 84804 115348 84856
rect 210424 84804 210476 84856
rect 245108 84804 245160 84856
rect 309784 84804 309836 84856
rect 441712 84804 441764 84856
rect 126796 84124 126848 84176
rect 167736 84124 167788 84176
rect 189816 84124 189868 84176
rect 428004 84124 428056 84176
rect 114376 84056 114428 84108
rect 203708 84056 203760 84108
rect 57888 83444 57940 83496
rect 98644 83444 98696 83496
rect 213276 83444 213328 83496
rect 252100 83444 252152 83496
rect 324964 83444 325016 83496
rect 441804 83444 441856 83496
rect 86868 82764 86920 82816
rect 164884 82764 164936 82816
rect 313924 82764 313976 82816
rect 435456 82764 435508 82816
rect 198096 82152 198148 82204
rect 232780 82152 232832 82204
rect 160836 82084 160888 82136
rect 213368 82084 213420 82136
rect 216128 82084 216180 82136
rect 249248 82084 249300 82136
rect 359464 82084 359516 82136
rect 441896 82084 441948 82136
rect 95148 81336 95200 81388
rect 173256 81336 173308 81388
rect 204996 81336 205048 81388
rect 281540 81336 281592 81388
rect 347044 81336 347096 81388
rect 408500 81336 408552 81388
rect 119988 81268 120040 81320
rect 170680 81268 170732 81320
rect 331220 80656 331272 80708
rect 340144 80656 340196 80708
rect 355324 80656 355376 80708
rect 111616 79976 111668 80028
rect 172060 79976 172112 80028
rect 200764 79976 200816 80028
rect 411904 79976 411956 80028
rect 125508 79908 125560 79960
rect 178868 79908 178920 79960
rect 337476 79296 337528 79348
rect 440424 79296 440476 79348
rect 124036 78616 124088 78668
rect 166264 78616 166316 78668
rect 270500 78616 270552 78668
rect 271052 78616 271104 78668
rect 438860 78616 438912 78668
rect 240968 78004 241020 78056
rect 271052 78004 271104 78056
rect 34428 77936 34480 77988
rect 241060 77936 241112 77988
rect 100024 77188 100076 77240
rect 170772 77188 170824 77240
rect 132408 77120 132460 77172
rect 176016 77120 176068 77172
rect 246396 76508 246448 76560
rect 404452 76508 404504 76560
rect 97264 75828 97316 75880
rect 170588 75828 170640 75880
rect 151544 75760 151596 75812
rect 181444 75760 181496 75812
rect 278688 75148 278740 75200
rect 448704 75148 448756 75200
rect 129648 74468 129700 74520
rect 210608 74468 210660 74520
rect 91008 74400 91060 74452
rect 160836 74400 160888 74452
rect 218704 73856 218756 73908
rect 239680 73856 239732 73908
rect 160744 73788 160796 73840
rect 218796 73788 218848 73840
rect 106924 73108 106976 73160
rect 214748 73108 214800 73160
rect 114468 73040 114520 73092
rect 174544 73040 174596 73092
rect 301504 72428 301556 72480
rect 398840 72428 398892 72480
rect 118608 71680 118660 71732
rect 195428 71680 195480 71732
rect 102048 71612 102100 71664
rect 178776 71612 178828 71664
rect 129004 70320 129056 70372
rect 171784 70320 171836 70372
rect 119988 69640 120040 69692
rect 251916 69640 251968 69692
rect 289084 69640 289136 69692
rect 383108 69640 383160 69692
rect 85488 68960 85540 69012
rect 169300 68960 169352 69012
rect 322940 68960 322992 69012
rect 323676 68960 323728 69012
rect 416872 68960 416924 69012
rect 126704 68892 126756 68944
rect 199384 68892 199436 68944
rect 67640 67532 67692 67584
rect 187056 67532 187108 67584
rect 93676 67464 93728 67516
rect 205088 67464 205140 67516
rect 330484 66852 330536 66904
rect 441620 66852 441672 66904
rect 115204 66172 115256 66224
rect 207664 66172 207716 66224
rect 122748 66104 122800 66156
rect 170404 66104 170456 66156
rect 332600 65492 332652 65544
rect 352656 65492 352708 65544
rect 104164 64812 104216 64864
rect 192484 64812 192536 64864
rect 331864 64812 331916 64864
rect 401600 64812 401652 64864
rect 121368 64744 121420 64796
rect 173164 64744 173216 64796
rect 318156 64132 318208 64184
rect 331864 64132 331916 64184
rect 108304 63452 108356 63504
rect 193864 63452 193916 63504
rect 355324 63452 355376 63504
rect 436100 63452 436152 63504
rect 68928 62772 68980 62824
rect 253204 62772 253256 62824
rect 308404 62772 308456 62824
rect 353944 62772 353996 62824
rect 111708 62024 111760 62076
rect 200856 62024 200908 62076
rect 73068 61344 73120 61396
rect 262956 61344 263008 61396
rect 288348 61344 288400 61396
rect 419724 61344 419776 61396
rect 99288 60664 99340 60716
rect 198004 60664 198056 60716
rect 271880 60664 271932 60716
rect 359556 60664 359608 60716
rect 269120 60256 269172 60308
rect 271880 60256 271932 60308
rect 70308 59984 70360 60036
rect 245016 59984 245068 60036
rect 3056 59304 3108 59356
rect 11704 59304 11756 59356
rect 103428 59304 103480 59356
rect 184296 59304 184348 59356
rect 66168 58624 66220 58676
rect 260288 58624 260340 58676
rect 271144 58624 271196 58676
rect 423680 58624 423732 58676
rect 104808 57876 104860 57928
rect 202328 57876 202380 57928
rect 91008 57196 91060 57248
rect 264428 57196 264480 57248
rect 112996 56516 113048 56568
rect 182824 56516 182876 56568
rect 97908 55836 97960 55888
rect 256056 55836 256108 55888
rect 260380 55836 260432 55888
rect 381544 55836 381596 55888
rect 381636 55836 381688 55888
rect 447324 55836 447376 55888
rect 107476 55156 107528 55208
rect 203616 55156 203668 55208
rect 311900 55156 311952 55208
rect 405832 55156 405884 55208
rect 244280 54544 244332 54596
rect 311900 54544 311952 54596
rect 102048 54476 102100 54528
rect 250536 54476 250588 54528
rect 125416 53728 125468 53780
rect 216036 53728 216088 53780
rect 89628 53048 89680 53100
rect 258816 53048 258868 53100
rect 115848 52368 115900 52420
rect 195336 52368 195388 52420
rect 104808 51688 104860 51740
rect 267740 51688 267792 51740
rect 339500 51688 339552 51740
rect 430672 51688 430724 51740
rect 110328 51008 110380 51060
rect 189724 51008 189776 51060
rect 241520 51008 241572 51060
rect 249800 51008 249852 51060
rect 433340 51008 433392 51060
rect 108948 50328 109000 50380
rect 242256 50328 242308 50380
rect 128268 49648 128320 49700
rect 180248 49648 180300 49700
rect 111708 48968 111760 49020
rect 243544 48968 243596 49020
rect 247684 48968 247736 49020
rect 414112 48968 414164 49020
rect 337384 48220 337436 48272
rect 437480 48220 437532 48272
rect 336004 48016 336056 48068
rect 337384 48016 337436 48068
rect 33048 47608 33100 47660
rect 240876 47608 240928 47660
rect 67180 47540 67232 47592
rect 280804 47540 280856 47592
rect 285680 47540 285732 47592
rect 334716 47540 334768 47592
rect 74448 46180 74500 46232
rect 262864 46180 262916 46232
rect 321560 46180 321612 46232
rect 408500 46180 408552 46232
rect 44088 44888 44140 44940
rect 211804 44888 211856 44940
rect 41328 44820 41380 44872
rect 225604 44820 225656 44872
rect 314660 44820 314712 44872
rect 444380 44820 444432 44872
rect 84108 43460 84160 43512
rect 253296 43460 253348 43512
rect 29644 43392 29696 43444
rect 265624 43392 265676 43444
rect 279424 43392 279476 43444
rect 415400 43392 415452 43444
rect 62028 42032 62080 42084
rect 264336 42032 264388 42084
rect 268384 42032 268436 42084
rect 449992 42032 450044 42084
rect 115848 40740 115900 40792
rect 249064 40740 249116 40792
rect 259368 40740 259420 40792
rect 430580 40740 430632 40792
rect 38568 40672 38620 40724
rect 269212 40672 269264 40724
rect 30288 39380 30340 39432
rect 181536 39380 181588 39432
rect 13728 39312 13780 39364
rect 244924 39312 244976 39364
rect 339408 38564 339460 38616
rect 418804 38564 418856 38616
rect 333980 37884 334032 37936
rect 338120 37884 338172 37936
rect 339408 37884 339460 37936
rect 209044 37204 209096 37256
rect 258080 37204 258132 37256
rect 259368 37204 259420 37256
rect 122748 36592 122800 36644
rect 206376 36592 206428 36644
rect 16488 36524 16540 36576
rect 235356 36524 235408 36576
rect 276664 36524 276716 36576
rect 414020 36524 414072 36576
rect 320824 35844 320876 35896
rect 395436 35844 395488 35896
rect 130384 35232 130436 35284
rect 213276 35232 213328 35284
rect 71044 35164 71096 35216
rect 239496 35164 239548 35216
rect 320180 34484 320232 34536
rect 320824 34484 320876 34536
rect 191196 33804 191248 33856
rect 280896 33804 280948 33856
rect 70216 33736 70268 33788
rect 218704 33736 218756 33788
rect 2872 33056 2924 33108
rect 40684 33056 40736 33108
rect 85488 32444 85540 32496
rect 246304 32444 246356 32496
rect 60648 32376 60700 32428
rect 275284 32376 275336 32428
rect 275284 31764 275336 31816
rect 276664 31764 276716 31816
rect 57244 31696 57296 31748
rect 278780 31696 278832 31748
rect 279424 31696 279476 31748
rect 112 31016 164 31068
rect 231308 31016 231360 31068
rect 278044 31016 278096 31068
rect 281540 31016 281592 31068
rect 388536 31016 388588 31068
rect 300860 30268 300912 30320
rect 301320 30268 301372 30320
rect 432604 30268 432656 30320
rect 118608 29656 118660 29708
rect 231216 29656 231268 29708
rect 56508 29588 56560 29640
rect 260104 29588 260156 29640
rect 277400 29588 277452 29640
rect 301320 29588 301372 29640
rect 99288 28296 99340 28348
rect 229744 28296 229796 28348
rect 49608 28228 49660 28280
rect 240784 28228 240836 28280
rect 271788 28228 271840 28280
rect 392768 28228 392820 28280
rect 52368 27548 52420 27600
rect 262220 27548 262272 27600
rect 262956 27548 263008 27600
rect 296720 27548 296772 27600
rect 374644 27548 374696 27600
rect 344284 27480 344336 27532
rect 405740 27480 405792 27532
rect 61936 26868 61988 26920
rect 160744 26868 160796 26920
rect 263600 26868 263652 26920
rect 296720 26868 296772 26920
rect 257344 25508 257396 25560
rect 445944 25508 445996 25560
rect 55128 24760 55180 24812
rect 307760 24760 307812 24812
rect 308404 24760 308456 24812
rect 92388 22788 92440 22840
rect 209136 22788 209188 22840
rect 45468 22720 45520 22772
rect 228364 22720 228416 22772
rect 250536 22720 250588 22772
rect 389916 22720 389968 22772
rect 346400 21428 346452 21480
rect 411444 21428 411496 21480
rect 95056 21360 95108 21412
rect 264244 21360 264296 21412
rect 284944 21360 284996 21412
rect 421564 21360 421616 21412
rect 224224 20612 224276 20664
rect 270500 20612 270552 20664
rect 271788 20612 271840 20664
rect 316040 20612 316092 20664
rect 316776 20612 316828 20664
rect 396724 20612 396776 20664
rect 305644 20544 305696 20596
rect 336740 20544 336792 20596
rect 337476 20544 337528 20596
rect 88248 20000 88300 20052
rect 216128 20000 216180 20052
rect 31668 19932 31720 19984
rect 224316 19932 224368 19984
rect 341524 19320 341576 19372
rect 346400 19320 346452 19372
rect 280804 19252 280856 19304
rect 284944 19252 284996 19304
rect 124128 18640 124180 18692
rect 210424 18640 210476 18692
rect 284944 18640 284996 18692
rect 370504 18640 370556 18692
rect 45376 18572 45428 18624
rect 198096 18572 198148 18624
rect 202144 18572 202196 18624
rect 288440 18572 288492 18624
rect 280896 17892 280948 17944
rect 363604 17892 363656 17944
rect 280160 17280 280212 17332
rect 280896 17280 280948 17332
rect 53656 17212 53708 17264
rect 242164 17212 242216 17264
rect 249156 16532 249208 16584
rect 249708 16532 249760 16584
rect 367836 16532 367888 16584
rect 39580 15920 39632 15972
rect 220176 15920 220228 15972
rect 9588 15852 9640 15904
rect 231124 15852 231176 15904
rect 343364 15852 343416 15904
rect 403624 15852 403676 15904
rect 255964 15104 256016 15156
rect 256608 15104 256660 15156
rect 310520 15104 310572 15156
rect 311440 14492 311492 14544
rect 360844 14492 360896 14544
rect 100668 14424 100720 14476
rect 258724 14424 258776 14476
rect 328736 14424 328788 14476
rect 382924 14424 382976 14476
rect 295340 13744 295392 13796
rect 295892 13744 295944 13796
rect 400312 13744 400364 13796
rect 96252 13132 96304 13184
rect 235264 13132 235316 13184
rect 54944 13064 54996 13116
rect 238116 13064 238168 13116
rect 299664 13064 299716 13116
rect 454040 13064 454092 13116
rect 264980 12452 265032 12504
rect 295340 12452 295392 12504
rect 251824 12384 251876 12436
rect 276112 12384 276164 12436
rect 277492 12384 277544 12436
rect 443000 12384 443052 12436
rect 385776 12316 385828 12368
rect 251180 11908 251232 11960
rect 251824 11908 251876 11960
rect 126888 11772 126940 11824
rect 217324 11772 217376 11824
rect 12164 11704 12216 11756
rect 233976 11704 234028 11756
rect 242900 11704 242952 11756
rect 244096 11704 244148 11756
rect 135260 11636 135312 11688
rect 136456 11636 136508 11688
rect 288440 10956 288492 11008
rect 288992 10956 289044 11008
rect 377496 10956 377548 11008
rect 81348 10344 81400 10396
rect 213184 10344 213236 10396
rect 24768 10276 24820 10328
rect 222936 10276 222988 10328
rect 261760 9596 261812 9648
rect 447140 9596 447192 9648
rect 85672 8984 85724 9036
rect 220084 8984 220136 9036
rect 59636 8916 59688 8968
rect 250444 8916 250496 8968
rect 345664 8236 345716 8288
rect 394148 8236 394200 8288
rect 114008 7624 114060 7676
rect 214564 7624 214616 7676
rect 66720 7556 66772 7608
rect 261484 7556 261536 7608
rect 342168 7556 342220 7608
rect 356704 7556 356756 7608
rect 325056 6808 325108 6860
rect 409880 6808 409932 6860
rect 318064 6740 318116 6792
rect 319444 6740 319496 6792
rect 121092 6196 121144 6248
rect 239404 6196 239456 6248
rect 58440 6128 58492 6180
rect 215944 6128 215996 6180
rect 298468 6128 298520 6180
rect 378876 6128 378928 6180
rect 324412 5516 324464 5568
rect 325056 5516 325108 5568
rect 316684 5448 316736 5500
rect 317328 5448 317380 5500
rect 425888 5448 425940 5500
rect 109316 4768 109368 4820
rect 238024 4768 238076 4820
rect 246212 4768 246264 4820
rect 407120 4768 407172 4820
rect 232504 4156 232556 4208
rect 235816 4156 235868 4208
rect 278688 4156 278740 4208
rect 283104 4156 283156 4208
rect 191104 4088 191156 4140
rect 247592 4088 247644 4140
rect 254676 4088 254728 4140
rect 258080 4088 258132 4140
rect 291844 4088 291896 4140
rect 301504 4088 301556 4140
rect 307116 4088 307168 4140
rect 307944 4088 307996 4140
rect 309876 4088 309928 4140
rect 289084 4020 289136 4072
rect 292580 4020 292632 4072
rect 306748 4020 306800 4072
rect 342904 4088 342956 4140
rect 348424 4088 348476 4140
rect 429844 4088 429896 4140
rect 332692 4020 332744 4072
rect 336004 4020 336056 4072
rect 312636 3952 312688 4004
rect 318156 3952 318208 4004
rect 291384 3680 291436 3732
rect 291844 3680 291896 3732
rect 11152 3544 11204 3596
rect 12256 3544 12308 3596
rect 27712 3544 27764 3596
rect 28908 3544 28960 3596
rect 44272 3544 44324 3596
rect 45376 3544 45428 3596
rect 64328 3544 64380 3596
rect 64788 3544 64840 3596
rect 8760 3476 8812 3528
rect 9588 3476 9640 3528
rect 9956 3476 10008 3528
rect 10968 3476 11020 3528
rect 15936 3476 15988 3528
rect 16488 3476 16540 3528
rect 17040 3476 17092 3528
rect 17868 3476 17920 3528
rect 18236 3476 18288 3528
rect 19248 3476 19300 3528
rect 24216 3476 24268 3528
rect 24768 3476 24820 3528
rect 20536 3408 20588 3460
rect 36544 3476 36596 3528
rect 40684 3476 40736 3528
rect 41328 3476 41380 3528
rect 41880 3476 41932 3528
rect 42708 3476 42760 3528
rect 43076 3476 43128 3528
rect 44088 3476 44140 3528
rect 48964 3476 49016 3528
rect 49608 3476 49660 3528
rect 50160 3476 50212 3528
rect 50988 3476 51040 3528
rect 52552 3476 52604 3528
rect 53656 3476 53708 3528
rect 56048 3476 56100 3528
rect 56508 3476 56560 3528
rect 57244 3476 57296 3528
rect 57888 3476 57940 3528
rect 63224 3476 63276 3528
rect 71044 3612 71096 3664
rect 351184 3612 351236 3664
rect 351644 3612 351696 3664
rect 69112 3544 69164 3596
rect 70216 3544 70268 3596
rect 119896 3544 119948 3596
rect 122104 3544 122156 3596
rect 276020 3544 276072 3596
rect 277124 3544 277176 3596
rect 65524 3476 65576 3528
rect 66168 3476 66220 3528
rect 67916 3476 67968 3528
rect 68928 3476 68980 3528
rect 72608 3476 72660 3528
rect 73068 3476 73120 3528
rect 73804 3476 73856 3528
rect 74448 3476 74500 3528
rect 75000 3476 75052 3528
rect 75828 3476 75880 3528
rect 76196 3476 76248 3528
rect 77208 3476 77260 3528
rect 80888 3476 80940 3528
rect 81348 3476 81400 3528
rect 90364 3476 90416 3528
rect 91008 3476 91060 3528
rect 91560 3476 91612 3528
rect 92388 3476 92440 3528
rect 92756 3476 92808 3528
rect 93768 3476 93820 3528
rect 93952 3476 94004 3528
rect 95056 3476 95108 3528
rect 97448 3476 97500 3528
rect 97908 3476 97960 3528
rect 98644 3476 98696 3528
rect 99288 3476 99340 3528
rect 99840 3476 99892 3528
rect 100668 3476 100720 3528
rect 101036 3476 101088 3528
rect 102048 3476 102100 3528
rect 105728 3476 105780 3528
rect 106188 3476 106240 3528
rect 106924 3476 106976 3528
rect 107568 3476 107620 3528
rect 108120 3476 108172 3528
rect 108948 3476 109000 3528
rect 110512 3476 110564 3528
rect 111708 3476 111760 3528
rect 115204 3476 115256 3528
rect 115848 3476 115900 3528
rect 116400 3476 116452 3528
rect 117228 3476 117280 3528
rect 117596 3476 117648 3528
rect 118608 3476 118660 3528
rect 118792 3476 118844 3528
rect 119988 3476 120040 3528
rect 122288 3476 122340 3528
rect 122748 3476 122800 3528
rect 123484 3476 123536 3528
rect 124128 3476 124180 3528
rect 124680 3476 124732 3528
rect 125508 3476 125560 3528
rect 125876 3476 125928 3528
rect 126888 3476 126940 3528
rect 140044 3476 140096 3528
rect 141424 3476 141476 3528
rect 143540 3476 143592 3528
rect 144828 3476 144880 3528
rect 240508 3476 240560 3528
rect 246396 3476 246448 3528
rect 248788 3476 248840 3528
rect 249708 3476 249760 3528
rect 252376 3476 252428 3528
rect 253204 3476 253256 3528
rect 266360 3476 266412 3528
rect 266544 3476 266596 3528
rect 271144 3476 271196 3528
rect 274824 3476 274876 3528
rect 275284 3476 275336 3528
rect 284300 3476 284352 3528
rect 285036 3476 285088 3528
rect 303528 3476 303580 3528
rect 305552 3476 305604 3528
rect 332600 3476 332652 3528
rect 333888 3476 333940 3528
rect 582196 3476 582248 3528
rect 583208 3476 583260 3528
rect 26516 3408 26568 3460
rect 27528 3408 27580 3460
rect 28908 3408 28960 3460
rect 29644 3408 29696 3460
rect 32404 3408 32456 3460
rect 33048 3408 33100 3460
rect 33600 3408 33652 3460
rect 34428 3408 34480 3460
rect 34796 3408 34848 3460
rect 35808 3408 35860 3460
rect 37096 3408 37148 3460
rect 87604 3408 87656 3460
rect 102232 3408 102284 3460
rect 130384 3408 130436 3460
rect 267740 3408 267792 3460
rect 268844 3408 268896 3460
rect 349252 3408 349304 3460
rect 357440 3408 357492 3460
rect 35992 3272 36044 3324
rect 37188 3272 37240 3324
rect 89168 3272 89220 3324
rect 89628 3272 89680 3324
rect 267740 3272 267792 3324
rect 281632 3272 281684 3324
rect 84476 3204 84528 3256
rect 85488 3204 85540 3256
rect 324964 3204 325016 3256
rect 325608 3204 325660 3256
rect 341524 3204 341576 3256
rect 344560 3204 344612 3256
rect 83280 3136 83332 3188
rect 84108 3136 84160 3188
rect 299388 3136 299440 3188
rect 301964 3136 302016 3188
rect 60832 3000 60884 3052
rect 61936 3000 61988 3052
rect 82084 3000 82136 3052
rect 82728 3000 82780 3052
rect 581000 3000 581052 3052
rect 582840 3000 582892 3052
rect 19432 2932 19484 2984
rect 20628 2932 20680 2984
rect 129372 2932 129424 2984
rect 133144 2932 133196 2984
rect 239312 2932 239364 2984
rect 240968 2932 241020 2984
rect 272432 2932 272484 2984
rect 273996 2932 274048 2984
rect 242900 2728 242952 2780
rect 412640 2728 412692 2780
rect 51356 2116 51408 2168
rect 58624 2116 58676 2168
rect 111616 2116 111668 2168
rect 222844 2116 222896 2168
rect 7656 2048 7708 2100
rect 54484 2048 54536 2100
rect 71504 2048 71556 2100
rect 233884 2048 233936 2100
rect 350448 2048 350500 2100
rect 381636 2048 381688 2100
rect 307760 552 307812 604
rect 309048 552 309100 604
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40052 703582 40356 703610
rect 8128 702506 8156 703520
rect 24320 702642 24348 703520
rect 24308 702636 24360 702642
rect 24308 702578 24360 702584
rect 8116 702500 8168 702506
rect 8116 702442 8168 702448
rect 3422 684312 3478 684321
rect 3422 684247 3478 684256
rect 3436 683194 3464 684247
rect 3424 683188 3476 683194
rect 3424 683130 3476 683136
rect 21364 683188 21416 683194
rect 21364 683130 21416 683136
rect 3514 671256 3570 671265
rect 3514 671191 3570 671200
rect 3528 670750 3556 671191
rect 3516 670744 3568 670750
rect 3516 670686 3568 670692
rect 3422 658200 3478 658209
rect 3422 658135 3478 658144
rect 3436 592686 3464 658135
rect 3516 632120 3568 632126
rect 3514 632088 3516 632097
rect 11704 632120 11756 632126
rect 3568 632088 3570 632097
rect 11704 632062 11756 632068
rect 3514 632023 3570 632032
rect 3514 619168 3570 619177
rect 3514 619103 3570 619112
rect 3528 618322 3556 619103
rect 3516 618316 3568 618322
rect 3516 618258 3568 618264
rect 3514 606112 3570 606121
rect 3514 606047 3570 606056
rect 3528 605878 3556 606047
rect 3516 605872 3568 605878
rect 3516 605814 3568 605820
rect 3424 592680 3476 592686
rect 3424 592622 3476 592628
rect 3424 589348 3476 589354
rect 3424 589290 3476 589296
rect 3436 580009 3464 589290
rect 3422 580000 3478 580009
rect 3422 579935 3478 579944
rect 11716 576162 11744 632062
rect 14464 618316 14516 618322
rect 14464 618258 14516 618264
rect 11704 576156 11756 576162
rect 11704 576098 11756 576104
rect 3422 566944 3478 566953
rect 3422 566879 3478 566888
rect 3330 553888 3386 553897
rect 3330 553823 3386 553832
rect 3344 553450 3372 553823
rect 3332 553444 3384 553450
rect 3332 553386 3384 553392
rect 3436 540258 3464 566879
rect 3424 540252 3476 540258
rect 3424 540194 3476 540200
rect 8208 537532 8260 537538
rect 8208 537474 8260 537480
rect 3424 532024 3476 532030
rect 3424 531966 3476 531972
rect 3436 527921 3464 531966
rect 3422 527912 3478 527921
rect 3422 527847 3478 527856
rect 3330 475688 3386 475697
rect 3330 475623 3386 475632
rect 3344 475386 3372 475623
rect 3332 475380 3384 475386
rect 3332 475322 3384 475328
rect 3436 451926 3464 527847
rect 3514 514856 3570 514865
rect 3514 514791 3516 514800
rect 3568 514791 3570 514800
rect 3516 514762 3568 514768
rect 3516 502308 3568 502314
rect 3516 502250 3568 502256
rect 3528 501809 3556 502250
rect 3514 501800 3570 501809
rect 3514 501735 3570 501744
rect 8220 475386 8248 537474
rect 14476 536081 14504 618258
rect 21376 543046 21404 683130
rect 22744 670744 22796 670750
rect 22744 670686 22796 670692
rect 21364 543040 21416 543046
rect 21364 542982 21416 542988
rect 22756 541686 22784 670686
rect 40052 594114 40080 703582
rect 40328 703474 40356 703582
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 412652 703582 413508 703610
rect 40512 703474 40540 703520
rect 40328 703446 40540 703474
rect 62028 702976 62080 702982
rect 62028 702918 62080 702924
rect 40040 594108 40092 594114
rect 40040 594050 40092 594056
rect 52276 587920 52328 587926
rect 52276 587862 52328 587868
rect 50988 582412 51040 582418
rect 50988 582354 51040 582360
rect 49608 571396 49660 571402
rect 49608 571338 49660 571344
rect 37188 561740 37240 561746
rect 37188 561682 37240 561688
rect 34520 543040 34572 543046
rect 34520 542982 34572 542988
rect 34532 542434 34560 542982
rect 34520 542428 34572 542434
rect 34520 542370 34572 542376
rect 35808 542428 35860 542434
rect 35808 542370 35860 542376
rect 22744 541680 22796 541686
rect 22744 541622 22796 541628
rect 17224 538892 17276 538898
rect 17224 538834 17276 538840
rect 14462 536072 14518 536081
rect 14462 536007 14518 536016
rect 14464 514820 14516 514826
rect 14464 514762 14516 514768
rect 8208 475380 8260 475386
rect 8208 475322 8260 475328
rect 3514 462632 3570 462641
rect 3514 462567 3570 462576
rect 3528 462398 3556 462567
rect 3516 462392 3568 462398
rect 3516 462334 3568 462340
rect 14476 459542 14504 514762
rect 15844 475380 15896 475386
rect 15844 475322 15896 475328
rect 14464 459536 14516 459542
rect 14464 459478 14516 459484
rect 3424 451920 3476 451926
rect 3424 451862 3476 451868
rect 3146 449576 3202 449585
rect 3146 449511 3202 449520
rect 3160 448594 3188 449511
rect 3148 448588 3200 448594
rect 3148 448530 3200 448536
rect 4804 444440 4856 444446
rect 4804 444382 4856 444388
rect 3146 423600 3202 423609
rect 3146 423535 3202 423544
rect 3160 422958 3188 423535
rect 3148 422952 3200 422958
rect 3148 422894 3200 422900
rect 3422 410544 3478 410553
rect 3422 410479 3478 410488
rect 2780 398744 2832 398750
rect 2780 398686 2832 398692
rect 2792 397497 2820 398686
rect 2778 397488 2834 397497
rect 2778 397423 2834 397432
rect 3436 391270 3464 410479
rect 4816 398750 4844 444382
rect 14464 428460 14516 428466
rect 14464 428402 14516 428408
rect 4804 398744 4856 398750
rect 4804 398686 4856 398692
rect 3424 391264 3476 391270
rect 3424 391206 3476 391212
rect 7562 387016 7618 387025
rect 7562 386951 7618 386960
rect 4802 385656 4858 385665
rect 4802 385591 4858 385600
rect 3516 380928 3568 380934
rect 3516 380870 3568 380876
rect 3240 371408 3292 371414
rect 3238 371376 3240 371385
rect 3292 371376 3294 371385
rect 3238 371311 3294 371320
rect 3330 359000 3386 359009
rect 3330 358935 3386 358944
rect 3344 354674 3372 358935
rect 3424 358624 3476 358630
rect 3424 358566 3476 358572
rect 3436 358465 3464 358566
rect 3422 358456 3478 358465
rect 3422 358391 3478 358400
rect 3344 354646 3464 354674
rect 20 336048 72 336054
rect 20 335990 72 335996
rect 32 6769 60 335990
rect 2780 254244 2832 254250
rect 2780 254186 2832 254192
rect 2792 254153 2820 254186
rect 2778 254144 2834 254153
rect 2778 254079 2834 254088
rect 3332 215280 3384 215286
rect 3332 215222 3384 215228
rect 3344 214985 3372 215222
rect 3330 214976 3386 214985
rect 3330 214911 3386 214920
rect 3056 202836 3108 202842
rect 3056 202778 3108 202784
rect 3068 201929 3096 202778
rect 3054 201920 3110 201929
rect 3054 201855 3110 201864
rect 2780 150340 2832 150346
rect 2780 150282 2832 150288
rect 2792 149841 2820 150282
rect 2778 149832 2834 149841
rect 2778 149767 2834 149776
rect 3148 111784 3200 111790
rect 3148 111726 3200 111732
rect 3160 110673 3188 111726
rect 3146 110664 3202 110673
rect 3146 110599 3202 110608
rect 3056 59356 3108 59362
rect 3056 59298 3108 59304
rect 3068 58585 3096 59298
rect 3054 58576 3110 58585
rect 3054 58511 3110 58520
rect 2872 33108 2924 33114
rect 2872 33050 2924 33056
rect 2884 32473 2912 33050
rect 2870 32464 2926 32473
rect 2870 32399 2926 32408
rect 112 31068 164 31074
rect 112 31010 164 31016
rect 18 6760 74 6769
rect 18 6695 74 6704
rect 124 490 152 31010
rect 3436 19417 3464 354646
rect 3528 345409 3556 380870
rect 4816 371414 4844 385591
rect 4804 371408 4856 371414
rect 4804 371350 4856 371356
rect 3514 345400 3570 345409
rect 3514 345335 3570 345344
rect 4816 321570 4844 371350
rect 7576 358630 7604 386951
rect 7564 358624 7616 358630
rect 7564 358566 7616 358572
rect 7564 329860 7616 329866
rect 7564 329802 7616 329808
rect 4804 321564 4856 321570
rect 4804 321506 4856 321512
rect 4066 319288 4122 319297
rect 4066 319223 4122 319232
rect 4080 318782 4108 319223
rect 4068 318776 4120 318782
rect 4068 318718 4120 318724
rect 3516 306332 3568 306338
rect 3516 306274 3568 306280
rect 3528 306241 3556 306274
rect 3514 306232 3570 306241
rect 3514 306167 3570 306176
rect 3514 293176 3570 293185
rect 3514 293111 3570 293120
rect 3528 292602 3556 293111
rect 3516 292596 3568 292602
rect 3516 292538 3568 292544
rect 4080 276690 4108 318718
rect 4804 310548 4856 310554
rect 4804 310490 4856 310496
rect 4068 276684 4120 276690
rect 4068 276626 4120 276632
rect 3514 267200 3570 267209
rect 3514 267135 3570 267144
rect 3528 267034 3556 267135
rect 3516 267028 3568 267034
rect 3516 266970 3568 266976
rect 4816 254250 4844 310490
rect 4804 254244 4856 254250
rect 4804 254186 4856 254192
rect 7576 241126 7604 329802
rect 11704 328500 11756 328506
rect 11704 328442 11756 328448
rect 3516 241120 3568 241126
rect 3514 241088 3516 241097
rect 7564 241120 7616 241126
rect 3568 241088 3570 241097
rect 7564 241062 7616 241068
rect 3514 241023 3570 241032
rect 4804 236020 4856 236026
rect 4804 235962 4856 235968
rect 3516 189032 3568 189038
rect 3516 188974 3568 188980
rect 3528 188873 3556 188974
rect 3514 188864 3570 188873
rect 3514 188799 3570 188808
rect 3516 164892 3568 164898
rect 3516 164834 3568 164840
rect 3528 162897 3556 164834
rect 3514 162888 3570 162897
rect 3514 162823 3570 162832
rect 4816 150346 4844 235962
rect 4804 150340 4856 150346
rect 4804 150282 4856 150288
rect 3516 137964 3568 137970
rect 3516 137906 3568 137912
rect 3528 136785 3556 137906
rect 3514 136776 3570 136785
rect 3514 136711 3570 136720
rect 3516 97980 3568 97986
rect 3516 97922 3568 97928
rect 3528 97617 3556 97922
rect 3514 97608 3570 97617
rect 3514 97543 3570 97552
rect 3516 87644 3568 87650
rect 3516 87586 3568 87592
rect 3528 84697 3556 87586
rect 3514 84688 3570 84697
rect 3514 84623 3570 84632
rect 5446 79520 5502 79529
rect 5446 79455 5502 79464
rect 4066 21312 4122 21321
rect 4066 21247 4122 21256
rect 3422 19408 3478 19417
rect 3422 19343 3478 19352
rect 1674 4856 1730 4865
rect 1674 4791 1730 4800
rect 400 598 612 626
rect 400 490 428 598
rect 124 462 428 490
rect 584 480 612 598
rect 1688 480 1716 4791
rect 2870 3360 2926 3369
rect 2870 3295 2926 3304
rect 2884 480 2912 3295
rect 4080 480 4108 21247
rect 5460 6914 5488 79455
rect 11716 59362 11744 328442
rect 14476 267034 14504 428402
rect 15856 389230 15884 475322
rect 17236 422958 17264 538834
rect 18604 534744 18656 534750
rect 18604 534686 18656 534692
rect 18616 502314 18644 534686
rect 34428 520940 34480 520946
rect 34428 520882 34480 520888
rect 18604 502308 18656 502314
rect 18604 502250 18656 502256
rect 25504 462392 25556 462398
rect 25504 462334 25556 462340
rect 25516 449886 25544 462334
rect 25504 449880 25556 449886
rect 25504 449822 25556 449828
rect 18604 448588 18656 448594
rect 18604 448530 18656 448536
rect 17224 422952 17276 422958
rect 17224 422894 17276 422900
rect 15844 389224 15896 389230
rect 15844 389166 15896 389172
rect 17236 383654 17264 422894
rect 17224 383648 17276 383654
rect 17224 383590 17276 383596
rect 18616 372609 18644 448530
rect 18602 372600 18658 372609
rect 18602 372535 18658 372544
rect 18616 371385 18644 372535
rect 18602 371376 18658 371385
rect 18602 371311 18658 371320
rect 19246 371376 19302 371385
rect 19246 371311 19302 371320
rect 16486 340096 16542 340105
rect 16486 340031 16542 340040
rect 14464 267028 14516 267034
rect 14464 266970 14516 266976
rect 14476 233238 14504 266970
rect 14464 233232 14516 233238
rect 14464 233174 14516 233180
rect 16500 193225 16528 340031
rect 17868 295384 17920 295390
rect 17868 295326 17920 295332
rect 17880 195090 17908 295326
rect 19260 293962 19288 371311
rect 22744 327752 22796 327758
rect 22744 327694 22796 327700
rect 19248 293956 19300 293962
rect 19248 293898 19300 293904
rect 18604 292596 18656 292602
rect 18604 292538 18656 292544
rect 18616 240786 18644 292538
rect 18604 240780 18656 240786
rect 18604 240722 18656 240728
rect 17224 195084 17276 195090
rect 17224 195026 17276 195032
rect 17868 195084 17920 195090
rect 17868 195026 17920 195032
rect 15842 193216 15898 193225
rect 15842 193151 15898 193160
rect 16486 193216 16542 193225
rect 16486 193151 16542 193160
rect 15856 97986 15884 193151
rect 17236 164898 17264 195026
rect 17880 194614 17908 195026
rect 17868 194608 17920 194614
rect 17868 194550 17920 194556
rect 17224 164892 17276 164898
rect 17224 164834 17276 164840
rect 22756 137970 22784 327694
rect 29644 316736 29696 316742
rect 29644 316678 29696 316684
rect 29656 189038 29684 316678
rect 32404 309800 32456 309806
rect 32404 309742 32456 309748
rect 29644 189032 29696 189038
rect 29644 188974 29696 188980
rect 22744 137964 22796 137970
rect 22744 137906 22796 137912
rect 15844 97980 15896 97986
rect 15844 97922 15896 97928
rect 12346 80744 12402 80753
rect 12346 80679 12402 80688
rect 11704 59356 11756 59362
rect 11704 59298 11756 59304
rect 10966 55856 11022 55865
rect 10966 55791 11022 55800
rect 6826 38040 6882 38049
rect 6826 37975 6882 37984
rect 6840 6914 6868 37975
rect 9588 15904 9640 15910
rect 9588 15846 9640 15852
rect 5276 6886 5488 6914
rect 6472 6886 6868 6914
rect 5276 480 5304 6886
rect 6472 480 6500 6886
rect 9600 3534 9628 15846
rect 10980 3534 11008 55791
rect 12164 11756 12216 11762
rect 12164 11698 12216 11704
rect 11152 3596 11204 3602
rect 11152 3538 11204 3544
rect 8760 3528 8812 3534
rect 8760 3470 8812 3476
rect 9588 3528 9640 3534
rect 9588 3470 9640 3476
rect 9956 3528 10008 3534
rect 9956 3470 10008 3476
rect 10968 3528 11020 3534
rect 10968 3470 11020 3476
rect 7656 2100 7708 2106
rect 7656 2042 7708 2048
rect 7668 480 7696 2042
rect 8772 480 8800 3470
rect 9968 480 9996 3470
rect 11164 480 11192 3538
rect 12176 3482 12204 11698
rect 12360 6914 12388 80679
rect 17866 77888 17922 77897
rect 17866 77823 17922 77832
rect 15106 69592 15162 69601
rect 15106 69527 15162 69536
rect 13728 39364 13780 39370
rect 13728 39306 13780 39312
rect 13740 6914 13768 39306
rect 15120 6914 15148 69527
rect 16488 36576 16540 36582
rect 16488 36518 16540 36524
rect 12268 6886 12388 6914
rect 13556 6886 13768 6914
rect 14752 6886 15148 6914
rect 12268 3602 12296 6886
rect 12256 3596 12308 3602
rect 12256 3538 12308 3544
rect 12176 3454 12388 3482
rect 12360 480 12388 3454
rect 13556 480 13584 6886
rect 14752 480 14780 6886
rect 16500 3534 16528 36518
rect 17880 3534 17908 77823
rect 19154 75168 19210 75177
rect 19154 75103 19210 75112
rect 19168 74534 19196 75103
rect 19168 74506 19288 74534
rect 19260 3534 19288 74506
rect 22006 72584 22062 72593
rect 22006 72519 22062 72528
rect 20626 25528 20682 25537
rect 20626 25463 20682 25472
rect 15936 3528 15988 3534
rect 15936 3470 15988 3476
rect 16488 3528 16540 3534
rect 16488 3470 16540 3476
rect 17040 3528 17092 3534
rect 17040 3470 17092 3476
rect 17868 3528 17920 3534
rect 17868 3470 17920 3476
rect 18236 3528 18288 3534
rect 18236 3470 18288 3476
rect 19248 3528 19300 3534
rect 19248 3470 19300 3476
rect 15948 480 15976 3470
rect 17052 480 17080 3470
rect 18248 480 18276 3470
rect 20536 3460 20588 3466
rect 20536 3402 20588 3408
rect 19432 2984 19484 2990
rect 19432 2926 19484 2932
rect 19444 480 19472 2926
rect 20548 1714 20576 3402
rect 20640 2990 20668 25463
rect 22020 6914 22048 72519
rect 32416 71777 32444 309742
rect 34336 280220 34388 280226
rect 34336 280162 34388 280168
rect 34348 191826 34376 280162
rect 34440 274650 34468 520882
rect 35820 396778 35848 542370
rect 37200 429146 37228 561682
rect 44088 560312 44140 560318
rect 44088 560254 44140 560260
rect 39948 558204 40000 558210
rect 39948 558146 40000 558152
rect 36728 429140 36780 429146
rect 36728 429082 36780 429088
rect 37188 429140 37240 429146
rect 37188 429082 37240 429088
rect 36740 428466 36768 429082
rect 36728 428460 36780 428466
rect 36728 428402 36780 428408
rect 39960 421598 39988 558146
rect 43444 553444 43496 553450
rect 43444 553386 43496 553392
rect 43456 536790 43484 553386
rect 43444 536784 43496 536790
rect 43444 536726 43496 536732
rect 44100 531282 44128 560254
rect 48228 543788 48280 543794
rect 48228 543730 48280 543736
rect 45466 536072 45522 536081
rect 45466 536007 45522 536016
rect 44088 531276 44140 531282
rect 44088 531218 44140 531224
rect 44100 528554 44128 531218
rect 44008 528526 44128 528554
rect 41328 511284 41380 511290
rect 41328 511226 41380 511232
rect 41236 435396 41288 435402
rect 41236 435338 41288 435344
rect 39948 421592 40000 421598
rect 39948 421534 40000 421540
rect 35808 396772 35860 396778
rect 35808 396714 35860 396720
rect 39304 380180 39356 380186
rect 39304 380122 39356 380128
rect 36544 330540 36596 330546
rect 36544 330482 36596 330488
rect 35162 329896 35218 329905
rect 35162 329831 35218 329840
rect 34428 274644 34480 274650
rect 34428 274586 34480 274592
rect 35176 215286 35204 329831
rect 36556 306338 36584 330482
rect 39316 318782 39344 380122
rect 41248 378078 41276 435338
rect 41236 378072 41288 378078
rect 41236 378014 41288 378020
rect 39304 318776 39356 318782
rect 39304 318718 39356 318724
rect 39948 311160 40000 311166
rect 39948 311102 40000 311108
rect 39960 310554 39988 311102
rect 39948 310548 40000 310554
rect 39948 310490 40000 310496
rect 36544 306332 36596 306338
rect 36544 306274 36596 306280
rect 39960 217977 39988 310490
rect 41248 298110 41276 378014
rect 41236 298104 41288 298110
rect 41236 298046 41288 298052
rect 41340 240145 41368 511226
rect 44008 427106 44036 528526
rect 44088 433356 44140 433362
rect 44088 433298 44140 433304
rect 43996 427100 44048 427106
rect 43996 427042 44048 427048
rect 43444 276684 43496 276690
rect 43444 276626 43496 276632
rect 43456 261526 43484 276626
rect 43444 261520 43496 261526
rect 43444 261462 43496 261468
rect 41326 240136 41382 240145
rect 41326 240071 41382 240080
rect 44100 232558 44128 433298
rect 45480 385014 45508 536007
rect 46848 507136 46900 507142
rect 46848 507078 46900 507084
rect 45468 385008 45520 385014
rect 45468 384950 45520 384956
rect 46860 285666 46888 507078
rect 48136 403640 48188 403646
rect 48136 403582 48188 403588
rect 48148 383654 48176 403582
rect 48240 398886 48268 543730
rect 49620 446418 49648 571338
rect 50896 545148 50948 545154
rect 50896 545090 50948 545096
rect 50908 527134 50936 545090
rect 50896 527128 50948 527134
rect 50896 527070 50948 527076
rect 50802 517576 50858 517585
rect 50802 517511 50858 517520
rect 50816 447817 50844 517511
rect 50802 447808 50858 447817
rect 50802 447743 50858 447752
rect 49608 446412 49660 446418
rect 49608 446354 49660 446360
rect 49608 440904 49660 440910
rect 49608 440846 49660 440852
rect 48228 398880 48280 398886
rect 48228 398822 48280 398828
rect 48148 383626 48268 383654
rect 48240 379574 48268 383626
rect 48228 379568 48280 379574
rect 48228 379510 48280 379516
rect 48136 300144 48188 300150
rect 48136 300086 48188 300092
rect 46848 285660 46900 285666
rect 46848 285602 46900 285608
rect 44088 232552 44140 232558
rect 44088 232494 44140 232500
rect 39946 217968 40002 217977
rect 39946 217903 40002 217912
rect 35164 215280 35216 215286
rect 35164 215222 35216 215228
rect 48148 208350 48176 300086
rect 48240 245614 48268 379510
rect 49620 331226 49648 440846
rect 50908 400246 50936 527070
rect 51000 518129 51028 582354
rect 50986 518120 51042 518129
rect 50986 518055 51042 518064
rect 51000 517585 51028 518055
rect 50986 517576 51042 517585
rect 50986 517511 51042 517520
rect 50988 462392 51040 462398
rect 50988 462334 51040 462340
rect 50896 400240 50948 400246
rect 50896 400182 50948 400188
rect 50896 398880 50948 398886
rect 50896 398822 50948 398828
rect 50908 378146 50936 398822
rect 50896 378140 50948 378146
rect 50896 378082 50948 378088
rect 49608 331220 49660 331226
rect 49608 331162 49660 331168
rect 49620 330546 49648 331162
rect 49608 330540 49660 330546
rect 49608 330482 49660 330488
rect 49608 295452 49660 295458
rect 49608 295394 49660 295400
rect 48228 245608 48280 245614
rect 48228 245550 48280 245556
rect 49620 214577 49648 295394
rect 50804 271924 50856 271930
rect 50804 271866 50856 271872
rect 49606 214568 49662 214577
rect 49606 214503 49662 214512
rect 48136 208344 48188 208350
rect 48136 208286 48188 208292
rect 40682 203552 40738 203561
rect 40682 203487 40738 203496
rect 33784 191820 33836 191826
rect 33784 191762 33836 191768
rect 34336 191820 34388 191826
rect 34336 191762 34388 191768
rect 33796 87650 33824 191762
rect 35162 178664 35218 178673
rect 35162 178599 35218 178608
rect 35176 111790 35204 178599
rect 35164 111784 35216 111790
rect 35164 111726 35216 111732
rect 33784 87644 33836 87650
rect 33784 87586 33836 87592
rect 36542 79384 36598 79393
rect 36542 79319 36598 79328
rect 34428 77988 34480 77994
rect 34428 77930 34480 77936
rect 32402 71768 32458 71777
rect 32402 71703 32458 71712
rect 23386 54496 23442 54505
rect 23386 54431 23442 54440
rect 23400 6914 23428 54431
rect 28906 50280 28962 50289
rect 28906 50215 28962 50224
rect 27526 48920 27582 48929
rect 27526 48855 27582 48864
rect 24768 10328 24820 10334
rect 24768 10270 24820 10276
rect 21836 6886 22048 6914
rect 23032 6886 23428 6914
rect 20628 2984 20680 2990
rect 20628 2926 20680 2932
rect 20548 1686 20668 1714
rect 20640 480 20668 1686
rect 21836 480 21864 6886
rect 23032 480 23060 6886
rect 24780 3534 24808 10270
rect 25318 6216 25374 6225
rect 25318 6151 25374 6160
rect 24216 3528 24268 3534
rect 24216 3470 24268 3476
rect 24768 3528 24820 3534
rect 24768 3470 24820 3476
rect 24228 480 24256 3470
rect 25332 480 25360 6151
rect 27540 3466 27568 48855
rect 28920 3602 28948 50215
rect 33048 47660 33100 47666
rect 33048 47602 33100 47608
rect 29644 43444 29696 43450
rect 29644 43386 29696 43392
rect 27712 3596 27764 3602
rect 27712 3538 27764 3544
rect 28908 3596 28960 3602
rect 28908 3538 28960 3544
rect 26516 3460 26568 3466
rect 26516 3402 26568 3408
rect 27528 3460 27580 3466
rect 27528 3402 27580 3408
rect 26528 480 26556 3402
rect 27724 480 27752 3538
rect 29656 3466 29684 43386
rect 30288 39432 30340 39438
rect 30288 39374 30340 39380
rect 30300 6914 30328 39374
rect 31668 19984 31720 19990
rect 31668 19926 31720 19932
rect 31680 6914 31708 19926
rect 30116 6886 30328 6914
rect 31312 6886 31708 6914
rect 28908 3460 28960 3466
rect 28908 3402 28960 3408
rect 29644 3460 29696 3466
rect 29644 3402 29696 3408
rect 28920 480 28948 3402
rect 30116 480 30144 6886
rect 31312 480 31340 6886
rect 33060 3466 33088 47602
rect 34440 3466 34468 77930
rect 35806 73808 35862 73817
rect 35806 73743 35862 73752
rect 35820 3466 35848 73743
rect 36556 3534 36584 79319
rect 37186 42120 37242 42129
rect 37186 42055 37242 42064
rect 36544 3528 36596 3534
rect 36544 3470 36596 3476
rect 32404 3460 32456 3466
rect 32404 3402 32456 3408
rect 33048 3460 33100 3466
rect 33048 3402 33100 3408
rect 33600 3460 33652 3466
rect 33600 3402 33652 3408
rect 34428 3460 34480 3466
rect 34428 3402 34480 3408
rect 34796 3460 34848 3466
rect 34796 3402 34848 3408
rect 35808 3460 35860 3466
rect 35808 3402 35860 3408
rect 37096 3460 37148 3466
rect 37096 3402 37148 3408
rect 32416 480 32444 3402
rect 33612 480 33640 3402
rect 34808 480 34836 3402
rect 35992 3324 36044 3330
rect 35992 3266 36044 3272
rect 36004 480 36032 3266
rect 37108 1714 37136 3402
rect 37200 3330 37228 42055
rect 38568 40724 38620 40730
rect 38568 40666 38620 40672
rect 38580 6914 38608 40666
rect 40696 33114 40724 203487
rect 50816 193934 50844 271866
rect 50908 235890 50936 378082
rect 51000 336054 51028 462334
rect 52288 457502 52316 587862
rect 55128 586560 55180 586566
rect 55128 586502 55180 586508
rect 53656 567248 53708 567254
rect 53656 567190 53708 567196
rect 52368 563100 52420 563106
rect 52368 563042 52420 563048
rect 52276 457496 52328 457502
rect 52276 457438 52328 457444
rect 52274 444680 52330 444689
rect 52274 444615 52330 444624
rect 52182 415440 52238 415449
rect 52182 415375 52238 415384
rect 50988 336048 51040 336054
rect 50988 335990 51040 335996
rect 50988 331356 51040 331362
rect 50988 331298 51040 331304
rect 50896 235884 50948 235890
rect 50896 235826 50948 235832
rect 50804 193928 50856 193934
rect 50804 193870 50856 193876
rect 47584 175976 47636 175982
rect 47584 175918 47636 175924
rect 42706 64152 42762 64161
rect 42706 64087 42762 64096
rect 41328 44872 41380 44878
rect 41328 44814 41380 44820
rect 40684 33108 40736 33114
rect 40684 33050 40736 33056
rect 39580 15972 39632 15978
rect 39580 15914 39632 15920
rect 38396 6886 38608 6914
rect 37188 3324 37240 3330
rect 37188 3266 37240 3272
rect 37108 1686 37228 1714
rect 37200 480 37228 1686
rect 38396 480 38424 6886
rect 39592 480 39620 15914
rect 41340 3534 41368 44814
rect 42720 3534 42748 64087
rect 44088 44940 44140 44946
rect 44088 44882 44140 44888
rect 44100 3534 44128 44882
rect 47596 44305 47624 175918
rect 51000 72457 51028 331298
rect 52196 291174 52224 415375
rect 52184 291168 52236 291174
rect 52184 291110 52236 291116
rect 52184 276072 52236 276078
rect 52184 276014 52236 276020
rect 52196 223553 52224 276014
rect 52288 253230 52316 444615
rect 52380 431254 52408 563042
rect 53668 438190 53696 567190
rect 54484 564460 54536 564466
rect 54484 564402 54536 564408
rect 53746 533352 53802 533361
rect 53746 533287 53802 533296
rect 53656 438184 53708 438190
rect 53656 438126 53708 438132
rect 52368 431248 52420 431254
rect 52368 431190 52420 431196
rect 52460 427100 52512 427106
rect 52460 427042 52512 427048
rect 52472 425746 52500 427042
rect 52460 425740 52512 425746
rect 52460 425682 52512 425688
rect 53656 425740 53708 425746
rect 53656 425682 53708 425688
rect 53668 378729 53696 425682
rect 53654 378720 53710 378729
rect 53654 378655 53710 378664
rect 53472 370524 53524 370530
rect 53472 370466 53524 370472
rect 52368 320204 52420 320210
rect 52368 320146 52420 320152
rect 52276 253224 52328 253230
rect 52276 253166 52328 253172
rect 52182 223544 52238 223553
rect 52182 223479 52238 223488
rect 51080 204944 51132 204950
rect 51080 204886 51132 204892
rect 51092 202842 51120 204886
rect 51080 202836 51132 202842
rect 51080 202778 51132 202784
rect 50986 72448 51042 72457
rect 50986 72383 51042 72392
rect 50986 71088 51042 71097
rect 50986 71023 51042 71032
rect 48226 65512 48282 65521
rect 48226 65447 48282 65456
rect 47582 44296 47638 44305
rect 47582 44231 47638 44240
rect 46846 35184 46902 35193
rect 46846 35119 46902 35128
rect 45468 22772 45520 22778
rect 45468 22714 45520 22720
rect 45376 18624 45428 18630
rect 45376 18566 45428 18572
rect 45388 16574 45416 18566
rect 45296 16546 45416 16574
rect 44272 3596 44324 3602
rect 44272 3538 44324 3544
rect 40684 3528 40736 3534
rect 40684 3470 40736 3476
rect 41328 3528 41380 3534
rect 41328 3470 41380 3476
rect 41880 3528 41932 3534
rect 41880 3470 41932 3476
rect 42708 3528 42760 3534
rect 42708 3470 42760 3476
rect 43076 3528 43128 3534
rect 43076 3470 43128 3476
rect 44088 3528 44140 3534
rect 44088 3470 44140 3476
rect 40696 480 40724 3470
rect 41892 480 41920 3470
rect 43088 480 43116 3470
rect 44284 480 44312 3538
rect 45296 3482 45324 16546
rect 45480 6914 45508 22714
rect 46860 6914 46888 35119
rect 48240 6914 48268 65447
rect 49608 28280 49660 28286
rect 49608 28222 49660 28228
rect 45388 6886 45508 6914
rect 46676 6886 46888 6914
rect 47872 6886 48268 6914
rect 45388 3602 45416 6886
rect 45376 3596 45428 3602
rect 45376 3538 45428 3544
rect 45296 3454 45508 3482
rect 45480 480 45508 3454
rect 46676 480 46704 6886
rect 47872 480 47900 6886
rect 49620 3534 49648 28222
rect 51000 3534 51028 71023
rect 52380 27606 52408 320146
rect 53484 302190 53512 370466
rect 53656 319456 53708 319462
rect 53656 319398 53708 319404
rect 53564 305040 53616 305046
rect 53564 304982 53616 304988
rect 53472 302184 53524 302190
rect 53472 302126 53524 302132
rect 53472 264988 53524 264994
rect 53472 264930 53524 264936
rect 53484 198694 53512 264930
rect 53576 216481 53604 304982
rect 53562 216472 53618 216481
rect 53562 216407 53618 216416
rect 53472 198688 53524 198694
rect 53472 198630 53524 198636
rect 53668 46209 53696 319398
rect 53760 258058 53788 533287
rect 54496 433362 54524 564402
rect 55140 519586 55168 586502
rect 57796 585200 57848 585206
rect 57796 585142 57848 585148
rect 56508 554804 56560 554810
rect 56508 554746 56560 554752
rect 55128 519580 55180 519586
rect 55128 519522 55180 519528
rect 54484 433356 54536 433362
rect 54484 433298 54536 433304
rect 56520 416673 56548 554746
rect 57704 547936 57756 547942
rect 57704 547878 57756 547884
rect 57612 453348 57664 453354
rect 57612 453290 57664 453296
rect 56506 416664 56562 416673
rect 56506 416599 56562 416608
rect 56520 415449 56548 416599
rect 56506 415440 56562 415449
rect 56506 415375 56562 415384
rect 56416 411324 56468 411330
rect 56416 411266 56468 411272
rect 55036 400240 55088 400246
rect 55036 400182 55088 400188
rect 54944 343664 54996 343670
rect 54944 343606 54996 343612
rect 54956 313274 54984 343606
rect 54944 313268 54996 313274
rect 54944 313210 54996 313216
rect 53748 258052 53800 258058
rect 53748 257994 53800 258000
rect 54944 253972 54996 253978
rect 54944 253914 54996 253920
rect 54956 227050 54984 253914
rect 55048 238678 55076 400182
rect 56324 358080 56376 358086
rect 56324 358022 56376 358028
rect 55128 325712 55180 325718
rect 55128 325654 55180 325660
rect 55036 238672 55088 238678
rect 55036 238614 55088 238620
rect 54944 227044 54996 227050
rect 54944 226986 54996 226992
rect 53746 51776 53802 51785
rect 53746 51711 53802 51720
rect 53654 46200 53710 46209
rect 53654 46135 53710 46144
rect 52368 27600 52420 27606
rect 52368 27542 52420 27548
rect 53656 17264 53708 17270
rect 53656 17206 53708 17212
rect 53668 3534 53696 17206
rect 48964 3528 49016 3534
rect 48964 3470 49016 3476
rect 49608 3528 49660 3534
rect 49608 3470 49660 3476
rect 50160 3528 50212 3534
rect 50160 3470 50212 3476
rect 50988 3528 51040 3534
rect 50988 3470 51040 3476
rect 52552 3528 52604 3534
rect 52552 3470 52604 3476
rect 53656 3528 53708 3534
rect 53656 3470 53708 3476
rect 48976 480 49004 3470
rect 50172 480 50200 3470
rect 51356 2168 51408 2174
rect 51356 2110 51408 2116
rect 51368 480 51396 2110
rect 52564 480 52592 3470
rect 53760 480 53788 51711
rect 54482 36544 54538 36553
rect 54482 36479 54538 36488
rect 54496 2106 54524 36479
rect 55140 24818 55168 325654
rect 56336 289814 56364 358022
rect 56428 340105 56456 411266
rect 57624 389026 57652 453290
rect 57716 405822 57744 547878
rect 57808 456074 57836 585142
rect 59268 581052 59320 581058
rect 59268 580994 59320 581000
rect 59084 565888 59136 565894
rect 59084 565830 59136 565836
rect 57888 460216 57940 460222
rect 57888 460158 57940 460164
rect 57796 456068 57848 456074
rect 57796 456010 57848 456016
rect 57796 414724 57848 414730
rect 57796 414666 57848 414672
rect 57704 405816 57756 405822
rect 57704 405758 57756 405764
rect 57612 389020 57664 389026
rect 57612 388962 57664 388968
rect 57702 382936 57758 382945
rect 57702 382871 57758 382880
rect 56506 366344 56562 366353
rect 56506 366279 56562 366288
rect 56414 340096 56470 340105
rect 56414 340031 56470 340040
rect 56416 291168 56468 291174
rect 56416 291110 56468 291116
rect 56428 289882 56456 291110
rect 56416 289876 56468 289882
rect 56416 289818 56468 289824
rect 56324 289808 56376 289814
rect 56324 289750 56376 289756
rect 56428 213897 56456 289818
rect 56520 271862 56548 366279
rect 56508 271856 56560 271862
rect 56508 271798 56560 271804
rect 57612 267028 57664 267034
rect 57612 266970 57664 266976
rect 56508 260908 56560 260914
rect 56508 260850 56560 260856
rect 56414 213888 56470 213897
rect 56414 213823 56470 213832
rect 56520 186998 56548 260850
rect 57244 258052 57296 258058
rect 57244 257994 57296 258000
rect 56508 186992 56560 186998
rect 56508 186934 56560 186940
rect 57256 31754 57284 257994
rect 57624 234598 57652 266970
rect 57716 262682 57744 382871
rect 57704 262676 57756 262682
rect 57704 262618 57756 262624
rect 57808 248414 57836 414666
rect 57716 248386 57836 248414
rect 57716 241398 57744 248386
rect 57796 241460 57848 241466
rect 57796 241402 57848 241408
rect 57704 241392 57756 241398
rect 57704 241334 57756 241340
rect 57808 240786 57836 241402
rect 57796 240780 57848 240786
rect 57796 240722 57848 240728
rect 57612 234592 57664 234598
rect 57612 234534 57664 234540
rect 57808 227633 57836 240722
rect 57794 227624 57850 227633
rect 57794 227559 57850 227568
rect 57900 83502 57928 460158
rect 59096 435402 59124 565830
rect 59280 529242 59308 580994
rect 61936 574116 61988 574122
rect 61936 574058 61988 574064
rect 60648 568608 60700 568614
rect 60648 568550 60700 568556
rect 60556 549296 60608 549302
rect 60556 549238 60608 549244
rect 59268 529236 59320 529242
rect 59268 529178 59320 529184
rect 59176 523728 59228 523734
rect 59176 523670 59228 523676
rect 59084 435396 59136 435402
rect 59084 435338 59136 435344
rect 59084 423700 59136 423706
rect 59084 423642 59136 423648
rect 59096 363662 59124 423642
rect 59188 389298 59216 523670
rect 60568 514758 60596 549238
rect 60556 514752 60608 514758
rect 60556 514694 60608 514700
rect 59268 444508 59320 444514
rect 59268 444450 59320 444456
rect 59176 389292 59228 389298
rect 59176 389234 59228 389240
rect 59084 363656 59136 363662
rect 59084 363598 59136 363604
rect 59174 355328 59230 355337
rect 59174 355263 59230 355272
rect 59084 345092 59136 345098
rect 59084 345034 59136 345040
rect 58624 337408 58676 337414
rect 58624 337350 58676 337356
rect 58636 241466 58664 337350
rect 59096 295322 59124 345034
rect 59084 295316 59136 295322
rect 59084 295258 59136 295264
rect 59084 263628 59136 263634
rect 59084 263570 59136 263576
rect 58624 241460 58676 241466
rect 58624 241402 58676 241408
rect 59096 230217 59124 263570
rect 59188 244254 59216 355263
rect 59280 263634 59308 444450
rect 60568 407153 60596 514694
rect 60660 456754 60688 568550
rect 60740 558680 60792 558686
rect 60740 558622 60792 558628
rect 60752 558210 60780 558622
rect 60740 558204 60792 558210
rect 60740 558146 60792 558152
rect 60648 456748 60700 456754
rect 60648 456690 60700 456696
rect 61842 453248 61898 453257
rect 61842 453183 61898 453192
rect 60646 445768 60702 445777
rect 60646 445703 60702 445712
rect 60554 407144 60610 407153
rect 60554 407079 60610 407088
rect 60660 383654 60688 445703
rect 60740 438184 60792 438190
rect 60740 438126 60792 438132
rect 60752 437510 60780 438126
rect 60740 437504 60792 437510
rect 60740 437446 60792 437452
rect 61856 388793 61884 453183
rect 61948 447846 61976 574058
rect 62040 558686 62068 702918
rect 67640 702704 67692 702710
rect 67640 702646 67692 702652
rect 66168 699712 66220 699718
rect 66168 699654 66220 699660
rect 63316 590776 63368 590782
rect 63316 590718 63368 590724
rect 62028 558680 62080 558686
rect 62028 558622 62080 558628
rect 62028 546508 62080 546514
rect 62028 546450 62080 546456
rect 62040 517478 62068 546450
rect 62028 517472 62080 517478
rect 62028 517414 62080 517420
rect 61936 447840 61988 447846
rect 61936 447782 61988 447788
rect 61936 437504 61988 437510
rect 61936 437446 61988 437452
rect 61842 388784 61898 388793
rect 61842 388719 61898 388728
rect 61842 388376 61898 388385
rect 61842 388311 61898 388320
rect 60568 383626 60688 383654
rect 60568 382401 60596 383626
rect 60554 382392 60610 382401
rect 60554 382327 60610 382336
rect 60462 346624 60518 346633
rect 60462 346559 60518 346568
rect 60476 314634 60504 346559
rect 60464 314628 60516 314634
rect 60464 314570 60516 314576
rect 60464 300892 60516 300898
rect 60464 300834 60516 300840
rect 59268 263628 59320 263634
rect 59268 263570 59320 263576
rect 59268 262676 59320 262682
rect 59268 262618 59320 262624
rect 59280 262274 59308 262618
rect 59268 262268 59320 262274
rect 59268 262210 59320 262216
rect 59176 244248 59228 244254
rect 59176 244190 59228 244196
rect 59082 230208 59138 230217
rect 59082 230143 59138 230152
rect 59280 202842 59308 262210
rect 60188 253224 60240 253230
rect 60188 253166 60240 253172
rect 60200 252618 60228 253166
rect 60188 252612 60240 252618
rect 60188 252554 60240 252560
rect 60476 233209 60504 300834
rect 60568 292534 60596 382327
rect 61752 342304 61804 342310
rect 61752 342246 61804 342252
rect 60646 331800 60702 331809
rect 60646 331735 60702 331744
rect 60556 292528 60608 292534
rect 60556 292470 60608 292476
rect 60556 252612 60608 252618
rect 60556 252554 60608 252560
rect 60462 233200 60518 233209
rect 60462 233135 60518 233144
rect 60568 222193 60596 252554
rect 60554 222184 60610 222193
rect 60554 222119 60610 222128
rect 59268 202836 59320 202842
rect 59268 202778 59320 202784
rect 57888 83496 57940 83502
rect 57888 83438 57940 83444
rect 57886 57216 57942 57225
rect 57886 57151 57942 57160
rect 57244 31748 57296 31754
rect 57244 31690 57296 31696
rect 56508 29640 56560 29646
rect 56508 29582 56560 29588
rect 55128 24812 55180 24818
rect 55128 24754 55180 24760
rect 54944 13116 54996 13122
rect 54944 13058 54996 13064
rect 54484 2100 54536 2106
rect 54484 2042 54536 2048
rect 54956 480 54984 13058
rect 56520 3534 56548 29582
rect 57242 17232 57298 17241
rect 57242 17167 57298 17176
rect 57256 6914 57284 17167
rect 57164 6886 57284 6914
rect 56048 3528 56100 3534
rect 56048 3470 56100 3476
rect 56508 3528 56560 3534
rect 56508 3470 56560 3476
rect 56060 480 56088 3470
rect 57164 3369 57192 6886
rect 57900 3534 57928 57151
rect 58622 53136 58678 53145
rect 58622 53071 58678 53080
rect 58440 6180 58492 6186
rect 58440 6122 58492 6128
rect 57244 3528 57296 3534
rect 57244 3470 57296 3476
rect 57888 3528 57940 3534
rect 57888 3470 57940 3476
rect 57150 3360 57206 3369
rect 57150 3295 57206 3304
rect 57256 480 57284 3470
rect 58452 480 58480 6122
rect 58636 2174 58664 53071
rect 60660 32434 60688 331735
rect 61764 309806 61792 342246
rect 61752 309800 61804 309806
rect 61752 309742 61804 309748
rect 61856 284306 61884 388311
rect 61948 384305 61976 437446
rect 62040 403646 62068 517414
rect 63328 454714 63356 590718
rect 64788 579692 64840 579698
rect 64788 579634 64840 579640
rect 64696 553444 64748 553450
rect 64696 553386 64748 553392
rect 63408 539640 63460 539646
rect 63408 539582 63460 539588
rect 63316 454708 63368 454714
rect 63316 454650 63368 454656
rect 63224 450560 63276 450566
rect 63224 450502 63276 450508
rect 62028 403640 62080 403646
rect 62028 403582 62080 403588
rect 63236 386374 63264 450502
rect 63420 393314 63448 539582
rect 64708 529854 64736 553386
rect 64800 530602 64828 579634
rect 65982 573472 66038 573481
rect 65982 573407 66038 573416
rect 65996 542337 66024 573407
rect 66074 559600 66130 559609
rect 66074 559535 66130 559544
rect 65982 542328 66038 542337
rect 65982 542263 66038 542272
rect 64788 530596 64840 530602
rect 64788 530538 64840 530544
rect 64696 529848 64748 529854
rect 64696 529790 64748 529796
rect 64708 528554 64736 529790
rect 64708 528526 64828 528554
rect 64696 449268 64748 449274
rect 64696 449210 64748 449216
rect 64602 416664 64658 416673
rect 64602 416599 64658 416608
rect 63328 393286 63448 393314
rect 63328 392018 63356 393286
rect 63316 392012 63368 392018
rect 63316 391954 63368 391960
rect 63224 386368 63276 386374
rect 63224 386310 63276 386316
rect 61934 384296 61990 384305
rect 61934 384231 61990 384240
rect 62026 374096 62082 374105
rect 62026 374031 62082 374040
rect 61936 335368 61988 335374
rect 61936 335310 61988 335316
rect 61948 317490 61976 335310
rect 61936 317484 61988 317490
rect 61936 317426 61988 317432
rect 61936 316056 61988 316062
rect 61936 315998 61988 316004
rect 61844 284300 61896 284306
rect 61844 284242 61896 284248
rect 61844 256760 61896 256766
rect 61844 256702 61896 256708
rect 61750 249928 61806 249937
rect 61750 249863 61806 249872
rect 61764 235958 61792 249863
rect 61752 235952 61804 235958
rect 61752 235894 61804 235900
rect 61856 228313 61884 256702
rect 61842 228304 61898 228313
rect 61842 228239 61898 228248
rect 61948 190369 61976 315998
rect 62040 247042 62068 374031
rect 63224 349172 63276 349178
rect 63224 349114 63276 349120
rect 63130 334656 63186 334665
rect 63130 334591 63186 334600
rect 63144 304978 63172 334591
rect 63236 318578 63264 349114
rect 63224 318572 63276 318578
rect 63224 318514 63276 318520
rect 63328 314974 63356 391954
rect 64616 389201 64644 416599
rect 64708 391377 64736 449210
rect 64800 414730 64828 528526
rect 65616 456748 65668 456754
rect 65616 456690 65668 456696
rect 65628 455462 65656 456690
rect 65616 455456 65668 455462
rect 65616 455398 65668 455404
rect 65892 455456 65944 455462
rect 65892 455398 65944 455404
rect 65904 439686 65932 455398
rect 65984 454028 66036 454034
rect 65984 453970 66036 453976
rect 65892 439680 65944 439686
rect 65892 439622 65944 439628
rect 65892 431248 65944 431254
rect 65892 431190 65944 431196
rect 64788 414724 64840 414730
rect 64788 414666 64840 414672
rect 64788 405816 64840 405822
rect 64788 405758 64840 405764
rect 64694 391368 64750 391377
rect 64694 391303 64750 391312
rect 64602 389192 64658 389201
rect 64602 389127 64658 389136
rect 63406 369064 63462 369073
rect 63406 368999 63462 369008
rect 63316 314968 63368 314974
rect 63316 314910 63368 314916
rect 63316 307828 63368 307834
rect 63316 307770 63368 307776
rect 63132 304972 63184 304978
rect 63132 304914 63184 304920
rect 62764 285728 62816 285734
rect 62764 285670 62816 285676
rect 62028 247036 62080 247042
rect 62028 246978 62080 246984
rect 62776 197985 62804 285670
rect 63224 273284 63276 273290
rect 63224 273226 63276 273232
rect 63236 240825 63264 273226
rect 63222 240816 63278 240825
rect 63222 240751 63278 240760
rect 63328 231849 63356 307770
rect 63420 284374 63448 368999
rect 64800 366382 64828 405758
rect 65522 381032 65578 381041
rect 65522 380967 65578 380976
rect 64788 366376 64840 366382
rect 64788 366318 64840 366324
rect 64694 362264 64750 362273
rect 64694 362199 64750 362208
rect 64602 336832 64658 336841
rect 64602 336767 64658 336776
rect 64512 334620 64564 334626
rect 64512 334562 64564 334568
rect 64524 316742 64552 334562
rect 64512 316736 64564 316742
rect 64512 316678 64564 316684
rect 64616 307766 64644 336767
rect 64604 307760 64656 307766
rect 64604 307702 64656 307708
rect 64708 298858 64736 362199
rect 64786 342952 64842 342961
rect 64786 342887 64842 342896
rect 64696 298852 64748 298858
rect 64696 298794 64748 298800
rect 63408 284368 63460 284374
rect 63406 284336 63408 284345
rect 63460 284336 63462 284345
rect 63406 284271 63462 284280
rect 64604 281580 64656 281586
rect 64604 281522 64656 281528
rect 63408 250504 63460 250510
rect 63408 250446 63460 250452
rect 63314 231840 63370 231849
rect 63314 231775 63370 231784
rect 63420 199442 63448 250446
rect 64512 249824 64564 249830
rect 64512 249766 64564 249772
rect 64524 212537 64552 249766
rect 64616 236609 64644 281522
rect 64696 278792 64748 278798
rect 64696 278734 64748 278740
rect 64602 236600 64658 236609
rect 64602 236535 64658 236544
rect 64708 229770 64736 278734
rect 64800 267850 64828 342887
rect 65536 316062 65564 380967
rect 65904 376689 65932 431190
rect 65996 389094 66024 453970
rect 66088 424289 66116 559535
rect 66180 536761 66208 699654
rect 67364 592748 67416 592754
rect 67364 592690 67416 592696
rect 66810 588432 66866 588441
rect 66810 588367 66866 588376
rect 66824 587926 66852 588367
rect 66812 587920 66864 587926
rect 66812 587862 66864 587868
rect 66260 586560 66312 586566
rect 66258 586528 66260 586537
rect 66312 586528 66314 586537
rect 66258 586463 66314 586472
rect 66810 585712 66866 585721
rect 66810 585647 66866 585656
rect 66824 585206 66852 585647
rect 66812 585200 66864 585206
rect 66812 585142 66864 585148
rect 66810 582992 66866 583001
rect 66810 582927 66866 582936
rect 66824 582418 66852 582927
rect 66812 582412 66864 582418
rect 66812 582354 66864 582360
rect 66718 581768 66774 581777
rect 66718 581703 66774 581712
rect 66732 581058 66760 581703
rect 66720 581052 66772 581058
rect 66720 580994 66772 581000
rect 66810 580272 66866 580281
rect 66810 580207 66866 580216
rect 66824 579698 66852 580207
rect 66812 579692 66864 579698
rect 66812 579634 66864 579640
rect 67376 574977 67404 592690
rect 67546 577552 67602 577561
rect 67546 577487 67602 577496
rect 67454 576192 67510 576201
rect 67454 576127 67456 576136
rect 67508 576127 67510 576136
rect 67456 576098 67508 576104
rect 67362 574968 67418 574977
rect 67362 574903 67418 574912
rect 67376 574122 67404 574903
rect 67364 574116 67416 574122
rect 67364 574058 67416 574064
rect 66810 572112 66866 572121
rect 66810 572047 66866 572056
rect 66824 571402 66852 572047
rect 66812 571396 66864 571402
rect 66812 571338 66864 571344
rect 67362 570752 67418 570761
rect 67362 570687 67418 570696
rect 66810 569392 66866 569401
rect 66810 569327 66866 569336
rect 66824 568614 66852 569327
rect 66812 568608 66864 568614
rect 66812 568550 66864 568556
rect 66810 568032 66866 568041
rect 66810 567967 66866 567976
rect 66824 567254 66852 567967
rect 66812 567248 66864 567254
rect 66812 567190 66864 567196
rect 66810 565040 66866 565049
rect 66810 564975 66866 564984
rect 66824 564466 66852 564975
rect 66812 564460 66864 564466
rect 66812 564402 66864 564408
rect 66810 563680 66866 563689
rect 66810 563615 66866 563624
rect 66824 563106 66852 563615
rect 66812 563100 66864 563106
rect 66812 563042 66864 563048
rect 66810 562320 66866 562329
rect 66810 562255 66866 562264
rect 66824 561746 66852 562255
rect 66812 561740 66864 561746
rect 66812 561682 66864 561688
rect 66810 560960 66866 560969
rect 66810 560895 66866 560904
rect 66824 560318 66852 560895
rect 66812 560312 66864 560318
rect 66812 560254 66864 560260
rect 66260 558680 66312 558686
rect 66260 558622 66312 558628
rect 66272 558385 66300 558622
rect 66258 558376 66314 558385
rect 66258 558311 66314 558320
rect 66810 555520 66866 555529
rect 66810 555455 66866 555464
rect 66824 554810 66852 555455
rect 66812 554804 66864 554810
rect 66812 554746 66864 554752
rect 66442 554160 66498 554169
rect 66442 554095 66498 554104
rect 66456 553450 66484 554095
rect 66444 553444 66496 553450
rect 66444 553386 66496 553392
rect 66810 550080 66866 550089
rect 66810 550015 66866 550024
rect 66824 549302 66852 550015
rect 66812 549296 66864 549302
rect 66812 549238 66864 549244
rect 66810 548720 66866 548729
rect 66810 548655 66866 548664
rect 66824 547942 66852 548655
rect 66812 547936 66864 547942
rect 66812 547878 66864 547884
rect 66902 547360 66958 547369
rect 66902 547295 66958 547304
rect 66916 546514 66944 547295
rect 66904 546508 66956 546514
rect 66904 546450 66956 546456
rect 66902 546000 66958 546009
rect 66902 545935 66958 545944
rect 66916 545154 66944 545935
rect 66904 545148 66956 545154
rect 66904 545090 66956 545096
rect 66902 544640 66958 544649
rect 66902 544575 66958 544584
rect 66916 543794 66944 544575
rect 66904 543788 66956 543794
rect 66904 543730 66956 543736
rect 66902 543280 66958 543289
rect 66902 543215 66958 543224
rect 66916 542434 66944 543215
rect 66904 542428 66956 542434
rect 66904 542370 66956 542376
rect 66994 541920 67050 541929
rect 66994 541855 67050 541864
rect 67008 541686 67036 541855
rect 66996 541680 67048 541686
rect 66996 541622 67048 541628
rect 67272 541680 67324 541686
rect 67272 541622 67324 541628
rect 67086 537432 67142 537441
rect 67086 537367 67142 537376
rect 66166 536752 66222 536761
rect 66166 536687 66222 536696
rect 66074 424280 66130 424289
rect 66074 424215 66130 424224
rect 66088 423706 66116 424215
rect 66076 423700 66128 423706
rect 66076 423642 66128 423648
rect 66076 421592 66128 421598
rect 66076 421534 66128 421540
rect 65984 389088 66036 389094
rect 65984 389030 66036 389036
rect 66088 381041 66116 421534
rect 66180 387802 66208 536687
rect 67100 523025 67128 537367
rect 67086 523016 67142 523025
rect 67086 522951 67142 522960
rect 66902 522880 66958 522889
rect 66902 522815 66958 522824
rect 66916 522306 66944 522815
rect 66904 522300 66956 522306
rect 66904 522242 66956 522248
rect 66350 439920 66406 439929
rect 66350 439855 66406 439864
rect 66364 439686 66392 439855
rect 66352 439680 66404 439686
rect 66352 439622 66404 439628
rect 66258 435432 66314 435441
rect 66258 435367 66260 435376
rect 66312 435367 66314 435376
rect 66260 435338 66312 435344
rect 66260 433288 66312 433294
rect 66258 433256 66260 433265
rect 66312 433256 66314 433265
rect 66258 433191 66314 433200
rect 66364 431954 66392 439622
rect 66810 437744 66866 437753
rect 66810 437679 66866 437688
rect 66824 437510 66852 437679
rect 66812 437504 66864 437510
rect 66812 437446 66864 437452
rect 66272 431926 66392 431954
rect 66168 387796 66220 387802
rect 66168 387738 66220 387744
rect 66074 381032 66130 381041
rect 66074 380967 66130 380976
rect 65890 376680 65946 376689
rect 65890 376615 65946 376624
rect 66168 369028 66220 369034
rect 66168 368970 66220 368976
rect 65982 357504 66038 357513
rect 65982 357439 66038 357448
rect 65890 332752 65946 332761
rect 65890 332687 65946 332696
rect 65524 316056 65576 316062
rect 65524 315998 65576 316004
rect 65904 303113 65932 332687
rect 65996 305289 66024 357439
rect 66180 322402 66208 368970
rect 66272 342310 66300 431926
rect 66536 431248 66588 431254
rect 66536 431190 66588 431196
rect 66548 431089 66576 431190
rect 66534 431080 66590 431089
rect 66534 431015 66590 431024
rect 66812 429140 66864 429146
rect 66812 429082 66864 429088
rect 66824 428641 66852 429082
rect 66810 428632 66866 428641
rect 66810 428567 66866 428576
rect 66810 426320 66866 426329
rect 66810 426255 66866 426264
rect 66824 425746 66852 426255
rect 66812 425740 66864 425746
rect 66812 425682 66864 425688
rect 66626 421968 66682 421977
rect 66626 421903 66682 421912
rect 66640 421598 66668 421903
rect 66628 421592 66680 421598
rect 66628 421534 66680 421540
rect 66810 415168 66866 415177
rect 66810 415103 66866 415112
rect 66824 414730 66852 415103
rect 66812 414724 66864 414730
rect 66812 414666 66864 414672
rect 66916 412634 66944 522242
rect 66732 412606 66944 412634
rect 66732 411330 66760 412606
rect 66720 411324 66772 411330
rect 66720 411266 66772 411272
rect 66732 410689 66760 411266
rect 66718 410680 66774 410689
rect 66718 410615 66774 410624
rect 66350 406192 66406 406201
rect 66350 406127 66406 406136
rect 66364 405822 66392 406127
rect 66352 405816 66404 405822
rect 66352 405758 66404 405764
rect 66350 403744 66406 403753
rect 66350 403679 66406 403688
rect 66364 403646 66392 403679
rect 66352 403640 66404 403646
rect 66352 403582 66404 403588
rect 66350 401568 66406 401577
rect 66350 401503 66406 401512
rect 66364 400246 66392 401503
rect 66352 400240 66404 400246
rect 66352 400182 66404 400188
rect 66350 399392 66406 399401
rect 66350 399327 66406 399336
rect 66364 398886 66392 399327
rect 66352 398880 66404 398886
rect 66352 398822 66404 398828
rect 66994 396944 67050 396953
rect 66994 396879 67050 396888
rect 67008 396778 67036 396879
rect 66996 396772 67048 396778
rect 66996 396714 67048 396720
rect 67284 396001 67312 541622
rect 67376 534070 67404 570687
rect 67468 562358 67496 576098
rect 67456 562352 67508 562358
rect 67456 562294 67508 562300
rect 67454 552800 67510 552809
rect 67454 552735 67510 552744
rect 67364 534064 67416 534070
rect 67364 534006 67416 534012
rect 67376 442241 67404 534006
rect 67362 442232 67418 442241
rect 67362 442167 67418 442176
rect 67468 412865 67496 552735
rect 67560 539782 67588 577487
rect 67652 566681 67680 702646
rect 72988 699718 73016 703520
rect 79324 702636 79376 702642
rect 79324 702578 79376 702584
rect 75184 700324 75236 700330
rect 75184 700266 75236 700272
rect 72976 699712 73028 699718
rect 72976 699654 73028 699660
rect 71780 605124 71832 605130
rect 71780 605066 71832 605072
rect 70308 596216 70360 596222
rect 70308 596158 70360 596164
rect 69112 592680 69164 592686
rect 69112 592622 69164 592628
rect 69124 589422 69152 592622
rect 70320 590753 70348 596158
rect 70306 590744 70362 590753
rect 70306 590679 70362 590688
rect 71134 590744 71190 590753
rect 71134 590679 71190 590688
rect 70306 589928 70362 589937
rect 70306 589863 70362 589872
rect 69112 589416 69164 589422
rect 69112 589358 69164 589364
rect 69124 589084 69152 589358
rect 70320 589098 70348 589863
rect 70150 589070 70348 589098
rect 71148 589084 71176 590679
rect 71792 589098 71820 605066
rect 75196 592754 75224 700266
rect 79336 595678 79364 702578
rect 88248 702568 88300 702574
rect 88248 702510 88300 702516
rect 86224 699712 86276 699718
rect 86224 699654 86276 699660
rect 86236 605130 86264 699654
rect 86224 605124 86276 605130
rect 86224 605066 86276 605072
rect 79324 595672 79376 595678
rect 79324 595614 79376 595620
rect 80336 595672 80388 595678
rect 80336 595614 80388 595620
rect 80348 594930 80376 595614
rect 80336 594924 80388 594930
rect 80336 594866 80388 594872
rect 75184 592748 75236 592754
rect 75184 592690 75236 592696
rect 78588 592136 78640 592142
rect 74906 592104 74962 592113
rect 78588 592078 78640 592084
rect 74906 592039 74962 592048
rect 73068 590844 73120 590850
rect 73068 590786 73120 590792
rect 71792 589084 72082 589098
rect 73080 589084 73108 590786
rect 73896 590776 73948 590782
rect 73896 590718 73948 590724
rect 73908 589084 73936 590718
rect 74920 589354 74948 592039
rect 77666 591016 77722 591025
rect 77666 590951 77722 590960
rect 74908 589348 74960 589354
rect 74908 589290 74960 589296
rect 76748 589348 76800 589354
rect 76748 589290 76800 589296
rect 74920 589084 74948 589290
rect 76760 589084 76788 589290
rect 77680 589084 77708 590951
rect 78600 589084 78628 592078
rect 79324 590844 79376 590850
rect 79324 590786 79376 590792
rect 71792 589070 72096 589084
rect 72068 588690 72096 589070
rect 72422 588704 72478 588713
rect 72068 588676 72422 588690
rect 72082 588662 72422 588676
rect 79336 588674 79364 590786
rect 80348 589084 80376 594866
rect 85948 594856 86000 594862
rect 85948 594798 86000 594804
rect 84108 592068 84160 592074
rect 84108 592010 84160 592016
rect 82266 590880 82322 590889
rect 82266 590815 82322 590824
rect 81346 589384 81402 589393
rect 81346 589319 81402 589328
rect 81360 589084 81388 589319
rect 82280 589084 82308 590815
rect 83186 589520 83242 589529
rect 83186 589455 83242 589464
rect 83200 589084 83228 589455
rect 84120 589084 84148 592010
rect 85028 592000 85080 592006
rect 85028 591942 85080 591948
rect 85040 589084 85068 591942
rect 85960 589084 85988 594798
rect 88260 593434 88288 702510
rect 88800 702500 88852 702506
rect 88800 702442 88852 702448
rect 88812 596174 88840 702442
rect 89180 699718 89208 703520
rect 95148 702636 95200 702642
rect 95148 702578 95200 702584
rect 89168 699712 89220 699718
rect 89168 699654 89220 699660
rect 90364 605872 90416 605878
rect 90364 605814 90416 605820
rect 88812 596146 89024 596174
rect 88248 593428 88300 593434
rect 88248 593370 88300 593376
rect 88260 592006 88288 593370
rect 88248 592000 88300 592006
rect 88248 591942 88300 591948
rect 86868 590708 86920 590714
rect 86868 590650 86920 590656
rect 86880 589084 86908 590650
rect 72422 588639 72478 588648
rect 79324 588668 79376 588674
rect 88734 588662 88932 588690
rect 79324 588610 79376 588616
rect 79784 588600 79836 588606
rect 75854 588526 75960 588554
rect 79534 588548 79784 588554
rect 88062 588568 88118 588577
rect 79534 588542 79836 588548
rect 79534 588526 79824 588542
rect 87814 588526 88062 588554
rect 75932 588470 75960 588526
rect 88062 588503 88118 588512
rect 75920 588464 75972 588470
rect 75920 588406 75972 588412
rect 88904 588402 88932 588662
rect 88892 588396 88944 588402
rect 88892 588338 88944 588344
rect 88996 588282 89024 596146
rect 90376 594318 90404 605814
rect 90364 594312 90416 594318
rect 90364 594254 90416 594260
rect 91100 594312 91152 594318
rect 91100 594254 91152 594260
rect 89812 594108 89864 594114
rect 89812 594050 89864 594056
rect 89076 589416 89128 589422
rect 89076 589358 89128 589364
rect 88812 588254 89024 588282
rect 67730 584352 67786 584361
rect 67730 584287 67786 584296
rect 67638 566672 67694 566681
rect 67638 566607 67694 566616
rect 67652 565894 67680 566607
rect 67640 565888 67692 565894
rect 67640 565830 67692 565836
rect 67548 539776 67600 539782
rect 67548 539718 67600 539724
rect 67548 539640 67600 539646
rect 67546 539608 67548 539617
rect 67600 539608 67602 539617
rect 67546 539543 67602 539552
rect 67744 462398 67772 584287
rect 67822 578912 67878 578921
rect 67822 578847 67878 578856
rect 67836 538286 67864 578847
rect 88812 576854 88840 588254
rect 88892 588192 88944 588198
rect 88892 588134 88944 588140
rect 88904 584526 88932 588134
rect 88984 587852 89036 587858
rect 88984 587794 89036 587800
rect 88996 586634 89024 587794
rect 88984 586628 89036 586634
rect 88984 586570 89036 586576
rect 89088 586514 89116 589358
rect 88996 586486 89116 586514
rect 88892 584520 88944 584526
rect 88892 584462 88944 584468
rect 88812 576826 88932 576854
rect 68284 562352 68336 562358
rect 68284 562294 68336 562300
rect 67824 538280 67876 538286
rect 67824 538222 67876 538228
rect 68296 476134 68324 562294
rect 88904 560153 88932 576826
rect 88890 560144 88946 560153
rect 88890 560079 88946 560088
rect 88892 541000 88944 541006
rect 88892 540942 88944 540948
rect 88798 540152 88854 540161
rect 88798 540087 88854 540096
rect 88812 539646 88840 540087
rect 69388 539640 69440 539646
rect 71872 539640 71924 539646
rect 69440 539588 69690 539594
rect 69388 539582 69690 539588
rect 71872 539582 71924 539588
rect 81164 539640 81216 539646
rect 81164 539582 81216 539588
rect 88800 539640 88852 539646
rect 88800 539582 88852 539588
rect 69400 539566 69690 539582
rect 68664 539294 68770 539322
rect 68664 536722 68692 539294
rect 68652 536716 68704 536722
rect 68652 536658 68704 536664
rect 68284 476128 68336 476134
rect 68284 476070 68336 476076
rect 67732 462392 67784 462398
rect 67732 462334 67784 462340
rect 68284 447228 68336 447234
rect 68284 447170 68336 447176
rect 67824 446412 67876 446418
rect 67824 446354 67876 446360
rect 67730 419656 67786 419665
rect 67730 419591 67786 419600
rect 67454 412856 67510 412865
rect 67454 412791 67510 412800
rect 67362 396944 67418 396953
rect 67362 396879 67418 396888
rect 67270 395992 67326 396001
rect 67270 395927 67326 395936
rect 66810 392592 66866 392601
rect 66810 392527 66866 392536
rect 66824 392018 66852 392527
rect 66812 392012 66864 392018
rect 66812 391954 66864 391960
rect 67376 365702 67404 396879
rect 66904 365696 66956 365702
rect 66904 365638 66956 365644
rect 67364 365696 67416 365702
rect 67364 365638 67416 365644
rect 66916 349178 66944 365638
rect 66904 349172 66956 349178
rect 66904 349114 66956 349120
rect 67364 349172 67416 349178
rect 67364 349114 67416 349120
rect 67376 348401 67404 349114
rect 67362 348392 67418 348401
rect 67362 348327 67418 348336
rect 67272 343732 67324 343738
rect 67272 343674 67324 343680
rect 66260 342304 66312 342310
rect 66260 342246 66312 342252
rect 66902 326768 66958 326777
rect 66902 326703 66958 326712
rect 66916 325718 66944 326703
rect 66904 325712 66956 325718
rect 66904 325654 66956 325660
rect 66258 322416 66314 322425
rect 66180 322374 66258 322402
rect 66180 316034 66208 322374
rect 66258 322351 66314 322360
rect 66904 321564 66956 321570
rect 66904 321506 66956 321512
rect 66810 321328 66866 321337
rect 66810 321263 66866 321272
rect 66824 320210 66852 321263
rect 66916 320249 66944 321506
rect 66902 320240 66958 320249
rect 66812 320204 66864 320210
rect 66902 320175 66958 320184
rect 66812 320146 66864 320152
rect 67284 319462 67312 343674
rect 67364 342304 67416 342310
rect 67364 342246 67416 342252
rect 67376 341465 67404 342246
rect 67362 341456 67418 341465
rect 67362 341391 67418 341400
rect 67364 331288 67416 331294
rect 67364 331230 67416 331236
rect 66996 319456 67048 319462
rect 66996 319398 67048 319404
rect 67272 319456 67324 319462
rect 67272 319398 67324 319404
rect 67008 319161 67036 319398
rect 66994 319152 67050 319161
rect 66994 319087 67050 319096
rect 66812 318572 66864 318578
rect 66812 318514 66864 318520
rect 66824 318073 66852 318514
rect 66810 318064 66866 318073
rect 66810 317999 66866 318008
rect 66720 317484 66772 317490
rect 66720 317426 66772 317432
rect 66088 316006 66208 316034
rect 66732 316034 66760 317426
rect 66810 316976 66866 316985
rect 66810 316911 66866 316920
rect 66824 316742 66852 316911
rect 66812 316736 66864 316742
rect 66812 316678 66864 316684
rect 66732 316006 66852 316034
rect 65982 305280 66038 305289
rect 65982 305215 66038 305224
rect 65890 303104 65946 303113
rect 65890 303039 65946 303048
rect 65984 274644 66036 274650
rect 65984 274586 66036 274592
rect 65996 274553 66024 274586
rect 65982 274544 66038 274553
rect 65982 274479 66038 274488
rect 65996 273737 66024 274479
rect 65982 273728 66038 273737
rect 65982 273663 66038 273672
rect 64788 267844 64840 267850
rect 64788 267786 64840 267792
rect 64696 229764 64748 229770
rect 64696 229706 64748 229712
rect 64800 219337 64828 267786
rect 65892 261520 65944 261526
rect 65892 261462 65944 261468
rect 65904 228993 65932 261462
rect 65982 255504 66038 255513
rect 65982 255439 66038 255448
rect 65890 228984 65946 228993
rect 65890 228919 65946 228928
rect 65996 222154 66024 255439
rect 66088 240786 66116 316006
rect 66628 315988 66680 315994
rect 66628 315930 66680 315936
rect 66534 315888 66590 315897
rect 66534 315823 66590 315832
rect 66548 314974 66576 315823
rect 66168 314968 66220 314974
rect 66168 314910 66220 314916
rect 66536 314968 66588 314974
rect 66536 314910 66588 314916
rect 66076 240780 66128 240786
rect 66076 240722 66128 240728
rect 65984 222148 66036 222154
rect 65984 222090 66036 222096
rect 64786 219328 64842 219337
rect 64786 219263 64842 219272
rect 66180 216617 66208 314910
rect 66640 314809 66668 315930
rect 66626 314800 66682 314809
rect 66626 314735 66682 314744
rect 66628 304972 66680 304978
rect 66628 304914 66680 304920
rect 66640 304201 66668 304914
rect 66626 304192 66682 304201
rect 66626 304127 66682 304136
rect 66720 302184 66772 302190
rect 66720 302126 66772 302132
rect 66732 300937 66760 302126
rect 66718 300928 66774 300937
rect 66718 300863 66774 300872
rect 66260 295316 66312 295322
rect 66260 295258 66312 295264
rect 66272 294409 66300 295258
rect 66258 294400 66314 294409
rect 66258 294335 66314 294344
rect 66628 289808 66680 289814
rect 66628 289750 66680 289756
rect 66640 288969 66668 289750
rect 66626 288960 66682 288969
rect 66626 288895 66682 288904
rect 66824 287054 66852 316006
rect 66904 314628 66956 314634
rect 66904 314570 66956 314576
rect 66916 313993 66944 314570
rect 66902 313984 66958 313993
rect 66902 313919 66958 313928
rect 66904 313268 66956 313274
rect 66904 313210 66956 313216
rect 66916 312905 66944 313210
rect 66902 312896 66958 312905
rect 66902 312831 66958 312840
rect 66994 311808 67050 311817
rect 66994 311743 67050 311752
rect 66904 309800 66956 309806
rect 66904 309742 66956 309748
rect 66916 309641 66944 309742
rect 66902 309632 66958 309641
rect 66902 309567 66958 309576
rect 66904 307760 66956 307766
rect 66904 307702 66956 307708
rect 66916 307465 66944 307702
rect 66902 307456 66958 307465
rect 66902 307391 66958 307400
rect 66902 306368 66958 306377
rect 66902 306303 66958 306312
rect 66916 305046 66944 306303
rect 66904 305040 66956 305046
rect 66904 304982 66956 304988
rect 66902 302016 66958 302025
rect 66902 301951 66958 301960
rect 66916 300898 66944 301951
rect 66904 300892 66956 300898
rect 66904 300834 66956 300840
rect 67008 300150 67036 311743
rect 67088 311160 67140 311166
rect 67088 311102 67140 311108
rect 67100 310729 67128 311102
rect 67086 310720 67142 310729
rect 67086 310655 67142 310664
rect 66996 300144 67048 300150
rect 66996 300086 67048 300092
rect 66904 298852 66956 298858
rect 66904 298794 66956 298800
rect 66916 298761 66944 298794
rect 66902 298752 66958 298761
rect 66902 298687 66958 298696
rect 66904 298104 66956 298110
rect 66904 298046 66956 298052
rect 66916 297673 66944 298046
rect 66902 297664 66958 297673
rect 66902 297599 66958 297608
rect 67178 296304 67234 296313
rect 67178 296239 67234 296248
rect 66902 295488 66958 295497
rect 66902 295423 66904 295432
rect 66956 295423 66958 295432
rect 66904 295394 66956 295400
rect 67192 295390 67220 296239
rect 67180 295384 67232 295390
rect 67180 295326 67232 295332
rect 66904 293956 66956 293962
rect 66904 293898 66956 293904
rect 66916 293321 66944 293898
rect 66902 293312 66958 293321
rect 66902 293247 66958 293256
rect 66904 292528 66956 292534
rect 66904 292470 66956 292476
rect 66916 292233 66944 292470
rect 66902 292224 66958 292233
rect 66902 292159 66958 292168
rect 66902 291136 66958 291145
rect 66902 291071 66958 291080
rect 66916 289882 66944 291071
rect 67376 290057 67404 331230
rect 67468 311166 67496 412791
rect 67546 395992 67602 396001
rect 67546 395927 67602 395936
rect 67560 394913 67588 395927
rect 67546 394904 67602 394913
rect 67546 394839 67602 394848
rect 67560 375426 67588 394839
rect 67640 389156 67692 389162
rect 67640 389098 67692 389104
rect 67548 375420 67600 375426
rect 67548 375362 67600 375368
rect 67456 311160 67508 311166
rect 67456 311102 67508 311108
rect 67560 299849 67588 375362
rect 67652 369034 67680 389098
rect 67744 378865 67772 419591
rect 67836 387122 67864 446354
rect 68296 440910 68324 447170
rect 68284 440904 68336 440910
rect 68284 440846 68336 440852
rect 68664 390402 68692 536658
rect 69584 535537 69612 539566
rect 70504 539294 70610 539322
rect 70780 539294 71530 539322
rect 70504 536790 70532 539294
rect 70492 536784 70544 536790
rect 70492 536726 70544 536732
rect 70504 535537 70532 536726
rect 69570 535528 69626 535537
rect 69570 535463 69626 535472
rect 70490 535528 70546 535537
rect 70490 535463 70546 535472
rect 70780 528554 70808 539294
rect 70412 528526 70808 528554
rect 70412 527542 70440 528526
rect 70400 527536 70452 527542
rect 70400 527478 70452 527484
rect 71044 527536 71096 527542
rect 71044 527478 71096 527484
rect 71056 527202 71084 527478
rect 71044 527196 71096 527202
rect 71044 527138 71096 527144
rect 68928 476128 68980 476134
rect 68928 476070 68980 476076
rect 68836 462392 68888 462398
rect 68836 462334 68888 462340
rect 68848 461650 68876 462334
rect 68836 461644 68888 461650
rect 68836 461586 68888 461592
rect 68940 447098 68968 476070
rect 69018 456920 69074 456929
rect 69018 456855 69074 456864
rect 68928 447092 68980 447098
rect 68928 447034 68980 447040
rect 68744 446412 68796 446418
rect 68744 446354 68796 446360
rect 68756 444380 68784 446354
rect 69032 444394 69060 456855
rect 71056 454034 71084 527138
rect 71044 454028 71096 454034
rect 71044 453970 71096 453976
rect 71780 449880 71832 449886
rect 71780 449822 71832 449828
rect 71792 449206 71820 449822
rect 71780 449200 71832 449206
rect 71780 449142 71832 449148
rect 71780 447840 71832 447846
rect 71780 447782 71832 447788
rect 71792 447166 71820 447782
rect 71884 447234 71912 539582
rect 72344 539294 72450 539322
rect 73172 539294 73370 539322
rect 73540 539294 74290 539322
rect 75104 539294 75210 539322
rect 75932 539294 76130 539322
rect 76760 539294 77050 539322
rect 78062 539294 78352 539322
rect 72344 536790 72372 539294
rect 72332 536784 72384 536790
rect 72332 536726 72384 536732
rect 72344 535537 72372 536726
rect 73172 536081 73200 539294
rect 73158 536072 73214 536081
rect 73158 536007 73214 536016
rect 72330 535528 72386 535537
rect 72330 535463 72386 535472
rect 73540 528554 73568 539294
rect 75104 538214 75132 539294
rect 75104 538186 75224 538214
rect 75196 536625 75224 538186
rect 75182 536616 75238 536625
rect 75182 536551 75238 536560
rect 73172 528526 73568 528554
rect 73172 453354 73200 528526
rect 73160 453348 73212 453354
rect 73160 453290 73212 453296
rect 75196 453257 75224 536551
rect 75182 453248 75238 453257
rect 75182 453183 75238 453192
rect 75932 450566 75960 539294
rect 76564 538280 76616 538286
rect 76564 538222 76616 538228
rect 76576 461514 76604 538222
rect 76760 536761 76788 539294
rect 76746 536752 76802 536761
rect 76746 536687 76802 536696
rect 78324 534818 78352 539294
rect 78692 539294 78890 539322
rect 79060 539294 79810 539322
rect 80822 539294 81112 539322
rect 78312 534812 78364 534818
rect 78312 534754 78364 534760
rect 77944 530596 77996 530602
rect 77944 530538 77996 530544
rect 76012 461508 76064 461514
rect 76012 461450 76064 461456
rect 76564 461508 76616 461514
rect 76564 461450 76616 461456
rect 75920 450560 75972 450566
rect 75920 450502 75972 450508
rect 72700 449200 72752 449206
rect 72700 449142 72752 449148
rect 72712 448633 72740 449142
rect 72698 448624 72754 448633
rect 72698 448559 72754 448568
rect 71872 447228 71924 447234
rect 71872 447170 71924 447176
rect 71780 447160 71832 447166
rect 71780 447102 71832 447108
rect 69032 444366 70242 444394
rect 71792 444380 71820 447102
rect 71884 446758 71912 447170
rect 73160 447092 73212 447098
rect 73160 447034 73212 447040
rect 71872 446752 71924 446758
rect 71872 446694 71924 446700
rect 73172 444380 73200 447034
rect 74816 446752 74868 446758
rect 74816 446694 74868 446700
rect 74828 444380 74856 446694
rect 76024 444394 76052 461450
rect 76576 460970 76604 461450
rect 76564 460964 76616 460970
rect 76564 460906 76616 460912
rect 77956 452674 77984 530538
rect 77944 452668 77996 452674
rect 77944 452610 77996 452616
rect 77956 444394 77984 452610
rect 78692 449274 78720 539294
rect 79060 528554 79088 539294
rect 80058 535664 80114 535673
rect 80058 535599 80114 535608
rect 80072 529802 80100 535599
rect 81084 532710 81112 539294
rect 81176 536790 81204 539582
rect 88156 539572 88208 539578
rect 88156 539514 88208 539520
rect 81452 539294 81650 539322
rect 82662 539294 82768 539322
rect 81164 536784 81216 536790
rect 81164 536726 81216 536732
rect 81072 532704 81124 532710
rect 81072 532646 81124 532652
rect 79980 529786 80100 529802
rect 79324 529780 79376 529786
rect 79324 529722 79376 529728
rect 79968 529780 80100 529786
rect 80020 529774 80100 529780
rect 79968 529722 80020 529728
rect 79336 529242 79364 529722
rect 79324 529236 79376 529242
rect 79324 529178 79376 529184
rect 78784 528526 79088 528554
rect 78784 523734 78812 528526
rect 78772 523728 78824 523734
rect 78772 523670 78824 523676
rect 79336 460934 79364 529178
rect 81452 464409 81480 539294
rect 82740 535498 82768 539294
rect 82832 539294 83490 539322
rect 84304 539294 84410 539322
rect 84580 539294 85330 539322
rect 86342 539294 86632 539322
rect 82728 535492 82780 535498
rect 82728 535434 82780 535440
rect 81438 464400 81494 464409
rect 81438 464335 81494 464344
rect 82832 462913 82860 539294
rect 84304 535537 84332 539294
rect 84290 535528 84346 535537
rect 84290 535463 84346 535472
rect 84580 528554 84608 539294
rect 86604 538214 86632 539294
rect 87064 539294 87354 539322
rect 86868 538214 86920 538218
rect 86604 538212 86920 538214
rect 86604 538186 86868 538212
rect 86868 538154 86920 538160
rect 86224 535492 86276 535498
rect 86224 535434 86276 535440
rect 84212 528526 84608 528554
rect 82818 462904 82874 462913
rect 82818 462839 82874 462848
rect 81440 461644 81492 461650
rect 81440 461586 81492 461592
rect 79336 460906 79456 460934
rect 78680 449268 78732 449274
rect 78680 449210 78732 449216
rect 79428 444514 79456 460906
rect 80886 447808 80942 447817
rect 80886 447743 80942 447752
rect 79416 444508 79468 444514
rect 79416 444450 79468 444456
rect 76024 444366 76314 444394
rect 77878 444366 77984 444394
rect 79428 444380 79456 444450
rect 80900 444380 80928 447743
rect 81452 444394 81480 461586
rect 82820 456068 82872 456074
rect 82820 456010 82872 456016
rect 82832 455433 82860 456010
rect 82818 455424 82874 455433
rect 82818 455359 82874 455368
rect 82832 444394 82860 455359
rect 84212 447817 84240 528526
rect 85580 519580 85632 519586
rect 85580 519522 85632 519528
rect 84198 447808 84254 447817
rect 84198 447743 84254 447752
rect 85592 445777 85620 519522
rect 86236 465769 86264 535434
rect 86222 465760 86278 465769
rect 86222 465695 86278 465704
rect 86880 453257 86908 538154
rect 87064 460934 87092 539294
rect 88168 536722 88196 539514
rect 88904 539458 88932 540942
rect 88366 539430 88932 539458
rect 88156 536716 88208 536722
rect 88156 536658 88208 536664
rect 88444 528554 88472 539430
rect 88352 528526 88472 528554
rect 87064 460906 87184 460934
rect 87052 457496 87104 457502
rect 87052 457438 87104 457444
rect 86866 453248 86922 453257
rect 86866 453183 86922 453192
rect 85578 445768 85634 445777
rect 85578 445703 85634 445712
rect 81452 444366 82386 444394
rect 82832 444366 83858 444394
rect 85592 444380 85620 445703
rect 87064 444553 87092 457438
rect 87156 456113 87184 460906
rect 88352 457473 88380 528526
rect 88338 457464 88394 457473
rect 88338 457399 88394 457408
rect 87142 456104 87198 456113
rect 87142 456039 87198 456048
rect 88996 454850 89024 586486
rect 89718 586256 89774 586265
rect 89718 586191 89774 586200
rect 89626 560144 89682 560153
rect 89626 560079 89682 560088
rect 89640 558958 89668 560079
rect 89628 558952 89680 558958
rect 89628 558894 89680 558900
rect 89732 532030 89760 586191
rect 89824 567361 89852 594050
rect 90362 589928 90418 589937
rect 90362 589863 90418 589872
rect 89810 567352 89866 567361
rect 89810 567287 89866 567296
rect 89720 532024 89772 532030
rect 89720 531966 89772 531972
rect 88340 454844 88392 454850
rect 88340 454786 88392 454792
rect 88984 454844 89036 454850
rect 88984 454786 89036 454792
rect 88352 454102 88380 454786
rect 88340 454096 88392 454102
rect 88340 454038 88392 454044
rect 87050 444544 87106 444553
rect 87050 444479 87106 444488
rect 87064 444380 87092 444479
rect 88352 444394 88380 454038
rect 90376 444961 90404 589863
rect 91112 576745 91140 594254
rect 93766 589384 93822 589393
rect 93766 589319 93822 589328
rect 93122 588704 93178 588713
rect 93122 588639 93178 588648
rect 91742 587616 91798 587625
rect 91742 587551 91798 587560
rect 91756 586566 91784 587551
rect 91744 586560 91796 586566
rect 91744 586502 91796 586508
rect 91374 584896 91430 584905
rect 91374 584831 91430 584840
rect 91388 584458 91416 584831
rect 91376 584452 91428 584458
rect 91376 584394 91428 584400
rect 91192 583704 91244 583710
rect 91190 583672 91192 583681
rect 91244 583672 91246 583681
rect 91190 583607 91246 583616
rect 91742 582176 91798 582185
rect 91742 582111 91798 582120
rect 91756 581058 91784 582111
rect 91744 581052 91796 581058
rect 91744 580994 91796 581000
rect 91742 580816 91798 580825
rect 91742 580751 91798 580760
rect 91756 579698 91784 580751
rect 91744 579692 91796 579698
rect 91744 579634 91796 579640
rect 91742 579456 91798 579465
rect 91742 579391 91798 579400
rect 91756 578270 91784 579391
rect 91744 578264 91796 578270
rect 91744 578206 91796 578212
rect 91098 576736 91154 576745
rect 91098 576671 91154 576680
rect 91112 576162 91140 576671
rect 91100 576156 91152 576162
rect 91100 576098 91152 576104
rect 91098 575376 91154 575385
rect 91098 575311 91154 575320
rect 91112 574122 91140 575311
rect 91100 574116 91152 574122
rect 91100 574058 91152 574064
rect 91098 574016 91154 574025
rect 91098 573951 91154 573960
rect 91112 572762 91140 573951
rect 91100 572756 91152 572762
rect 91100 572698 91152 572704
rect 91190 572656 91246 572665
rect 91190 572591 91246 572600
rect 91098 571432 91154 571441
rect 91098 571367 91100 571376
rect 91152 571367 91154 571376
rect 91100 571338 91152 571344
rect 91204 570654 91232 572591
rect 91192 570648 91244 570654
rect 91192 570590 91244 570596
rect 91098 570072 91154 570081
rect 91098 570007 91154 570016
rect 91112 569974 91140 570007
rect 91100 569968 91152 569974
rect 91100 569910 91152 569916
rect 91098 568712 91154 568721
rect 91098 568647 91154 568656
rect 91112 568614 91140 568647
rect 91100 568608 91152 568614
rect 91100 568550 91152 568556
rect 91466 567352 91522 567361
rect 91466 567287 91522 567296
rect 91376 565888 91428 565894
rect 91374 565856 91376 565865
rect 91428 565856 91430 565865
rect 91374 565791 91430 565800
rect 91480 565146 91508 567287
rect 91468 565140 91520 565146
rect 91468 565082 91520 565088
rect 91374 564496 91430 564505
rect 91374 564431 91376 564440
rect 91428 564431 91430 564440
rect 91376 564402 91428 564408
rect 91374 563136 91430 563145
rect 91374 563071 91376 563080
rect 91428 563071 91430 563080
rect 91376 563042 91428 563048
rect 91098 561504 91154 561513
rect 91098 561439 91154 561448
rect 91112 557410 91140 561439
rect 91190 558784 91246 558793
rect 91190 558719 91246 558728
rect 91204 557598 91232 558719
rect 91192 557592 91244 557598
rect 91192 557534 91244 557540
rect 91282 557424 91338 557433
rect 91112 557382 91232 557410
rect 91098 556064 91154 556073
rect 91098 555999 91154 556008
rect 91112 554849 91140 555999
rect 91098 554840 91154 554849
rect 91098 554775 91154 554784
rect 91098 554704 91154 554713
rect 91098 554639 91154 554648
rect 91112 553450 91140 554639
rect 91100 553444 91152 553450
rect 91100 553386 91152 553392
rect 91100 552152 91152 552158
rect 91098 552120 91100 552129
rect 91152 552120 91154 552129
rect 91098 552055 91154 552064
rect 91098 550760 91154 550769
rect 91098 550695 91100 550704
rect 91152 550695 91154 550704
rect 91100 550666 91152 550672
rect 91098 549400 91154 549409
rect 91098 549335 91154 549344
rect 91112 547913 91140 549335
rect 91098 547904 91154 547913
rect 91098 547839 91154 547848
rect 91098 545184 91154 545193
rect 91098 545119 91100 545128
rect 91152 545119 91154 545128
rect 91100 545090 91152 545096
rect 91098 542464 91154 542473
rect 91098 542399 91100 542408
rect 91152 542399 91154 542408
rect 91100 542370 91152 542376
rect 91100 541680 91152 541686
rect 91100 541622 91152 541628
rect 91112 541249 91140 541622
rect 91098 541240 91154 541249
rect 91098 541175 91154 541184
rect 91098 539744 91154 539753
rect 91098 539679 91100 539688
rect 91152 539679 91154 539688
rect 91100 539650 91152 539656
rect 91204 538898 91232 557382
rect 91282 557359 91338 557368
rect 91296 556306 91324 557359
rect 91284 556300 91336 556306
rect 91284 556242 91336 556248
rect 92110 553344 92166 553353
rect 92110 553279 92166 553288
rect 92124 552090 92152 553279
rect 92112 552084 92164 552090
rect 92112 552026 92164 552032
rect 91374 548040 91430 548049
rect 91374 547975 91430 547984
rect 91388 547942 91416 547975
rect 91376 547936 91428 547942
rect 91376 547878 91428 547884
rect 91282 546544 91338 546553
rect 91282 546479 91338 546488
rect 91192 538892 91244 538898
rect 91192 538834 91244 538840
rect 91296 538778 91324 546479
rect 91204 538750 91324 538778
rect 90454 535528 90510 535537
rect 90454 535463 90510 535472
rect 90468 459649 90496 535463
rect 91204 534750 91232 538750
rect 91388 538642 91416 547878
rect 91558 546544 91614 546553
rect 91558 546479 91560 546488
rect 91612 546479 91614 546488
rect 91560 546450 91612 546456
rect 92386 542328 92442 542337
rect 92386 542263 92442 542272
rect 91296 538614 91416 538642
rect 91296 537538 91324 538614
rect 91284 537532 91336 537538
rect 91284 537474 91336 537480
rect 91192 534744 91244 534750
rect 91192 534686 91244 534692
rect 90454 459640 90510 459649
rect 90454 459575 90510 459584
rect 91558 450528 91614 450537
rect 91558 450463 91614 450472
rect 90362 444952 90418 444961
rect 90362 444887 90418 444896
rect 90376 444394 90404 444887
rect 88352 444366 88458 444394
rect 90206 444366 90404 444394
rect 91572 444380 91600 450463
rect 92400 449177 92428 542263
rect 93136 451274 93164 588639
rect 93780 465730 93808 589319
rect 94504 588668 94556 588674
rect 94504 588610 94556 588616
rect 93768 465724 93820 465730
rect 93768 465666 93820 465672
rect 93044 451246 93164 451274
rect 92386 449168 92442 449177
rect 92386 449103 92442 449112
rect 93044 447137 93072 451246
rect 94516 448526 94544 588610
rect 95160 584458 95188 702578
rect 99288 702500 99340 702506
rect 99288 702442 99340 702448
rect 96618 592104 96674 592113
rect 96618 592039 96674 592048
rect 95882 590880 95938 590889
rect 95882 590815 95938 590824
rect 95240 586560 95292 586566
rect 95240 586502 95292 586508
rect 95148 584452 95200 584458
rect 95148 584394 95200 584400
rect 95148 571396 95200 571402
rect 95148 571338 95200 571344
rect 95160 569226 95188 571338
rect 95148 569220 95200 569226
rect 95148 569162 95200 569168
rect 95146 547904 95202 547913
rect 95146 547839 95202 547848
rect 94596 545148 94648 545154
rect 94596 545090 94648 545096
rect 94608 464409 94636 545090
rect 94594 464400 94650 464409
rect 94594 464335 94650 464344
rect 95160 460193 95188 547839
rect 95252 460222 95280 586502
rect 95896 577522 95924 590815
rect 95884 577516 95936 577522
rect 95884 577458 95936 577464
rect 95884 542428 95936 542434
rect 95884 542370 95936 542376
rect 95896 469849 95924 542370
rect 95882 469840 95938 469849
rect 95882 469775 95938 469784
rect 95240 460216 95292 460222
rect 95146 460184 95202 460193
rect 95240 460158 95292 460164
rect 95146 460119 95202 460128
rect 95884 454708 95936 454714
rect 95884 454650 95936 454656
rect 95896 451246 95924 454650
rect 95884 451240 95936 451246
rect 95884 451182 95936 451188
rect 94504 448520 94556 448526
rect 94504 448462 94556 448468
rect 93030 447128 93086 447137
rect 93030 447063 93086 447072
rect 93044 444689 93072 447063
rect 94516 444689 94544 448462
rect 93030 444680 93086 444689
rect 93030 444615 93086 444624
rect 94502 444680 94558 444689
rect 94502 444615 94558 444624
rect 93044 444380 93072 444615
rect 94516 444394 94544 444615
rect 95896 444394 95924 451182
rect 96632 445777 96660 592039
rect 97262 591016 97318 591025
rect 97262 590951 97318 590960
rect 97276 454034 97304 590951
rect 98644 586628 98696 586634
rect 98644 586570 98696 586576
rect 97906 543824 97962 543833
rect 97906 543759 97962 543768
rect 97920 471209 97948 543759
rect 98000 532704 98052 532710
rect 98000 532646 98052 532652
rect 98012 531457 98040 532646
rect 97998 531448 98054 531457
rect 97998 531383 98054 531392
rect 98012 531350 98040 531383
rect 98000 531344 98052 531350
rect 98000 531286 98052 531292
rect 97906 471200 97962 471209
rect 97906 471135 97962 471144
rect 97264 454028 97316 454034
rect 97264 453970 97316 453976
rect 98656 451353 98684 586570
rect 99300 583710 99328 702442
rect 105464 700330 105492 703520
rect 137848 700398 137876 703520
rect 154132 702545 154160 703520
rect 170324 702710 170352 703520
rect 202800 702914 202828 703520
rect 202788 702908 202840 702914
rect 202788 702850 202840 702856
rect 170312 702704 170364 702710
rect 170312 702646 170364 702652
rect 191748 702704 191800 702710
rect 191748 702646 191800 702652
rect 154118 702536 154174 702545
rect 154118 702471 154174 702480
rect 124864 700392 124916 700398
rect 124864 700334 124916 700340
rect 137836 700392 137888 700398
rect 137836 700334 137888 700340
rect 105452 700324 105504 700330
rect 105452 700266 105504 700272
rect 106924 594924 106976 594930
rect 106924 594866 106976 594872
rect 103520 592136 103572 592142
rect 103520 592078 103572 592084
rect 101404 589348 101456 589354
rect 101404 589290 101456 589296
rect 99288 583704 99340 583710
rect 99288 583646 99340 583652
rect 99300 583030 99328 583646
rect 99288 583024 99340 583030
rect 99288 582966 99340 582972
rect 100024 568608 100076 568614
rect 100024 568550 100076 568556
rect 98642 451344 98698 451353
rect 98642 451279 98698 451288
rect 96618 445768 96674 445777
rect 96618 445703 96674 445712
rect 97630 445768 97686 445777
rect 97630 445703 97686 445712
rect 94516 444366 94714 444394
rect 95896 444366 96186 444394
rect 97644 444380 97672 445703
rect 98656 444394 98684 451279
rect 100036 449274 100064 568550
rect 100024 449268 100076 449274
rect 100024 449210 100076 449216
rect 101416 444514 101444 589290
rect 101496 569968 101548 569974
rect 101496 569910 101548 569916
rect 101508 566506 101536 569910
rect 101496 566500 101548 566506
rect 101496 566442 101548 566448
rect 102784 565888 102836 565894
rect 102784 565830 102836 565836
rect 101496 564460 101548 564466
rect 101496 564402 101548 564408
rect 101508 479505 101536 564402
rect 101588 539708 101640 539714
rect 101588 539650 101640 539656
rect 101494 479496 101550 479505
rect 101494 479431 101550 479440
rect 101600 456113 101628 539650
rect 101586 456104 101642 456113
rect 101586 456039 101642 456048
rect 102140 454028 102192 454034
rect 102140 453970 102192 453976
rect 102152 445777 102180 453970
rect 102796 453354 102824 565830
rect 102784 453348 102836 453354
rect 102784 453290 102836 453296
rect 103532 449206 103560 592078
rect 105544 588600 105596 588606
rect 105544 588542 105596 588548
rect 104256 552152 104308 552158
rect 104256 552094 104308 552100
rect 104164 546508 104216 546514
rect 104164 546450 104216 546456
rect 104176 457065 104204 546450
rect 104268 468489 104296 552094
rect 104254 468480 104310 468489
rect 104254 468415 104310 468424
rect 105556 467838 105584 588542
rect 106186 554840 106242 554849
rect 106186 554775 106242 554784
rect 105544 467832 105596 467838
rect 105544 467774 105596 467780
rect 105556 466478 105584 467774
rect 104900 466472 104952 466478
rect 104900 466414 104952 466420
rect 105544 466472 105596 466478
rect 105544 466414 105596 466420
rect 104162 457056 104218 457065
rect 104162 456991 104218 457000
rect 103520 449200 103572 449206
rect 103520 449142 103572 449148
rect 103704 449200 103756 449206
rect 103704 449142 103756 449148
rect 102138 445768 102194 445777
rect 102138 445703 102194 445712
rect 101404 444508 101456 444514
rect 101404 444450 101456 444456
rect 101416 444394 101444 444450
rect 98656 444366 99130 444394
rect 100878 444366 101444 444394
rect 102152 444394 102180 445703
rect 102152 444366 102258 444394
rect 103716 444380 103744 449142
rect 104912 444394 104940 466414
rect 106200 463010 106228 554775
rect 106188 463004 106240 463010
rect 106188 462946 106240 462952
rect 106936 451178 106964 594866
rect 113180 593428 113232 593434
rect 113180 593370 113232 593376
rect 112444 592068 112496 592074
rect 112444 592010 112496 592016
rect 111062 589520 111118 589529
rect 111062 589455 111118 589464
rect 108304 583024 108356 583030
rect 108304 582966 108356 582972
rect 107660 465724 107712 465730
rect 107660 465666 107712 465672
rect 106924 451172 106976 451178
rect 106924 451114 106976 451120
rect 104912 444366 105386 444394
rect 106936 444380 106964 451114
rect 107672 444394 107700 465666
rect 108316 447817 108344 582966
rect 109040 577516 109092 577522
rect 109040 577458 109092 577464
rect 108396 552084 108448 552090
rect 108396 552026 108448 552032
rect 108408 464409 108436 552026
rect 108394 464400 108450 464409
rect 108394 464335 108450 464344
rect 108302 447808 108358 447817
rect 108302 447743 108358 447752
rect 109052 447098 109080 577458
rect 111076 561746 111104 589455
rect 111064 561740 111116 561746
rect 111064 561682 111116 561688
rect 111708 561740 111760 561746
rect 111708 561682 111760 561688
rect 109040 447092 109092 447098
rect 109040 447034 109092 447040
rect 109776 447092 109828 447098
rect 109776 447034 109828 447040
rect 109498 444544 109554 444553
rect 109498 444479 109554 444488
rect 109512 444394 109540 444479
rect 109788 444394 109816 447034
rect 111522 444544 111578 444553
rect 111522 444479 111578 444488
rect 107672 444366 108330 444394
rect 109512 444380 109816 444394
rect 111536 444394 111564 444479
rect 111720 444394 111748 561682
rect 112456 556238 112484 592010
rect 112444 556232 112496 556238
rect 112444 556174 112496 556180
rect 112456 459542 112484 556174
rect 112536 553444 112588 553450
rect 112536 553386 112588 553392
rect 112444 459536 112496 459542
rect 112444 459478 112496 459484
rect 112456 445806 112484 459478
rect 112548 458833 112576 553386
rect 112534 458824 112590 458833
rect 112534 458759 112590 458768
rect 112444 445800 112496 445806
rect 112444 445742 112496 445748
rect 112904 445800 112956 445806
rect 113192 445777 113220 593370
rect 115296 590708 115348 590714
rect 115296 590650 115348 590656
rect 115204 572756 115256 572762
rect 115204 572698 115256 572704
rect 115216 445777 115244 572698
rect 115308 562562 115336 590650
rect 119342 585712 119398 585721
rect 119342 585647 119398 585656
rect 116584 584520 116636 584526
rect 116584 584462 116636 584468
rect 115296 562556 115348 562562
rect 115296 562498 115348 562504
rect 116596 451994 116624 584462
rect 117964 562556 118016 562562
rect 117964 562498 118016 562504
rect 117976 552022 118004 562498
rect 117964 552016 118016 552022
rect 117964 551958 118016 551964
rect 118608 552016 118660 552022
rect 118608 551958 118660 551964
rect 118620 550662 118648 551958
rect 118608 550656 118660 550662
rect 118608 550598 118660 550604
rect 116584 451988 116636 451994
rect 116584 451930 116636 451936
rect 116122 446448 116178 446457
rect 116122 446383 116178 446392
rect 112904 445742 112956 445748
rect 113178 445768 113234 445777
rect 111536 444380 111748 444394
rect 112916 444380 112944 445742
rect 113178 445703 113234 445712
rect 114374 445768 114430 445777
rect 114374 445703 114430 445712
rect 115202 445768 115258 445777
rect 115202 445703 115258 445712
rect 114388 444553 114416 445703
rect 114374 444544 114430 444553
rect 114374 444479 114430 444488
rect 114388 444380 114416 444479
rect 116136 444380 116164 446383
rect 118620 445777 118648 550598
rect 119356 448594 119384 585647
rect 120724 578264 120776 578270
rect 120724 578206 120776 578212
rect 120736 568546 120764 578206
rect 123116 576156 123168 576162
rect 123116 576098 123168 576104
rect 122196 574116 122248 574122
rect 122196 574058 122248 574064
rect 121552 570648 121604 570654
rect 121552 570590 121604 570596
rect 120724 568540 120776 568546
rect 120724 568482 120776 568488
rect 121368 568540 121420 568546
rect 121368 568482 121420 568488
rect 121380 567254 121408 568482
rect 121368 567248 121420 567254
rect 121368 567190 121420 567196
rect 120816 463004 120868 463010
rect 120816 462946 120868 462952
rect 119344 448588 119396 448594
rect 119344 448530 119396 448536
rect 117594 445768 117650 445777
rect 117594 445703 117650 445712
rect 118606 445768 118662 445777
rect 118606 445703 118662 445712
rect 117608 444380 117636 445703
rect 118700 444440 118752 444446
rect 119356 444394 119384 448530
rect 120078 444680 120134 444689
rect 120078 444615 120134 444624
rect 120092 444446 120120 444615
rect 118752 444388 119384 444394
rect 118700 444382 119384 444388
rect 120080 444440 120132 444446
rect 120080 444382 120132 444388
rect 120724 444440 120776 444446
rect 120724 444382 120776 444388
rect 109512 444366 109802 444380
rect 111550 444366 111748 444380
rect 118712 444366 119384 444382
rect 120630 417072 120686 417081
rect 120630 417007 120686 417016
rect 85670 391096 85726 391105
rect 73344 391060 73396 391066
rect 85670 391031 85726 391040
rect 92754 391096 92810 391105
rect 92810 391068 93058 391082
rect 103822 391068 104112 391082
rect 92810 391054 93072 391068
rect 92754 391031 92810 391040
rect 73344 391002 73396 391008
rect 71870 390688 71926 390697
rect 71806 390660 71870 390674
rect 71792 390646 71870 390660
rect 69938 390416 69994 390425
rect 68480 390374 68770 390402
rect 68480 389162 68508 390374
rect 69994 390388 70334 390402
rect 69994 390374 70348 390388
rect 69938 390351 69994 390360
rect 68468 389156 68520 389162
rect 68468 389098 68520 389104
rect 67824 387116 67876 387122
rect 67824 387058 67876 387064
rect 67730 378856 67786 378865
rect 67730 378791 67786 378800
rect 70320 373318 70348 390374
rect 70308 373312 70360 373318
rect 70308 373254 70360 373260
rect 71688 371272 71740 371278
rect 71688 371214 71740 371220
rect 67732 369164 67784 369170
rect 67732 369106 67784 369112
rect 67640 369028 67692 369034
rect 67640 368970 67692 368976
rect 67744 354674 67772 369106
rect 69662 363760 69718 363769
rect 69662 363695 69718 363704
rect 67652 354646 67772 354674
rect 67546 299840 67602 299849
rect 67546 299775 67602 299784
rect 67362 290048 67418 290057
rect 67362 289983 67418 289992
rect 66904 289876 66956 289882
rect 66904 289818 66956 289824
rect 66824 287026 66944 287054
rect 66810 286784 66866 286793
rect 66810 286719 66866 286728
rect 66824 285734 66852 286719
rect 66812 285728 66864 285734
rect 66916 285705 66944 287026
rect 66812 285670 66864 285676
rect 66902 285696 66958 285705
rect 66902 285631 66958 285640
rect 66258 284608 66314 284617
rect 66258 284543 66314 284552
rect 66272 284374 66300 284543
rect 66260 284368 66312 284374
rect 66260 284310 66312 284316
rect 66996 284300 67048 284306
rect 66996 284242 67048 284248
rect 66810 282432 66866 282441
rect 66810 282367 66866 282376
rect 66824 281586 66852 282367
rect 66812 281580 66864 281586
rect 66812 281522 66864 281528
rect 66810 279168 66866 279177
rect 66810 279103 66866 279112
rect 66824 278798 66852 279103
rect 66812 278792 66864 278798
rect 66812 278734 66864 278740
rect 66902 278080 66958 278089
rect 66902 278015 66958 278024
rect 66350 276176 66406 276185
rect 66350 276111 66406 276120
rect 66364 276078 66392 276111
rect 66352 276072 66404 276078
rect 66352 276014 66404 276020
rect 66810 274000 66866 274009
rect 66810 273935 66866 273944
rect 66824 273290 66852 273935
rect 66812 273284 66864 273290
rect 66812 273226 66864 273232
rect 66718 272912 66774 272921
rect 66718 272847 66774 272856
rect 66732 271930 66760 272847
rect 66720 271924 66772 271930
rect 66720 271866 66772 271872
rect 66812 271856 66864 271862
rect 66810 271824 66812 271833
rect 66864 271824 66866 271833
rect 66810 271759 66866 271768
rect 66810 268560 66866 268569
rect 66810 268495 66866 268504
rect 66824 267850 66852 268495
rect 66812 267844 66864 267850
rect 66812 267786 66864 267792
rect 66916 267034 66944 278015
rect 67008 277273 67036 284242
rect 67546 283520 67602 283529
rect 67546 283455 67602 283464
rect 67454 281344 67510 281353
rect 67454 281279 67510 281288
rect 67178 280256 67234 280265
rect 67178 280191 67180 280200
rect 67232 280191 67234 280200
rect 67180 280162 67232 280168
rect 66994 277264 67050 277273
rect 66994 277199 67050 277208
rect 66904 267028 66956 267034
rect 66904 266970 66956 266976
rect 67178 266384 67234 266393
rect 67178 266319 67234 266328
rect 66902 265296 66958 265305
rect 66902 265231 66958 265240
rect 66916 264994 66944 265231
rect 66904 264988 66956 264994
rect 66904 264930 66956 264936
rect 66442 264208 66498 264217
rect 66442 264143 66498 264152
rect 66456 263634 66484 264143
rect 66444 263628 66496 263634
rect 66444 263570 66496 263576
rect 66902 263120 66958 263129
rect 66902 263055 66958 263064
rect 66916 262274 66944 263055
rect 66904 262268 66956 262274
rect 66904 262210 66956 262216
rect 66534 262032 66590 262041
rect 66534 261967 66590 261976
rect 66548 261526 66576 261967
rect 66536 261520 66588 261526
rect 66536 261462 66588 261468
rect 66350 260944 66406 260953
rect 66350 260879 66352 260888
rect 66404 260879 66406 260888
rect 66352 260850 66404 260856
rect 66260 258120 66312 258126
rect 66258 258088 66260 258097
rect 66312 258088 66314 258097
rect 66258 258023 66314 258032
rect 66810 257680 66866 257689
rect 66810 257615 66866 257624
rect 66824 256766 66852 257615
rect 66812 256760 66864 256766
rect 66812 256702 66864 256708
rect 66626 254416 66682 254425
rect 66626 254351 66682 254360
rect 66640 253978 66668 254351
rect 66628 253972 66680 253978
rect 66628 253914 66680 253920
rect 66810 253328 66866 253337
rect 66810 253263 66866 253272
rect 66824 252618 66852 253263
rect 66812 252612 66864 252618
rect 66812 252554 66864 252560
rect 66810 251152 66866 251161
rect 66810 251087 66866 251096
rect 66824 249830 66852 251087
rect 66812 249824 66864 249830
rect 66812 249766 66864 249772
rect 66812 247036 66864 247042
rect 66812 246978 66864 246984
rect 66824 246809 66852 246978
rect 66810 246800 66866 246809
rect 66810 246735 66866 246744
rect 66812 245608 66864 245614
rect 66812 245550 66864 245556
rect 66824 244633 66852 245550
rect 66810 244624 66866 244633
rect 66810 244559 66866 244568
rect 66812 244248 66864 244254
rect 66812 244190 66864 244196
rect 66824 243545 66852 244190
rect 66810 243536 66866 243545
rect 66810 243471 66866 243480
rect 66166 216608 66222 216617
rect 66166 216543 66222 216552
rect 64510 212528 64566 212537
rect 64510 212463 64566 212472
rect 63408 199436 63460 199442
rect 63408 199378 63460 199384
rect 62762 197976 62818 197985
rect 62762 197911 62818 197920
rect 61934 190360 61990 190369
rect 61934 190295 61990 190304
rect 66074 129296 66130 129305
rect 66074 129231 66130 129240
rect 65522 128072 65578 128081
rect 65522 128007 65578 128016
rect 65536 127022 65564 128007
rect 62028 127016 62080 127022
rect 62028 126958 62080 126964
rect 65524 127016 65576 127022
rect 65524 126958 65576 126964
rect 62040 77217 62068 126958
rect 64970 126304 65026 126313
rect 64970 126239 65026 126248
rect 64984 125633 65012 126239
rect 64786 125624 64842 125633
rect 64786 125559 64842 125568
rect 64970 125624 65026 125633
rect 64970 125559 65026 125568
rect 63408 121508 63460 121514
rect 63408 121450 63460 121456
rect 63420 84862 63448 121450
rect 63408 84856 63460 84862
rect 63408 84798 63460 84804
rect 64800 81433 64828 125559
rect 65982 122632 66038 122641
rect 65982 122567 66038 122576
rect 65996 121514 66024 122567
rect 65984 121508 66036 121514
rect 65984 121450 66036 121456
rect 66088 94518 66116 129231
rect 66166 125216 66222 125225
rect 66166 125151 66222 125160
rect 66076 94512 66128 94518
rect 66076 94454 66128 94460
rect 66180 82793 66208 125151
rect 66166 82784 66222 82793
rect 66166 82719 66222 82728
rect 64786 81424 64842 81433
rect 64786 81359 64842 81368
rect 62026 77208 62082 77217
rect 62026 77143 62082 77152
rect 64786 65648 64842 65657
rect 64786 65583 64842 65592
rect 62028 42084 62080 42090
rect 62028 42026 62080 42032
rect 60648 32428 60700 32434
rect 60648 32370 60700 32376
rect 61936 26920 61988 26926
rect 61936 26862 61988 26868
rect 59636 8968 59688 8974
rect 59636 8910 59688 8916
rect 58624 2168 58676 2174
rect 58624 2110 58676 2116
rect 59648 480 59676 8910
rect 61948 3058 61976 26862
rect 60832 3052 60884 3058
rect 60832 2994 60884 3000
rect 61936 3052 61988 3058
rect 61936 2994 61988 3000
rect 60844 480 60872 2994
rect 62040 480 62068 42026
rect 64800 3602 64828 65583
rect 66168 58676 66220 58682
rect 66168 58618 66220 58624
rect 64328 3596 64380 3602
rect 64328 3538 64380 3544
rect 64788 3596 64840 3602
rect 64788 3538 64840 3544
rect 63224 3528 63276 3534
rect 63224 3470 63276 3476
rect 63236 480 63264 3470
rect 64340 480 64368 3538
rect 66180 3534 66208 58618
rect 67192 47598 67220 266319
rect 67362 256592 67418 256601
rect 67362 256527 67418 256536
rect 67270 252240 67326 252249
rect 67270 252175 67326 252184
rect 67284 235793 67312 252175
rect 67270 235784 67326 235793
rect 67270 235719 67326 235728
rect 67376 224913 67404 256527
rect 67468 240038 67496 281279
rect 67560 262954 67588 283455
rect 67652 269657 67680 354646
rect 67732 354000 67784 354006
rect 67732 353942 67784 353948
rect 67744 324601 67772 353942
rect 69676 335354 69704 363695
rect 70308 362228 70360 362234
rect 70308 362170 70360 362176
rect 70320 335354 70348 362170
rect 71596 349852 71648 349858
rect 71596 349794 71648 349800
rect 71608 345014 71636 349794
rect 69308 335326 69704 335354
rect 70136 335326 70348 335354
rect 71516 344986 71636 345014
rect 67824 332648 67876 332654
rect 67824 332590 67876 332596
rect 67730 324592 67786 324601
rect 67730 324527 67786 324536
rect 67836 308553 67864 332590
rect 69308 331362 69336 335326
rect 69296 331356 69348 331362
rect 69296 331298 69348 331304
rect 69308 329474 69336 331298
rect 69388 329588 69440 329594
rect 69388 329530 69440 329536
rect 69400 329497 69428 329530
rect 69000 329446 69336 329474
rect 69386 329488 69442 329497
rect 70136 329474 70164 335326
rect 71516 331906 71544 344986
rect 71700 335354 71728 371214
rect 71608 335326 71728 335354
rect 70768 331900 70820 331906
rect 70768 331842 70820 331848
rect 71504 331900 71556 331906
rect 71504 331842 71556 331848
rect 70780 329474 70808 331842
rect 71608 329474 71636 335326
rect 71792 332654 71820 390646
rect 71870 390623 71926 390632
rect 73172 389094 73200 390388
rect 73160 389088 73212 389094
rect 73356 389065 73384 391002
rect 85684 390833 85712 391031
rect 85670 390824 85726 390833
rect 85606 390796 85670 390810
rect 85592 390782 85670 390796
rect 74552 390374 74842 390402
rect 76406 390374 76604 390402
rect 73804 389088 73856 389094
rect 73160 389030 73212 389036
rect 73342 389056 73398 389065
rect 73804 389030 73856 389036
rect 73342 388991 73398 389000
rect 73816 383722 73844 389030
rect 74552 388385 74580 390374
rect 74538 388376 74594 388385
rect 74538 388311 74594 388320
rect 76576 385014 76604 390374
rect 77864 389026 77892 390388
rect 77852 389020 77904 389026
rect 77852 388962 77904 388968
rect 77864 388385 77892 388962
rect 79520 388793 79548 390388
rect 79506 388784 79562 388793
rect 79506 388719 79562 388728
rect 79520 388550 79548 388719
rect 79508 388544 79560 388550
rect 79508 388486 79560 388492
rect 77850 388376 77906 388385
rect 77850 388311 77906 388320
rect 80900 386374 80928 390388
rect 82096 390374 82386 390402
rect 82096 387802 82124 390374
rect 82084 387796 82136 387802
rect 82084 387738 82136 387744
rect 80060 386368 80112 386374
rect 80060 386310 80112 386316
rect 80888 386368 80940 386374
rect 80888 386310 80940 386316
rect 76564 385008 76616 385014
rect 76564 384950 76616 384956
rect 73804 383716 73856 383722
rect 73804 383658 73856 383664
rect 73158 371920 73214 371929
rect 73158 371855 73214 371864
rect 72424 354068 72476 354074
rect 72424 354010 72476 354016
rect 72436 337414 72464 354010
rect 73066 345128 73122 345137
rect 73066 345063 73122 345072
rect 72424 337408 72476 337414
rect 72424 337350 72476 337356
rect 71780 332648 71832 332654
rect 71780 332590 71832 332596
rect 72240 331356 72292 331362
rect 72240 331298 72292 331304
rect 72252 329474 72280 331298
rect 73080 329474 73108 345063
rect 69736 329446 70164 329474
rect 70472 329446 70808 329474
rect 71208 329446 71636 329474
rect 71944 329446 72280 329474
rect 72680 329446 73108 329474
rect 73172 329474 73200 371855
rect 73816 371278 73844 383658
rect 76576 373289 76604 384950
rect 80072 381546 80100 386310
rect 80060 381540 80112 381546
rect 80060 381482 80112 381488
rect 81348 376032 81400 376038
rect 81348 375974 81400 375980
rect 77944 374672 77996 374678
rect 77944 374614 77996 374620
rect 76562 373280 76618 373289
rect 76562 373215 76618 373224
rect 73804 371272 73856 371278
rect 73804 371214 73856 371220
rect 75826 364984 75882 364993
rect 75826 364919 75882 364928
rect 75734 360224 75790 360233
rect 75734 360159 75790 360168
rect 74448 351280 74500 351286
rect 74448 351222 74500 351228
rect 74460 329474 74488 351222
rect 75644 333260 75696 333266
rect 75644 333202 75696 333208
rect 75656 331362 75684 333202
rect 75644 331356 75696 331362
rect 75644 331298 75696 331304
rect 75182 331256 75238 331265
rect 75182 331191 75238 331200
rect 75196 329474 75224 331191
rect 75748 329474 75776 360159
rect 75840 331265 75868 364919
rect 76564 356720 76616 356726
rect 76564 356662 76616 356668
rect 75826 331256 75882 331265
rect 75826 331191 75882 331200
rect 76576 329594 76604 356662
rect 77208 352640 77260 352646
rect 77208 352582 77260 352588
rect 77116 341556 77168 341562
rect 77116 341498 77168 341504
rect 77128 332178 77156 341498
rect 76656 332172 76708 332178
rect 76656 332114 76708 332120
rect 77116 332172 77168 332178
rect 77116 332114 77168 332120
rect 76564 329588 76616 329594
rect 76564 329530 76616 329536
rect 76668 329474 76696 332114
rect 77220 329474 77248 352582
rect 73172 329446 73416 329474
rect 74152 329446 74488 329474
rect 74888 329446 75224 329474
rect 75624 329446 75776 329474
rect 76360 329446 76696 329474
rect 77096 329446 77248 329474
rect 77482 329488 77538 329497
rect 69386 329423 69442 329432
rect 77956 329474 77984 374614
rect 79968 367804 80020 367810
rect 79968 367746 80020 367752
rect 79874 352744 79930 352753
rect 79874 352679 79930 352688
rect 78588 340264 78640 340270
rect 78588 340206 78640 340212
rect 78600 329746 78628 340206
rect 79888 335354 79916 352679
rect 77538 329446 77984 329474
rect 78554 329718 78628 329746
rect 79704 335326 79916 335354
rect 78554 329460 78582 329718
rect 79704 329474 79732 335326
rect 79980 331809 80008 367746
rect 81360 349178 81388 375974
rect 82096 360874 82124 387738
rect 83936 384985 83964 390388
rect 83922 384976 83978 384985
rect 83922 384911 83978 384920
rect 85592 370734 85620 390782
rect 85670 390759 85726 390768
rect 89810 390416 89866 390425
rect 87064 389298 87092 390388
rect 87052 389292 87104 389298
rect 87052 389234 87104 389240
rect 86224 388544 86276 388550
rect 86224 388486 86276 388492
rect 85580 370728 85632 370734
rect 85580 370670 85632 370676
rect 81624 360868 81676 360874
rect 81624 360810 81676 360816
rect 82084 360868 82136 360874
rect 82084 360810 82136 360816
rect 80152 349172 80204 349178
rect 80152 349114 80204 349120
rect 81348 349172 81400 349178
rect 81348 349114 81400 349120
rect 80164 345014 80192 349114
rect 81348 347064 81400 347070
rect 81348 347006 81400 347012
rect 80164 344986 80376 345014
rect 79966 331800 80022 331809
rect 79966 331735 79968 331744
rect 80020 331735 80022 331744
rect 79968 331706 80020 331712
rect 79980 331675 80008 331706
rect 80244 331628 80296 331634
rect 80244 331570 80296 331576
rect 80256 329474 80284 331570
rect 79304 329446 79732 329474
rect 80040 329446 80284 329474
rect 80348 329474 80376 344986
rect 81360 331634 81388 347006
rect 81636 345014 81664 360810
rect 84108 355360 84160 355366
rect 84108 355302 84160 355308
rect 81636 344986 81848 345014
rect 81438 342408 81494 342417
rect 81438 342343 81494 342352
rect 81348 331628 81400 331634
rect 81348 331570 81400 331576
rect 81452 329746 81480 342343
rect 81452 329718 81526 329746
rect 80348 329446 80776 329474
rect 81498 329460 81526 329718
rect 81820 329474 81848 344986
rect 83830 336016 83886 336025
rect 83830 335951 83886 335960
rect 83096 332172 83148 332178
rect 83096 332114 83148 332120
rect 83108 329474 83136 332114
rect 83844 329474 83872 335951
rect 84120 332178 84148 355302
rect 86236 351121 86264 388486
rect 86316 371204 86368 371210
rect 86316 371146 86368 371152
rect 86328 370734 86356 371146
rect 86316 370728 86368 370734
rect 86316 370670 86368 370676
rect 86222 351112 86278 351121
rect 86222 351047 86278 351056
rect 86328 349761 86356 370670
rect 86958 367296 87014 367305
rect 86958 367231 87014 367240
rect 86868 352572 86920 352578
rect 86868 352514 86920 352520
rect 86314 349752 86370 349761
rect 86314 349687 86370 349696
rect 85580 340944 85632 340950
rect 85580 340886 85632 340892
rect 85396 338428 85448 338434
rect 85396 338370 85448 338376
rect 84108 332172 84160 332178
rect 84108 332114 84160 332120
rect 84384 331764 84436 331770
rect 84384 331706 84436 331712
rect 81820 329446 82248 329474
rect 82800 329446 83136 329474
rect 83536 329446 83872 329474
rect 77482 329423 77538 329432
rect 84396 329202 84424 331706
rect 85408 329474 85436 338370
rect 85008 329446 85436 329474
rect 85592 329474 85620 340886
rect 86880 329474 86908 352514
rect 85592 329446 85744 329474
rect 86480 329446 86908 329474
rect 86972 329474 87000 367231
rect 87064 354074 87092 389234
rect 88536 388686 88564 390388
rect 91282 390416 91338 390425
rect 89866 390374 90404 390402
rect 89810 390351 89866 390360
rect 90376 389065 90404 390374
rect 91338 390374 92060 390402
rect 91282 390351 91338 390360
rect 90362 389056 90418 389065
rect 90362 388991 90418 389000
rect 88524 388680 88576 388686
rect 88524 388622 88576 388628
rect 89626 370560 89682 370569
rect 89626 370495 89682 370504
rect 89534 358048 89590 358057
rect 89534 357983 89590 357992
rect 87052 354068 87104 354074
rect 87052 354010 87104 354016
rect 87602 353968 87658 353977
rect 87602 353903 87658 353912
rect 87616 341562 87644 353903
rect 87604 341556 87656 341562
rect 87604 341498 87656 341504
rect 88248 331764 88300 331770
rect 88248 331706 88300 331712
rect 88260 329474 88288 331706
rect 88984 331492 89036 331498
rect 88984 331434 89036 331440
rect 88996 329474 89024 331434
rect 89548 329474 89576 357983
rect 89640 331498 89668 370495
rect 90376 364334 90404 388991
rect 91006 386472 91062 386481
rect 91006 386407 91062 386416
rect 90376 364306 90496 364334
rect 90468 351218 90496 364306
rect 90456 351212 90508 351218
rect 90456 351154 90508 351160
rect 90364 347812 90416 347818
rect 90364 347754 90416 347760
rect 90376 331770 90404 347754
rect 90468 338434 90496 351154
rect 90456 338428 90508 338434
rect 90456 338370 90508 338376
rect 90364 331764 90416 331770
rect 90364 331706 90416 331712
rect 89628 331492 89680 331498
rect 89628 331434 89680 331440
rect 90456 331492 90508 331498
rect 90456 331434 90508 331440
rect 90468 329474 90496 331434
rect 91020 329474 91048 386407
rect 92032 383654 92060 390374
rect 92480 388680 92532 388686
rect 92478 388648 92480 388657
rect 92532 388648 92534 388657
rect 92478 388583 92534 388592
rect 93044 388482 93072 391054
rect 103808 391066 104112 391068
rect 103808 391060 104124 391066
rect 103808 391054 104072 391060
rect 102138 390552 102194 390561
rect 102194 390524 102258 390538
rect 102194 390510 102272 390524
rect 102138 390487 102194 390496
rect 94226 390416 94282 390425
rect 97354 390416 97410 390425
rect 94282 390374 95004 390402
rect 94226 390351 94282 390360
rect 93766 388648 93822 388657
rect 93766 388583 93822 388592
rect 93032 388476 93084 388482
rect 93032 388418 93084 388424
rect 92032 383626 92244 383654
rect 91098 365800 91154 365809
rect 91098 365735 91154 365744
rect 91112 345014 91140 365735
rect 92216 360942 92244 383626
rect 92294 377360 92350 377369
rect 92294 377295 92350 377304
rect 92308 365809 92336 377295
rect 93122 367568 93178 367577
rect 93122 367503 93178 367512
rect 92294 365800 92350 365809
rect 92294 365735 92350 365744
rect 92204 360936 92256 360942
rect 92204 360878 92256 360884
rect 92386 345808 92442 345817
rect 92386 345743 92442 345752
rect 91112 344986 92060 345014
rect 91928 332172 91980 332178
rect 91928 332114 91980 332120
rect 91940 329474 91968 332114
rect 86972 329446 87216 329474
rect 87952 329446 88288 329474
rect 88688 329446 89024 329474
rect 89424 329446 89576 329474
rect 90160 329446 90496 329474
rect 90896 329446 91048 329474
rect 91632 329446 91968 329474
rect 92032 329474 92060 344986
rect 92400 332178 92428 345743
rect 92388 332172 92440 332178
rect 92388 332114 92440 332120
rect 93136 331498 93164 367503
rect 93780 357406 93808 388583
rect 94976 383654 95004 390374
rect 96172 389162 96200 390388
rect 98826 390416 98882 390425
rect 97410 390374 97856 390402
rect 97354 390351 97410 390360
rect 96160 389156 96212 389162
rect 96160 389098 96212 389104
rect 96172 389065 96200 389098
rect 96158 389056 96214 389065
rect 96158 388991 96214 389000
rect 95238 388512 95294 388521
rect 95238 388447 95294 388456
rect 94976 383626 95188 383654
rect 95160 379545 95188 383626
rect 95146 379536 95202 379545
rect 95146 379471 95202 379480
rect 93768 357400 93820 357406
rect 93768 357342 93820 357348
rect 95160 343777 95188 379471
rect 95252 376038 95280 388447
rect 95240 376032 95292 376038
rect 95240 375974 95292 375980
rect 96528 355428 96580 355434
rect 96528 355370 96580 355376
rect 95146 343768 95202 343777
rect 95146 343703 95202 343712
rect 95160 340270 95188 343703
rect 95148 340264 95200 340270
rect 95148 340206 95200 340212
rect 93492 340196 93544 340202
rect 93492 340138 93544 340144
rect 93124 331492 93176 331498
rect 93124 331434 93176 331440
rect 93504 329474 93532 340138
rect 95148 339516 95200 339522
rect 95148 339458 95200 339464
rect 94228 336048 94280 336054
rect 94228 335990 94280 335996
rect 94136 331492 94188 331498
rect 94136 331434 94188 331440
rect 94148 329474 94176 331434
rect 94240 331265 94268 335990
rect 95160 331498 95188 339458
rect 96342 338736 96398 338745
rect 96342 338671 96398 338680
rect 96356 332178 96384 338671
rect 96540 335354 96568 355370
rect 97828 341601 97856 390374
rect 98882 390374 99328 390402
rect 98826 390351 98882 390360
rect 98644 388476 98696 388482
rect 98644 388418 98696 388424
rect 98656 369238 98684 388418
rect 99196 385756 99248 385762
rect 99196 385698 99248 385704
rect 98644 369232 98696 369238
rect 98644 369174 98696 369180
rect 99208 355473 99236 385698
rect 99300 385665 99328 390374
rect 100772 390289 100800 390388
rect 100758 390280 100814 390289
rect 100758 390215 100814 390224
rect 99286 385656 99342 385665
rect 99286 385591 99342 385600
rect 99286 371376 99342 371385
rect 99286 371311 99342 371320
rect 99194 355464 99250 355473
rect 99194 355399 99196 355408
rect 99248 355399 99250 355408
rect 99196 355370 99248 355376
rect 99208 355339 99236 355370
rect 99194 349752 99250 349761
rect 99194 349687 99250 349696
rect 97814 341592 97870 341601
rect 97814 341527 97870 341536
rect 97080 337408 97132 337414
rect 97080 337350 97132 337356
rect 96448 335326 96568 335354
rect 95608 332172 95660 332178
rect 95608 332114 95660 332120
rect 96344 332172 96396 332178
rect 96344 332114 96396 332120
rect 95148 331492 95200 331498
rect 95148 331434 95200 331440
rect 94226 331256 94282 331265
rect 94226 331191 94282 331200
rect 94870 331256 94926 331265
rect 94870 331191 94926 331200
rect 94884 329474 94912 331191
rect 95620 329474 95648 332114
rect 96448 329474 96476 335326
rect 97092 329474 97120 337350
rect 97814 335744 97870 335753
rect 97814 335679 97870 335688
rect 97828 329474 97856 335679
rect 98552 331492 98604 331498
rect 98552 331434 98604 331440
rect 98564 329474 98592 331434
rect 99208 329474 99236 349687
rect 99300 331498 99328 371311
rect 100772 360233 100800 390215
rect 102244 389337 102272 390510
rect 102230 389328 102286 389337
rect 102230 389263 102286 389272
rect 103808 389094 103836 391054
rect 104072 391002 104124 391008
rect 104990 390416 105046 390425
rect 106554 390416 106610 390425
rect 105046 390374 105386 390402
rect 104990 390351 105046 390360
rect 108026 390416 108082 390425
rect 106610 390374 107332 390402
rect 106554 390351 106610 390360
rect 101404 389088 101456 389094
rect 101404 389030 101456 389036
rect 103796 389088 103848 389094
rect 103796 389030 103848 389036
rect 100758 360224 100814 360233
rect 100758 360159 100814 360168
rect 101126 360224 101182 360233
rect 101126 360159 101182 360168
rect 101140 359582 101168 360159
rect 101128 359576 101180 359582
rect 101128 359518 101180 359524
rect 99378 353560 99434 353569
rect 99378 353495 99434 353504
rect 99392 352578 99420 353495
rect 100666 352608 100722 352617
rect 99380 352572 99432 352578
rect 100666 352543 100722 352552
rect 99380 352514 99432 352520
rect 100574 345672 100630 345681
rect 100574 345607 100630 345616
rect 100588 332178 100616 345607
rect 100024 332172 100076 332178
rect 100024 332114 100076 332120
rect 100576 332172 100628 332178
rect 100576 332114 100628 332120
rect 99288 331492 99340 331498
rect 99288 331434 99340 331440
rect 100036 329474 100064 332114
rect 100680 329474 100708 352543
rect 100758 340096 100814 340105
rect 100758 340031 100814 340040
rect 92032 329446 92368 329474
rect 93104 329446 93532 329474
rect 93840 329446 94176 329474
rect 94576 329446 94912 329474
rect 95312 329446 95648 329474
rect 96048 329446 96476 329474
rect 96784 329446 97120 329474
rect 97520 329446 97856 329474
rect 98256 329446 98592 329474
rect 98992 329446 99236 329474
rect 99728 329446 100064 329474
rect 100464 329446 100708 329474
rect 100772 329474 100800 340031
rect 101416 331809 101444 389030
rect 105004 380934 105032 390351
rect 107304 390266 107332 390374
rect 109498 390416 109554 390425
rect 108082 390388 108422 390402
rect 108082 390374 108436 390388
rect 108026 390351 108082 390360
rect 107304 390238 107608 390266
rect 107474 388512 107530 388521
rect 107474 388447 107530 388456
rect 104992 380928 105044 380934
rect 104992 380870 105044 380876
rect 105544 380928 105596 380934
rect 105544 380870 105596 380876
rect 104164 375488 104216 375494
rect 104164 375430 104216 375436
rect 103426 360904 103482 360913
rect 103426 360839 103482 360848
rect 102048 354748 102100 354754
rect 102048 354690 102100 354696
rect 101402 331800 101458 331809
rect 101402 331735 101458 331744
rect 102060 329474 102088 354690
rect 103440 332178 103468 360839
rect 104176 337385 104204 375430
rect 104900 364404 104952 364410
rect 104900 364346 104952 364352
rect 104162 337376 104218 337385
rect 104162 337311 104218 337320
rect 104440 334008 104492 334014
rect 104440 333950 104492 333956
rect 102968 332172 103020 332178
rect 102968 332114 103020 332120
rect 103428 332172 103480 332178
rect 103428 332114 103480 332120
rect 102980 329474 103008 332114
rect 103242 331800 103298 331809
rect 103242 331735 103298 331744
rect 100772 329446 101200 329474
rect 101936 329446 102088 329474
rect 102672 329446 103008 329474
rect 84272 329174 84424 329202
rect 103256 329202 103284 331735
rect 104452 329474 104480 333950
rect 104912 329746 104940 364346
rect 105556 352578 105584 380870
rect 105544 352572 105596 352578
rect 105544 352514 105596 352520
rect 107488 351937 107516 388447
rect 106922 351928 106978 351937
rect 106922 351863 106978 351872
rect 107474 351928 107530 351937
rect 107474 351863 107530 351872
rect 104990 349072 105046 349081
rect 104990 349007 105046 349016
rect 105004 345014 105032 349007
rect 105004 344986 105216 345014
rect 104144 329446 104480 329474
rect 104866 329718 104940 329746
rect 104866 329460 104894 329718
rect 105188 329474 105216 344986
rect 106280 338156 106332 338162
rect 106280 338098 106332 338104
rect 106292 329746 106320 338098
rect 106936 336025 106964 351863
rect 107580 343058 107608 390238
rect 108408 389473 108436 390374
rect 115938 390416 115994 390425
rect 109554 390374 110276 390402
rect 109498 390351 109554 390360
rect 108394 389464 108450 389473
rect 108394 389399 108450 389408
rect 109684 380928 109736 380934
rect 109684 380870 109736 380876
rect 107752 366376 107804 366382
rect 107752 366318 107804 366324
rect 107764 357474 107792 366318
rect 108762 361720 108818 361729
rect 108762 361655 108818 361664
rect 107752 357468 107804 357474
rect 107752 357410 107804 357416
rect 107764 345014 107792 357410
rect 108776 355366 108804 361655
rect 109696 358086 109724 380870
rect 110248 378826 110276 390374
rect 111444 389230 111472 390388
rect 111432 389224 111484 389230
rect 111432 389166 111484 389172
rect 111444 385694 111472 389166
rect 112916 389065 112944 390388
rect 113088 389836 113140 389842
rect 113088 389778 113140 389784
rect 112902 389056 112958 389065
rect 112902 388991 112958 389000
rect 111432 385688 111484 385694
rect 111432 385630 111484 385636
rect 110236 378820 110288 378826
rect 110236 378762 110288 378768
rect 110328 362976 110380 362982
rect 110328 362918 110380 362924
rect 109684 358080 109736 358086
rect 109684 358022 109736 358028
rect 108764 355360 108816 355366
rect 108764 355302 108816 355308
rect 108304 347132 108356 347138
rect 108304 347074 108356 347080
rect 107764 344986 107976 345014
rect 107568 343052 107620 343058
rect 107568 342994 107620 343000
rect 107476 342916 107528 342922
rect 107476 342858 107528 342864
rect 106922 336016 106978 336025
rect 106922 335951 106978 335960
rect 106292 329718 106366 329746
rect 105188 329446 105616 329474
rect 106338 329460 106366 329718
rect 107488 329474 107516 342858
rect 107844 336796 107896 336802
rect 107844 336738 107896 336744
rect 107856 329474 107884 336738
rect 107088 329446 107516 329474
rect 107640 329446 107884 329474
rect 107948 329474 107976 344986
rect 108316 334626 108344 347074
rect 110234 339688 110290 339697
rect 110234 339623 110290 339632
rect 108304 334620 108356 334626
rect 108304 334562 108356 334568
rect 109408 331560 109460 331566
rect 109408 331502 109460 331508
rect 109420 329474 109448 331502
rect 110248 329474 110276 339623
rect 110340 331566 110368 362918
rect 113100 361622 113128 389778
rect 114480 387802 114508 390388
rect 118790 390416 118846 390425
rect 115994 390388 116150 390402
rect 115994 390374 116164 390388
rect 115938 390351 115994 390360
rect 116136 389065 116164 390374
rect 117608 389065 117636 390388
rect 118846 390388 119002 390402
rect 118846 390374 119016 390388
rect 118790 390351 118846 390360
rect 116122 389056 116178 389065
rect 116122 388991 116178 389000
rect 117134 389056 117190 389065
rect 117134 388991 117190 389000
rect 117594 389056 117650 389065
rect 117594 388991 117650 389000
rect 118606 389056 118662 389065
rect 118606 388991 118662 389000
rect 114468 387796 114520 387802
rect 114468 387738 114520 387744
rect 114480 367946 114508 387738
rect 117148 378049 117176 388991
rect 118620 382974 118648 388991
rect 118988 388482 119016 390374
rect 120460 390318 120488 390388
rect 120448 390312 120500 390318
rect 120448 390254 120500 390260
rect 120460 388521 120488 390254
rect 120644 389842 120672 417007
rect 120632 389836 120684 389842
rect 120632 389778 120684 389784
rect 120446 388512 120502 388521
rect 118976 388476 119028 388482
rect 120446 388447 120502 388456
rect 118976 388418 119028 388424
rect 118988 387025 119016 388418
rect 118974 387016 119030 387025
rect 118974 386951 119030 386960
rect 118608 382968 118660 382974
rect 118608 382910 118660 382916
rect 116582 378040 116638 378049
rect 116582 377975 116638 377984
rect 117134 378040 117190 378049
rect 117134 377975 117190 377984
rect 116596 376825 116624 377975
rect 116582 376816 116638 376825
rect 116582 376751 116638 376760
rect 114558 372736 114614 372745
rect 114558 372671 114614 372680
rect 113824 367940 113876 367946
rect 113824 367882 113876 367888
rect 114468 367940 114520 367946
rect 114468 367882 114520 367888
rect 113836 367130 113864 367882
rect 113824 367124 113876 367130
rect 113824 367066 113876 367072
rect 111800 361616 111852 361622
rect 111800 361558 111852 361564
rect 113088 361616 113140 361622
rect 113088 361558 113140 361564
rect 111062 357640 111118 357649
rect 111062 357575 111118 357584
rect 111076 352753 111104 357575
rect 111708 355360 111760 355366
rect 111708 355302 111760 355308
rect 111062 352744 111118 352753
rect 111062 352679 111118 352688
rect 111614 342272 111670 342281
rect 111614 342207 111670 342216
rect 110328 331560 110380 331566
rect 110328 331502 110380 331508
rect 110880 331356 110932 331362
rect 110880 331298 110932 331304
rect 110892 329474 110920 331298
rect 111628 329474 111656 342207
rect 111720 331362 111748 355302
rect 111708 331356 111760 331362
rect 111708 331298 111760 331304
rect 107948 329446 108376 329474
rect 109112 329446 109448 329474
rect 109848 329446 110276 329474
rect 110584 329446 110920 329474
rect 111320 329446 111656 329474
rect 111812 329474 111840 361558
rect 113836 351286 113864 367066
rect 114468 353320 114520 353326
rect 114468 353262 114520 353268
rect 113824 351280 113876 351286
rect 113824 351222 113876 351228
rect 114374 350568 114430 350577
rect 114374 350503 114430 350512
rect 112352 338224 112404 338230
rect 112352 338166 112404 338172
rect 112364 329474 112392 338166
rect 114388 332178 114416 350503
rect 113824 332172 113876 332178
rect 113824 332114 113876 332120
rect 114376 332172 114428 332178
rect 114376 332114 114428 332120
rect 113836 329474 113864 332114
rect 114480 329474 114508 353262
rect 111812 329446 112056 329474
rect 112364 329446 112792 329474
rect 113528 329446 113864 329474
rect 114264 329446 114508 329474
rect 114572 329474 114600 372671
rect 114650 339960 114706 339969
rect 114650 339895 114706 339904
rect 114664 329730 114692 339895
rect 116596 338881 116624 376751
rect 119986 375320 120042 375329
rect 119986 375255 120042 375264
rect 120000 374066 120028 375255
rect 119988 374060 120040 374066
rect 119988 374002 120040 374008
rect 117964 371340 118016 371346
rect 117964 371282 118016 371288
rect 117976 354006 118004 371282
rect 117964 354000 118016 354006
rect 117964 353942 118016 353948
rect 118882 349208 118938 349217
rect 118882 349143 118938 349152
rect 118896 345014 118924 349143
rect 119894 346488 119950 346497
rect 119894 346423 119950 346432
rect 118896 344986 119016 345014
rect 117228 341012 117280 341018
rect 117228 340954 117280 340960
rect 116582 338872 116638 338881
rect 116582 338807 116638 338816
rect 117042 334112 117098 334121
rect 117042 334047 117098 334056
rect 116768 332172 116820 332178
rect 116768 332114 116820 332120
rect 114652 329724 114704 329730
rect 114652 329666 114704 329672
rect 115710 329724 115762 329730
rect 115710 329666 115762 329672
rect 115722 329474 115750 329666
rect 116780 329474 116808 332114
rect 114572 329446 115000 329474
rect 115400 329460 115750 329474
rect 115400 329446 115736 329460
rect 116472 329446 116808 329474
rect 103256 329174 103408 329202
rect 115400 329118 115428 329446
rect 117056 329338 117084 334047
rect 117240 332178 117268 340954
rect 118240 336048 118292 336054
rect 118240 335990 118292 335996
rect 117228 332172 117280 332178
rect 117228 332114 117280 332120
rect 118252 329474 118280 335990
rect 118884 331628 118936 331634
rect 118884 331570 118936 331576
rect 118896 329474 118924 331570
rect 117944 329446 118280 329474
rect 118680 329446 118924 329474
rect 118988 329474 119016 344986
rect 119908 331634 119936 346423
rect 119896 331628 119948 331634
rect 119896 331570 119948 331576
rect 120000 331362 120028 374002
rect 120736 353977 120764 444382
rect 120828 390318 120856 462946
rect 121380 429214 121408 567190
rect 121460 556300 121512 556306
rect 121460 556242 121512 556248
rect 121368 429208 121420 429214
rect 121368 429150 121420 429156
rect 121472 392601 121500 556242
rect 121564 417489 121592 570590
rect 122208 558958 122236 574058
rect 122104 558952 122156 558958
rect 122104 558894 122156 558900
rect 122196 558952 122248 558958
rect 122196 558894 122248 558900
rect 122932 558952 122984 558958
rect 122932 558894 122984 558900
rect 121644 451920 121696 451926
rect 121644 451862 121696 451868
rect 121656 440230 121684 451862
rect 121644 440224 121696 440230
rect 121644 440166 121696 440172
rect 121656 440065 121684 440166
rect 121642 440056 121698 440065
rect 121642 439991 121698 440000
rect 121644 429208 121696 429214
rect 121644 429150 121696 429156
rect 121656 428505 121684 429150
rect 121642 428496 121698 428505
rect 121642 428431 121698 428440
rect 121550 417480 121606 417489
rect 121550 417415 121606 417424
rect 122116 397361 122144 558894
rect 122746 428496 122802 428505
rect 122746 428431 122802 428440
rect 122102 397352 122158 397361
rect 122102 397287 122158 397296
rect 121552 396024 121604 396030
rect 121552 395966 121604 395972
rect 121564 394913 121592 395966
rect 121550 394904 121606 394913
rect 121550 394839 121606 394848
rect 121458 392592 121514 392601
rect 121458 392527 121514 392536
rect 121472 392018 121500 392527
rect 121460 392012 121512 392018
rect 121460 391954 121512 391960
rect 120816 390312 120868 390318
rect 120816 390254 120868 390260
rect 121564 382945 121592 394839
rect 121550 382936 121606 382945
rect 121550 382871 121606 382880
rect 122760 368529 122788 428431
rect 122944 421977 122972 558894
rect 123022 447808 123078 447817
rect 123022 447743 123078 447752
rect 123036 435305 123064 447743
rect 123022 435296 123078 435305
rect 123022 435231 123078 435240
rect 123022 426048 123078 426057
rect 123022 425983 123078 425992
rect 122930 421968 122986 421977
rect 122930 421903 122986 421912
rect 122944 421598 122972 421903
rect 122932 421592 122984 421598
rect 122932 421534 122984 421540
rect 122932 415200 122984 415206
rect 122930 415168 122932 415177
rect 122984 415168 122986 415177
rect 122930 415103 122986 415112
rect 122944 385762 122972 415103
rect 122932 385756 122984 385762
rect 122932 385698 122984 385704
rect 122102 368520 122158 368529
rect 122102 368455 122158 368464
rect 122746 368520 122802 368529
rect 122746 368455 122802 368464
rect 120816 360936 120868 360942
rect 120816 360878 120868 360884
rect 120722 353968 120778 353977
rect 120722 353903 120778 353912
rect 120828 350606 120856 360878
rect 121460 353388 121512 353394
rect 121460 353330 121512 353336
rect 120080 350600 120132 350606
rect 120080 350542 120132 350548
rect 120816 350600 120868 350606
rect 120816 350542 120868 350548
rect 119988 331356 120040 331362
rect 119988 331298 120040 331304
rect 120092 329746 120120 350542
rect 121472 349858 121500 353330
rect 121552 349920 121604 349926
rect 121552 349862 121604 349868
rect 121460 349852 121512 349858
rect 121460 349794 121512 349800
rect 121564 335354 121592 349862
rect 121736 348424 121788 348430
rect 121736 348366 121788 348372
rect 121748 345014 121776 348366
rect 122116 347138 122144 368455
rect 123036 356726 123064 425983
rect 123128 424153 123156 576098
rect 124876 541686 124904 700334
rect 129004 700324 129056 700330
rect 129004 700266 129056 700272
rect 127440 566500 127492 566506
rect 127440 566442 127492 566448
rect 127452 565894 127480 566442
rect 126980 565888 127032 565894
rect 126980 565830 127032 565836
rect 127440 565888 127492 565894
rect 127440 565830 127492 565836
rect 124956 552084 125008 552090
rect 124956 552026 125008 552032
rect 124864 541680 124916 541686
rect 124864 541622 124916 541628
rect 124862 538792 124918 538801
rect 124862 538727 124918 538736
rect 124220 534812 124272 534818
rect 124220 534754 124272 534760
rect 123576 449268 123628 449274
rect 123576 449210 123628 449216
rect 123114 424144 123170 424153
rect 123114 424079 123170 424088
rect 123482 424144 123538 424153
rect 123482 424079 123538 424088
rect 123496 385082 123524 424079
rect 123588 411369 123616 449210
rect 124128 444372 124180 444378
rect 124128 444314 124180 444320
rect 124140 444281 124168 444314
rect 124126 444272 124182 444281
rect 124126 444207 124182 444216
rect 124126 442096 124182 442105
rect 124126 442031 124182 442040
rect 124140 441658 124168 442031
rect 124128 441652 124180 441658
rect 124128 441594 124180 441600
rect 124128 438864 124180 438870
rect 124128 438806 124180 438812
rect 124140 437889 124168 438806
rect 124126 437880 124182 437889
rect 124126 437815 124182 437824
rect 124128 433356 124180 433362
rect 124128 433298 124180 433304
rect 124140 433265 124168 433298
rect 124126 433256 124182 433265
rect 124126 433191 124182 433200
rect 124036 431928 124088 431934
rect 124036 431870 124088 431876
rect 124048 431089 124076 431870
rect 124034 431080 124090 431089
rect 124034 431015 124090 431024
rect 124128 412752 124180 412758
rect 124126 412720 124128 412729
rect 124180 412720 124182 412729
rect 124126 412655 124182 412664
rect 123574 411360 123630 411369
rect 123574 411295 123630 411304
rect 124126 408368 124182 408377
rect 124126 408303 124182 408312
rect 124140 407794 124168 408303
rect 124128 407788 124180 407794
rect 124128 407730 124180 407736
rect 124128 406224 124180 406230
rect 124126 406192 124128 406201
rect 124180 406192 124182 406201
rect 124126 406127 124182 406136
rect 123850 403744 123906 403753
rect 123850 403679 123906 403688
rect 123864 403374 123892 403679
rect 123852 403368 123904 403374
rect 123852 403310 123904 403316
rect 123942 401568 123998 401577
rect 123942 401503 123998 401512
rect 123956 400926 123984 401503
rect 123944 400920 123996 400926
rect 123944 400862 123996 400868
rect 124126 399392 124182 399401
rect 124126 399327 124182 399336
rect 124140 398886 124168 399327
rect 124128 398880 124180 398886
rect 124128 398822 124180 398828
rect 123758 397352 123814 397361
rect 123758 397287 123814 397296
rect 123772 393990 123800 397287
rect 123760 393984 123812 393990
rect 123760 393926 123812 393932
rect 123484 385076 123536 385082
rect 123484 385018 123536 385024
rect 123496 369170 123524 385018
rect 124232 384985 124260 534754
rect 124876 529922 124904 538727
rect 124864 529916 124916 529922
rect 124864 529858 124916 529864
rect 124968 529854 124996 552026
rect 126886 549400 126942 549409
rect 126886 549335 126942 549344
rect 125048 534812 125100 534818
rect 125048 534754 125100 534760
rect 125060 534138 125088 534754
rect 125048 534132 125100 534138
rect 125048 534074 125100 534080
rect 124956 529848 125008 529854
rect 124956 529790 125008 529796
rect 124864 477556 124916 477562
rect 124864 477498 124916 477504
rect 124312 451988 124364 451994
rect 124312 451930 124364 451936
rect 124324 444378 124352 451930
rect 124876 451246 124904 477498
rect 125600 453348 125652 453354
rect 125600 453290 125652 453296
rect 124864 451240 124916 451246
rect 124864 451182 124916 451188
rect 124864 447160 124916 447166
rect 124864 447102 124916 447108
rect 124312 444372 124364 444378
rect 124312 444314 124364 444320
rect 124312 420912 124364 420918
rect 124310 420880 124312 420889
rect 124364 420880 124366 420889
rect 124310 420815 124366 420824
rect 124324 419665 124352 420815
rect 124310 419656 124366 419665
rect 124310 419591 124366 419600
rect 124218 384976 124274 384985
rect 124218 384911 124274 384920
rect 124402 382528 124458 382537
rect 124402 382463 124458 382472
rect 124416 378078 124444 382463
rect 124404 378072 124456 378078
rect 124404 378014 124456 378020
rect 123484 369164 123536 369170
rect 123484 369106 123536 369112
rect 124126 364440 124182 364449
rect 124126 364375 124182 364384
rect 123024 356720 123076 356726
rect 124036 356720 124088 356726
rect 123024 356662 123076 356668
rect 124034 356688 124036 356697
rect 124088 356688 124090 356697
rect 124034 356623 124090 356632
rect 122194 356280 122250 356289
rect 122194 356215 122250 356224
rect 122104 347132 122156 347138
rect 122104 347074 122156 347080
rect 121748 344986 121960 345014
rect 121472 335326 121592 335354
rect 120540 331356 120592 331362
rect 120540 331298 120592 331304
rect 120092 329718 120166 329746
rect 118988 329446 119416 329474
rect 120138 329460 120166 329718
rect 120552 329474 120580 331298
rect 121472 329474 121500 335326
rect 121932 329474 121960 344986
rect 122208 340202 122236 356215
rect 122196 340196 122248 340202
rect 122196 340138 122248 340144
rect 124140 331634 124168 364375
rect 124876 345710 124904 447102
rect 124956 445800 125008 445806
rect 124956 445742 125008 445748
rect 124968 436762 124996 445742
rect 124956 436756 125008 436762
rect 124956 436698 125008 436704
rect 125612 406994 125640 453290
rect 125692 413976 125744 413982
rect 125692 413918 125744 413924
rect 125704 412758 125732 413918
rect 125692 412752 125744 412758
rect 125692 412694 125744 412700
rect 125520 406966 125640 406994
rect 125520 406230 125548 406966
rect 125508 406224 125560 406230
rect 125508 406166 125560 406172
rect 124956 403368 125008 403374
rect 124956 403310 125008 403316
rect 124968 378078 124996 403310
rect 125520 402354 125548 406166
rect 125508 402348 125560 402354
rect 125508 402290 125560 402296
rect 125600 398880 125652 398886
rect 125600 398822 125652 398828
rect 125048 397520 125100 397526
rect 125048 397462 125100 397468
rect 125060 389162 125088 397462
rect 125048 389156 125100 389162
rect 125048 389098 125100 389104
rect 125612 383654 125640 398822
rect 125600 383648 125652 383654
rect 125600 383590 125652 383596
rect 125704 380186 125732 412694
rect 125692 380180 125744 380186
rect 125692 380122 125744 380128
rect 124956 378072 125008 378078
rect 124956 378014 125008 378020
rect 126244 365832 126296 365838
rect 126244 365774 126296 365780
rect 125506 360224 125562 360233
rect 125506 360159 125562 360168
rect 124954 351112 125010 351121
rect 124954 351047 125010 351056
rect 124864 345704 124916 345710
rect 124864 345646 124916 345652
rect 123392 331628 123444 331634
rect 123392 331570 123444 331576
rect 124128 331628 124180 331634
rect 124128 331570 124180 331576
rect 123404 329474 123432 331570
rect 124876 331498 124904 345646
rect 124968 338337 124996 351047
rect 124954 338328 125010 338337
rect 124954 338263 125010 338272
rect 124128 331492 124180 331498
rect 124128 331434 124180 331440
rect 124864 331492 124916 331498
rect 124864 331434 124916 331440
rect 124140 329474 124168 331434
rect 124678 331392 124734 331401
rect 124678 331327 124734 331336
rect 120552 329446 120888 329474
rect 121472 329446 121624 329474
rect 121932 329446 122360 329474
rect 123096 329446 123432 329474
rect 123832 329446 124168 329474
rect 124692 329338 124720 331327
rect 124968 329905 124996 338263
rect 125520 331401 125548 360159
rect 126256 349926 126284 365774
rect 126244 349920 126296 349926
rect 126244 349862 126296 349868
rect 126796 349240 126848 349246
rect 126796 349182 126848 349188
rect 126808 348945 126836 349182
rect 125598 348936 125654 348945
rect 125598 348871 125654 348880
rect 126794 348936 126850 348945
rect 126794 348871 126850 348880
rect 125506 331392 125562 331401
rect 125506 331327 125562 331336
rect 124954 329896 125010 329905
rect 125612 329866 125640 348871
rect 126900 340241 126928 549335
rect 126992 413982 127020 565830
rect 128360 550724 128412 550730
rect 128360 550666 128412 550672
rect 127624 488572 127676 488578
rect 127624 488514 127676 488520
rect 126980 413976 127032 413982
rect 126980 413918 127032 413924
rect 127636 396030 127664 488514
rect 127716 458244 127768 458250
rect 127716 458186 127768 458192
rect 127728 451178 127756 458186
rect 127716 451172 127768 451178
rect 127716 451114 127768 451120
rect 127716 444508 127768 444514
rect 127716 444450 127768 444456
rect 127624 396024 127676 396030
rect 127624 395966 127676 395972
rect 127728 359514 127756 444450
rect 127808 402348 127860 402354
rect 127808 402290 127860 402296
rect 126980 359508 127032 359514
rect 126980 359450 127032 359456
rect 127716 359508 127768 359514
rect 127716 359450 127768 359456
rect 126992 345014 127020 359450
rect 126992 344986 127112 345014
rect 126334 340232 126390 340241
rect 126334 340167 126390 340176
rect 126886 340232 126942 340241
rect 126886 340167 126942 340176
rect 124954 329831 125010 329840
rect 125600 329860 125652 329866
rect 124968 329474 124996 329831
rect 125600 329802 125652 329808
rect 125612 329474 125640 329802
rect 126348 329474 126376 340167
rect 127084 329474 127112 344986
rect 127820 342553 127848 402290
rect 128372 387802 128400 550666
rect 129016 538218 129044 700266
rect 141424 594856 141476 594862
rect 141424 594798 141476 594804
rect 132500 584452 132552 584458
rect 132500 584394 132552 584400
rect 129740 569220 129792 569226
rect 129740 569162 129792 569168
rect 129752 568614 129780 569162
rect 129740 568608 129792 568614
rect 129740 568550 129792 568556
rect 129004 538212 129056 538218
rect 129004 538154 129056 538160
rect 129648 536852 129700 536858
rect 129648 536794 129700 536800
rect 128452 452668 128504 452674
rect 128452 452610 128504 452616
rect 128360 387796 128412 387802
rect 128360 387738 128412 387744
rect 127806 342544 127862 342553
rect 127806 342479 127862 342488
rect 127820 329474 127848 342479
rect 128464 337414 128492 452610
rect 129660 343913 129688 536794
rect 129752 415206 129780 568550
rect 131580 541680 131632 541686
rect 131580 541622 131632 541628
rect 131592 541074 131620 541622
rect 131120 541068 131172 541074
rect 131120 541010 131172 541016
rect 131580 541068 131632 541074
rect 131580 541010 131632 541016
rect 130384 445052 130436 445058
rect 130384 444994 130436 445000
rect 129740 415200 129792 415206
rect 129740 415142 129792 415148
rect 130396 369073 130424 444994
rect 130476 444440 130528 444446
rect 130476 444382 130528 444388
rect 130488 409834 130516 444382
rect 130476 409828 130528 409834
rect 130476 409770 130528 409776
rect 131132 391270 131160 541010
rect 131764 465112 131816 465118
rect 131764 465054 131816 465060
rect 131776 440230 131804 465054
rect 131764 440224 131816 440230
rect 131764 440166 131816 440172
rect 132512 438870 132540 584394
rect 134524 565140 134576 565146
rect 134524 565082 134576 565088
rect 134536 553450 134564 565082
rect 134524 553444 134576 553450
rect 134524 553386 134576 553392
rect 133144 542428 133196 542434
rect 133144 542370 133196 542376
rect 133156 536625 133184 542370
rect 133142 536616 133198 536625
rect 133142 536551 133198 536560
rect 133880 454096 133932 454102
rect 133880 454038 133932 454044
rect 133144 439544 133196 439550
rect 133144 439486 133196 439492
rect 132500 438864 132552 438870
rect 132500 438806 132552 438812
rect 131120 391264 131172 391270
rect 131120 391206 131172 391212
rect 131304 378208 131356 378214
rect 131304 378150 131356 378156
rect 130476 378072 130528 378078
rect 130476 378014 130528 378020
rect 130488 370705 130516 378014
rect 130474 370696 130530 370705
rect 130474 370631 130530 370640
rect 130382 369064 130438 369073
rect 130382 368999 130438 369008
rect 131026 367432 131082 367441
rect 131026 367367 131082 367376
rect 130384 363656 130436 363662
rect 130384 363598 130436 363604
rect 130396 350713 130424 363598
rect 131040 357406 131068 367367
rect 131028 357400 131080 357406
rect 131080 357348 131160 357354
rect 131028 357342 131160 357348
rect 131040 357326 131160 357342
rect 131040 357277 131068 357326
rect 130382 350704 130438 350713
rect 130382 350639 130438 350648
rect 131026 350704 131082 350713
rect 131026 350639 131082 350648
rect 129002 343904 129058 343913
rect 129002 343839 129058 343848
rect 129646 343904 129702 343913
rect 129646 343839 129702 343848
rect 128452 337408 128504 337414
rect 128452 337350 128504 337356
rect 129016 331809 129044 343839
rect 130750 332480 130806 332489
rect 130750 332415 130806 332424
rect 129002 331800 129058 331809
rect 129002 331735 129058 331744
rect 129280 331560 129332 331566
rect 129280 331502 129332 331508
rect 129292 329474 129320 331502
rect 130016 331492 130068 331498
rect 130016 331434 130068 331440
rect 130028 329474 130056 331434
rect 130764 329474 130792 332415
rect 131040 331498 131068 350639
rect 131028 331492 131080 331498
rect 131028 331434 131080 331440
rect 131132 329746 131160 357326
rect 131316 345014 131344 378150
rect 133156 367810 133184 439486
rect 133788 438864 133840 438870
rect 133788 438806 133840 438812
rect 133800 438190 133828 438806
rect 133788 438184 133840 438190
rect 133788 438126 133840 438132
rect 133144 367804 133196 367810
rect 133144 367746 133196 367752
rect 133786 361720 133842 361729
rect 133786 361655 133842 361664
rect 133694 347848 133750 347857
rect 133694 347783 133750 347792
rect 131316 344986 131528 345014
rect 131132 329718 131206 329746
rect 124968 329446 125304 329474
rect 125612 329446 126040 329474
rect 126348 329446 126776 329474
rect 127084 329446 127512 329474
rect 127820 329446 128248 329474
rect 128984 329446 129320 329474
rect 129720 329446 130056 329474
rect 130456 329446 130792 329474
rect 131178 329460 131206 329718
rect 131500 329474 131528 344986
rect 132500 335368 132552 335374
rect 133708 335354 133736 347783
rect 132500 335310 132552 335316
rect 133616 335326 133736 335354
rect 132512 333305 132540 335310
rect 132498 333296 132554 333305
rect 132498 333231 132554 333240
rect 132776 331696 132828 331702
rect 132776 331638 132828 331644
rect 132788 329474 132816 331638
rect 133616 329474 133644 335326
rect 133800 331702 133828 361655
rect 133892 347070 133920 454038
rect 134536 407794 134564 553386
rect 137926 546544 137982 546553
rect 137926 546479 137982 546488
rect 137284 473408 137336 473414
rect 137284 473350 137336 473356
rect 134524 407788 134576 407794
rect 134524 407730 134576 407736
rect 134536 371550 134564 407730
rect 137296 391377 137324 473350
rect 137376 448588 137428 448594
rect 137376 448530 137428 448536
rect 137282 391368 137338 391377
rect 137282 391303 137338 391312
rect 134524 371544 134576 371550
rect 134524 371486 134576 371492
rect 135168 371544 135220 371550
rect 135168 371486 135220 371492
rect 135180 371278 135208 371486
rect 135168 371272 135220 371278
rect 135168 371214 135220 371220
rect 134984 347744 135036 347750
rect 134984 347686 135036 347692
rect 134996 347070 135024 347686
rect 133880 347064 133932 347070
rect 133880 347006 133932 347012
rect 134984 347064 135036 347070
rect 134984 347006 135036 347012
rect 134522 344312 134578 344321
rect 134522 344247 134578 344256
rect 133970 336968 134026 336977
rect 133970 336903 134026 336912
rect 133984 336054 134012 336903
rect 133972 336048 134024 336054
rect 133972 335990 134024 335996
rect 134536 332489 134564 344247
rect 134800 343664 134852 343670
rect 134800 343606 134852 343612
rect 134812 336734 134840 343606
rect 135180 340202 135208 371214
rect 137388 369073 137416 448530
rect 137374 369064 137430 369073
rect 137374 368999 137430 369008
rect 137284 343664 137336 343670
rect 137284 343606 137336 343612
rect 137190 340912 137246 340921
rect 137190 340847 137246 340856
rect 135168 340196 135220 340202
rect 135168 340138 135220 340144
rect 134800 336728 134852 336734
rect 134800 336670 134852 336676
rect 134890 335608 134946 335617
rect 134890 335543 134946 335552
rect 134522 332480 134578 332489
rect 134522 332415 134578 332424
rect 133788 331696 133840 331702
rect 133788 331638 133840 331644
rect 134246 331392 134302 331401
rect 134246 331327 134302 331336
rect 134260 329474 134288 331327
rect 134904 329474 134932 335543
rect 135168 334076 135220 334082
rect 135168 334018 135220 334024
rect 135180 331566 135208 334018
rect 135718 331800 135774 331809
rect 135718 331735 135774 331744
rect 135168 331560 135220 331566
rect 135168 331502 135220 331508
rect 135732 329474 135760 331735
rect 137008 331220 137060 331226
rect 137008 331162 137060 331168
rect 136454 330032 136510 330041
rect 136454 329967 136510 329976
rect 136468 329474 136496 329967
rect 131500 329446 131928 329474
rect 132480 329446 132816 329474
rect 133216 329446 133644 329474
rect 133952 329446 134288 329474
rect 134688 329446 134932 329474
rect 135424 329446 135760 329474
rect 136160 329446 136496 329474
rect 137020 329338 137048 331162
rect 137204 329474 137232 340847
rect 137296 331226 137324 343606
rect 137940 340921 137968 546479
rect 140780 534132 140832 534138
rect 140780 534074 140832 534080
rect 140792 532710 140820 534074
rect 140780 532704 140832 532710
rect 140780 532646 140832 532652
rect 141436 513369 141464 594798
rect 148416 581052 148468 581058
rect 148416 580994 148468 581000
rect 142804 579692 142856 579698
rect 142804 579634 142856 579640
rect 142816 574802 142844 579634
rect 142804 574796 142856 574802
rect 142804 574738 142856 574744
rect 141516 527196 141568 527202
rect 141516 527138 141568 527144
rect 141422 513360 141478 513369
rect 141422 513295 141478 513304
rect 141528 510610 141556 527138
rect 142066 513360 142122 513369
rect 142066 513295 142122 513304
rect 141516 510604 141568 510610
rect 141516 510546 141568 510552
rect 138664 492720 138716 492726
rect 138664 492662 138716 492668
rect 138676 374678 138704 492662
rect 142080 446826 142108 513295
rect 140780 446820 140832 446826
rect 140780 446762 140832 446768
rect 142068 446820 142120 446826
rect 142068 446762 142120 446768
rect 140792 446457 140820 446762
rect 140778 446448 140834 446457
rect 140778 446383 140834 446392
rect 141422 444952 141478 444961
rect 141422 444887 141478 444896
rect 140044 426488 140096 426494
rect 140044 426430 140096 426436
rect 138664 374672 138716 374678
rect 138664 374614 138716 374620
rect 139308 363044 139360 363050
rect 139308 362986 139360 362992
rect 137926 340912 137982 340921
rect 137926 340847 137982 340856
rect 139320 331498 139348 362986
rect 140056 347041 140084 426430
rect 140688 376780 140740 376786
rect 140688 376722 140740 376728
rect 140042 347032 140098 347041
rect 140042 346967 140098 346976
rect 140136 346452 140188 346458
rect 140136 346394 140188 346400
rect 139492 340196 139544 340202
rect 139492 340138 139544 340144
rect 139398 339688 139454 339697
rect 139398 339623 139454 339632
rect 139412 339590 139440 339623
rect 139400 339584 139452 339590
rect 139400 339526 139452 339532
rect 139504 335354 139532 340138
rect 140044 336048 140096 336054
rect 140044 335990 140096 335996
rect 139412 335326 139532 335354
rect 138664 331492 138716 331498
rect 138664 331434 138716 331440
rect 139308 331492 139360 331498
rect 139308 331434 139360 331440
rect 137284 331220 137336 331226
rect 137284 331162 137336 331168
rect 138676 329474 138704 331434
rect 137204 329446 137632 329474
rect 138368 329446 138704 329474
rect 139412 329474 139440 335326
rect 140056 334665 140084 335990
rect 140042 334656 140098 334665
rect 140042 334591 140098 334600
rect 140148 333266 140176 346394
rect 140136 333260 140188 333266
rect 140136 333202 140188 333208
rect 140700 329474 140728 376722
rect 141436 356794 141464 444887
rect 142816 431934 142844 574738
rect 144828 539708 144880 539714
rect 144828 539650 144880 539656
rect 142894 537024 142950 537033
rect 142894 536959 142950 536968
rect 142908 447137 142936 536959
rect 142894 447128 142950 447137
rect 142894 447063 142950 447072
rect 142988 446820 143040 446826
rect 142988 446762 143040 446768
rect 142804 431928 142856 431934
rect 142804 431870 142856 431876
rect 143000 380225 143028 446762
rect 143448 421592 143500 421598
rect 143448 421534 143500 421540
rect 143356 394732 143408 394738
rect 143356 394674 143408 394680
rect 142986 380216 143042 380225
rect 142986 380151 143042 380160
rect 143368 363633 143396 394674
rect 143354 363624 143410 363633
rect 143354 363559 143410 363568
rect 143368 363050 143396 363559
rect 143356 363044 143408 363050
rect 143356 362986 143408 362992
rect 140780 356788 140832 356794
rect 140780 356730 140832 356736
rect 141424 356788 141476 356794
rect 141424 356730 141476 356736
rect 140792 345014 140820 356730
rect 140792 344986 140912 345014
rect 139412 329446 139840 329474
rect 140576 329446 140728 329474
rect 140884 329474 140912 344986
rect 143460 340241 143488 421534
rect 143540 374128 143592 374134
rect 143540 374070 143592 374076
rect 143552 370530 143580 374070
rect 143540 370524 143592 370530
rect 143540 370466 143592 370472
rect 144736 365764 144788 365770
rect 144736 365706 144788 365712
rect 143446 340232 143502 340241
rect 143446 340167 143502 340176
rect 141882 334248 141938 334257
rect 141882 334183 141938 334192
rect 140884 329446 141312 329474
rect 117056 329310 117208 329338
rect 124324 329310 124720 329338
rect 136896 329310 137048 329338
rect 124324 329118 124352 329310
rect 141896 329202 141924 334183
rect 144550 332208 144606 332217
rect 144550 332143 144606 332152
rect 143080 331424 143132 331430
rect 143080 331366 143132 331372
rect 143092 329474 143120 331366
rect 143816 331356 143868 331362
rect 143816 331298 143868 331304
rect 143828 329474 143856 331298
rect 144564 329474 144592 332143
rect 144748 331362 144776 365706
rect 144840 331809 144868 539650
rect 148324 535560 148376 535566
rect 148324 535502 148376 535508
rect 147588 521688 147640 521694
rect 147588 521630 147640 521636
rect 147496 476060 147548 476066
rect 147496 476002 147548 476008
rect 147508 444310 147536 476002
rect 147496 444304 147548 444310
rect 147496 444246 147548 444252
rect 147496 434716 147548 434722
rect 147496 434658 147548 434664
rect 147508 433362 147536 434658
rect 147496 433356 147548 433362
rect 147496 433298 147548 433304
rect 147508 387122 147536 433298
rect 146944 387116 146996 387122
rect 146944 387058 146996 387064
rect 147496 387116 147548 387122
rect 147496 387058 147548 387064
rect 146208 369912 146260 369918
rect 146208 369854 146260 369860
rect 145564 369164 145616 369170
rect 145564 369106 145616 369112
rect 145576 332217 145604 369106
rect 146116 360256 146168 360262
rect 146116 360198 146168 360204
rect 146128 358057 146156 360198
rect 146114 358048 146170 358057
rect 146114 357983 146170 357992
rect 146220 335354 146248 369854
rect 146956 358766 146984 387058
rect 147600 363089 147628 521630
rect 148336 447098 148364 535502
rect 148428 535401 148456 580994
rect 184204 565956 184256 565962
rect 184204 565898 184256 565904
rect 162768 564460 162820 564466
rect 162768 564402 162820 564408
rect 153108 560380 153160 560386
rect 153108 560322 153160 560328
rect 151820 557592 151872 557598
rect 151820 557534 151872 557540
rect 148414 535392 148470 535401
rect 148414 535327 148470 535336
rect 148966 535392 149022 535401
rect 148966 535327 149022 535336
rect 148980 460222 149008 535327
rect 151832 488578 151860 557534
rect 151820 488572 151872 488578
rect 151820 488514 151872 488520
rect 148968 460216 149020 460222
rect 148968 460158 149020 460164
rect 148980 459610 149008 460158
rect 148416 459604 148468 459610
rect 148416 459546 148468 459552
rect 148968 459604 149020 459610
rect 148968 459546 149020 459552
rect 148324 447092 148376 447098
rect 148324 447034 148376 447040
rect 148324 444304 148376 444310
rect 148324 444246 148376 444252
rect 147586 363080 147642 363089
rect 147586 363015 147642 363024
rect 147600 360913 147628 363015
rect 147586 360904 147642 360913
rect 147586 360839 147642 360848
rect 146944 358760 146996 358766
rect 146944 358702 146996 358708
rect 147588 358760 147640 358766
rect 147588 358702 147640 358708
rect 147600 358086 147628 358702
rect 147588 358080 147640 358086
rect 147588 358022 147640 358028
rect 146128 335326 146248 335354
rect 145562 332208 145618 332217
rect 145562 332143 145618 332152
rect 144826 331800 144882 331809
rect 144826 331735 144882 331744
rect 144920 331424 144972 331430
rect 144920 331366 144972 331372
rect 144736 331356 144788 331362
rect 144736 331298 144788 331304
rect 144932 331226 144960 331366
rect 145286 331256 145342 331265
rect 144920 331220 144972 331226
rect 145286 331191 145342 331200
rect 144920 331162 144972 331168
rect 145300 329474 145328 331191
rect 146128 329474 146156 335326
rect 146760 331832 146812 331838
rect 146760 331774 146812 331780
rect 146772 329474 146800 331774
rect 147600 329474 147628 358022
rect 147678 353560 147734 353569
rect 147678 353495 147734 353504
rect 147692 349761 147720 353495
rect 148336 350849 148364 444246
rect 148428 434722 148456 459546
rect 151084 438184 151136 438190
rect 151084 438126 151136 438132
rect 148416 434716 148468 434722
rect 148416 434658 148468 434664
rect 148416 388476 148468 388482
rect 148416 388418 148468 388424
rect 147770 350840 147826 350849
rect 147770 350775 147826 350784
rect 148322 350840 148378 350849
rect 148322 350775 148378 350784
rect 147678 349752 147734 349761
rect 147678 349687 147734 349696
rect 147784 345014 147812 350775
rect 147784 344986 148272 345014
rect 148140 332648 148192 332654
rect 148140 332590 148192 332596
rect 148152 329474 148180 332590
rect 142784 329446 143120 329474
rect 143520 329446 143856 329474
rect 144256 329446 144592 329474
rect 144992 329446 145328 329474
rect 145728 329446 146156 329474
rect 146464 329446 146800 329474
rect 147200 329446 147628 329474
rect 147936 329446 148180 329474
rect 148244 329474 148272 344986
rect 148428 336025 148456 388418
rect 148506 378176 148562 378185
rect 148506 378111 148562 378120
rect 148520 371210 148548 378111
rect 148508 371204 148560 371210
rect 148508 371146 148560 371152
rect 151096 369209 151124 438126
rect 151820 369232 151872 369238
rect 151082 369200 151138 369209
rect 151820 369174 151872 369180
rect 151082 369135 151138 369144
rect 151726 360224 151782 360233
rect 151726 360159 151782 360168
rect 149426 356144 149482 356153
rect 149426 356079 149482 356088
rect 149440 350441 149468 356079
rect 149426 350432 149482 350441
rect 149426 350367 149482 350376
rect 150346 347032 150402 347041
rect 150346 346967 150402 346976
rect 150360 345014 150388 346967
rect 150268 344986 150388 345014
rect 149244 337408 149296 337414
rect 149244 337350 149296 337356
rect 148414 336016 148470 336025
rect 148414 335951 148470 335960
rect 149256 329798 149284 337350
rect 150268 331401 150296 344986
rect 150348 336864 150400 336870
rect 150348 336806 150400 336812
rect 150360 331838 150388 336806
rect 150348 331832 150400 331838
rect 150348 331774 150400 331780
rect 149702 331392 149758 331401
rect 149702 331327 149758 331336
rect 150254 331392 150310 331401
rect 150254 331327 150310 331336
rect 151176 331356 151228 331362
rect 149244 329792 149296 329798
rect 149244 329734 149296 329740
rect 149716 329474 149744 331327
rect 151176 331298 151228 331304
rect 150438 331256 150494 331265
rect 150438 331191 150494 331200
rect 150348 330608 150400 330614
rect 150348 330550 150400 330556
rect 150360 329474 150388 330550
rect 150452 329730 150480 331191
rect 150440 329724 150492 329730
rect 150440 329666 150492 329672
rect 151188 329474 151216 331298
rect 151740 329474 151768 360159
rect 151832 359009 151860 369174
rect 153120 359281 153148 560322
rect 160834 559056 160890 559065
rect 160834 558991 160890 559000
rect 156604 552152 156656 552158
rect 156604 552094 156656 552100
rect 155224 531344 155276 531350
rect 155224 531286 155276 531292
rect 155236 500954 155264 531286
rect 155224 500948 155276 500954
rect 155224 500890 155276 500896
rect 155868 498840 155920 498846
rect 155868 498782 155920 498788
rect 155222 456920 155278 456929
rect 155222 456855 155278 456864
rect 153842 451344 153898 451353
rect 153842 451279 153898 451288
rect 153856 369238 153884 451279
rect 153936 392012 153988 392018
rect 153936 391954 153988 391960
rect 153948 372638 153976 391954
rect 153936 372632 153988 372638
rect 153934 372600 153936 372609
rect 153988 372600 153990 372609
rect 153934 372535 153990 372544
rect 153844 369232 153896 369238
rect 153844 369174 153896 369180
rect 152462 359272 152518 359281
rect 152462 359207 152518 359216
rect 153106 359272 153162 359281
rect 153106 359207 153162 359216
rect 151818 359000 151874 359009
rect 151818 358935 151874 358944
rect 152476 352646 152504 359207
rect 152646 359000 152702 359009
rect 152646 358935 152702 358944
rect 152660 352646 152688 358935
rect 153120 358873 153148 359207
rect 153106 358864 153162 358873
rect 153106 358799 153162 358808
rect 153844 353320 153896 353326
rect 153844 353262 153896 353268
rect 154672 353320 154724 353326
rect 154672 353262 154724 353268
rect 152464 352640 152516 352646
rect 152464 352582 152516 352588
rect 152648 352640 152700 352646
rect 152648 352582 152700 352588
rect 152660 351966 152688 352582
rect 152648 351960 152700 351966
rect 152648 351902 152700 351908
rect 153108 351960 153160 351966
rect 153108 351902 153160 351908
rect 152464 339584 152516 339590
rect 152464 339526 152516 339532
rect 152476 334665 152504 339526
rect 152462 334656 152518 334665
rect 152462 334591 152518 334600
rect 153014 332888 153070 332897
rect 153014 332823 153070 332832
rect 152924 331356 152976 331362
rect 152924 331298 152976 331304
rect 152646 331256 152702 331265
rect 152646 331191 152702 331200
rect 152660 329474 152688 331191
rect 152936 331158 152964 331298
rect 153028 331226 153056 332823
rect 153016 331220 153068 331226
rect 153016 331162 153068 331168
rect 152924 331152 152976 331158
rect 152924 331094 152976 331100
rect 153120 329746 153148 351902
rect 153856 336054 153884 353262
rect 154684 345014 154712 353262
rect 154684 344986 154896 345014
rect 154210 338192 154266 338201
rect 154210 338127 154266 338136
rect 154224 336734 154252 338127
rect 154762 336968 154818 336977
rect 154762 336903 154818 336912
rect 154212 336728 154264 336734
rect 154212 336670 154264 336676
rect 153844 336048 153896 336054
rect 153844 335990 153896 335996
rect 154672 335776 154724 335782
rect 154672 335718 154724 335724
rect 154120 331356 154172 331362
rect 154120 331298 154172 331304
rect 148244 329446 148672 329474
rect 149408 329446 149744 329474
rect 150144 329446 150388 329474
rect 150880 329446 151216 329474
rect 151616 329446 151768 329474
rect 152352 329446 152688 329474
rect 153074 329718 153148 329746
rect 153074 329460 153102 329718
rect 154132 329474 154160 331298
rect 154684 329474 154712 335718
rect 154776 333334 154804 336903
rect 154764 333328 154816 333334
rect 154764 333270 154816 333276
rect 153824 329446 154160 329474
rect 154560 329446 154712 329474
rect 154868 329474 154896 344986
rect 155236 338065 155264 456855
rect 155314 389328 155370 389337
rect 155314 389263 155370 389272
rect 155328 353326 155356 389263
rect 155316 353320 155368 353326
rect 155316 353262 155368 353268
rect 155222 338056 155278 338065
rect 155222 337991 155278 338000
rect 155880 335782 155908 498782
rect 156616 386481 156644 552094
rect 160742 535800 160798 535809
rect 160742 535735 160798 535744
rect 159364 460964 159416 460970
rect 159364 460906 159416 460912
rect 157984 436756 158036 436762
rect 157984 436698 158036 436704
rect 156602 386472 156658 386481
rect 156602 386407 156658 386416
rect 156510 344992 156566 345001
rect 156510 344927 156566 344936
rect 156524 343738 156552 344927
rect 156512 343732 156564 343738
rect 156512 343674 156564 343680
rect 156510 340096 156566 340105
rect 156510 340031 156566 340040
rect 156524 339930 156552 340031
rect 156512 339924 156564 339930
rect 156512 339866 156564 339872
rect 155868 335776 155920 335782
rect 155868 335718 155920 335724
rect 156616 331906 156644 386407
rect 156696 385688 156748 385694
rect 156696 385630 156748 385636
rect 156708 343738 156736 385630
rect 156788 350600 156840 350606
rect 156788 350542 156840 350548
rect 156696 343732 156748 343738
rect 156696 343674 156748 343680
rect 156800 337385 156828 350542
rect 157340 343052 157392 343058
rect 157340 342994 157392 343000
rect 157246 338056 157302 338065
rect 157246 337991 157302 338000
rect 156786 337376 156842 337385
rect 156786 337311 156842 337320
rect 156604 331900 156656 331906
rect 156604 331842 156656 331848
rect 157260 331242 157288 337991
rect 157352 331537 157380 342994
rect 157338 331528 157394 331537
rect 157338 331463 157394 331472
rect 157260 331214 157380 331242
rect 156052 331152 156104 331158
rect 156052 331094 156104 331100
rect 155868 330608 155920 330614
rect 155868 330550 155920 330556
rect 155880 329866 155908 330550
rect 155868 329860 155920 329866
rect 155868 329802 155920 329808
rect 156064 329798 156092 331094
rect 156970 329896 157026 329905
rect 156970 329831 157026 329840
rect 155960 329792 156012 329798
rect 155958 329760 155960 329769
rect 156052 329792 156104 329798
rect 156012 329760 156014 329769
rect 156052 329734 156104 329740
rect 155958 329695 156014 329704
rect 156696 329724 156748 329730
rect 156696 329666 156748 329672
rect 156708 329633 156736 329666
rect 156694 329624 156750 329633
rect 156694 329559 156750 329568
rect 154868 329446 155296 329474
rect 152646 329216 152702 329225
rect 141896 329174 142048 329202
rect 152646 329151 152702 329160
rect 152660 329118 152688 329151
rect 115388 329112 115440 329118
rect 115388 329054 115440 329060
rect 124312 329112 124364 329118
rect 139308 329112 139360 329118
rect 124312 329054 124364 329060
rect 139104 329060 139308 329066
rect 139104 329054 139360 329060
rect 152648 329112 152700 329118
rect 156328 329112 156380 329118
rect 152648 329054 152700 329060
rect 156032 329060 156328 329066
rect 156032 329054 156380 329060
rect 139104 329038 139348 329054
rect 156032 329038 156368 329054
rect 156584 328902 156920 328930
rect 156696 328840 156748 328846
rect 156696 328782 156748 328788
rect 67822 308544 67878 308553
rect 67822 308479 67878 308488
rect 67836 307834 67864 308479
rect 67824 307828 67876 307834
rect 67824 307770 67876 307776
rect 67730 270736 67786 270745
rect 67730 270671 67786 270680
rect 67638 269648 67694 269657
rect 67638 269583 67694 269592
rect 67548 262948 67600 262954
rect 67548 262890 67600 262896
rect 67546 259856 67602 259865
rect 67546 259791 67602 259800
rect 67560 253230 67588 259791
rect 67548 253224 67600 253230
rect 67548 253166 67600 253172
rect 67744 250510 67772 270671
rect 68284 262948 68336 262954
rect 68284 262890 68336 262896
rect 67732 250504 67784 250510
rect 67732 250446 67784 250452
rect 67638 245712 67694 245721
rect 67638 245647 67694 245656
rect 67456 240032 67508 240038
rect 67456 239974 67508 239980
rect 67362 224904 67418 224913
rect 67362 224839 67418 224848
rect 67652 200870 67680 245647
rect 67732 240168 67784 240174
rect 67732 240110 67784 240116
rect 67744 238513 67772 240110
rect 67730 238504 67786 238513
rect 67730 238439 67786 238448
rect 68296 225622 68324 262890
rect 156708 254658 156736 328782
rect 156892 328506 156920 328902
rect 156880 328500 156932 328506
rect 156880 328442 156932 328448
rect 156880 328364 156932 328370
rect 156880 328306 156932 328312
rect 156788 328296 156840 328302
rect 156788 328238 156840 328244
rect 156800 327321 156828 328238
rect 156892 327729 156920 328306
rect 156878 327720 156934 327729
rect 156878 327655 156934 327664
rect 156984 327350 157012 329831
rect 156972 327344 157024 327350
rect 156786 327312 156842 327321
rect 156972 327286 157024 327292
rect 156786 327247 156842 327256
rect 157352 310457 157380 331214
rect 157432 331220 157484 331226
rect 157432 331162 157484 331168
rect 157444 329089 157472 331162
rect 157430 329080 157486 329089
rect 157430 329015 157486 329024
rect 157338 310448 157394 310457
rect 157338 310383 157394 310392
rect 156880 278044 156932 278050
rect 156880 277986 156932 277992
rect 156696 254652 156748 254658
rect 156696 254594 156748 254600
rect 68376 253224 68428 253230
rect 68376 253166 68428 253172
rect 68388 239601 68416 253166
rect 156788 252476 156840 252482
rect 156788 252418 156840 252424
rect 155316 242072 155368 242078
rect 80978 242040 81034 242049
rect 154670 242040 154726 242049
rect 81034 241998 81296 242026
rect 80978 241975 81034 241984
rect 69662 241904 69718 241913
rect 69662 241839 69718 241848
rect 68480 241590 68816 241618
rect 69368 241590 69612 241618
rect 68480 240174 68508 241590
rect 68468 240168 68520 240174
rect 68468 240110 68520 240116
rect 69584 240106 69612 241590
rect 69572 240100 69624 240106
rect 69572 240042 69624 240048
rect 68374 239592 68430 239601
rect 68374 239527 68430 239536
rect 68284 225616 68336 225622
rect 68284 225558 68336 225564
rect 69676 206961 69704 241839
rect 70104 241590 70348 241618
rect 69756 240032 69808 240038
rect 69756 239974 69808 239980
rect 69768 231810 69796 239974
rect 70320 239494 70348 241590
rect 70412 241590 70840 241618
rect 71576 241590 71728 241618
rect 70308 239488 70360 239494
rect 70308 239430 70360 239436
rect 69756 231804 69808 231810
rect 69756 231746 69808 231752
rect 70412 211818 70440 241590
rect 71700 238785 71728 241590
rect 71792 241590 72312 241618
rect 72712 241590 73048 241618
rect 73172 241590 73784 241618
rect 74520 241590 74580 241618
rect 71686 238776 71742 238785
rect 71686 238711 71742 238720
rect 71792 226302 71820 241590
rect 72712 240145 72740 241590
rect 72422 240136 72478 240145
rect 72698 240136 72754 240145
rect 72422 240071 72478 240080
rect 72516 240100 72568 240106
rect 71780 226296 71832 226302
rect 71780 226238 71832 226244
rect 70400 211812 70452 211818
rect 70400 211754 70452 211760
rect 69662 206952 69718 206961
rect 69662 206887 69718 206896
rect 67640 200864 67692 200870
rect 67640 200806 67692 200812
rect 72436 196625 72464 240071
rect 72698 240071 72754 240080
rect 72516 240042 72568 240048
rect 72528 202774 72556 240042
rect 73172 238746 73200 241590
rect 73802 241496 73858 241505
rect 73802 241431 73858 241440
rect 73160 238740 73212 238746
rect 73160 238682 73212 238688
rect 73816 210361 73844 241431
rect 74552 220561 74580 241590
rect 74644 241590 75256 241618
rect 75932 241590 75992 241618
rect 76728 241590 77064 241618
rect 74644 234569 74672 241590
rect 75932 240106 75960 241590
rect 75184 240100 75236 240106
rect 75184 240042 75236 240048
rect 75920 240100 75972 240106
rect 75920 240042 75972 240048
rect 75196 238678 75224 240042
rect 77036 239465 77064 241590
rect 77404 241590 77464 241618
rect 77864 241590 78200 241618
rect 78692 241590 78936 241618
rect 79672 241590 80008 241618
rect 80408 241590 80744 241618
rect 77300 240168 77352 240174
rect 77300 240110 77352 240116
rect 77022 239456 77078 239465
rect 77022 239391 77078 239400
rect 76562 238776 76618 238785
rect 76562 238711 76618 238720
rect 75184 238672 75236 238678
rect 75184 238614 75236 238620
rect 74630 234560 74686 234569
rect 74630 234495 74686 234504
rect 75196 220833 75224 238614
rect 76576 223417 76604 238711
rect 76562 223408 76618 223417
rect 76562 223343 76618 223352
rect 75182 220824 75238 220833
rect 75182 220759 75238 220768
rect 74538 220552 74594 220561
rect 74538 220487 74594 220496
rect 77312 211138 77340 240110
rect 77404 235890 77432 241590
rect 77864 240174 77892 241590
rect 77852 240168 77904 240174
rect 77852 240110 77904 240116
rect 77392 235884 77444 235890
rect 77392 235826 77444 235832
rect 77300 211132 77352 211138
rect 77300 211074 77352 211080
rect 73802 210352 73858 210361
rect 73802 210287 73858 210296
rect 72516 202768 72568 202774
rect 72516 202710 72568 202716
rect 78692 200025 78720 241590
rect 79980 223582 80008 241590
rect 80716 239290 80744 241590
rect 80704 239284 80756 239290
rect 80704 239226 80756 239232
rect 81268 224777 81296 241998
rect 154726 241998 155264 242026
rect 155316 242014 155368 242020
rect 156694 242040 156750 242049
rect 154670 241975 154726 241984
rect 81880 241590 82216 241618
rect 82616 241590 82768 241618
rect 82188 239834 82216 241590
rect 82740 240106 82768 241590
rect 83338 241466 83366 241604
rect 83752 241590 84088 241618
rect 84824 241590 85160 241618
rect 85560 241590 85620 241618
rect 83326 241460 83378 241466
rect 83326 241402 83378 241408
rect 83338 241346 83366 241402
rect 83338 241318 83412 241346
rect 82912 240168 82964 240174
rect 82912 240110 82964 240116
rect 82728 240100 82780 240106
rect 82728 240042 82780 240048
rect 82176 239828 82228 239834
rect 82176 239770 82228 239776
rect 82728 239828 82780 239834
rect 82728 239770 82780 239776
rect 81348 239284 81400 239290
rect 81348 239226 81400 239232
rect 81254 224768 81310 224777
rect 81254 224703 81310 224712
rect 79968 223576 80020 223582
rect 79968 223518 80020 223524
rect 81360 209545 81388 239226
rect 82740 218754 82768 239770
rect 82728 218748 82780 218754
rect 82728 218690 82780 218696
rect 81346 209536 81402 209545
rect 81346 209471 81402 209480
rect 82924 206825 82952 240110
rect 83384 238754 83412 241318
rect 83752 240174 83780 241590
rect 83740 240168 83792 240174
rect 83740 240110 83792 240116
rect 85132 240106 85160 241590
rect 83556 240100 83608 240106
rect 83556 240042 83608 240048
rect 85120 240100 85172 240106
rect 85120 240042 85172 240048
rect 83384 238726 83504 238754
rect 83476 208321 83504 238726
rect 83568 217326 83596 240042
rect 83646 239592 83702 239601
rect 83646 239527 83702 239536
rect 83660 229838 83688 239527
rect 83648 229832 83700 229838
rect 83648 229774 83700 229780
rect 83556 217320 83608 217326
rect 83556 217262 83608 217268
rect 83462 208312 83518 208321
rect 83462 208247 83518 208256
rect 82910 206816 82966 206825
rect 82910 206751 82966 206760
rect 78678 200016 78734 200025
rect 78678 199951 78734 199960
rect 72422 196616 72478 196625
rect 72422 196551 72478 196560
rect 85592 192545 85620 241590
rect 85684 241590 86296 241618
rect 86972 241590 87032 241618
rect 87156 241590 87768 241618
rect 88504 241590 88840 241618
rect 89240 241590 89668 241618
rect 85684 225049 85712 241590
rect 86224 240780 86276 240786
rect 86224 240722 86276 240728
rect 85670 225040 85726 225049
rect 85670 224975 85726 224984
rect 86236 220697 86264 240722
rect 86866 226128 86922 226137
rect 86866 226063 86922 226072
rect 86880 225049 86908 226063
rect 86866 225040 86922 225049
rect 86866 224975 86922 224984
rect 86222 220688 86278 220697
rect 86222 220623 86278 220632
rect 86880 200705 86908 224975
rect 86972 205630 87000 241590
rect 87156 215286 87184 241590
rect 88812 239426 88840 241590
rect 88800 239420 88852 239426
rect 88800 239362 88852 239368
rect 89536 239420 89588 239426
rect 89536 239362 89588 239368
rect 89548 222057 89576 239362
rect 89534 222048 89590 222057
rect 89534 221983 89590 221992
rect 87144 215280 87196 215286
rect 87144 215222 87196 215228
rect 86960 205624 87012 205630
rect 86960 205566 87012 205572
rect 86866 200696 86922 200705
rect 86866 200631 86922 200640
rect 89640 193866 89668 241590
rect 89732 241590 89976 241618
rect 90376 241590 90712 241618
rect 91204 241590 91448 241618
rect 91848 241590 92184 241618
rect 92492 241590 92920 241618
rect 93136 241590 93472 241618
rect 93964 241590 94208 241618
rect 89732 209030 89760 241590
rect 90376 238754 90404 241590
rect 91100 240168 91152 240174
rect 91100 240110 91152 240116
rect 89824 238726 90404 238754
rect 89824 226409 89852 238726
rect 91006 227488 91062 227497
rect 91006 227423 91062 227432
rect 91020 226409 91048 227423
rect 89810 226400 89866 226409
rect 89810 226335 89866 226344
rect 91006 226400 91062 226409
rect 91006 226335 91062 226344
rect 90916 209704 90968 209710
rect 90916 209646 90968 209652
rect 90928 209030 90956 209646
rect 89720 209024 89772 209030
rect 89720 208966 89772 208972
rect 90916 209024 90968 209030
rect 90916 208966 90968 208972
rect 89628 193860 89680 193866
rect 89628 193802 89680 193808
rect 85578 192536 85634 192545
rect 85578 192471 85634 192480
rect 90928 186969 90956 208966
rect 91020 202337 91048 226335
rect 91112 204270 91140 240110
rect 91204 233073 91232 241590
rect 91848 240174 91876 241590
rect 91836 240168 91888 240174
rect 91836 240110 91888 240116
rect 91190 233064 91246 233073
rect 91190 232999 91246 233008
rect 92492 206689 92520 241590
rect 92572 240100 92624 240106
rect 92572 240042 92624 240048
rect 92584 238241 92612 240042
rect 93136 238754 93164 241590
rect 93858 241496 93914 241505
rect 93858 241431 93914 241440
rect 92676 238726 93164 238754
rect 92570 238232 92626 238241
rect 92570 238167 92626 238176
rect 92676 233238 92704 238726
rect 93872 236026 93900 241431
rect 93860 236020 93912 236026
rect 93860 235962 93912 235968
rect 92664 233232 92716 233238
rect 92664 233174 92716 233180
rect 92676 232762 92704 233174
rect 92664 232756 92716 232762
rect 92664 232698 92716 232704
rect 93124 232756 93176 232762
rect 93124 232698 93176 232704
rect 92478 206680 92534 206689
rect 92478 206615 92534 206624
rect 91100 204264 91152 204270
rect 91100 204206 91152 204212
rect 91006 202328 91062 202337
rect 91006 202263 91062 202272
rect 93136 193186 93164 232698
rect 93964 209681 93992 241590
rect 94930 241505 94958 241604
rect 95252 241590 95680 241618
rect 95896 241590 96416 241618
rect 97152 241590 97488 241618
rect 97888 241590 97948 241618
rect 98624 241590 99144 241618
rect 99360 241590 99420 241618
rect 100096 241590 100708 241618
rect 94916 241496 94972 241505
rect 94916 241431 94972 241440
rect 94504 236020 94556 236026
rect 94504 235962 94556 235968
rect 94516 229022 94544 235962
rect 94504 229016 94556 229022
rect 94504 228958 94556 228964
rect 95252 212401 95280 241590
rect 95896 238754 95924 241590
rect 97460 239494 97488 241590
rect 97264 239488 97316 239494
rect 97264 239430 97316 239436
rect 97448 239488 97500 239494
rect 97448 239430 97500 239436
rect 95344 238726 95924 238754
rect 95344 224262 95372 238726
rect 95332 224256 95384 224262
rect 95332 224198 95384 224204
rect 97276 213926 97304 239430
rect 97264 213920 97316 213926
rect 97264 213862 97316 213868
rect 95238 212392 95294 212401
rect 95238 212327 95294 212336
rect 96526 212392 96582 212401
rect 96526 212327 96582 212336
rect 93950 209672 94006 209681
rect 93950 209607 94006 209616
rect 95146 209672 95202 209681
rect 95146 209607 95202 209616
rect 93766 206680 93822 206689
rect 93766 206615 93822 206624
rect 93124 193180 93176 193186
rect 93124 193122 93176 193128
rect 90914 186960 90970 186969
rect 90914 186895 90970 186904
rect 93780 185609 93808 206615
rect 95160 188465 95188 209607
rect 96540 191049 96568 212327
rect 97920 199889 97948 241590
rect 99116 238754 99144 241590
rect 99116 238726 99328 238754
rect 99300 215937 99328 238726
rect 99286 215928 99342 215937
rect 99286 215863 99342 215872
rect 99392 207806 99420 241590
rect 100680 217705 100708 241590
rect 100772 241590 100832 241618
rect 101568 241590 102088 241618
rect 100666 217696 100722 217705
rect 100666 217631 100722 217640
rect 100668 208276 100720 208282
rect 100668 208218 100720 208224
rect 100680 207806 100708 208218
rect 99380 207800 99432 207806
rect 99380 207742 99432 207748
rect 100668 207800 100720 207806
rect 100668 207742 100720 207748
rect 97906 199880 97962 199889
rect 97906 199815 97962 199824
rect 96526 191040 96582 191049
rect 96526 190975 96582 190984
rect 95146 188456 95202 188465
rect 95146 188391 95202 188400
rect 100680 187105 100708 207742
rect 100772 204202 100800 241590
rect 101956 239420 102008 239426
rect 101956 239362 102008 239368
rect 101968 237289 101996 239362
rect 101954 237280 102010 237289
rect 101954 237215 102010 237224
rect 101968 236065 101996 237215
rect 101402 236056 101458 236065
rect 101402 235991 101458 236000
rect 101954 236056 102010 236065
rect 101954 235991 102010 236000
rect 101416 226273 101444 235991
rect 101402 226264 101458 226273
rect 101402 226199 101458 226208
rect 102060 210905 102088 241590
rect 102244 241590 102304 241618
rect 102704 241590 103040 241618
rect 103776 241590 104112 241618
rect 104512 241590 104848 241618
rect 105248 241590 105584 241618
rect 102244 237289 102272 241590
rect 102704 239426 102732 241590
rect 103612 240236 103664 240242
rect 103612 240178 103664 240184
rect 102692 239420 102744 239426
rect 102692 239362 102744 239368
rect 102230 237280 102286 237289
rect 102230 237215 102286 237224
rect 103624 234433 103652 240178
rect 104084 239222 104112 241590
rect 104820 240242 104848 241590
rect 104808 240236 104860 240242
rect 104808 240178 104860 240184
rect 105556 239290 105584 241590
rect 105648 241590 105984 241618
rect 106292 241590 106720 241618
rect 107456 241590 107608 241618
rect 105544 239284 105596 239290
rect 105544 239226 105596 239232
rect 104072 239216 104124 239222
rect 104072 239158 104124 239164
rect 104808 239216 104860 239222
rect 104808 239158 104860 239164
rect 103610 234424 103666 234433
rect 103610 234359 103666 234368
rect 104164 225616 104216 225622
rect 104164 225558 104216 225564
rect 102046 210896 102102 210905
rect 102046 210831 102102 210840
rect 104176 209778 104204 225558
rect 104164 209772 104216 209778
rect 104164 209714 104216 209720
rect 100760 204196 100812 204202
rect 100760 204138 100812 204144
rect 104820 195265 104848 239158
rect 105648 238754 105676 241590
rect 106188 239284 106240 239290
rect 106188 239226 106240 239232
rect 104912 238726 105676 238754
rect 104912 220794 104940 238726
rect 104900 220788 104952 220794
rect 104900 220730 104952 220736
rect 106200 218822 106228 239226
rect 106292 222086 106320 241590
rect 106280 222080 106332 222086
rect 106280 222022 106332 222028
rect 106188 218816 106240 218822
rect 106188 218758 106240 218764
rect 104806 195256 104862 195265
rect 104806 195191 104862 195200
rect 107580 194449 107608 241590
rect 107764 241590 108192 241618
rect 108592 241590 108928 241618
rect 109664 241590 110276 241618
rect 110400 241590 110736 241618
rect 111136 241590 111748 241618
rect 107660 240168 107712 240174
rect 107660 240110 107712 240116
rect 107672 216646 107700 240110
rect 107764 235249 107792 241590
rect 108592 240174 108620 241590
rect 108580 240168 108632 240174
rect 108580 240110 108632 240116
rect 110248 238754 110276 241590
rect 110708 239873 110736 241590
rect 110694 239864 110750 239873
rect 110694 239799 110750 239808
rect 110248 238726 110368 238754
rect 107750 235240 107806 235249
rect 107750 235175 107806 235184
rect 110340 230353 110368 238726
rect 110326 230344 110382 230353
rect 110326 230279 110382 230288
rect 111720 224942 111748 241590
rect 111812 241590 111872 241618
rect 112608 241590 113128 241618
rect 113344 241590 113680 241618
rect 114080 241590 114508 241618
rect 111708 224936 111760 224942
rect 111708 224878 111760 224884
rect 107660 216640 107712 216646
rect 107660 216582 107712 216588
rect 111812 215121 111840 241590
rect 111890 239456 111946 239465
rect 111890 239391 111946 239400
rect 111904 233918 111932 239391
rect 111892 233912 111944 233918
rect 111892 233854 111944 233860
rect 111798 215112 111854 215121
rect 111798 215047 111854 215056
rect 112994 215112 113050 215121
rect 112994 215047 113050 215056
rect 113008 196654 113036 215047
rect 113100 205057 113128 241590
rect 113652 240038 113680 241590
rect 113640 240032 113692 240038
rect 113640 239974 113692 239980
rect 114480 206990 114508 241590
rect 114664 241590 114816 241618
rect 115552 241590 115888 241618
rect 116288 241590 116624 241618
rect 117024 241590 117268 241618
rect 117760 241590 117912 241618
rect 114664 235890 114692 241590
rect 115204 240168 115256 240174
rect 115204 240110 115256 240116
rect 114652 235884 114704 235890
rect 114652 235826 114704 235832
rect 115216 226001 115244 240110
rect 115860 239465 115888 241590
rect 115846 239456 115902 239465
rect 115846 239391 115902 239400
rect 116596 239358 116624 241590
rect 116584 239352 116636 239358
rect 116584 239294 116636 239300
rect 117136 239352 117188 239358
rect 117136 239294 117188 239300
rect 115202 225992 115258 226001
rect 115202 225927 115258 225936
rect 117148 213761 117176 239294
rect 117134 213752 117190 213761
rect 117134 213687 117190 213696
rect 114468 206984 114520 206990
rect 114468 206926 114520 206932
rect 113086 205048 113142 205057
rect 113086 204983 113142 204992
rect 117240 200841 117268 241590
rect 117884 240106 117912 241590
rect 117976 241590 118312 241618
rect 119048 241590 119384 241618
rect 117872 240100 117924 240106
rect 117872 240042 117924 240048
rect 117976 238754 118004 241590
rect 119356 240106 119384 241590
rect 119448 241590 119784 241618
rect 120520 241590 120856 241618
rect 118608 240100 118660 240106
rect 118608 240042 118660 240048
rect 119344 240100 119396 240106
rect 119344 240042 119396 240048
rect 118516 240032 118568 240038
rect 118516 239974 118568 239980
rect 117332 238726 118004 238754
rect 117332 229090 117360 238726
rect 118528 238678 118556 239974
rect 118516 238672 118568 238678
rect 118516 238614 118568 238620
rect 117320 229084 117372 229090
rect 117320 229026 117372 229032
rect 117226 200832 117282 200841
rect 117226 200767 117282 200776
rect 118620 197334 118648 240042
rect 119448 238754 119476 241590
rect 119988 240100 120040 240106
rect 119988 240042 120040 240048
rect 118712 238726 119476 238754
rect 118712 213858 118740 238726
rect 120000 219065 120028 240042
rect 120828 239358 120856 241590
rect 120920 241590 121256 241618
rect 121992 241590 122328 241618
rect 122728 241590 122788 241618
rect 123464 241590 124076 241618
rect 124200 241590 124260 241618
rect 120816 239352 120868 239358
rect 120816 239294 120868 239300
rect 120920 238754 120948 241590
rect 122300 239494 122328 241590
rect 122288 239488 122340 239494
rect 122288 239430 122340 239436
rect 121368 239352 121420 239358
rect 121368 239294 121420 239300
rect 120092 238726 120948 238754
rect 119986 219056 120042 219065
rect 119986 218991 120042 219000
rect 118700 213852 118752 213858
rect 118700 213794 118752 213800
rect 120092 198626 120120 238726
rect 121380 202881 121408 239294
rect 121366 202872 121422 202881
rect 121366 202807 121422 202816
rect 120080 198620 120132 198626
rect 120080 198562 120132 198568
rect 122760 198121 122788 241590
rect 124048 238754 124076 241590
rect 124048 238726 124168 238754
rect 124140 212498 124168 238726
rect 124232 222902 124260 241590
rect 124324 241590 124936 241618
rect 125612 241590 125672 241618
rect 126408 241590 126928 241618
rect 124324 231742 124352 241590
rect 125612 237386 125640 241590
rect 125600 237380 125652 237386
rect 125600 237322 125652 237328
rect 124312 231736 124364 231742
rect 124312 231678 124364 231684
rect 124220 222896 124272 222902
rect 124220 222838 124272 222844
rect 124128 212492 124180 212498
rect 124128 212434 124180 212440
rect 126900 200802 126928 241590
rect 126992 241590 127144 241618
rect 127268 241590 127880 241618
rect 128616 241590 128676 241618
rect 126992 218006 127020 241590
rect 127268 220114 127296 241590
rect 128648 240106 128676 241590
rect 128740 241590 129352 241618
rect 129844 241590 130088 241618
rect 130824 241590 131068 241618
rect 131560 241590 131896 241618
rect 128636 240100 128688 240106
rect 128636 240042 128688 240048
rect 128740 239986 128768 241590
rect 128820 240780 128872 240786
rect 128820 240722 128872 240728
rect 128372 239958 128768 239986
rect 127256 220108 127308 220114
rect 127256 220050 127308 220056
rect 128372 219201 128400 239958
rect 128832 238754 128860 240722
rect 129648 240100 129700 240106
rect 129648 240042 129700 240048
rect 128740 238726 128860 238754
rect 128740 234598 128768 238726
rect 128728 234592 128780 234598
rect 128728 234534 128780 234540
rect 128358 219192 128414 219201
rect 128358 219127 128414 219136
rect 126980 218000 127032 218006
rect 126980 217942 127032 217948
rect 129660 205601 129688 240042
rect 129844 234433 129872 241590
rect 130106 240952 130162 240961
rect 130106 240887 130162 240896
rect 130120 235958 130148 240887
rect 130108 235952 130160 235958
rect 130108 235894 130160 235900
rect 129830 234424 129886 234433
rect 129830 234359 129886 234368
rect 131040 211041 131068 241590
rect 131868 240106 131896 241590
rect 131960 241590 132296 241618
rect 133032 241590 133368 241618
rect 131856 240100 131908 240106
rect 131856 240042 131908 240048
rect 131960 239290 131988 241590
rect 133340 240106 133368 241590
rect 133708 241590 133768 241618
rect 134504 241590 134932 241618
rect 135240 241590 135392 241618
rect 132408 240100 132460 240106
rect 132408 240042 132460 240048
rect 133328 240100 133380 240106
rect 133328 240042 133380 240048
rect 131212 239284 131264 239290
rect 131212 239226 131264 239232
rect 131948 239284 132000 239290
rect 131948 239226 132000 239232
rect 131224 235278 131252 239226
rect 131212 235272 131264 235278
rect 131212 235214 131264 235220
rect 132420 216578 132448 240042
rect 133144 233980 133196 233986
rect 133144 233922 133196 233928
rect 133156 223553 133184 233922
rect 133142 223544 133198 223553
rect 133142 223479 133198 223488
rect 133708 223281 133736 241590
rect 133788 240100 133840 240106
rect 133788 240042 133840 240048
rect 133694 223272 133750 223281
rect 133694 223207 133750 223216
rect 133144 218816 133196 218822
rect 133144 218758 133196 218764
rect 132408 216572 132460 216578
rect 132408 216514 132460 216520
rect 131026 211032 131082 211041
rect 131026 210967 131082 210976
rect 133156 208049 133184 218758
rect 133142 208040 133198 208049
rect 133142 207975 133198 207984
rect 133800 206922 133828 240042
rect 134904 238754 134932 241590
rect 135364 240106 135392 241590
rect 135456 241590 135976 241618
rect 136652 241590 136712 241618
rect 137296 241590 137448 241618
rect 138184 241590 138520 241618
rect 135352 240100 135404 240106
rect 135352 240042 135404 240048
rect 134904 238726 135208 238754
rect 135180 224369 135208 238726
rect 135456 232937 135484 241590
rect 136548 240100 136600 240106
rect 136548 240042 136600 240048
rect 135442 232928 135498 232937
rect 135442 232863 135498 232872
rect 136560 228857 136588 240042
rect 136546 228848 136602 228857
rect 136546 228783 136602 228792
rect 135166 224360 135222 224369
rect 135166 224295 135222 224304
rect 136652 218822 136680 241590
rect 137296 237153 137324 241590
rect 138492 240106 138520 241590
rect 138584 241590 138920 241618
rect 139412 241590 139656 241618
rect 140056 241590 140392 241618
rect 140792 241590 141128 241618
rect 141864 241590 142108 241618
rect 142600 241590 142936 241618
rect 138480 240100 138532 240106
rect 138480 240042 138532 240048
rect 138584 239290 138612 241590
rect 139308 240100 139360 240106
rect 139308 240042 139360 240048
rect 138020 239284 138072 239290
rect 138020 239226 138072 239232
rect 138572 239284 138624 239290
rect 138572 239226 138624 239232
rect 137282 237144 137338 237153
rect 137282 237079 137338 237088
rect 136640 218816 136692 218822
rect 136640 218758 136692 218764
rect 133788 206916 133840 206922
rect 133788 206858 133840 206864
rect 129646 205592 129702 205601
rect 129646 205527 129702 205536
rect 137296 204950 137324 237079
rect 137928 229764 137980 229770
rect 137928 229706 137980 229712
rect 137940 227730 137968 229706
rect 137928 227724 137980 227730
rect 137928 227666 137980 227672
rect 138032 227633 138060 239226
rect 139320 230382 139348 240042
rect 139308 230376 139360 230382
rect 139308 230318 139360 230324
rect 138018 227624 138074 227633
rect 138018 227559 138074 227568
rect 138032 221921 138060 227559
rect 139412 226234 139440 241590
rect 140056 238754 140084 241590
rect 139504 238726 140084 238754
rect 139504 227361 139532 238726
rect 140792 235634 140820 241590
rect 140792 235606 140912 235634
rect 140778 235240 140834 235249
rect 140778 235175 140834 235184
rect 140792 234297 140820 235175
rect 140778 234288 140834 234297
rect 140778 234223 140834 234232
rect 139584 233912 139636 233918
rect 139584 233854 139636 233860
rect 139596 231713 139624 233854
rect 140884 232626 140912 235606
rect 140872 232620 140924 232626
rect 140872 232562 140924 232568
rect 139582 231704 139638 231713
rect 139582 231639 139638 231648
rect 141424 229832 141476 229838
rect 141424 229774 141476 229780
rect 139490 227352 139546 227361
rect 139490 227287 139546 227296
rect 139400 226228 139452 226234
rect 139400 226170 139452 226176
rect 138018 221912 138074 221921
rect 138018 221847 138074 221856
rect 141436 213625 141464 229774
rect 141422 213616 141478 213625
rect 141422 213551 141478 213560
rect 137284 204944 137336 204950
rect 137284 204886 137336 204892
rect 126888 200796 126940 200802
rect 126888 200738 126940 200744
rect 122746 198112 122802 198121
rect 122746 198047 122802 198056
rect 118608 197328 118660 197334
rect 118608 197270 118660 197276
rect 112996 196648 113048 196654
rect 112996 196590 113048 196596
rect 133144 195288 133196 195294
rect 133144 195230 133196 195236
rect 107566 194440 107622 194449
rect 107566 194375 107622 194384
rect 129002 193896 129058 193905
rect 129002 193831 129058 193840
rect 110328 189100 110380 189106
rect 110328 189042 110380 189048
rect 100666 187096 100722 187105
rect 100666 187031 100722 187040
rect 93766 185600 93822 185609
rect 93766 185535 93822 185544
rect 100668 184952 100720 184958
rect 100668 184894 100720 184900
rect 98458 180840 98514 180849
rect 98458 180775 98514 180784
rect 97446 179480 97502 179489
rect 97446 179415 97502 179424
rect 97460 176905 97488 179415
rect 98472 177585 98500 180775
rect 98458 177576 98514 177585
rect 98458 177511 98514 177520
rect 97446 176896 97502 176905
rect 97446 176831 97502 176840
rect 100680 176769 100708 184894
rect 101954 183696 102010 183705
rect 101954 183631 102010 183640
rect 101968 177585 101996 183631
rect 108948 183592 109000 183598
rect 108948 183534 109000 183540
rect 103334 182200 103390 182209
rect 103334 182135 103390 182144
rect 102048 178016 102100 178022
rect 102048 177958 102100 177964
rect 101954 177576 102010 177585
rect 101954 177511 102010 177520
rect 102060 176769 102088 177958
rect 103348 176769 103376 182135
rect 105726 180976 105782 180985
rect 105726 180911 105782 180920
rect 105740 177585 105768 180911
rect 107014 179616 107070 179625
rect 107014 179551 107070 179560
rect 105726 177576 105782 177585
rect 105726 177511 105782 177520
rect 107028 177041 107056 179551
rect 108960 177585 108988 183534
rect 110340 177585 110368 189042
rect 114468 185020 114520 185026
rect 114468 184962 114520 184968
rect 112258 182336 112314 182345
rect 112258 182271 112314 182280
rect 108946 177576 109002 177585
rect 108946 177511 109002 177520
rect 110326 177576 110382 177585
rect 110326 177511 110382 177520
rect 112272 177449 112300 182271
rect 114480 177585 114508 184962
rect 117228 183660 117280 183666
rect 117228 183602 117280 183608
rect 115848 180872 115900 180878
rect 115848 180814 115900 180820
rect 115860 177585 115888 180814
rect 117240 177585 117268 183602
rect 123484 182232 123536 182238
rect 123484 182174 123536 182180
rect 119804 179512 119856 179518
rect 119804 179454 119856 179460
rect 114466 177576 114522 177585
rect 114466 177511 114522 177520
rect 115846 177576 115902 177585
rect 115846 177511 115902 177520
rect 117226 177576 117282 177585
rect 117226 177511 117282 177520
rect 112258 177440 112314 177449
rect 112258 177375 112314 177384
rect 119816 177041 119844 179454
rect 123496 177585 123524 182174
rect 128176 179444 128228 179450
rect 128176 179386 128228 179392
rect 125048 178084 125100 178090
rect 125048 178026 125100 178032
rect 123482 177576 123538 177585
rect 123482 177511 123538 177520
rect 107014 177032 107070 177041
rect 107014 176967 107070 176976
rect 119802 177032 119858 177041
rect 119802 176967 119858 176976
rect 125060 176769 125088 178026
rect 128188 176769 128216 179386
rect 100666 176760 100722 176769
rect 100666 176695 100722 176704
rect 102046 176760 102102 176769
rect 102046 176695 102102 176704
rect 103334 176760 103390 176769
rect 103334 176695 103390 176704
rect 125046 176760 125102 176769
rect 125046 176695 125102 176704
rect 128174 176760 128230 176769
rect 128174 176695 128230 176704
rect 129016 175982 129044 193831
rect 129096 187740 129148 187746
rect 129096 187682 129148 187688
rect 129108 178022 129136 187682
rect 133156 178673 133184 195230
rect 142080 194585 142108 241590
rect 142908 240106 142936 241590
rect 143000 241590 143152 241618
rect 143644 241590 143888 241618
rect 144288 241590 144624 241618
rect 145360 241590 145696 241618
rect 146096 241590 146248 241618
rect 146832 241590 147444 241618
rect 147568 241590 147628 241618
rect 148304 241590 148916 241618
rect 149040 241590 149100 241618
rect 149776 241590 150112 241618
rect 142896 240100 142948 240106
rect 142896 240042 142948 240048
rect 143000 240038 143028 241590
rect 143356 240100 143408 240106
rect 143356 240042 143408 240048
rect 142252 240032 142304 240038
rect 142252 239974 142304 239980
rect 142988 240032 143040 240038
rect 142988 239974 143040 239980
rect 142264 235929 142292 239974
rect 142250 235920 142306 235929
rect 142250 235855 142306 235864
rect 143368 230450 143396 240042
rect 143540 239352 143592 239358
rect 143540 239294 143592 239300
rect 143552 232558 143580 239294
rect 143644 233238 143672 241590
rect 144288 239358 144316 241590
rect 145668 240106 145696 241590
rect 145656 240100 145708 240106
rect 145656 240042 145708 240048
rect 146116 240100 146168 240106
rect 146116 240042 146168 240048
rect 144276 239352 144328 239358
rect 144276 239294 144328 239300
rect 143632 233232 143684 233238
rect 143632 233174 143684 233180
rect 143540 232552 143592 232558
rect 143460 232500 143540 232506
rect 143460 232494 143592 232500
rect 143460 232478 143580 232494
rect 143356 230444 143408 230450
rect 143356 230386 143408 230392
rect 143460 219434 143488 232478
rect 146128 227633 146156 240042
rect 146114 227624 146170 227633
rect 146114 227559 146170 227568
rect 146220 223553 146248 241590
rect 147416 238754 147444 241590
rect 147416 238726 147536 238754
rect 147508 231577 147536 238726
rect 147494 231568 147550 231577
rect 147494 231503 147550 231512
rect 146206 223544 146262 223553
rect 146206 223479 146262 223488
rect 143368 219406 143488 219434
rect 142804 218748 142856 218754
rect 142804 218690 142856 218696
rect 142816 205562 142844 218690
rect 143368 217841 143396 219406
rect 143446 219056 143502 219065
rect 143446 218991 143502 219000
rect 143460 218074 143488 218991
rect 143448 218068 143500 218074
rect 143448 218010 143500 218016
rect 143354 217832 143410 217841
rect 143354 217767 143410 217776
rect 142804 205556 142856 205562
rect 142804 205498 142856 205504
rect 147600 199510 147628 241590
rect 148888 238754 148916 241590
rect 148888 238726 149008 238754
rect 148980 204241 149008 238726
rect 149072 237318 149100 241590
rect 150084 241233 150112 241590
rect 150452 241590 150512 241618
rect 150636 241590 151248 241618
rect 151984 241590 152044 241618
rect 150070 241224 150126 241233
rect 150070 241159 150126 241168
rect 149060 237312 149112 237318
rect 149060 237254 149112 237260
rect 150452 234598 150480 241590
rect 150636 235657 150664 241590
rect 151726 241224 151782 241233
rect 151726 241159 151782 241168
rect 150622 235648 150678 235657
rect 150622 235583 150678 235592
rect 150440 234592 150492 234598
rect 150440 234534 150492 234540
rect 148966 204232 149022 204241
rect 148966 204167 149022 204176
rect 151740 202201 151768 241159
rect 152016 240145 152044 241590
rect 152108 241590 152720 241618
rect 153456 241590 153516 241618
rect 152002 240136 152058 240145
rect 152002 240071 152058 240080
rect 152108 234530 152136 241590
rect 153106 240136 153162 240145
rect 153488 240106 153516 241590
rect 153580 241590 154192 241618
rect 153106 240071 153162 240080
rect 153476 240100 153528 240106
rect 152738 237416 152794 237425
rect 152738 237351 152794 237360
rect 152752 235890 152780 237351
rect 152464 235884 152516 235890
rect 152464 235826 152516 235832
rect 152740 235884 152792 235890
rect 152740 235826 152792 235832
rect 152370 235784 152426 235793
rect 152370 235719 152372 235728
rect 152424 235719 152426 235728
rect 152372 235690 152424 235696
rect 152096 234524 152148 234530
rect 152096 234466 152148 234472
rect 152476 219065 152504 235826
rect 152922 235784 152978 235793
rect 152922 235719 152978 235728
rect 152936 233986 152964 235719
rect 152924 233980 152976 233986
rect 152924 233922 152976 233928
rect 152462 219056 152518 219065
rect 152462 218991 152518 219000
rect 153120 204921 153148 240071
rect 153476 240042 153528 240048
rect 153382 238640 153438 238649
rect 153382 238575 153438 238584
rect 153396 235929 153424 238575
rect 153580 235929 153608 241590
rect 154488 240100 154540 240106
rect 154488 240042 154540 240048
rect 153382 235920 153438 235929
rect 153382 235855 153438 235864
rect 153566 235920 153622 235929
rect 153566 235855 153622 235864
rect 153106 204912 153162 204921
rect 153106 204847 153162 204856
rect 151726 202192 151782 202201
rect 151726 202127 151782 202136
rect 147588 199504 147640 199510
rect 147588 199446 147640 199452
rect 154500 195401 154528 240042
rect 155236 240009 155264 241998
rect 155222 240000 155278 240009
rect 155222 239935 155278 239944
rect 155224 233912 155276 233918
rect 155224 233854 155276 233860
rect 155236 223417 155264 233854
rect 155328 231713 155356 242014
rect 156694 241975 156750 241984
rect 155664 241590 155724 241618
rect 155500 240440 155552 240446
rect 155500 240382 155552 240388
rect 155512 234569 155540 240382
rect 155696 240145 155724 241590
rect 156386 241398 156414 241604
rect 156374 241392 156426 241398
rect 156374 241334 156426 241340
rect 156708 240446 156736 241975
rect 156696 240440 156748 240446
rect 156696 240382 156748 240388
rect 155682 240136 155738 240145
rect 155682 240071 155738 240080
rect 155774 240000 155830 240009
rect 155774 239935 155830 239944
rect 155498 234560 155554 234569
rect 155498 234495 155554 234504
rect 155682 234560 155738 234569
rect 155682 234495 155684 234504
rect 155736 234495 155738 234504
rect 155684 234466 155736 234472
rect 155788 231713 155816 239935
rect 155960 235748 156012 235754
rect 155960 235690 156012 235696
rect 155972 235249 156000 235690
rect 155958 235240 156014 235249
rect 155958 235175 156014 235184
rect 155868 233164 155920 233170
rect 155868 233106 155920 233112
rect 155880 232626 155908 233106
rect 156604 232756 156656 232762
rect 156604 232698 156656 232704
rect 155868 232620 155920 232626
rect 155868 232562 155920 232568
rect 155314 231704 155370 231713
rect 155314 231639 155370 231648
rect 155774 231704 155830 231713
rect 155774 231639 155830 231648
rect 155222 223408 155278 223417
rect 155222 223343 155278 223352
rect 154486 195392 154542 195401
rect 154486 195327 154542 195336
rect 142066 194576 142122 194585
rect 142066 194511 142122 194520
rect 139400 193928 139452 193934
rect 139400 193870 139452 193876
rect 139412 193118 139440 193870
rect 139400 193112 139452 193118
rect 139400 193054 139452 193060
rect 155880 189786 155908 232562
rect 156616 193905 156644 232698
rect 156800 198626 156828 252418
rect 156892 233238 156920 277986
rect 157996 255241 158024 436698
rect 158074 385656 158130 385665
rect 158074 385591 158130 385600
rect 158088 291825 158116 385591
rect 159376 374649 159404 460906
rect 160756 420918 160784 535735
rect 160848 527134 160876 558991
rect 160836 527128 160888 527134
rect 160836 527070 160888 527076
rect 162216 436144 162268 436150
rect 162216 436086 162268 436092
rect 160744 420912 160796 420918
rect 160744 420854 160796 420860
rect 160744 393984 160796 393990
rect 160744 393926 160796 393932
rect 159454 389464 159510 389473
rect 159454 389399 159510 389408
rect 159362 374640 159418 374649
rect 159362 374575 159418 374584
rect 158720 373312 158772 373318
rect 158720 373254 158772 373260
rect 158260 332648 158312 332654
rect 158260 332590 158312 332596
rect 158272 325446 158300 332590
rect 158260 325440 158312 325446
rect 158260 325382 158312 325388
rect 158166 324456 158222 324465
rect 158732 324442 158760 373254
rect 159362 369200 159418 369209
rect 159362 369135 159418 369144
rect 158812 339924 158864 339930
rect 158812 339866 158864 339872
rect 158824 339697 158852 339866
rect 158810 339688 158866 339697
rect 158810 339623 158866 339632
rect 159376 338065 159404 369135
rect 159468 342145 159496 389399
rect 160756 380186 160784 393926
rect 160744 380180 160796 380186
rect 160744 380122 160796 380128
rect 160836 378820 160888 378826
rect 160836 378762 160888 378768
rect 160098 378720 160154 378729
rect 160098 378655 160154 378664
rect 159454 342136 159510 342145
rect 159454 342071 159510 342080
rect 159362 338056 159418 338065
rect 159362 337991 159418 338000
rect 158810 336016 158866 336025
rect 158810 335951 158866 335960
rect 158824 324850 158852 335951
rect 158904 335776 158956 335782
rect 158904 335718 158956 335724
rect 158916 335481 158944 335718
rect 158902 335472 158958 335481
rect 158902 335407 158958 335416
rect 158904 334076 158956 334082
rect 158904 334018 158956 334024
rect 158916 329186 158944 334018
rect 158996 331356 159048 331362
rect 158996 331298 159048 331304
rect 158904 329180 158956 329186
rect 158904 329122 158956 329128
rect 158904 327888 158956 327894
rect 158904 327830 158956 327836
rect 158916 327593 158944 327830
rect 158902 327584 158958 327593
rect 158902 327519 158958 327528
rect 158902 326496 158958 326505
rect 158902 326431 158958 326440
rect 158916 325718 158944 326431
rect 159008 326369 159036 331298
rect 159456 329792 159508 329798
rect 159456 329734 159508 329740
rect 158994 326360 159050 326369
rect 158994 326295 159050 326304
rect 158904 325712 158956 325718
rect 158904 325654 158956 325660
rect 158824 324822 159128 324850
rect 158732 324414 158852 324442
rect 158166 324391 158222 324400
rect 158180 309913 158208 324391
rect 158718 324320 158774 324329
rect 158718 324255 158774 324264
rect 158732 323066 158760 324255
rect 158720 323060 158772 323066
rect 158720 323002 158772 323008
rect 158718 322144 158774 322153
rect 158718 322079 158774 322088
rect 158732 321638 158760 322079
rect 158720 321632 158772 321638
rect 158720 321574 158772 321580
rect 158718 321056 158774 321065
rect 158718 320991 158774 321000
rect 158732 320210 158760 320991
rect 158720 320204 158772 320210
rect 158720 320146 158772 320152
rect 158720 319456 158772 319462
rect 158720 319398 158772 319404
rect 158732 318889 158760 319398
rect 158718 318880 158774 318889
rect 158718 318815 158774 318824
rect 158718 317792 158774 317801
rect 158718 317727 158774 317736
rect 158732 317490 158760 317727
rect 158720 317484 158772 317490
rect 158720 317426 158772 317432
rect 158824 317422 158852 324414
rect 158904 324216 158956 324222
rect 158904 324158 158956 324164
rect 158916 323241 158944 324158
rect 158902 323232 158958 323241
rect 158902 323167 158958 323176
rect 158812 317416 158864 317422
rect 158812 317358 158864 317364
rect 158824 316713 158852 317358
rect 158810 316704 158866 316713
rect 158810 316639 158866 316648
rect 159100 316034 159128 324822
rect 159362 319424 159418 319433
rect 159362 319359 159418 319368
rect 158824 316006 159128 316034
rect 158718 315616 158774 315625
rect 158718 315551 158774 315560
rect 158732 314770 158760 315551
rect 158720 314764 158772 314770
rect 158720 314706 158772 314712
rect 158720 314628 158772 314634
rect 158720 314570 158772 314576
rect 158732 314537 158760 314570
rect 158718 314528 158774 314537
rect 158718 314463 158774 314472
rect 158718 313440 158774 313449
rect 158718 313375 158774 313384
rect 158732 313342 158760 313375
rect 158720 313336 158772 313342
rect 158720 313278 158772 313284
rect 158166 309904 158222 309913
rect 158166 309839 158222 309848
rect 158718 306912 158774 306921
rect 158718 306847 158774 306856
rect 158732 306406 158760 306847
rect 158720 306400 158772 306406
rect 158720 306342 158772 306348
rect 158824 306374 158852 316006
rect 158824 306346 158944 306374
rect 158810 305824 158866 305833
rect 158810 305759 158866 305768
rect 158824 305046 158852 305759
rect 158812 305040 158864 305046
rect 158812 304982 158864 304988
rect 158718 304736 158774 304745
rect 158718 304671 158774 304680
rect 158260 301504 158312 301510
rect 158260 301446 158312 301452
rect 158074 291816 158130 291825
rect 158130 291774 158208 291802
rect 158074 291751 158130 291760
rect 158074 287736 158130 287745
rect 158074 287671 158130 287680
rect 157982 255232 158038 255241
rect 157982 255167 158038 255176
rect 157984 243568 158036 243574
rect 157984 243510 158036 243516
rect 156972 241528 157024 241534
rect 156972 241470 157024 241476
rect 156880 233232 156932 233238
rect 156880 233174 156932 233180
rect 156984 231810 157012 241470
rect 157338 233064 157394 233073
rect 157338 232999 157394 233008
rect 157352 232558 157380 232999
rect 157340 232552 157392 232558
rect 157340 232494 157392 232500
rect 156972 231804 157024 231810
rect 156972 231746 157024 231752
rect 157338 224768 157394 224777
rect 157338 224703 157394 224712
rect 157352 224262 157380 224703
rect 157340 224256 157392 224262
rect 157340 224198 157392 224204
rect 157996 199889 158024 243510
rect 158088 226302 158116 287671
rect 158180 242185 158208 291774
rect 158272 268025 158300 301446
rect 158732 298790 158760 304671
rect 158916 300121 158944 306346
rect 158902 300112 158958 300121
rect 158902 300047 158958 300056
rect 158720 298784 158772 298790
rect 158720 298726 158772 298732
rect 158720 297424 158772 297430
rect 158720 297366 158772 297372
rect 158732 297129 158760 297366
rect 158718 297120 158774 297129
rect 158718 297055 158774 297064
rect 158720 295316 158772 295322
rect 158720 295258 158772 295264
rect 158732 294953 158760 295258
rect 158718 294944 158774 294953
rect 158718 294879 158774 294888
rect 158810 293856 158866 293865
rect 158810 293791 158866 293800
rect 158718 293040 158774 293049
rect 158718 292975 158774 292984
rect 158732 292670 158760 292975
rect 158720 292664 158772 292670
rect 158720 292606 158772 292612
rect 158824 292602 158852 293791
rect 158812 292596 158864 292602
rect 158812 292538 158864 292544
rect 158718 291952 158774 291961
rect 158718 291887 158774 291896
rect 158732 291310 158760 291887
rect 158720 291304 158772 291310
rect 158720 291246 158772 291252
rect 158718 290864 158774 290873
rect 158718 290799 158774 290808
rect 158732 289882 158760 290799
rect 159272 290216 159324 290222
rect 159272 290158 159324 290164
rect 158720 289876 158772 289882
rect 158720 289818 158772 289824
rect 158810 289776 158866 289785
rect 158810 289711 158866 289720
rect 158824 288454 158852 289711
rect 159284 288697 159312 290158
rect 159270 288688 159326 288697
rect 159270 288623 159326 288632
rect 158812 288448 158864 288454
rect 158812 288390 158864 288396
rect 158718 287600 158774 287609
rect 158718 287535 158774 287544
rect 158732 287094 158760 287535
rect 158720 287088 158772 287094
rect 158720 287030 158772 287036
rect 158812 287020 158864 287026
rect 158812 286962 158864 286968
rect 158824 286521 158852 286962
rect 158810 286512 158866 286521
rect 158810 286447 158866 286456
rect 158720 286340 158772 286346
rect 158720 286282 158772 286288
rect 158732 285433 158760 286282
rect 158718 285424 158774 285433
rect 158718 285359 158774 285368
rect 158720 284368 158772 284374
rect 158718 284336 158720 284345
rect 158772 284336 158774 284345
rect 158718 284271 158774 284280
rect 158720 282600 158772 282606
rect 158720 282542 158772 282548
rect 158732 282169 158760 282542
rect 158718 282160 158774 282169
rect 158718 282095 158774 282104
rect 158718 281072 158774 281081
rect 158718 281007 158774 281016
rect 158732 280294 158760 281007
rect 158720 280288 158772 280294
rect 158720 280230 158772 280236
rect 158720 280152 158772 280158
rect 158720 280094 158772 280100
rect 158732 279993 158760 280094
rect 158718 279984 158774 279993
rect 158718 279919 158774 279928
rect 158718 278896 158774 278905
rect 158718 278831 158720 278840
rect 158772 278831 158774 278840
rect 158720 278802 158772 278808
rect 158720 277296 158772 277302
rect 158720 277238 158772 277244
rect 158732 276729 158760 277238
rect 158718 276720 158774 276729
rect 158718 276655 158774 276664
rect 158718 275632 158774 275641
rect 158718 275567 158774 275576
rect 158732 274922 158760 275567
rect 158720 274916 158772 274922
rect 158720 274858 158772 274864
rect 158720 274644 158772 274650
rect 158720 274586 158772 274592
rect 158732 274553 158760 274586
rect 158718 274544 158774 274553
rect 158718 274479 158774 274488
rect 158810 273456 158866 273465
rect 158810 273391 158866 273400
rect 158718 271280 158774 271289
rect 158718 271215 158774 271224
rect 158732 270570 158760 271215
rect 158824 271182 158852 273391
rect 158812 271176 158864 271182
rect 158812 271118 158864 271124
rect 158720 270564 158772 270570
rect 158720 270506 158772 270512
rect 158718 269104 158774 269113
rect 158718 269039 158720 269048
rect 158772 269039 158774 269048
rect 158720 269010 158772 269016
rect 158258 268016 158314 268025
rect 158258 267951 158314 267960
rect 158718 265840 158774 265849
rect 158718 265775 158774 265784
rect 158732 264994 158760 265775
rect 158720 264988 158772 264994
rect 158720 264930 158772 264936
rect 158720 262676 158772 262682
rect 158720 262618 158772 262624
rect 158732 262585 158760 262618
rect 158718 262576 158774 262585
rect 158718 262511 158774 262520
rect 158996 261588 159048 261594
rect 158996 261530 159048 261536
rect 159008 261497 159036 261530
rect 158994 261488 159050 261497
rect 158994 261423 159050 261432
rect 158810 258224 158866 258233
rect 158810 258159 158866 258168
rect 158824 258126 158852 258159
rect 158812 258120 158864 258126
rect 158812 258062 158864 258068
rect 158720 258052 158772 258058
rect 158720 257994 158772 258000
rect 158732 257145 158760 257994
rect 158718 257136 158774 257145
rect 158718 257071 158774 257080
rect 158718 256320 158774 256329
rect 158718 256255 158774 256264
rect 158536 255332 158588 255338
rect 158536 255274 158588 255280
rect 158548 255241 158576 255274
rect 158534 255232 158590 255241
rect 158534 255167 158590 255176
rect 158260 254584 158312 254590
rect 158260 254526 158312 254532
rect 158166 242176 158222 242185
rect 158166 242111 158222 242120
rect 158272 233170 158300 254526
rect 158732 253230 158760 256255
rect 158720 253224 158772 253230
rect 158720 253166 158772 253172
rect 158718 253056 158774 253065
rect 158718 252991 158774 253000
rect 158732 252618 158760 252991
rect 158720 252612 158772 252618
rect 158720 252554 158772 252560
rect 158904 251252 158956 251258
rect 158904 251194 158956 251200
rect 158718 250880 158774 250889
rect 158718 250815 158774 250824
rect 158732 249830 158760 250815
rect 158720 249824 158772 249830
rect 158720 249766 158772 249772
rect 158810 249792 158866 249801
rect 158810 249727 158866 249736
rect 158824 248470 158852 249727
rect 158916 248713 158944 251194
rect 158902 248704 158958 248713
rect 158902 248639 158958 248648
rect 158812 248464 158864 248470
rect 158812 248406 158864 248412
rect 158718 244352 158774 244361
rect 158718 244287 158720 244296
rect 158772 244287 158774 244296
rect 158720 244258 158772 244264
rect 158718 243264 158774 243273
rect 158718 243199 158774 243208
rect 158732 242962 158760 243199
rect 158720 242956 158772 242962
rect 158720 242898 158772 242904
rect 158718 233200 158774 233209
rect 158260 233164 158312 233170
rect 158718 233135 158774 233144
rect 158260 233106 158312 233112
rect 158732 231878 158760 233135
rect 159376 232801 159404 319359
rect 159468 304298 159496 329734
rect 159546 311264 159602 311273
rect 159546 311199 159602 311208
rect 159560 305697 159588 311199
rect 160006 308000 160062 308009
rect 160112 307986 160140 378655
rect 160744 356720 160796 356726
rect 160744 356662 160796 356668
rect 160190 329624 160246 329633
rect 160190 329559 160246 329568
rect 160204 326505 160232 329559
rect 160190 326496 160246 326505
rect 160190 326431 160246 326440
rect 160756 324222 160784 356662
rect 160744 324216 160796 324222
rect 160744 324158 160796 324164
rect 160742 316704 160798 316713
rect 160742 316639 160798 316648
rect 160062 307958 160140 307986
rect 160006 307935 160062 307944
rect 159546 305688 159602 305697
rect 159546 305623 159602 305632
rect 159456 304292 159508 304298
rect 159456 304234 159508 304240
rect 160112 302938 160140 307958
rect 160100 302932 160152 302938
rect 160100 302874 160152 302880
rect 159456 302252 159508 302258
rect 159456 302194 159508 302200
rect 159468 283257 159496 302194
rect 159914 299296 159970 299305
rect 159914 299231 159970 299240
rect 159928 296177 159956 299231
rect 160008 296744 160060 296750
rect 160008 296686 160060 296692
rect 159914 296168 159970 296177
rect 159914 296103 159970 296112
rect 160020 296041 160048 296686
rect 160006 296032 160062 296041
rect 160006 295967 160062 295976
rect 159548 294636 159600 294642
rect 159548 294578 159600 294584
rect 159454 283248 159510 283257
rect 159454 283183 159510 283192
rect 159456 261588 159508 261594
rect 159456 261530 159508 261536
rect 159178 232792 159234 232801
rect 159178 232727 159180 232736
rect 159232 232727 159234 232736
rect 159362 232792 159418 232801
rect 159362 232727 159418 232736
rect 159180 232698 159232 232704
rect 158720 231872 158772 231878
rect 158720 231814 158772 231820
rect 158076 226296 158128 226302
rect 158076 226238 158128 226244
rect 157982 199880 158038 199889
rect 157982 199815 158038 199824
rect 158088 199481 158116 226238
rect 158168 224188 158220 224194
rect 158168 224130 158220 224136
rect 158180 211070 158208 224130
rect 158168 211064 158220 211070
rect 158168 211006 158220 211012
rect 159468 200114 159496 261530
rect 159560 247625 159588 294578
rect 159638 271824 159694 271833
rect 159638 271759 159694 271768
rect 159652 270201 159680 271759
rect 159638 270192 159694 270201
rect 159638 270127 159694 270136
rect 159652 269822 159680 270127
rect 159640 269816 159692 269822
rect 159640 269758 159692 269764
rect 160098 260808 160154 260817
rect 160098 260743 160154 260752
rect 159730 249112 159786 249121
rect 159730 249047 159786 249056
rect 159546 247616 159602 247625
rect 159546 247551 159602 247560
rect 159744 238754 159772 249047
rect 160006 244896 160062 244905
rect 160006 244831 160062 244840
rect 159652 238726 159772 238754
rect 159652 222154 159680 238726
rect 160020 224233 160048 244831
rect 160006 224224 160062 224233
rect 160006 224159 160062 224168
rect 159640 222148 159692 222154
rect 159640 222090 159692 222096
rect 160112 202881 160140 260743
rect 160192 241392 160244 241398
rect 160192 241334 160244 241340
rect 160204 241097 160232 241334
rect 160190 241088 160246 241097
rect 160190 241023 160246 241032
rect 160756 206689 160784 316639
rect 160848 296857 160876 378762
rect 162122 370696 162178 370705
rect 162122 370631 162178 370640
rect 161480 343732 161532 343738
rect 161480 343674 161532 343680
rect 161492 327894 161520 343674
rect 161480 327888 161532 327894
rect 161480 327830 161532 327836
rect 161480 327344 161532 327350
rect 161480 327286 161532 327292
rect 161492 324970 161520 327286
rect 161480 324964 161532 324970
rect 161480 324906 161532 324912
rect 160834 296848 160890 296857
rect 160834 296783 160890 296792
rect 160848 262682 160876 296783
rect 161020 274916 161072 274922
rect 161020 274858 161072 274864
rect 160928 262880 160980 262886
rect 160928 262822 160980 262828
rect 160836 262676 160888 262682
rect 160836 262618 160888 262624
rect 160834 251832 160890 251841
rect 160834 251767 160890 251776
rect 160742 206680 160798 206689
rect 160742 206615 160798 206624
rect 160098 202872 160154 202881
rect 160098 202807 160154 202816
rect 160848 200114 160876 251767
rect 160940 226137 160968 262822
rect 161032 261526 161060 274858
rect 161020 261520 161072 261526
rect 161020 261462 161072 261468
rect 161572 244928 161624 244934
rect 161572 244870 161624 244876
rect 161584 240961 161612 244870
rect 161570 240952 161626 240961
rect 161570 240887 161626 240896
rect 160926 226128 160982 226137
rect 160926 226063 160982 226072
rect 162136 211041 162164 370631
rect 162228 290222 162256 436086
rect 162780 344321 162808 564402
rect 166356 561808 166408 561814
rect 166356 561750 166408 561756
rect 166264 538280 166316 538286
rect 166264 538222 166316 538228
rect 164884 504416 164936 504422
rect 164884 504358 164936 504364
rect 163504 441652 163556 441658
rect 163504 441594 163556 441600
rect 162952 346452 163004 346458
rect 162952 346394 163004 346400
rect 162766 344312 162822 344321
rect 162766 344247 162822 344256
rect 162858 342136 162914 342145
rect 162858 342071 162914 342080
rect 162308 338224 162360 338230
rect 162308 338166 162360 338172
rect 162216 290216 162268 290222
rect 162216 290158 162268 290164
rect 162216 283892 162268 283898
rect 162216 283834 162268 283840
rect 162228 237318 162256 283834
rect 162320 279478 162348 338166
rect 162768 284368 162820 284374
rect 162768 284310 162820 284316
rect 162780 282198 162808 284310
rect 162768 282192 162820 282198
rect 162768 282134 162820 282140
rect 162308 279472 162360 279478
rect 162308 279414 162360 279420
rect 162400 278860 162452 278866
rect 162400 278802 162452 278808
rect 162412 247790 162440 278802
rect 162768 260840 162820 260846
rect 162768 260782 162820 260788
rect 162780 260681 162808 260782
rect 162766 260672 162822 260681
rect 162766 260607 162822 260616
rect 162492 250504 162544 250510
rect 162492 250446 162544 250452
rect 162400 247784 162452 247790
rect 162400 247726 162452 247732
rect 162216 237312 162268 237318
rect 162216 237254 162268 237260
rect 162504 234297 162532 250446
rect 162872 238754 162900 342071
rect 162964 340202 162992 346394
rect 162952 340196 163004 340202
rect 162952 340138 163004 340144
rect 162952 336116 163004 336122
rect 162952 336058 163004 336064
rect 162964 330886 162992 336058
rect 162952 330880 163004 330886
rect 162952 330822 163004 330828
rect 162950 327720 163006 327729
rect 162950 327655 163006 327664
rect 162964 324902 162992 327655
rect 162952 324896 163004 324902
rect 162952 324838 163004 324844
rect 162950 288552 163006 288561
rect 162950 288487 163006 288496
rect 162964 282606 162992 288487
rect 162952 282600 163004 282606
rect 162952 282542 163004 282548
rect 163516 262177 163544 441594
rect 164148 411324 164200 411330
rect 164148 411266 164200 411272
rect 163596 325440 163648 325446
rect 163596 325382 163648 325388
rect 163608 282266 163636 325382
rect 164160 314702 164188 411266
rect 164896 374134 164924 504358
rect 165528 467900 165580 467906
rect 165528 467842 165580 467848
rect 164884 374128 164936 374134
rect 164884 374070 164936 374076
rect 164148 314696 164200 314702
rect 164148 314638 164200 314644
rect 164896 313313 164924 374070
rect 164974 339552 165030 339561
rect 164974 339487 165030 339496
rect 164988 322153 165016 339487
rect 165158 337376 165214 337385
rect 165158 337311 165214 337320
rect 165172 329118 165200 337311
rect 165160 329112 165212 329118
rect 165160 329054 165212 329060
rect 165160 328500 165212 328506
rect 165160 328442 165212 328448
rect 165172 325009 165200 328442
rect 165158 325000 165214 325009
rect 165158 324935 165214 324944
rect 165068 324896 165120 324902
rect 165068 324838 165120 324844
rect 165080 323649 165108 324838
rect 165066 323640 165122 323649
rect 165066 323575 165122 323584
rect 164974 322144 165030 322153
rect 164974 322079 165030 322088
rect 164976 320204 165028 320210
rect 164976 320146 165028 320152
rect 164882 313304 164938 313313
rect 164882 313239 164938 313248
rect 164988 311846 165016 320146
rect 165434 313304 165490 313313
rect 165434 313239 165490 313248
rect 164976 311840 165028 311846
rect 164976 311782 165028 311788
rect 164976 304292 165028 304298
rect 164976 304234 165028 304240
rect 164882 303648 164938 303657
rect 164882 303583 164938 303592
rect 164896 286346 164924 303583
rect 164884 286340 164936 286346
rect 164884 286282 164936 286288
rect 164884 284980 164936 284986
rect 164884 284922 164936 284928
rect 163596 282260 163648 282266
rect 163596 282202 163648 282208
rect 163688 280220 163740 280226
rect 163688 280162 163740 280168
rect 163596 275324 163648 275330
rect 163596 275266 163648 275272
rect 163502 262168 163558 262177
rect 163502 262103 163558 262112
rect 163502 254552 163558 254561
rect 163502 254487 163558 254496
rect 162780 238726 162900 238754
rect 162490 234288 162546 234297
rect 162490 234223 162546 234232
rect 162780 233753 162808 238726
rect 162214 233744 162270 233753
rect 162214 233679 162270 233688
rect 162766 233744 162822 233753
rect 162766 233679 162822 233688
rect 162122 211032 162178 211041
rect 162122 210967 162178 210976
rect 162228 205601 162256 233679
rect 162780 233345 162808 233679
rect 162766 233336 162822 233345
rect 162766 233271 162822 233280
rect 163516 223281 163544 254487
rect 163608 230353 163636 275266
rect 163700 258058 163728 280162
rect 163778 261488 163834 261497
rect 163778 261423 163834 261432
rect 163688 258052 163740 258058
rect 163688 257994 163740 258000
rect 163792 252482 163820 261423
rect 164148 256760 164200 256766
rect 164148 256702 164200 256708
rect 164160 254153 164188 256702
rect 164146 254144 164202 254153
rect 164146 254079 164202 254088
rect 163780 252476 163832 252482
rect 163780 252418 163832 252424
rect 163686 250472 163742 250481
rect 163686 250407 163742 250416
rect 163700 234569 163728 250407
rect 163686 234560 163742 234569
rect 163686 234495 163742 234504
rect 163594 230344 163650 230353
rect 163594 230279 163650 230288
rect 164896 228993 164924 284922
rect 164988 258738 165016 304234
rect 165448 289814 165476 313239
rect 165540 303657 165568 467842
rect 166276 363769 166304 538222
rect 166368 444378 166396 561750
rect 173806 557560 173862 557569
rect 173806 557495 173862 557504
rect 172428 538892 172480 538898
rect 172428 538834 172480 538840
rect 169022 526416 169078 526425
rect 169022 526351 169078 526360
rect 166356 444372 166408 444378
rect 166356 444314 166408 444320
rect 166262 363760 166318 363769
rect 166262 363695 166318 363704
rect 165894 332752 165950 332761
rect 165894 332687 165950 332696
rect 165620 330880 165672 330886
rect 165620 330822 165672 330828
rect 165632 326398 165660 330822
rect 165908 330614 165936 332687
rect 166368 332246 166396 444314
rect 169036 439550 169064 526351
rect 170404 524476 170456 524482
rect 170404 524418 170456 524424
rect 169024 439544 169076 439550
rect 169024 439486 169076 439492
rect 169024 427848 169076 427854
rect 169024 427790 169076 427796
rect 167644 423700 167696 423706
rect 167644 423642 167696 423648
rect 167184 388476 167236 388482
rect 167184 388418 167236 388424
rect 167196 388385 167224 388418
rect 167182 388376 167238 388385
rect 167182 388311 167238 388320
rect 167000 381540 167052 381546
rect 167000 381482 167052 381488
rect 167012 381002 167040 381482
rect 167000 380996 167052 381002
rect 167000 380938 167052 380944
rect 166908 363656 166960 363662
rect 166908 363598 166960 363604
rect 166356 332240 166408 332246
rect 166356 332182 166408 332188
rect 166264 331900 166316 331906
rect 166264 331842 166316 331848
rect 165896 330608 165948 330614
rect 165896 330550 165948 330556
rect 165620 326392 165672 326398
rect 165620 326334 165672 326340
rect 165526 303648 165582 303657
rect 165526 303583 165582 303592
rect 166276 290494 166304 331842
rect 166448 329180 166500 329186
rect 166448 329122 166500 329128
rect 166356 321632 166408 321638
rect 166356 321574 166408 321580
rect 166368 298761 166396 321574
rect 166460 320890 166488 329122
rect 166920 325694 166948 363598
rect 166736 325666 166948 325694
rect 166448 320884 166500 320890
rect 166448 320826 166500 320832
rect 166736 317422 166764 325666
rect 167012 319462 167040 380938
rect 167656 358086 167684 423642
rect 168288 388476 168340 388482
rect 168288 388418 168340 388424
rect 167736 358148 167788 358154
rect 167736 358090 167788 358096
rect 167092 358080 167144 358086
rect 167092 358022 167144 358028
rect 167644 358080 167696 358086
rect 167644 358022 167696 358028
rect 167104 356862 167132 358022
rect 167092 356856 167144 356862
rect 167092 356798 167144 356804
rect 167748 356794 167776 358090
rect 167736 356788 167788 356794
rect 167736 356730 167788 356736
rect 167642 343768 167698 343777
rect 167642 343703 167698 343712
rect 167656 331906 167684 343703
rect 167644 331900 167696 331906
rect 167644 331842 167696 331848
rect 167748 331022 167776 356730
rect 167736 331016 167788 331022
rect 167736 330958 167788 330964
rect 167644 329860 167696 329866
rect 167644 329802 167696 329808
rect 167000 319456 167052 319462
rect 167000 319398 167052 319404
rect 167012 318730 167040 319398
rect 166828 318702 167040 318730
rect 166448 317416 166500 317422
rect 166448 317358 166500 317364
rect 166724 317416 166776 317422
rect 166724 317358 166776 317364
rect 166460 316742 166488 317358
rect 166448 316736 166500 316742
rect 166448 316678 166500 316684
rect 166354 298752 166410 298761
rect 166354 298687 166410 298696
rect 166264 290488 166316 290494
rect 166264 290430 166316 290436
rect 165436 289808 165488 289814
rect 165436 289750 165488 289756
rect 166356 289808 166408 289814
rect 166356 289750 166408 289756
rect 165068 287700 165120 287706
rect 165068 287642 165120 287648
rect 165080 262886 165108 287642
rect 166264 287088 166316 287094
rect 166264 287030 166316 287036
rect 165068 262880 165120 262886
rect 165068 262822 165120 262828
rect 165436 262880 165488 262886
rect 165436 262822 165488 262828
rect 165066 262168 165122 262177
rect 165066 262103 165122 262112
rect 164976 258732 165028 258738
rect 164976 258674 165028 258680
rect 165080 242865 165108 262103
rect 165066 242856 165122 242865
rect 165066 242791 165122 242800
rect 165448 230382 165476 262822
rect 165526 253192 165582 253201
rect 165526 253127 165582 253136
rect 165436 230376 165488 230382
rect 165436 230318 165488 230324
rect 165448 229634 165476 230318
rect 165436 229628 165488 229634
rect 165436 229570 165488 229576
rect 164882 228984 164938 228993
rect 164882 228919 164938 228928
rect 163502 223272 163558 223281
rect 163502 223207 163558 223216
rect 162766 211032 162822 211041
rect 162766 210967 162822 210976
rect 162780 210769 162808 210967
rect 162766 210760 162822 210769
rect 162766 210695 162822 210704
rect 162214 205592 162270 205601
rect 162214 205527 162270 205536
rect 159376 200086 159496 200114
rect 160756 200086 160876 200114
rect 158074 199472 158130 199481
rect 158074 199407 158130 199416
rect 156788 198620 156840 198626
rect 156788 198562 156840 198568
rect 156800 196897 156828 198562
rect 156786 196888 156842 196897
rect 156786 196823 156842 196832
rect 159376 195906 159404 200086
rect 160756 198694 160784 200086
rect 160744 198688 160796 198694
rect 160744 198630 160796 198636
rect 158720 195900 158772 195906
rect 158720 195842 158772 195848
rect 159364 195900 159416 195906
rect 159364 195842 159416 195848
rect 158732 195294 158760 195842
rect 158720 195288 158772 195294
rect 158720 195230 158772 195236
rect 156602 193896 156658 193905
rect 156602 193831 156658 193840
rect 155868 189780 155920 189786
rect 155868 189722 155920 189728
rect 133788 186380 133840 186386
rect 133788 186322 133840 186328
rect 133142 178664 133198 178673
rect 133142 178599 133198 178608
rect 132408 178152 132460 178158
rect 132408 178094 132460 178100
rect 129096 178016 129148 178022
rect 129096 177958 129148 177964
rect 132420 176769 132448 178094
rect 133800 177585 133828 186322
rect 134800 182300 134852 182306
rect 134800 182242 134852 182248
rect 134812 177585 134840 182242
rect 148232 180940 148284 180946
rect 148232 180882 148284 180888
rect 148244 177585 148272 180882
rect 160756 178809 160784 198630
rect 163516 187241 163544 223207
rect 165540 191826 165568 253127
rect 166276 240854 166304 287030
rect 166368 276185 166396 289750
rect 166724 284368 166776 284374
rect 166724 284310 166776 284316
rect 166354 276176 166410 276185
rect 166354 276111 166410 276120
rect 166448 267096 166500 267102
rect 166448 267038 166500 267044
rect 166460 266393 166488 267038
rect 166446 266384 166502 266393
rect 166446 266319 166502 266328
rect 166356 252612 166408 252618
rect 166356 252554 166408 252560
rect 166264 240848 166316 240854
rect 166264 240790 166316 240796
rect 166368 230382 166396 252554
rect 166736 237425 166764 284310
rect 166828 255513 166856 318702
rect 167656 274038 167684 329802
rect 168102 328400 168158 328409
rect 168102 328335 168158 328344
rect 168116 327758 168144 328335
rect 168104 327752 168156 327758
rect 168104 327694 168156 327700
rect 167644 274032 167696 274038
rect 167644 273974 167696 273980
rect 167736 271176 167788 271182
rect 167736 271118 167788 271124
rect 167644 268388 167696 268394
rect 167644 268330 167696 268336
rect 166906 266384 166962 266393
rect 166906 266319 166962 266328
rect 166814 255504 166870 255513
rect 166814 255439 166870 255448
rect 166722 237416 166778 237425
rect 166722 237351 166778 237360
rect 166356 230376 166408 230382
rect 166356 230318 166408 230324
rect 166264 229628 166316 229634
rect 166264 229570 166316 229576
rect 165528 191820 165580 191826
rect 165528 191762 165580 191768
rect 164884 189780 164936 189786
rect 164884 189722 164936 189728
rect 163502 187232 163558 187241
rect 163502 187167 163558 187176
rect 162860 182300 162912 182306
rect 162860 182242 162912 182248
rect 160742 178800 160798 178809
rect 160742 178735 160798 178744
rect 133786 177576 133842 177585
rect 133786 177511 133842 177520
rect 134798 177576 134854 177585
rect 134798 177511 134854 177520
rect 148230 177576 148286 177585
rect 148230 177511 148286 177520
rect 136088 176792 136140 176798
rect 130750 176760 130806 176769
rect 130750 176695 130752 176704
rect 130804 176695 130806 176704
rect 132406 176760 132462 176769
rect 132406 176695 132462 176704
rect 136086 176760 136088 176769
rect 140780 176792 140832 176798
rect 136140 176760 136142 176769
rect 158996 176792 159048 176798
rect 140780 176734 140832 176740
rect 158994 176760 158996 176769
rect 159048 176760 159050 176769
rect 136086 176695 136142 176704
rect 130752 176666 130804 176672
rect 140792 176662 140820 176734
rect 158994 176695 159050 176704
rect 140780 176656 140832 176662
rect 140780 176598 140832 176604
rect 129004 175976 129056 175982
rect 129004 175918 129056 175924
rect 129464 175976 129516 175982
rect 129464 175918 129516 175924
rect 129476 175681 129504 175918
rect 129462 175672 129518 175681
rect 129462 175607 129518 175616
rect 162872 175234 162900 182242
rect 164896 175273 164924 189722
rect 165528 178152 165580 178158
rect 165528 178094 165580 178100
rect 164974 177032 165030 177041
rect 164974 176967 165030 176976
rect 164882 175264 164938 175273
rect 162860 175228 162912 175234
rect 164882 175199 164938 175208
rect 162860 175170 162912 175176
rect 164988 171018 165016 176967
rect 165158 175672 165214 175681
rect 165158 175607 165214 175616
rect 165172 171086 165200 175607
rect 165540 173874 165568 178094
rect 165528 173868 165580 173874
rect 165528 173810 165580 173816
rect 165160 171080 165212 171086
rect 165160 171022 165212 171028
rect 164976 171012 165028 171018
rect 164976 170954 165028 170960
rect 67638 123584 67694 123593
rect 67638 123519 67694 123528
rect 67454 120864 67510 120873
rect 67454 120799 67510 120808
rect 67362 100736 67418 100745
rect 67362 100671 67418 100680
rect 67376 90370 67404 100671
rect 67468 91798 67496 120799
rect 67546 102368 67602 102377
rect 67546 102303 67602 102312
rect 67560 95033 67588 102303
rect 67546 95024 67602 95033
rect 67546 94959 67602 94968
rect 67456 91792 67508 91798
rect 67456 91734 67508 91740
rect 67364 90364 67416 90370
rect 67364 90306 67416 90312
rect 67652 67590 67680 123519
rect 166276 106865 166304 229570
rect 166354 183696 166410 183705
rect 166354 183631 166410 183640
rect 166368 157350 166396 183631
rect 166920 182073 166948 266319
rect 167656 231577 167684 268330
rect 167748 249082 167776 271118
rect 168116 269793 168144 327694
rect 168196 270632 168248 270638
rect 168196 270574 168248 270580
rect 168102 269784 168158 269793
rect 168102 269719 168158 269728
rect 167826 249248 167882 249257
rect 167826 249183 167882 249192
rect 167736 249076 167788 249082
rect 167736 249018 167788 249024
rect 167840 240786 167868 249183
rect 167918 242856 167974 242865
rect 167918 242791 167974 242800
rect 167932 241641 167960 242791
rect 167918 241632 167974 241641
rect 167918 241567 167974 241576
rect 167828 240780 167880 240786
rect 167828 240722 167880 240728
rect 167734 237416 167790 237425
rect 167734 237351 167790 237360
rect 167642 231568 167698 231577
rect 167642 231503 167698 231512
rect 167000 221468 167052 221474
rect 167000 221410 167052 221416
rect 167012 220561 167040 221410
rect 166998 220552 167054 220561
rect 166998 220487 167054 220496
rect 167656 199345 167684 231503
rect 167748 221474 167776 237351
rect 167932 237153 167960 241567
rect 167918 237144 167974 237153
rect 167918 237079 167974 237088
rect 168208 234666 168236 270574
rect 168300 242865 168328 388418
rect 168380 332240 168432 332246
rect 168380 332182 168432 332188
rect 168286 242856 168342 242865
rect 168286 242791 168342 242800
rect 168392 237425 168420 332182
rect 169036 284374 169064 427790
rect 169116 371340 169168 371346
rect 169116 371282 169168 371288
rect 169128 337521 169156 371282
rect 169208 369232 169260 369238
rect 169208 369174 169260 369180
rect 169114 337512 169170 337521
rect 169114 337447 169170 337456
rect 169116 331016 169168 331022
rect 169116 330958 169168 330964
rect 169024 284368 169076 284374
rect 169024 284310 169076 284316
rect 169024 280288 169076 280294
rect 169024 280230 169076 280236
rect 169036 277370 169064 280230
rect 169024 277364 169076 277370
rect 169024 277306 169076 277312
rect 169128 269890 169156 330958
rect 169220 329798 169248 369174
rect 170416 336841 170444 524418
rect 171048 477556 171100 477562
rect 171048 477498 171100 477504
rect 170494 356824 170550 356833
rect 170494 356759 170550 356768
rect 170402 336832 170458 336841
rect 170402 336767 170458 336776
rect 169208 329792 169260 329798
rect 169208 329734 169260 329740
rect 169668 317552 169720 317558
rect 169668 317494 169720 317500
rect 169208 302932 169260 302938
rect 169208 302874 169260 302880
rect 169220 280537 169248 302874
rect 169680 302433 169708 317494
rect 170416 307086 170444 336767
rect 170404 307080 170456 307086
rect 170404 307022 170456 307028
rect 169666 302424 169722 302433
rect 169666 302359 169722 302368
rect 170402 284336 170458 284345
rect 170402 284271 170458 284280
rect 169206 280528 169262 280537
rect 169206 280463 169262 280472
rect 169668 275596 169720 275602
rect 169668 275538 169720 275544
rect 169116 269884 169168 269890
rect 169116 269826 169168 269832
rect 169024 256012 169076 256018
rect 169024 255954 169076 255960
rect 168472 247716 168524 247722
rect 168472 247658 168524 247664
rect 168484 242049 168512 247658
rect 168470 242040 168526 242049
rect 168470 241975 168526 241984
rect 168378 237416 168434 237425
rect 168378 237351 168434 237360
rect 168196 234660 168248 234666
rect 168196 234602 168248 234608
rect 167736 221468 167788 221474
rect 167736 221410 167788 221416
rect 169036 213858 169064 255954
rect 169680 247081 169708 275538
rect 170416 274650 170444 284271
rect 170404 274644 170456 274650
rect 170404 274586 170456 274592
rect 170404 269816 170456 269822
rect 170404 269758 170456 269764
rect 169666 247072 169722 247081
rect 169666 247007 169722 247016
rect 169024 213852 169076 213858
rect 169024 213794 169076 213800
rect 167826 199472 167882 199481
rect 167826 199407 167882 199416
rect 168380 199436 168432 199442
rect 167642 199336 167698 199345
rect 167642 199271 167698 199280
rect 167000 198076 167052 198082
rect 167000 198018 167052 198024
rect 167012 193186 167040 198018
rect 167000 193180 167052 193186
rect 167000 193122 167052 193128
rect 166906 182064 166962 182073
rect 166906 181999 166962 182008
rect 166448 180872 166500 180878
rect 166448 180814 166500 180820
rect 166460 165578 166488 180814
rect 167736 179512 167788 179518
rect 167736 179454 167788 179460
rect 167642 178256 167698 178265
rect 167642 178191 167698 178200
rect 166538 175400 166594 175409
rect 166538 175335 166594 175344
rect 166448 165572 166500 165578
rect 166448 165514 166500 165520
rect 166552 165510 166580 175335
rect 166540 165504 166592 165510
rect 166540 165446 166592 165452
rect 167656 162858 167684 178191
rect 167748 167006 167776 179454
rect 167840 173466 167868 199407
rect 168380 199378 168432 199384
rect 168392 198694 168420 199378
rect 168380 198688 168432 198694
rect 168380 198630 168432 198636
rect 169036 192681 169064 213794
rect 169760 200864 169812 200870
rect 169760 200806 169812 200812
rect 169772 200122 169800 200806
rect 169760 200116 169812 200122
rect 169760 200058 169812 200064
rect 169022 192672 169078 192681
rect 169022 192607 169078 192616
rect 169022 186960 169078 186969
rect 169022 186895 169078 186904
rect 167918 175536 167974 175545
rect 167918 175471 167974 175480
rect 167828 173460 167880 173466
rect 167828 173402 167880 173408
rect 167826 171592 167882 171601
rect 167826 171527 167882 171536
rect 167736 167000 167788 167006
rect 167736 166942 167788 166948
rect 167644 162852 167696 162858
rect 167644 162794 167696 162800
rect 167840 159390 167868 171527
rect 167932 168366 167960 175471
rect 167920 168360 167972 168366
rect 167920 168302 167972 168308
rect 167828 159384 167880 159390
rect 167828 159326 167880 159332
rect 166356 157344 166408 157350
rect 166356 157286 166408 157292
rect 166356 153264 166408 153270
rect 166356 153206 166408 153212
rect 166262 106856 166318 106865
rect 166262 106791 166318 106800
rect 166264 104168 166316 104174
rect 166264 104110 166316 104116
rect 164974 101416 165030 101425
rect 164974 101351 165030 101360
rect 164884 98048 164936 98054
rect 164884 97990 164936 97996
rect 113178 94752 113234 94761
rect 113178 94687 113234 94696
rect 130750 94752 130806 94761
rect 130750 94687 130806 94696
rect 97264 94512 97316 94518
rect 97264 94454 97316 94460
rect 74814 92440 74870 92449
rect 74814 92375 74870 92384
rect 74828 91118 74856 92375
rect 88062 92168 88118 92177
rect 88062 92103 88118 92112
rect 86866 91352 86922 91361
rect 86866 91287 86922 91296
rect 85486 91216 85542 91225
rect 85486 91151 85542 91160
rect 86774 91216 86830 91225
rect 86774 91151 86830 91160
rect 74816 91112 74868 91118
rect 74816 91054 74868 91060
rect 85500 69018 85528 91151
rect 86788 84153 86816 91151
rect 86774 84144 86830 84153
rect 86774 84079 86830 84088
rect 86880 82822 86908 91287
rect 88076 90409 88104 92103
rect 91650 92032 91706 92041
rect 91650 91967 91706 91976
rect 89074 91216 89130 91225
rect 89074 91151 89130 91160
rect 91006 91216 91062 91225
rect 91006 91151 91062 91160
rect 88062 90400 88118 90409
rect 88062 90335 88118 90344
rect 89088 85513 89116 91151
rect 89720 91112 89772 91118
rect 89720 91054 89772 91060
rect 89732 86873 89760 91054
rect 89718 86864 89774 86873
rect 89718 86799 89774 86808
rect 89074 85504 89130 85513
rect 89074 85439 89130 85448
rect 86868 82816 86920 82822
rect 86868 82758 86920 82764
rect 86866 76528 86922 76537
rect 86866 76463 86922 76472
rect 85488 69012 85540 69018
rect 85488 68954 85540 68960
rect 67640 67584 67692 67590
rect 67640 67526 67692 67532
rect 77206 64288 77262 64297
rect 77206 64223 77262 64232
rect 68928 62824 68980 62830
rect 68928 62766 68980 62772
rect 67180 47592 67232 47598
rect 67180 47534 67232 47540
rect 66720 7608 66772 7614
rect 66720 7550 66772 7556
rect 65524 3528 65576 3534
rect 65524 3470 65576 3476
rect 66168 3528 66220 3534
rect 66168 3470 66220 3476
rect 65536 480 65564 3470
rect 66732 480 66760 7550
rect 68940 3534 68968 62766
rect 75826 61432 75882 61441
rect 73068 61396 73120 61402
rect 75826 61367 75882 61376
rect 73068 61338 73120 61344
rect 70308 60036 70360 60042
rect 70308 59978 70360 59984
rect 70216 33788 70268 33794
rect 70216 33730 70268 33736
rect 70228 16574 70256 33730
rect 70136 16546 70256 16574
rect 69112 3596 69164 3602
rect 69112 3538 69164 3544
rect 67916 3528 67968 3534
rect 67916 3470 67968 3476
rect 68928 3528 68980 3534
rect 68928 3470 68980 3476
rect 67928 480 67956 3470
rect 69124 480 69152 3538
rect 70136 3482 70164 16546
rect 70320 6914 70348 59978
rect 71044 35216 71096 35222
rect 71044 35158 71096 35164
rect 70228 6886 70348 6914
rect 70228 3602 70256 6886
rect 71056 3670 71084 35158
rect 71044 3664 71096 3670
rect 71044 3606 71096 3612
rect 70216 3596 70268 3602
rect 70216 3538 70268 3544
rect 73080 3534 73108 61338
rect 74448 46232 74500 46238
rect 74448 46174 74500 46180
rect 74460 3534 74488 46174
rect 75840 3534 75868 61367
rect 77220 3534 77248 64223
rect 79966 62792 80022 62801
rect 79966 62727 80022 62736
rect 78586 58576 78642 58585
rect 78586 58511 78642 58520
rect 72608 3528 72660 3534
rect 70136 3454 70348 3482
rect 72608 3470 72660 3476
rect 73068 3528 73120 3534
rect 73068 3470 73120 3476
rect 73804 3528 73856 3534
rect 73804 3470 73856 3476
rect 74448 3528 74500 3534
rect 74448 3470 74500 3476
rect 75000 3528 75052 3534
rect 75000 3470 75052 3476
rect 75828 3528 75880 3534
rect 75828 3470 75880 3476
rect 76196 3528 76248 3534
rect 76196 3470 76248 3476
rect 77208 3528 77260 3534
rect 77208 3470 77260 3476
rect 70320 480 70348 3454
rect 71504 2100 71556 2106
rect 71504 2042 71556 2048
rect 71516 480 71544 2042
rect 72620 480 72648 3470
rect 73816 480 73844 3470
rect 75012 480 75040 3470
rect 76208 480 76236 3470
rect 77390 3360 77446 3369
rect 77390 3295 77446 3304
rect 77404 480 77432 3295
rect 78600 480 78628 58511
rect 79980 6914 80008 62727
rect 82726 59936 82782 59945
rect 82726 59871 82782 59880
rect 81348 10396 81400 10402
rect 81348 10338 81400 10344
rect 79704 6886 80008 6914
rect 79704 480 79732 6886
rect 81360 3534 81388 10338
rect 80888 3528 80940 3534
rect 80888 3470 80940 3476
rect 81348 3528 81400 3534
rect 81348 3470 81400 3476
rect 80900 480 80928 3470
rect 82740 3058 82768 59871
rect 84108 43512 84160 43518
rect 84108 43454 84160 43460
rect 84120 3194 84148 43454
rect 85488 32496 85540 32502
rect 85488 32438 85540 32444
rect 85500 3262 85528 32438
rect 85672 9036 85724 9042
rect 85672 8978 85724 8984
rect 84476 3256 84528 3262
rect 84476 3198 84528 3204
rect 85488 3256 85540 3262
rect 85488 3198 85540 3204
rect 83280 3188 83332 3194
rect 83280 3130 83332 3136
rect 84108 3188 84160 3194
rect 84108 3130 84160 3136
rect 82084 3052 82136 3058
rect 82084 2994 82136 3000
rect 82728 3052 82780 3058
rect 82728 2994 82780 3000
rect 82096 480 82124 2994
rect 83292 480 83320 3130
rect 84488 480 84516 3198
rect 85684 480 85712 8978
rect 86880 480 86908 76463
rect 87602 75304 87658 75313
rect 87602 75239 87658 75248
rect 87616 3466 87644 75239
rect 91020 74458 91048 91151
rect 91664 89593 91692 91967
rect 95054 91352 95110 91361
rect 95054 91287 95110 91296
rect 93674 91216 93730 91225
rect 93674 91151 93730 91160
rect 91650 89584 91706 89593
rect 91650 89519 91706 89528
rect 91008 74452 91060 74458
rect 91008 74394 91060 74400
rect 93688 67522 93716 91151
rect 95068 87650 95096 91287
rect 95146 91216 95202 91225
rect 95146 91151 95202 91160
rect 96526 91216 96582 91225
rect 96526 91151 96582 91160
rect 95056 87644 95108 87650
rect 95056 87586 95108 87592
rect 95160 81394 95188 91151
rect 96540 84017 96568 91151
rect 96526 84008 96582 84017
rect 96526 83943 96582 83952
rect 95148 81388 95200 81394
rect 95148 81330 95200 81336
rect 97276 75886 97304 94454
rect 113192 93906 113220 94687
rect 130764 93974 130792 94687
rect 162124 94512 162176 94518
rect 162124 94454 162176 94460
rect 162858 94480 162914 94489
rect 130752 93968 130804 93974
rect 130752 93910 130804 93916
rect 113180 93900 113232 93906
rect 113180 93842 113232 93848
rect 153200 93900 153252 93906
rect 162136 93854 162164 94454
rect 162858 94415 162914 94424
rect 153200 93842 153252 93848
rect 119710 93392 119766 93401
rect 119710 93327 119766 93336
rect 123022 93392 123078 93401
rect 123022 93327 123078 93336
rect 103426 93256 103482 93265
rect 103426 93191 103482 93200
rect 97354 92440 97410 92449
rect 97354 92375 97410 92384
rect 100114 92440 100170 92449
rect 100114 92375 100170 92384
rect 103150 92440 103206 92449
rect 103150 92375 103206 92384
rect 97368 91186 97396 92375
rect 100024 91792 100076 91798
rect 100024 91734 100076 91740
rect 98734 91352 98790 91361
rect 98734 91287 98790 91296
rect 97814 91216 97870 91225
rect 97356 91180 97408 91186
rect 97814 91151 97870 91160
rect 97356 91122 97408 91128
rect 97828 80073 97856 91151
rect 98748 86737 98776 91287
rect 99286 91216 99342 91225
rect 99286 91151 99342 91160
rect 98734 86728 98790 86737
rect 98734 86663 98790 86672
rect 98644 83496 98696 83502
rect 98644 83438 98696 83444
rect 97814 80064 97870 80073
rect 97814 79999 97870 80008
rect 97264 75880 97316 75886
rect 97264 75822 97316 75828
rect 93766 69728 93822 69737
rect 93766 69663 93822 69672
rect 93676 67516 93728 67522
rect 93676 67458 93728 67464
rect 91008 57248 91060 57254
rect 91008 57190 91060 57196
rect 89628 53100 89680 53106
rect 89628 53042 89680 53048
rect 88248 20052 88300 20058
rect 88248 19994 88300 20000
rect 88260 6914 88288 19994
rect 87984 6886 88288 6914
rect 87604 3460 87656 3466
rect 87604 3402 87656 3408
rect 87984 480 88012 6886
rect 89640 3330 89668 53042
rect 91020 3534 91048 57190
rect 92388 22840 92440 22846
rect 92388 22782 92440 22788
rect 92400 3534 92428 22782
rect 93780 3534 93808 69663
rect 95146 68232 95202 68241
rect 95146 68167 95202 68176
rect 95056 21412 95108 21418
rect 95056 21354 95108 21360
rect 95068 3534 95096 21354
rect 90364 3528 90416 3534
rect 90364 3470 90416 3476
rect 91008 3528 91060 3534
rect 91008 3470 91060 3476
rect 91560 3528 91612 3534
rect 91560 3470 91612 3476
rect 92388 3528 92440 3534
rect 92388 3470 92440 3476
rect 92756 3528 92808 3534
rect 92756 3470 92808 3476
rect 93768 3528 93820 3534
rect 93768 3470 93820 3476
rect 93952 3528 94004 3534
rect 93952 3470 94004 3476
rect 95056 3528 95108 3534
rect 95056 3470 95108 3476
rect 89168 3324 89220 3330
rect 89168 3266 89220 3272
rect 89628 3324 89680 3330
rect 89628 3266 89680 3272
rect 89180 480 89208 3266
rect 90376 480 90404 3470
rect 91572 480 91600 3470
rect 92768 480 92796 3470
rect 93964 480 93992 3470
rect 95160 480 95188 68167
rect 97908 55888 97960 55894
rect 97908 55830 97960 55836
rect 96252 13184 96304 13190
rect 96252 13126 96304 13132
rect 96264 480 96292 13126
rect 97920 3534 97948 55830
rect 98656 18601 98684 83438
rect 99300 60722 99328 91151
rect 100036 77246 100064 91734
rect 100128 91118 100156 92375
rect 100574 91216 100630 91225
rect 100574 91151 100630 91160
rect 102046 91216 102102 91225
rect 102046 91151 102102 91160
rect 100116 91112 100168 91118
rect 100116 91054 100168 91060
rect 100588 85241 100616 91151
rect 100574 85232 100630 85241
rect 100574 85167 100630 85176
rect 100024 77240 100076 77246
rect 100024 77182 100076 77188
rect 102060 71670 102088 91151
rect 103164 91050 103192 92375
rect 103152 91044 103204 91050
rect 103152 90986 103204 90992
rect 102048 71664 102100 71670
rect 102048 71606 102100 71612
rect 99288 60716 99340 60722
rect 99288 60658 99340 60664
rect 103440 59362 103468 93191
rect 119724 93158 119752 93327
rect 123036 93226 123064 93327
rect 123024 93220 123076 93226
rect 123024 93162 123076 93168
rect 119712 93152 119764 93158
rect 119712 93094 119764 93100
rect 134432 92472 134484 92478
rect 108578 92440 108634 92449
rect 108578 92375 108634 92384
rect 116766 92440 116822 92449
rect 116766 92375 116822 92384
rect 124126 92440 124182 92449
rect 124126 92375 124182 92384
rect 134430 92440 134432 92449
rect 134484 92440 134486 92449
rect 134430 92375 134486 92384
rect 151358 92440 151414 92449
rect 151358 92375 151414 92384
rect 104254 91216 104310 91225
rect 104164 91180 104216 91186
rect 104254 91151 104310 91160
rect 104806 91216 104862 91225
rect 104806 91151 104862 91160
rect 105542 91216 105598 91225
rect 105542 91151 105598 91160
rect 106186 91216 106242 91225
rect 106186 91151 106242 91160
rect 107474 91216 107530 91225
rect 107474 91151 107530 91160
rect 108486 91216 108542 91225
rect 108486 91151 108542 91160
rect 104164 91122 104216 91128
rect 104176 64870 104204 91122
rect 104268 88233 104296 91151
rect 104254 88224 104310 88233
rect 104254 88159 104310 88168
rect 104164 64864 104216 64870
rect 104164 64806 104216 64812
rect 103428 59356 103480 59362
rect 103428 59298 103480 59304
rect 104820 57934 104848 91151
rect 105556 85377 105584 91151
rect 105542 85368 105598 85377
rect 105542 85303 105598 85312
rect 106200 82657 106228 91151
rect 106924 90364 106976 90370
rect 106924 90306 106976 90312
rect 106186 82648 106242 82657
rect 106186 82583 106242 82592
rect 106186 82104 106242 82113
rect 106186 82039 106242 82048
rect 104808 57928 104860 57934
rect 104808 57870 104860 57876
rect 102048 54528 102100 54534
rect 102048 54470 102100 54476
rect 99288 28348 99340 28354
rect 99288 28290 99340 28296
rect 98642 18592 98698 18601
rect 98642 18527 98698 18536
rect 99300 3534 99328 28290
rect 100668 14476 100720 14482
rect 100668 14418 100720 14424
rect 100680 3534 100708 14418
rect 102060 3534 102088 54470
rect 104808 51740 104860 51746
rect 104808 51682 104860 51688
rect 103426 24168 103482 24177
rect 103426 24103 103482 24112
rect 103440 6914 103468 24103
rect 104820 6914 104848 51682
rect 103348 6886 103468 6914
rect 104544 6886 104848 6914
rect 97448 3528 97500 3534
rect 97448 3470 97500 3476
rect 97908 3528 97960 3534
rect 97908 3470 97960 3476
rect 98644 3528 98696 3534
rect 98644 3470 98696 3476
rect 99288 3528 99340 3534
rect 99288 3470 99340 3476
rect 99840 3528 99892 3534
rect 99840 3470 99892 3476
rect 100668 3528 100720 3534
rect 100668 3470 100720 3476
rect 101036 3528 101088 3534
rect 101036 3470 101088 3476
rect 102048 3528 102100 3534
rect 102048 3470 102100 3476
rect 97460 480 97488 3470
rect 98656 480 98684 3470
rect 99852 480 99880 3470
rect 101048 480 101076 3470
rect 102232 3460 102284 3466
rect 102232 3402 102284 3408
rect 102244 480 102272 3402
rect 103348 480 103376 6886
rect 104544 480 104572 6886
rect 106200 3534 106228 82039
rect 106936 73166 106964 90306
rect 106924 73160 106976 73166
rect 106924 73102 106976 73108
rect 107488 55214 107516 91151
rect 108304 91112 108356 91118
rect 108304 91054 108356 91060
rect 107566 78024 107622 78033
rect 107566 77959 107622 77968
rect 107476 55208 107528 55214
rect 107476 55150 107528 55156
rect 107580 3534 107608 77959
rect 108316 63510 108344 91054
rect 108500 86970 108528 91151
rect 108592 91118 108620 92375
rect 110142 91760 110198 91769
rect 110142 91695 110198 91704
rect 108580 91112 108632 91118
rect 108580 91054 108632 91060
rect 110156 89729 110184 91695
rect 111706 91352 111762 91361
rect 111706 91287 111762 91296
rect 114374 91352 114430 91361
rect 114374 91287 114430 91296
rect 115478 91352 115534 91361
rect 115478 91287 115534 91296
rect 115754 91352 115810 91361
rect 115754 91287 115810 91296
rect 110326 91216 110382 91225
rect 110326 91151 110382 91160
rect 111614 91216 111670 91225
rect 111614 91151 111670 91160
rect 110142 89720 110198 89729
rect 110142 89655 110198 89664
rect 108488 86964 108540 86970
rect 108488 86906 108540 86912
rect 108304 63504 108356 63510
rect 108304 63446 108356 63452
rect 110340 51066 110368 91151
rect 111628 80034 111656 91151
rect 111616 80028 111668 80034
rect 111616 79970 111668 79976
rect 111720 62082 111748 91287
rect 112994 91216 113050 91225
rect 112994 91151 113050 91160
rect 111708 62076 111760 62082
rect 111708 62018 111760 62024
rect 113008 56574 113036 91151
rect 114388 84114 114416 91287
rect 114466 91216 114522 91225
rect 114466 91151 114522 91160
rect 114376 84108 114428 84114
rect 114376 84050 114428 84056
rect 113086 80880 113142 80889
rect 113086 80815 113142 80824
rect 112996 56568 113048 56574
rect 112996 56510 113048 56516
rect 110328 51060 110380 51066
rect 110328 51002 110380 51008
rect 108948 50380 109000 50386
rect 108948 50322 109000 50328
rect 108960 3534 108988 50322
rect 111708 49020 111760 49026
rect 111708 48962 111760 48968
rect 109316 4820 109368 4826
rect 109316 4762 109368 4768
rect 105728 3528 105780 3534
rect 105728 3470 105780 3476
rect 106188 3528 106240 3534
rect 106188 3470 106240 3476
rect 106924 3528 106976 3534
rect 106924 3470 106976 3476
rect 107568 3528 107620 3534
rect 107568 3470 107620 3476
rect 108120 3528 108172 3534
rect 108120 3470 108172 3476
rect 108948 3528 109000 3534
rect 108948 3470 109000 3476
rect 105740 480 105768 3470
rect 106936 480 106964 3470
rect 108132 480 108160 3470
rect 109328 480 109356 4762
rect 111720 3534 111748 48962
rect 113100 6914 113128 80815
rect 114480 73098 114508 91151
rect 115492 87961 115520 91287
rect 115478 87952 115534 87961
rect 115478 87887 115534 87896
rect 115204 87644 115256 87650
rect 115204 87586 115256 87592
rect 114468 73092 114520 73098
rect 114468 73034 114520 73040
rect 115216 66230 115244 87586
rect 115768 85542 115796 91287
rect 115846 91216 115902 91225
rect 115846 91151 115902 91160
rect 115756 85536 115808 85542
rect 115756 85478 115808 85484
rect 115296 84856 115348 84862
rect 115296 84798 115348 84804
rect 115308 74497 115336 84798
rect 115294 74488 115350 74497
rect 115294 74423 115350 74432
rect 115204 66224 115256 66230
rect 115204 66166 115256 66172
rect 115860 52426 115888 91151
rect 116780 91118 116808 92375
rect 121182 91760 121238 91769
rect 121182 91695 121238 91704
rect 117134 91216 117190 91225
rect 117134 91151 117190 91160
rect 118606 91216 118662 91225
rect 118606 91151 118662 91160
rect 119986 91216 120042 91225
rect 119986 91151 120042 91160
rect 116584 91112 116636 91118
rect 116584 91054 116636 91060
rect 116768 91112 116820 91118
rect 116768 91054 116820 91060
rect 116596 67561 116624 91054
rect 117148 88330 117176 91151
rect 117136 88324 117188 88330
rect 117136 88266 117188 88272
rect 117226 76664 117282 76673
rect 117226 76599 117282 76608
rect 116582 67552 116638 67561
rect 116582 67487 116638 67496
rect 115848 52420 115900 52426
rect 115848 52362 115900 52368
rect 115848 40792 115900 40798
rect 115848 40734 115900 40740
rect 114008 7676 114060 7682
rect 114008 7618 114060 7624
rect 112824 6886 113128 6914
rect 110512 3528 110564 3534
rect 110512 3470 110564 3476
rect 111708 3528 111760 3534
rect 111708 3470 111760 3476
rect 110524 480 110552 3470
rect 111616 2168 111668 2174
rect 111616 2110 111668 2116
rect 111628 480 111656 2110
rect 112824 480 112852 6886
rect 114020 480 114048 7618
rect 115860 3534 115888 40734
rect 117240 3534 117268 76599
rect 118620 71738 118648 91151
rect 120000 81326 120028 91151
rect 121196 89690 121224 91695
rect 121366 91216 121422 91225
rect 121366 91151 121422 91160
rect 121826 91216 121882 91225
rect 121826 91151 121882 91160
rect 122746 91216 122802 91225
rect 122746 91151 122802 91160
rect 124034 91216 124090 91225
rect 124034 91151 124090 91160
rect 121184 89684 121236 89690
rect 121184 89626 121236 89632
rect 119988 81320 120040 81326
rect 119988 81262 120040 81268
rect 118608 71732 118660 71738
rect 118608 71674 118660 71680
rect 119988 69692 120040 69698
rect 119988 69634 120040 69640
rect 118608 29708 118660 29714
rect 118608 29650 118660 29656
rect 118620 3534 118648 29650
rect 119896 3596 119948 3602
rect 119896 3538 119948 3544
rect 115204 3528 115256 3534
rect 115204 3470 115256 3476
rect 115848 3528 115900 3534
rect 115848 3470 115900 3476
rect 116400 3528 116452 3534
rect 116400 3470 116452 3476
rect 117228 3528 117280 3534
rect 117228 3470 117280 3476
rect 117596 3528 117648 3534
rect 117596 3470 117648 3476
rect 118608 3528 118660 3534
rect 118608 3470 118660 3476
rect 118792 3528 118844 3534
rect 118792 3470 118844 3476
rect 115216 480 115244 3470
rect 116412 480 116440 3470
rect 117608 480 117636 3470
rect 118804 480 118832 3470
rect 119908 480 119936 3538
rect 120000 3534 120028 69634
rect 121380 64802 121408 91151
rect 121840 88262 121868 91151
rect 121828 88256 121880 88262
rect 121828 88198 121880 88204
rect 122102 66872 122158 66881
rect 122102 66807 122158 66816
rect 121368 64796 121420 64802
rect 121368 64738 121420 64744
rect 121092 6248 121144 6254
rect 121092 6190 121144 6196
rect 119988 3528 120040 3534
rect 119988 3470 120040 3476
rect 121104 480 121132 6190
rect 122116 3602 122144 66807
rect 122760 66162 122788 91151
rect 124048 78674 124076 91151
rect 124140 90982 124168 92375
rect 136454 91760 136510 91769
rect 136454 91695 136510 91704
rect 126702 91488 126758 91497
rect 126702 91423 126704 91432
rect 126756 91423 126758 91432
rect 129004 91452 129056 91458
rect 126704 91394 126756 91400
rect 129004 91394 129056 91400
rect 125506 91352 125562 91361
rect 125506 91287 125562 91296
rect 126702 91352 126758 91361
rect 126702 91287 126758 91296
rect 125414 91216 125470 91225
rect 125414 91151 125470 91160
rect 124128 90976 124180 90982
rect 124128 90918 124180 90924
rect 124036 78668 124088 78674
rect 124036 78610 124088 78616
rect 122748 66156 122800 66162
rect 122748 66098 122800 66104
rect 125428 53786 125456 91151
rect 125520 79966 125548 91287
rect 125508 79960 125560 79966
rect 125508 79902 125560 79908
rect 126716 68950 126744 91287
rect 126794 91216 126850 91225
rect 126794 91151 126850 91160
rect 128266 91216 128322 91225
rect 128266 91151 128322 91160
rect 126808 84182 126836 91151
rect 126796 84176 126848 84182
rect 126796 84118 126848 84124
rect 126704 68944 126756 68950
rect 126704 68886 126756 68892
rect 125506 68368 125562 68377
rect 125506 68303 125562 68312
rect 125416 53780 125468 53786
rect 125416 53722 125468 53728
rect 122748 36644 122800 36650
rect 122748 36586 122800 36592
rect 122104 3596 122156 3602
rect 122104 3538 122156 3544
rect 122760 3534 122788 36586
rect 124128 18692 124180 18698
rect 124128 18634 124180 18640
rect 124140 3534 124168 18634
rect 125520 3534 125548 68303
rect 128280 49706 128308 91151
rect 129016 70378 129044 91394
rect 129646 91216 129702 91225
rect 129646 91151 129702 91160
rect 132406 91216 132462 91225
rect 132406 91151 132462 91160
rect 133788 91180 133840 91186
rect 129660 74526 129688 91151
rect 132420 77178 132448 91151
rect 133788 91122 133840 91128
rect 133800 86601 133828 91122
rect 136468 89457 136496 91695
rect 151372 91118 151400 92375
rect 151542 91352 151598 91361
rect 151542 91287 151598 91296
rect 151360 91112 151412 91118
rect 151360 91054 151412 91060
rect 136454 89448 136510 89457
rect 136454 89383 136510 89392
rect 133786 86592 133842 86601
rect 133786 86527 133842 86536
rect 132408 77172 132460 77178
rect 132408 77114 132460 77120
rect 151556 75818 151584 91287
rect 151726 91216 151782 91225
rect 151726 91151 151782 91160
rect 152462 91216 152518 91225
rect 152462 91151 152518 91160
rect 151740 85474 151768 91151
rect 152476 86902 152504 91151
rect 153212 90953 153240 93842
rect 162044 93826 162164 93854
rect 158720 91112 158772 91118
rect 158720 91054 158772 91060
rect 153198 90944 153254 90953
rect 153198 90879 153254 90888
rect 158732 89622 158760 91054
rect 161938 90400 161994 90409
rect 161938 90335 161994 90344
rect 158720 89616 158772 89622
rect 158720 89558 158772 89564
rect 161952 88097 161980 90335
rect 161938 88088 161994 88097
rect 161938 88023 161994 88032
rect 152464 86896 152516 86902
rect 152464 86838 152516 86844
rect 151728 85468 151780 85474
rect 151728 85410 151780 85416
rect 162044 85241 162072 93826
rect 162124 91384 162176 91390
rect 162124 91326 162176 91332
rect 162136 89457 162164 91326
rect 162872 90953 162900 94415
rect 162858 90944 162914 90953
rect 162858 90879 162914 90888
rect 162122 89448 162178 89457
rect 162122 89383 162178 89392
rect 162030 85232 162086 85241
rect 162030 85167 162086 85176
rect 164896 82822 164924 97990
rect 164988 87961 165016 101351
rect 165528 96688 165580 96694
rect 165528 96630 165580 96636
rect 165540 95033 165568 96630
rect 165526 95024 165582 95033
rect 165526 94959 165582 94968
rect 164974 87952 165030 87961
rect 164974 87887 165030 87896
rect 164884 82816 164936 82822
rect 164884 82758 164936 82764
rect 160836 82136 160888 82142
rect 160836 82078 160888 82084
rect 151544 75812 151596 75818
rect 151544 75754 151596 75760
rect 129648 74520 129700 74526
rect 129648 74462 129700 74468
rect 160848 74458 160876 82078
rect 166276 78674 166304 104110
rect 166368 85474 166396 153206
rect 167644 144968 167696 144974
rect 167644 144910 167696 144916
rect 166448 126268 166500 126274
rect 166448 126210 166500 126216
rect 166460 92478 166488 126210
rect 166540 110492 166592 110498
rect 166540 110434 166592 110440
rect 166448 92472 166500 92478
rect 166448 92414 166500 92420
rect 166552 86737 166580 110434
rect 167656 93974 167684 144910
rect 167736 135924 167788 135930
rect 167736 135866 167788 135872
rect 167748 108769 167776 135866
rect 169036 131753 169064 186895
rect 170416 184249 170444 269758
rect 170508 261594 170536 356759
rect 170588 334008 170640 334014
rect 170588 333950 170640 333956
rect 170600 319462 170628 333950
rect 170588 319456 170640 319462
rect 170588 319398 170640 319404
rect 170586 294536 170642 294545
rect 170586 294471 170642 294480
rect 170600 268433 170628 294471
rect 170586 268424 170642 268433
rect 170586 268359 170642 268368
rect 170496 261588 170548 261594
rect 170496 261530 170548 261536
rect 170956 259480 171008 259486
rect 170956 259422 171008 259428
rect 170588 254652 170640 254658
rect 170588 254594 170640 254600
rect 170494 254008 170550 254017
rect 170494 253943 170550 253952
rect 170508 197334 170536 253943
rect 170600 240174 170628 254594
rect 170968 240961 170996 259422
rect 171060 254017 171088 477498
rect 172242 455424 172298 455433
rect 172440 455394 172468 538834
rect 173164 525088 173216 525094
rect 173164 525030 173216 525036
rect 172242 455359 172244 455368
rect 172296 455359 172298 455368
rect 172428 455388 172480 455394
rect 172244 455330 172296 455336
rect 172428 455330 172480 455336
rect 171782 450120 171838 450129
rect 171782 450055 171838 450064
rect 171140 380928 171192 380934
rect 171140 380870 171192 380876
rect 171152 259486 171180 380870
rect 171796 306513 171824 450055
rect 171876 387184 171928 387190
rect 171876 387126 171928 387132
rect 171888 380934 171916 387126
rect 171876 380928 171928 380934
rect 171876 380870 171928 380876
rect 172518 373280 172574 373289
rect 172518 373215 172574 373224
rect 171874 349752 171930 349761
rect 171874 349687 171930 349696
rect 171782 306504 171838 306513
rect 171782 306439 171838 306448
rect 171796 280158 171824 306439
rect 171784 280152 171836 280158
rect 171784 280094 171836 280100
rect 171230 275224 171286 275233
rect 171230 275159 171286 275168
rect 171244 267734 171272 275159
rect 171244 267706 171364 267734
rect 171140 259480 171192 259486
rect 171140 259422 171192 259428
rect 171046 254008 171102 254017
rect 171046 253943 171102 253952
rect 171138 247072 171194 247081
rect 171138 247007 171194 247016
rect 170954 240952 171010 240961
rect 170954 240887 171010 240896
rect 170588 240168 170640 240174
rect 170588 240110 170640 240116
rect 171152 227361 171180 247007
rect 171336 243574 171364 267706
rect 171888 245041 171916 349687
rect 172532 275913 172560 373215
rect 172612 329792 172664 329798
rect 172612 329734 172664 329740
rect 172624 314673 172652 329734
rect 173176 317558 173204 525030
rect 173256 455388 173308 455394
rect 173256 455330 173308 455336
rect 173268 329798 173296 455330
rect 173820 353297 173848 557495
rect 180248 550724 180300 550730
rect 180248 550666 180300 550672
rect 182088 550724 182140 550730
rect 182088 550666 182140 550672
rect 177394 549536 177450 549545
rect 177394 549471 177450 549480
rect 175924 542496 175976 542502
rect 175924 542438 175976 542444
rect 175094 532536 175150 532545
rect 175094 532471 175150 532480
rect 175002 384296 175058 384305
rect 175002 384231 175058 384240
rect 175016 383761 175044 384231
rect 175002 383752 175058 383761
rect 175002 383687 175058 383696
rect 174542 353424 174598 353433
rect 174542 353359 174598 353368
rect 173806 353288 173862 353297
rect 173806 353223 173862 353232
rect 173820 352617 173848 353223
rect 173806 352608 173862 352617
rect 173806 352543 173862 352552
rect 173346 350840 173402 350849
rect 173346 350775 173402 350784
rect 173256 329792 173308 329798
rect 173256 329734 173308 329740
rect 173164 317552 173216 317558
rect 173164 317494 173216 317500
rect 172610 314664 172666 314673
rect 172610 314599 172666 314608
rect 173162 285832 173218 285841
rect 173162 285767 173218 285776
rect 172518 275904 172574 275913
rect 172518 275839 172574 275848
rect 172532 275602 172560 275839
rect 172520 275596 172572 275602
rect 172520 275538 172572 275544
rect 172428 269816 172480 269822
rect 172428 269758 172480 269764
rect 172336 258052 172388 258058
rect 172336 257994 172388 258000
rect 172348 250481 172376 257994
rect 172334 250472 172390 250481
rect 172334 250407 172390 250416
rect 171874 245032 171930 245041
rect 171874 244967 171930 244976
rect 172334 244896 172390 244905
rect 172334 244831 172390 244840
rect 171324 243568 171376 243574
rect 171324 243510 171376 243516
rect 171692 243568 171744 243574
rect 171692 243510 171744 243516
rect 171784 243568 171836 243574
rect 172348 243545 172376 244831
rect 171784 243510 171836 243516
rect 172334 243536 172390 243545
rect 171704 243001 171732 243510
rect 171690 242992 171746 243001
rect 171690 242927 171746 242936
rect 171138 227352 171194 227361
rect 171138 227287 171194 227296
rect 171796 222086 171824 243510
rect 172334 243471 172390 243480
rect 172058 227352 172114 227361
rect 172058 227287 172114 227296
rect 171784 222080 171836 222086
rect 171784 222022 171836 222028
rect 170496 197328 170548 197334
rect 170496 197270 170548 197276
rect 170402 184240 170458 184249
rect 170402 184175 170458 184184
rect 169392 183660 169444 183666
rect 169392 183602 169444 183608
rect 169114 180840 169170 180849
rect 169114 180775 169170 180784
rect 169128 155922 169156 180775
rect 169404 177313 169432 183602
rect 170508 182850 170536 197270
rect 170496 182844 170548 182850
rect 170496 182786 170548 182792
rect 170496 182232 170548 182238
rect 170496 182174 170548 182180
rect 169390 177304 169446 177313
rect 169390 177239 169446 177248
rect 169206 176896 169262 176905
rect 169206 176831 169262 176840
rect 169220 168298 169248 176831
rect 170404 176792 170456 176798
rect 170404 176734 170456 176740
rect 169760 175976 169812 175982
rect 169760 175918 169812 175924
rect 169772 172514 169800 175918
rect 169760 172508 169812 172514
rect 169760 172450 169812 172456
rect 169208 168292 169260 168298
rect 169208 168234 169260 168240
rect 170416 158030 170444 176734
rect 170508 169726 170536 182174
rect 171796 173913 171824 222022
rect 171874 210352 171930 210361
rect 171874 210287 171930 210296
rect 171888 200977 171916 210287
rect 171874 200968 171930 200977
rect 171874 200903 171930 200912
rect 172072 198121 172100 227287
rect 172440 217297 172468 269758
rect 173176 227730 173204 285767
rect 173254 279712 173310 279721
rect 173254 279647 173310 279656
rect 173268 250510 173296 279647
rect 173360 267034 173388 350775
rect 173438 273320 173494 273329
rect 173438 273255 173494 273264
rect 173348 267028 173400 267034
rect 173348 266970 173400 266976
rect 173348 265668 173400 265674
rect 173348 265610 173400 265616
rect 173256 250504 173308 250510
rect 173256 250446 173308 250452
rect 173360 243574 173388 265610
rect 173452 258058 173480 273255
rect 174556 262993 174584 353359
rect 175016 318889 175044 383687
rect 175108 362234 175136 532471
rect 175188 514820 175240 514826
rect 175188 514762 175240 514768
rect 175096 362228 175148 362234
rect 175096 362170 175148 362176
rect 175002 318880 175058 318889
rect 175002 318815 175058 318824
rect 175016 316034 175044 318815
rect 174648 316006 175044 316034
rect 174648 305833 174676 316006
rect 175096 314764 175148 314770
rect 175096 314706 175148 314712
rect 174634 305824 174690 305833
rect 174634 305759 174690 305768
rect 174636 291236 174688 291242
rect 174636 291178 174688 291184
rect 174542 262984 174598 262993
rect 174542 262919 174598 262928
rect 173440 258052 173492 258058
rect 173440 257994 173492 258000
rect 173440 249824 173492 249830
rect 173440 249766 173492 249772
rect 173348 243568 173400 243574
rect 173348 243510 173400 243516
rect 173452 229809 173480 249766
rect 174544 234660 174596 234666
rect 174544 234602 174596 234608
rect 173438 229800 173494 229809
rect 173438 229735 173494 229744
rect 173164 227724 173216 227730
rect 173164 227666 173216 227672
rect 172426 217288 172482 217297
rect 172426 217223 172482 217232
rect 171874 198112 171930 198121
rect 171874 198047 171930 198056
rect 172058 198112 172114 198121
rect 172058 198047 172114 198056
rect 171782 173904 171838 173913
rect 171782 173839 171838 173848
rect 170496 169720 170548 169726
rect 170496 169662 170548 169668
rect 170404 158024 170456 158030
rect 170404 157966 170456 157972
rect 169116 155916 169168 155922
rect 169116 155858 169168 155864
rect 171888 151094 171916 198047
rect 171968 183592 172020 183598
rect 171968 183534 172020 183540
rect 171980 161430 172008 183534
rect 173176 172446 173204 227666
rect 173254 200696 173310 200705
rect 173254 200631 173310 200640
rect 173164 172440 173216 172446
rect 173164 172382 173216 172388
rect 171968 161424 172020 161430
rect 171968 161366 172020 161372
rect 171876 151088 171928 151094
rect 171876 151030 171928 151036
rect 173268 148374 173296 200631
rect 174556 186289 174584 234602
rect 174648 229022 174676 291178
rect 174818 257272 174874 257281
rect 174818 257207 174874 257216
rect 174832 249257 174860 257207
rect 174818 249248 174874 249257
rect 174818 249183 174874 249192
rect 174636 229016 174688 229022
rect 174636 228958 174688 228964
rect 174542 186280 174598 186289
rect 174542 186215 174598 186224
rect 174544 180940 174596 180946
rect 174544 180882 174596 180888
rect 173346 179616 173402 179625
rect 173346 179551 173402 179560
rect 173360 161362 173388 179551
rect 173440 173460 173492 173466
rect 173440 173402 173492 173408
rect 173348 161356 173400 161362
rect 173348 161298 173400 161304
rect 173256 148368 173308 148374
rect 173256 148310 173308 148316
rect 171784 142180 171836 142186
rect 171784 142122 171836 142128
rect 170404 139460 170456 139466
rect 170404 139402 170456 139408
rect 169116 138712 169168 138718
rect 169116 138654 169168 138660
rect 169022 131744 169078 131753
rect 169022 131679 169078 131688
rect 167828 116612 167880 116618
rect 167828 116554 167880 116560
rect 167840 111761 167868 116554
rect 167826 111752 167882 111761
rect 167826 111687 167882 111696
rect 167828 110424 167880 110430
rect 167828 110366 167880 110372
rect 167840 110129 167868 110366
rect 167826 110120 167882 110129
rect 167826 110055 167882 110064
rect 167734 108760 167790 108769
rect 167734 108695 167790 108704
rect 167828 106344 167880 106350
rect 167828 106286 167880 106292
rect 167736 105596 167788 105602
rect 167736 105538 167788 105544
rect 167644 93968 167696 93974
rect 167644 93910 167696 93916
rect 166538 86728 166594 86737
rect 166538 86663 166594 86672
rect 166356 85468 166408 85474
rect 166356 85410 166408 85416
rect 167748 84182 167776 105538
rect 167840 89593 167868 106286
rect 169024 102196 169076 102202
rect 169024 102138 169076 102144
rect 168288 96008 168340 96014
rect 168288 95950 168340 95956
rect 168300 91390 168328 95950
rect 168288 91384 168340 91390
rect 168288 91326 168340 91332
rect 167826 89584 167882 89593
rect 167826 89519 167882 89528
rect 167736 84176 167788 84182
rect 167736 84118 167788 84124
rect 166264 78668 166316 78674
rect 166264 78610 166316 78616
rect 169036 74497 169064 102138
rect 169128 86902 169156 138654
rect 169208 134564 169260 134570
rect 169208 134506 169260 134512
rect 169116 86896 169168 86902
rect 169116 86838 169168 86844
rect 169220 86601 169248 134506
rect 169300 117360 169352 117366
rect 169300 117302 169352 117308
rect 169312 93537 169340 117302
rect 169298 93528 169354 93537
rect 169298 93463 169354 93472
rect 169298 89176 169354 89185
rect 169298 89111 169354 89120
rect 169206 86592 169262 86601
rect 169206 86527 169262 86536
rect 169022 74488 169078 74497
rect 160836 74452 160888 74458
rect 169022 74423 169078 74432
rect 160836 74394 160888 74400
rect 160744 73840 160796 73846
rect 160744 73782 160796 73788
rect 129004 70372 129056 70378
rect 129004 70314 129056 70320
rect 128268 49700 128320 49706
rect 128268 49642 128320 49648
rect 141422 44840 141478 44849
rect 141422 44775 141478 44784
rect 130384 35284 130436 35290
rect 130384 35226 130436 35232
rect 126888 11824 126940 11830
rect 126888 11766 126940 11772
rect 126900 3534 126928 11766
rect 122288 3528 122340 3534
rect 122288 3470 122340 3476
rect 122748 3528 122800 3534
rect 122748 3470 122800 3476
rect 123484 3528 123536 3534
rect 123484 3470 123536 3476
rect 124128 3528 124180 3534
rect 124128 3470 124180 3476
rect 124680 3528 124732 3534
rect 124680 3470 124732 3476
rect 125508 3528 125560 3534
rect 125508 3470 125560 3476
rect 125876 3528 125928 3534
rect 125876 3470 125928 3476
rect 126888 3528 126940 3534
rect 126888 3470 126940 3476
rect 122300 480 122328 3470
rect 123496 480 123524 3470
rect 124692 480 124720 3470
rect 125888 480 125916 3470
rect 130396 3466 130424 35226
rect 135258 18592 135314 18601
rect 135258 18527 135314 18536
rect 133142 15872 133198 15881
rect 133142 15807 133198 15816
rect 132958 3496 133014 3505
rect 130384 3460 130436 3466
rect 132958 3431 133014 3440
rect 130384 3402 130436 3408
rect 129372 2984 129424 2990
rect 129372 2926 129424 2932
rect 129384 480 129412 2926
rect 132972 480 133000 3431
rect 133156 2990 133184 15807
rect 135272 11694 135300 18527
rect 135260 11688 135312 11694
rect 135260 11630 135312 11636
rect 136456 11688 136508 11694
rect 136456 11630 136508 11636
rect 133144 2984 133196 2990
rect 133144 2926 133196 2932
rect 136468 480 136496 11630
rect 141436 3534 141464 44775
rect 144826 39264 144882 39273
rect 144826 39199 144882 39208
rect 144840 3534 144868 39199
rect 160756 26926 160784 73782
rect 169312 69018 169340 89111
rect 169300 69012 169352 69018
rect 169300 68954 169352 68960
rect 170416 66162 170444 139402
rect 170496 120148 170548 120154
rect 170496 120090 170548 120096
rect 170508 88330 170536 120090
rect 170586 105224 170642 105233
rect 170586 105159 170642 105168
rect 170496 88324 170548 88330
rect 170496 88266 170548 88272
rect 170600 75886 170628 105159
rect 170680 101516 170732 101522
rect 170680 101458 170732 101464
rect 170692 81326 170720 101458
rect 170772 87712 170824 87718
rect 170772 87654 170824 87660
rect 170680 81320 170732 81326
rect 170680 81262 170732 81268
rect 170784 77246 170812 87654
rect 170772 77240 170824 77246
rect 170772 77182 170824 77188
rect 170588 75880 170640 75886
rect 170588 75822 170640 75828
rect 171796 70378 171824 142122
rect 171968 124228 172020 124234
rect 171968 124170 172020 124176
rect 171876 122868 171928 122874
rect 171876 122810 171928 122816
rect 171888 88262 171916 122810
rect 171980 93226 172008 124170
rect 173348 111852 173400 111858
rect 173348 111794 173400 111800
rect 173256 107704 173308 107710
rect 173256 107646 173308 107652
rect 172060 104236 172112 104242
rect 172060 104178 172112 104184
rect 171968 93220 172020 93226
rect 171968 93162 172020 93168
rect 171876 88256 171928 88262
rect 171876 88198 171928 88204
rect 172072 80034 172100 104178
rect 173164 95940 173216 95946
rect 173164 95882 173216 95888
rect 172060 80028 172112 80034
rect 172060 79970 172112 79976
rect 171784 70372 171836 70378
rect 171784 70314 171836 70320
rect 170404 66156 170456 66162
rect 170404 66098 170456 66104
rect 173176 64802 173204 95882
rect 173268 81394 173296 107646
rect 173360 94518 173388 111794
rect 173452 100065 173480 173402
rect 174556 150414 174584 180882
rect 174544 150408 174596 150414
rect 174544 150350 174596 150356
rect 174542 119368 174598 119377
rect 174542 119303 174598 119312
rect 173438 100056 173494 100065
rect 173438 99991 173494 100000
rect 173440 98116 173492 98122
rect 173440 98058 173492 98064
rect 173348 94512 173400 94518
rect 173348 94454 173400 94460
rect 173452 84153 173480 98058
rect 173438 84144 173494 84153
rect 173438 84079 173494 84088
rect 173256 81388 173308 81394
rect 173256 81330 173308 81336
rect 174556 73098 174584 119303
rect 174544 73092 174596 73098
rect 174544 73034 174596 73040
rect 173164 64796 173216 64802
rect 173164 64738 173216 64744
rect 160744 26920 160796 26926
rect 160744 26862 160796 26868
rect 175108 19281 175136 314706
rect 175200 210905 175228 514762
rect 175280 329792 175332 329798
rect 175280 329734 175332 329740
rect 175292 297430 175320 329734
rect 175280 297424 175332 297430
rect 175280 297366 175332 297372
rect 175292 297226 175320 297366
rect 175280 297220 175332 297226
rect 175280 297162 175332 297168
rect 175936 267102 175964 542438
rect 177304 534812 177356 534818
rect 177304 534754 177356 534760
rect 176016 530596 176068 530602
rect 176016 530538 176068 530544
rect 176028 345137 176056 530538
rect 177316 353394 177344 534754
rect 177408 522306 177436 549471
rect 180154 545320 180210 545329
rect 180154 545255 180210 545264
rect 178774 537160 178830 537169
rect 178774 537095 178830 537104
rect 177396 522300 177448 522306
rect 177396 522242 177448 522248
rect 178684 495508 178736 495514
rect 178684 495450 178736 495456
rect 177396 474768 177448 474774
rect 177396 474710 177448 474716
rect 177408 391241 177436 474710
rect 177856 396092 177908 396098
rect 177856 396034 177908 396040
rect 177394 391232 177450 391241
rect 177394 391167 177450 391176
rect 177396 359576 177448 359582
rect 177396 359518 177448 359524
rect 177304 353388 177356 353394
rect 177304 353330 177356 353336
rect 176200 349240 176252 349246
rect 176200 349182 176252 349188
rect 176014 345128 176070 345137
rect 176014 345063 176070 345072
rect 176028 319530 176056 345063
rect 176108 336796 176160 336802
rect 176108 336738 176160 336744
rect 176016 319524 176068 319530
rect 176016 319466 176068 319472
rect 176016 297220 176068 297226
rect 176016 297162 176068 297168
rect 175924 267096 175976 267102
rect 175924 267038 175976 267044
rect 175924 261520 175976 261526
rect 175924 261462 175976 261468
rect 175936 229022 175964 261462
rect 175924 229016 175976 229022
rect 175924 228958 175976 228964
rect 176028 227361 176056 297162
rect 176120 273970 176148 336738
rect 176212 329186 176240 349182
rect 176658 345944 176714 345953
rect 176658 345879 176714 345888
rect 176672 345681 176700 345879
rect 176658 345672 176714 345681
rect 176658 345607 176714 345616
rect 176200 329180 176252 329186
rect 176200 329122 176252 329128
rect 177316 311137 177344 353330
rect 177408 331974 177436 359518
rect 177868 345953 177896 396034
rect 178040 387116 178092 387122
rect 178040 387058 178092 387064
rect 177946 373280 178002 373289
rect 177946 373215 178002 373224
rect 177854 345944 177910 345953
rect 177854 345879 177910 345888
rect 177486 338328 177542 338337
rect 177486 338263 177542 338272
rect 177396 331968 177448 331974
rect 177396 331910 177448 331916
rect 177302 311128 177358 311137
rect 177302 311063 177358 311072
rect 177500 310593 177528 338263
rect 177486 310584 177542 310593
rect 177486 310519 177542 310528
rect 177854 310584 177910 310593
rect 177854 310519 177910 310528
rect 177304 309800 177356 309806
rect 177304 309742 177356 309748
rect 176934 309088 176990 309097
rect 176934 309023 176990 309032
rect 176948 308417 176976 309023
rect 176934 308408 176990 308417
rect 176934 308343 176990 308352
rect 176200 279472 176252 279478
rect 176200 279414 176252 279420
rect 176108 273964 176160 273970
rect 176108 273906 176160 273912
rect 176212 233986 176240 279414
rect 176566 272504 176622 272513
rect 176566 272439 176622 272448
rect 176580 271969 176608 272439
rect 176566 271960 176622 271969
rect 176566 271895 176622 271904
rect 176200 233980 176252 233986
rect 176200 233922 176252 233928
rect 176014 227352 176070 227361
rect 176014 227287 176070 227296
rect 175186 210896 175242 210905
rect 175186 210831 175242 210840
rect 175924 189100 175976 189106
rect 175924 189042 175976 189048
rect 175936 162790 175964 189042
rect 176016 186380 176068 186386
rect 176016 186322 176068 186328
rect 176028 175166 176056 186322
rect 176016 175160 176068 175166
rect 176016 175102 176068 175108
rect 175924 162784 175976 162790
rect 175924 162726 175976 162732
rect 175924 121508 175976 121514
rect 175924 121450 175976 121456
rect 175936 93158 175964 121450
rect 176016 100768 176068 100774
rect 176016 100710 176068 100716
rect 175924 93152 175976 93158
rect 175924 93094 175976 93100
rect 176028 77178 176056 100710
rect 176016 77172 176068 77178
rect 176016 77114 176068 77120
rect 176580 30297 176608 271895
rect 177316 254561 177344 309742
rect 177486 269784 177542 269793
rect 177486 269719 177542 269728
rect 177396 255332 177448 255338
rect 177396 255274 177448 255280
rect 177302 254552 177358 254561
rect 177302 254487 177358 254496
rect 177304 250980 177356 250986
rect 177304 250922 177356 250928
rect 177316 234433 177344 250922
rect 177302 234424 177358 234433
rect 177302 234359 177358 234368
rect 176658 234288 176714 234297
rect 176658 234223 176714 234232
rect 176672 233918 176700 234223
rect 176660 233912 176712 233918
rect 176660 233854 176712 233860
rect 177316 189854 177344 234359
rect 177408 223417 177436 255274
rect 177500 243574 177528 269719
rect 177868 265033 177896 310519
rect 177960 308417 177988 373215
rect 177946 308408 178002 308417
rect 177946 308343 178002 308352
rect 177948 297424 178000 297430
rect 177948 297366 178000 297372
rect 177854 265024 177910 265033
rect 177854 264959 177910 264968
rect 177488 243568 177540 243574
rect 177488 243510 177540 243516
rect 177960 234297 177988 297366
rect 178052 295089 178080 387058
rect 178132 380180 178184 380186
rect 178132 380122 178184 380128
rect 178144 379642 178172 380122
rect 178132 379636 178184 379642
rect 178132 379578 178184 379584
rect 178696 347041 178724 495450
rect 178788 421598 178816 537095
rect 180064 534744 180116 534750
rect 180064 534686 180116 534692
rect 180076 476066 180104 534686
rect 180168 511290 180196 545255
rect 180260 528562 180288 550666
rect 180248 528556 180300 528562
rect 180248 528498 180300 528504
rect 180248 516180 180300 516186
rect 180248 516122 180300 516128
rect 180156 511284 180208 511290
rect 180156 511226 180208 511232
rect 180260 498846 180288 516122
rect 180248 498840 180300 498846
rect 180248 498782 180300 498788
rect 180156 496868 180208 496874
rect 180156 496810 180208 496816
rect 180064 476060 180116 476066
rect 180064 476002 180116 476008
rect 180064 438932 180116 438938
rect 180064 438874 180116 438880
rect 178776 421592 178828 421598
rect 178776 421534 178828 421540
rect 178776 379636 178828 379642
rect 178776 379578 178828 379584
rect 178682 347032 178738 347041
rect 178682 346967 178738 346976
rect 178682 345672 178738 345681
rect 178682 345607 178738 345616
rect 178696 314770 178724 345607
rect 178684 314764 178736 314770
rect 178684 314706 178736 314712
rect 178684 313948 178736 313954
rect 178684 313890 178736 313896
rect 178038 295080 178094 295089
rect 178038 295015 178094 295024
rect 178052 294642 178080 295015
rect 178040 294636 178092 294642
rect 178040 294578 178092 294584
rect 178696 273329 178724 313890
rect 178682 273320 178738 273329
rect 178682 273255 178738 273264
rect 178684 269884 178736 269890
rect 178684 269826 178736 269832
rect 178696 269142 178724 269826
rect 178684 269136 178736 269142
rect 178684 269078 178736 269084
rect 178040 269000 178092 269006
rect 178040 268942 178092 268948
rect 178052 268394 178080 268942
rect 178040 268388 178092 268394
rect 178040 268330 178092 268336
rect 177946 234288 178002 234297
rect 177946 234223 178002 234232
rect 177946 224360 178002 224369
rect 177946 224295 178002 224304
rect 177394 223408 177450 223417
rect 177394 223343 177450 223352
rect 177856 217184 177908 217190
rect 177856 217126 177908 217132
rect 177304 189848 177356 189854
rect 177304 189790 177356 189796
rect 177304 187740 177356 187746
rect 177304 187682 177356 187688
rect 177316 173194 177344 187682
rect 177868 184278 177896 217126
rect 177960 187066 177988 224295
rect 178040 224256 178092 224262
rect 178040 224198 178092 224204
rect 178052 223689 178080 224198
rect 178038 223680 178094 223689
rect 178038 223615 178094 223624
rect 178696 203561 178724 269078
rect 178788 269006 178816 379578
rect 178866 278760 178922 278769
rect 178866 278695 178922 278704
rect 178776 269000 178828 269006
rect 178776 268942 178828 268948
rect 178776 249824 178828 249830
rect 178776 249766 178828 249772
rect 178788 217190 178816 249766
rect 178880 232937 178908 278695
rect 179328 267096 179380 267102
rect 179328 267038 179380 267044
rect 179340 241913 179368 267038
rect 179420 253224 179472 253230
rect 179420 253166 179472 253172
rect 179432 252550 179460 253166
rect 179420 252544 179472 252550
rect 179420 252486 179472 252492
rect 180076 250986 180104 438874
rect 180168 317393 180196 496810
rect 181628 483676 181680 483682
rect 181628 483618 181680 483624
rect 180248 480276 180300 480282
rect 180248 480218 180300 480224
rect 180260 388482 180288 480218
rect 181444 418192 181496 418198
rect 181444 418134 181496 418140
rect 180248 388476 180300 388482
rect 180248 388418 180300 388424
rect 180340 387116 180392 387122
rect 180340 387058 180392 387064
rect 180246 352608 180302 352617
rect 180246 352543 180302 352552
rect 180154 317384 180210 317393
rect 180154 317319 180210 317328
rect 180156 313336 180208 313342
rect 180156 313278 180208 313284
rect 180168 278118 180196 313278
rect 180156 278112 180208 278118
rect 180156 278054 180208 278060
rect 180156 274712 180208 274718
rect 180156 274654 180208 274660
rect 180168 262886 180196 274654
rect 180156 262880 180208 262886
rect 180156 262822 180208 262828
rect 180260 259457 180288 352543
rect 180352 347857 180380 387058
rect 180338 347848 180394 347857
rect 180338 347783 180394 347792
rect 180352 305017 180380 347783
rect 180338 305008 180394 305017
rect 180338 304943 180394 304952
rect 180706 305008 180762 305017
rect 180706 304943 180762 304952
rect 180720 273222 180748 304943
rect 180708 273216 180760 273222
rect 180708 273158 180760 273164
rect 180340 264988 180392 264994
rect 180340 264930 180392 264936
rect 180246 259448 180302 259457
rect 180246 259383 180302 259392
rect 180246 257952 180302 257961
rect 180246 257887 180302 257896
rect 180064 250980 180116 250986
rect 180064 250922 180116 250928
rect 180156 249960 180208 249966
rect 180156 249902 180208 249908
rect 179420 247784 179472 247790
rect 179420 247726 179472 247732
rect 179432 246362 179460 247726
rect 179420 246356 179472 246362
rect 179420 246298 179472 246304
rect 178958 241904 179014 241913
rect 178958 241839 179014 241848
rect 179326 241904 179382 241913
rect 179326 241839 179382 241848
rect 178972 238513 179000 241839
rect 179418 239456 179474 239465
rect 179418 239391 179474 239400
rect 179432 238513 179460 239391
rect 178958 238504 179014 238513
rect 178958 238439 179014 238448
rect 179418 238504 179474 238513
rect 179418 238439 179474 238448
rect 178866 232928 178922 232937
rect 178866 232863 178922 232872
rect 180168 229094 180196 249902
rect 180076 229066 180196 229094
rect 180076 226001 180104 229066
rect 180062 225992 180118 226001
rect 180062 225927 180118 225936
rect 178776 217184 178828 217190
rect 178776 217126 178828 217132
rect 178774 210896 178830 210905
rect 178774 210831 178830 210840
rect 178682 203552 178738 203561
rect 178682 203487 178738 203496
rect 177948 187060 178000 187066
rect 177948 187002 178000 187008
rect 178684 184952 178736 184958
rect 178684 184894 178736 184900
rect 177856 184272 177908 184278
rect 177856 184214 177908 184220
rect 177394 178120 177450 178129
rect 177394 178055 177450 178064
rect 177304 173188 177356 173194
rect 177304 173130 177356 173136
rect 177408 166938 177436 178055
rect 177396 166932 177448 166938
rect 177396 166874 177448 166880
rect 178696 157282 178724 184894
rect 178788 181558 178816 210831
rect 180076 210361 180104 225927
rect 180260 220794 180288 257887
rect 180352 254658 180380 264930
rect 180340 254652 180392 254658
rect 180340 254594 180392 254600
rect 180340 251864 180392 251870
rect 180340 251806 180392 251812
rect 180352 251258 180380 251806
rect 180340 251252 180392 251258
rect 180340 251194 180392 251200
rect 180708 251252 180760 251258
rect 180708 251194 180760 251200
rect 180248 220788 180300 220794
rect 180248 220730 180300 220736
rect 180062 210352 180118 210361
rect 180062 210287 180118 210296
rect 180062 205048 180118 205057
rect 180062 204983 180118 204992
rect 178776 181552 178828 181558
rect 178776 181494 178828 181500
rect 178684 157276 178736 157282
rect 178684 157218 178736 157224
rect 177304 151836 177356 151842
rect 177304 151778 177356 151784
rect 177316 89622 177344 151778
rect 178684 146328 178736 146334
rect 178684 146270 178736 146276
rect 177396 145036 177448 145042
rect 177396 144978 177448 144984
rect 177408 100774 177436 144978
rect 177488 101448 177540 101454
rect 177488 101390 177540 101396
rect 177396 100768 177448 100774
rect 177396 100710 177448 100716
rect 177394 90536 177450 90545
rect 177394 90471 177450 90480
rect 177304 89616 177356 89622
rect 177304 89558 177356 89564
rect 177302 87544 177358 87553
rect 177302 87479 177358 87488
rect 177316 35193 177344 87479
rect 177408 82793 177436 90471
rect 177500 89690 177528 101390
rect 178696 92177 178724 146270
rect 178776 111920 178828 111926
rect 178776 111862 178828 111868
rect 178682 92168 178738 92177
rect 178682 92103 178738 92112
rect 177488 89684 177540 89690
rect 177488 89626 177540 89632
rect 177394 82784 177450 82793
rect 177394 82719 177450 82728
rect 178788 71670 178816 111862
rect 178868 106956 178920 106962
rect 178868 106898 178920 106904
rect 178880 79966 178908 106898
rect 178868 79960 178920 79966
rect 178868 79902 178920 79908
rect 178776 71664 178828 71670
rect 178776 71606 178828 71612
rect 177302 35184 177358 35193
rect 177302 35119 177358 35128
rect 176566 30288 176622 30297
rect 176566 30223 176622 30232
rect 175094 19272 175150 19281
rect 175094 19207 175150 19216
rect 180076 10305 180104 204983
rect 180154 202464 180210 202473
rect 180154 202399 180210 202408
rect 180168 44849 180196 202399
rect 180260 178673 180288 220730
rect 180720 188358 180748 251194
rect 181456 246537 181484 418134
rect 181640 387190 181668 483618
rect 182100 467838 182128 550666
rect 182824 543788 182876 543794
rect 182824 543730 182876 543736
rect 182088 467832 182140 467838
rect 182088 467774 182140 467780
rect 181628 387184 181680 387190
rect 181628 387126 181680 387132
rect 181536 386436 181588 386442
rect 181536 386378 181588 386384
rect 181442 246528 181498 246537
rect 181442 246463 181498 246472
rect 181444 245676 181496 245682
rect 181444 245618 181496 245624
rect 181456 216578 181484 245618
rect 181548 237386 181576 386378
rect 181628 352572 181680 352578
rect 181628 352514 181680 352520
rect 181640 285054 181668 352514
rect 181718 335744 181774 335753
rect 181718 335679 181774 335688
rect 181628 285048 181680 285054
rect 181628 284990 181680 284996
rect 181628 283960 181680 283966
rect 181628 283902 181680 283908
rect 181640 265674 181668 283902
rect 181732 279478 181760 335679
rect 181720 279472 181772 279478
rect 181720 279414 181772 279420
rect 182088 274032 182140 274038
rect 182088 273974 182140 273980
rect 182100 273290 182128 273974
rect 182088 273284 182140 273290
rect 182088 273226 182140 273232
rect 181628 265668 181680 265674
rect 181628 265610 181680 265616
rect 181628 262676 181680 262682
rect 181628 262618 181680 262624
rect 181536 237380 181588 237386
rect 181536 237322 181588 237328
rect 181444 216572 181496 216578
rect 181444 216514 181496 216520
rect 180708 188352 180760 188358
rect 180708 188294 180760 188300
rect 180338 182200 180394 182209
rect 180338 182135 180394 182144
rect 180246 178664 180302 178673
rect 180246 178599 180302 178608
rect 180352 158710 180380 182135
rect 181456 181490 181484 216514
rect 181640 208282 181668 262618
rect 182100 260846 182128 273226
rect 182088 260840 182140 260846
rect 182088 260782 182140 260788
rect 182836 260778 182864 543730
rect 183468 430636 183520 430642
rect 183468 430578 183520 430584
rect 182914 368384 182970 368393
rect 182914 368319 182970 368328
rect 182928 287706 182956 368319
rect 183008 341012 183060 341018
rect 183008 340954 183060 340960
rect 183020 304298 183048 340954
rect 183008 304292 183060 304298
rect 183008 304234 183060 304240
rect 182916 287700 182968 287706
rect 182916 287642 182968 287648
rect 182916 285728 182968 285734
rect 182916 285670 182968 285676
rect 182928 277302 182956 285670
rect 182916 277296 182968 277302
rect 182916 277238 182968 277244
rect 183376 276684 183428 276690
rect 183376 276626 183428 276632
rect 182916 260840 182968 260846
rect 182916 260782 182968 260788
rect 182824 260772 182876 260778
rect 182824 260714 182876 260720
rect 181720 258732 181772 258738
rect 181720 258674 181772 258680
rect 181732 227730 181760 258674
rect 182454 249928 182510 249937
rect 182454 249863 182510 249872
rect 182468 249121 182496 249863
rect 182454 249112 182510 249121
rect 182454 249047 182510 249056
rect 182824 248464 182876 248470
rect 182824 248406 182876 248412
rect 182088 237380 182140 237386
rect 182088 237322 182140 237328
rect 182100 234433 182128 237322
rect 182086 234424 182142 234433
rect 182086 234359 182142 234368
rect 182086 233336 182142 233345
rect 182086 233271 182142 233280
rect 182100 230489 182128 233271
rect 182836 233073 182864 248406
rect 182822 233064 182878 233073
rect 182822 232999 182878 233008
rect 182086 230480 182142 230489
rect 182086 230415 182142 230424
rect 181720 227724 181772 227730
rect 181720 227666 181772 227672
rect 182272 218816 182324 218822
rect 182272 218758 182324 218764
rect 182284 214606 182312 218758
rect 182272 214600 182324 214606
rect 182272 214542 182324 214548
rect 181628 208276 181680 208282
rect 181628 208218 181680 208224
rect 181628 207052 181680 207058
rect 181628 206994 181680 207000
rect 181640 202774 181668 206994
rect 181628 202768 181680 202774
rect 181628 202710 181680 202716
rect 181536 194608 181588 194614
rect 181536 194550 181588 194556
rect 181548 183569 181576 194550
rect 181534 183560 181590 183569
rect 181534 183495 181590 183504
rect 181444 181484 181496 181490
rect 181444 181426 181496 181432
rect 181534 180976 181590 180985
rect 181534 180911 181590 180920
rect 181548 160070 181576 180911
rect 182928 180810 182956 260782
rect 183008 259480 183060 259486
rect 183008 259422 183060 259428
rect 183020 258097 183048 259422
rect 183006 258088 183062 258097
rect 183006 258023 183062 258032
rect 183388 243137 183416 276626
rect 183480 249937 183508 430578
rect 184216 378214 184244 565898
rect 188526 560416 188582 560425
rect 188526 560351 188582 560360
rect 187056 554872 187108 554878
rect 187056 554814 187108 554820
rect 186226 553480 186282 553489
rect 186226 553415 186282 553424
rect 184846 541104 184902 541113
rect 184846 541039 184902 541048
rect 184756 448588 184808 448594
rect 184756 448530 184808 448536
rect 184296 383716 184348 383722
rect 184296 383658 184348 383664
rect 184204 378208 184256 378214
rect 184204 378150 184256 378156
rect 184216 320958 184244 378150
rect 184308 371890 184336 383658
rect 184296 371884 184348 371890
rect 184296 371826 184348 371832
rect 184480 329180 184532 329186
rect 184480 329122 184532 329128
rect 184204 320952 184256 320958
rect 184204 320894 184256 320900
rect 184296 316736 184348 316742
rect 184296 316678 184348 316684
rect 184308 267889 184336 316678
rect 184386 287872 184442 287881
rect 184386 287807 184442 287816
rect 184294 267880 184350 267889
rect 184294 267815 184350 267824
rect 184400 262682 184428 287807
rect 184388 262676 184440 262682
rect 184388 262618 184440 262624
rect 184296 257372 184348 257378
rect 184296 257314 184348 257320
rect 183466 249928 183522 249937
rect 183466 249863 183522 249872
rect 184308 245682 184336 257314
rect 184296 245676 184348 245682
rect 184296 245618 184348 245624
rect 183098 243128 183154 243137
rect 183098 243063 183154 243072
rect 183374 243128 183430 243137
rect 183374 243063 183430 243072
rect 183112 242214 183140 243063
rect 184296 242956 184348 242962
rect 184296 242898 184348 242904
rect 183100 242208 183152 242214
rect 183100 242150 183152 242156
rect 184308 233918 184336 242898
rect 184296 233912 184348 233918
rect 184296 233854 184348 233860
rect 184294 233200 184350 233209
rect 184294 233135 184350 233144
rect 184308 231878 184336 233135
rect 184296 231872 184348 231878
rect 184296 231814 184348 231820
rect 183466 228304 183522 228313
rect 183466 228239 183522 228248
rect 183480 226137 183508 228239
rect 183466 226128 183522 226137
rect 183466 226063 183522 226072
rect 184202 207632 184258 207641
rect 184202 207567 184258 207576
rect 182916 180804 182968 180810
rect 182916 180746 182968 180752
rect 181536 160064 181588 160070
rect 181536 160006 181588 160012
rect 181444 159384 181496 159390
rect 181444 159326 181496 159332
rect 180340 158704 180392 158710
rect 180340 158646 180392 158652
rect 181456 150346 181484 159326
rect 181444 150340 181496 150346
rect 181444 150282 181496 150288
rect 180248 143608 180300 143614
rect 180248 143550 180300 143556
rect 180260 49706 180288 143550
rect 181536 141432 181588 141438
rect 181536 141374 181588 141380
rect 181444 131776 181496 131782
rect 181444 131718 181496 131724
rect 180340 109064 180392 109070
rect 180340 109006 180392 109012
rect 180352 84017 180380 109006
rect 180338 84008 180394 84017
rect 180338 83943 180394 83952
rect 181456 75818 181484 131718
rect 181548 110430 181576 141374
rect 182916 127628 182968 127634
rect 182916 127570 182968 127576
rect 181628 113212 181680 113218
rect 181628 113154 181680 113160
rect 181536 110424 181588 110430
rect 181536 110366 181588 110372
rect 181640 88233 181668 113154
rect 181720 99408 181772 99414
rect 181720 99350 181772 99356
rect 181626 88224 181682 88233
rect 181626 88159 181682 88168
rect 181536 86284 181588 86290
rect 181536 86226 181588 86232
rect 181444 75812 181496 75818
rect 181444 75754 181496 75760
rect 180248 49700 180300 49706
rect 180248 49642 180300 49648
rect 180154 44840 180210 44849
rect 180154 44775 180210 44784
rect 181548 39438 181576 86226
rect 181732 85513 181760 99350
rect 182824 97300 182876 97306
rect 182824 97242 182876 97248
rect 181718 85504 181774 85513
rect 181718 85439 181774 85448
rect 182836 56574 182864 97242
rect 182928 91089 182956 127570
rect 182914 91080 182970 91089
rect 182914 91015 182970 91024
rect 182824 56568 182876 56574
rect 182824 56510 182876 56516
rect 181536 39432 181588 39438
rect 181536 39374 181588 39380
rect 180062 10296 180118 10305
rect 180062 10231 180118 10240
rect 140044 3528 140096 3534
rect 140044 3470 140096 3476
rect 141424 3528 141476 3534
rect 141424 3470 141476 3476
rect 143540 3528 143592 3534
rect 143540 3470 143592 3476
rect 144828 3528 144880 3534
rect 144828 3470 144880 3476
rect 140056 480 140084 3470
rect 143552 480 143580 3470
rect 184216 2689 184244 207567
rect 184308 201113 184336 231814
rect 184492 217938 184520 329122
rect 184768 273329 184796 448530
rect 184860 313177 184888 541039
rect 185582 382528 185638 382537
rect 185582 382463 185638 382472
rect 185596 347070 185624 382463
rect 185584 347064 185636 347070
rect 185584 347006 185636 347012
rect 185582 339688 185638 339697
rect 185582 339623 185638 339632
rect 185596 315353 185624 339623
rect 185582 315344 185638 315353
rect 185582 315279 185638 315288
rect 184846 313168 184902 313177
rect 184846 313103 184902 313112
rect 185582 312624 185638 312633
rect 185582 312559 185638 312568
rect 184754 273320 184810 273329
rect 184754 273255 184810 273264
rect 184848 267028 184900 267034
rect 184848 266970 184900 266976
rect 184860 266422 184888 266970
rect 184848 266416 184900 266422
rect 184848 266358 184900 266364
rect 184756 245676 184808 245682
rect 184756 245618 184808 245624
rect 184768 244905 184796 245618
rect 184754 244896 184810 244905
rect 184754 244831 184810 244840
rect 184756 235272 184808 235278
rect 184756 235214 184808 235220
rect 184480 217932 184532 217938
rect 184480 217874 184532 217880
rect 184294 201104 184350 201113
rect 184294 201039 184350 201048
rect 184294 187232 184350 187241
rect 184294 187167 184350 187176
rect 184308 123457 184336 187167
rect 184768 184210 184796 235214
rect 184756 184204 184808 184210
rect 184756 184146 184808 184152
rect 184860 182918 184888 266358
rect 185596 253230 185624 312559
rect 186240 300898 186268 553415
rect 186964 545148 187016 545154
rect 186964 545090 187016 545096
rect 186976 517478 187004 545090
rect 186964 517472 187016 517478
rect 186964 517414 187016 517420
rect 186964 465112 187016 465118
rect 186964 465054 187016 465060
rect 185768 300892 185820 300898
rect 185768 300834 185820 300840
rect 186228 300892 186280 300898
rect 186228 300834 186280 300840
rect 185674 293992 185730 294001
rect 185674 293927 185730 293936
rect 185688 284986 185716 293927
rect 185676 284980 185728 284986
rect 185676 284922 185728 284928
rect 185676 278112 185728 278118
rect 185676 278054 185728 278060
rect 185584 253224 185636 253230
rect 185584 253166 185636 253172
rect 185584 247104 185636 247110
rect 185584 247046 185636 247052
rect 185596 235278 185624 247046
rect 185688 235890 185716 278054
rect 185780 275330 185808 300834
rect 185768 275324 185820 275330
rect 185768 275266 185820 275272
rect 185766 273320 185822 273329
rect 185766 273255 185822 273264
rect 186226 273320 186282 273329
rect 186226 273255 186282 273264
rect 185780 262138 185808 273255
rect 185768 262132 185820 262138
rect 185768 262074 185820 262080
rect 186240 259418 186268 273255
rect 186976 262206 187004 465054
rect 187068 360262 187096 554814
rect 187608 549296 187660 549302
rect 187608 549238 187660 549244
rect 187148 462392 187200 462398
rect 187148 462334 187200 462340
rect 187160 448526 187188 462334
rect 187148 448520 187200 448526
rect 187148 448462 187200 448468
rect 187146 369064 187202 369073
rect 187146 368999 187202 369008
rect 187056 360256 187108 360262
rect 187056 360198 187108 360204
rect 187068 323610 187096 360198
rect 187056 323604 187108 323610
rect 187056 323546 187108 323552
rect 187160 295322 187188 368999
rect 187620 350441 187648 549238
rect 188436 546508 188488 546514
rect 188436 546450 188488 546456
rect 188342 534984 188398 534993
rect 188342 534919 188398 534928
rect 187698 378312 187754 378321
rect 187698 378247 187754 378256
rect 187712 378146 187740 378247
rect 187700 378140 187752 378146
rect 187700 378082 187752 378088
rect 187606 350432 187662 350441
rect 187606 350367 187662 350376
rect 187620 350033 187648 350367
rect 187606 350024 187662 350033
rect 187606 349959 187662 349968
rect 188356 309806 188384 534919
rect 188448 514758 188476 546450
rect 188540 531282 188568 560351
rect 191104 557592 191156 557598
rect 191104 557534 191156 557540
rect 188620 553512 188672 553518
rect 188620 553454 188672 553460
rect 188632 534070 188660 553454
rect 188620 534064 188672 534070
rect 188620 534006 188672 534012
rect 188528 531276 188580 531282
rect 188528 531218 188580 531224
rect 188436 514752 188488 514758
rect 188436 514694 188488 514700
rect 188436 467832 188488 467838
rect 188436 467774 188488 467780
rect 188448 316062 188476 467774
rect 189724 405748 189776 405754
rect 189724 405690 189776 405696
rect 188988 400444 189040 400450
rect 188988 400386 189040 400392
rect 188528 379568 188580 379574
rect 188528 379510 188580 379516
rect 188540 370530 188568 379510
rect 189000 378321 189028 400386
rect 189080 385076 189132 385082
rect 189080 385018 189132 385024
rect 188986 378312 189042 378321
rect 188986 378247 189042 378256
rect 189092 377466 189120 385018
rect 189170 381032 189226 381041
rect 189170 380967 189226 380976
rect 189080 377460 189132 377466
rect 189080 377402 189132 377408
rect 189184 375193 189212 380967
rect 189170 375184 189226 375193
rect 189170 375119 189226 375128
rect 188528 370524 188580 370530
rect 188528 370466 188580 370472
rect 189078 360360 189134 360369
rect 189078 360295 189134 360304
rect 188526 350024 188582 350033
rect 188526 349959 188582 349968
rect 188540 325106 188568 349959
rect 188528 325100 188580 325106
rect 188528 325042 188580 325048
rect 188436 316056 188488 316062
rect 188436 315998 188488 316004
rect 188448 313954 188476 315998
rect 188436 313948 188488 313954
rect 188436 313890 188488 313896
rect 188528 312588 188580 312594
rect 188528 312530 188580 312536
rect 188344 309800 188396 309806
rect 188344 309742 188396 309748
rect 187608 307080 187660 307086
rect 187608 307022 187660 307028
rect 187620 302433 187648 307022
rect 187606 302424 187662 302433
rect 187606 302359 187662 302368
rect 187148 295316 187200 295322
rect 187148 295258 187200 295264
rect 187240 294024 187292 294030
rect 187240 293966 187292 293972
rect 187056 287088 187108 287094
rect 187056 287030 187108 287036
rect 187068 269074 187096 287030
rect 187252 285734 187280 293966
rect 187240 285728 187292 285734
rect 187240 285670 187292 285676
rect 187620 283121 187648 302359
rect 188436 302320 188488 302326
rect 188436 302262 188488 302268
rect 188344 298852 188396 298858
rect 188344 298794 188396 298800
rect 187606 283112 187662 283121
rect 187606 283047 187662 283056
rect 187514 281480 187570 281489
rect 187514 281415 187570 281424
rect 187056 269068 187108 269074
rect 187056 269010 187108 269016
rect 187056 263628 187108 263634
rect 187056 263570 187108 263576
rect 186320 262200 186372 262206
rect 186320 262142 186372 262148
rect 186964 262200 187016 262206
rect 186964 262142 187016 262148
rect 186332 261497 186360 262142
rect 186318 261488 186374 261497
rect 186318 261423 186374 261432
rect 186228 259412 186280 259418
rect 186228 259354 186280 259360
rect 186228 259276 186280 259282
rect 186228 259218 186280 259224
rect 186240 258126 186268 259218
rect 186228 258120 186280 258126
rect 186228 258062 186280 258068
rect 186136 253224 186188 253230
rect 186136 253166 186188 253172
rect 185676 235884 185728 235890
rect 185676 235826 185728 235832
rect 185584 235272 185636 235278
rect 185584 235214 185636 235220
rect 185582 230344 185638 230353
rect 185582 230279 185638 230288
rect 185596 209001 185624 230279
rect 186148 214713 186176 253166
rect 186240 249762 186268 258062
rect 187068 251870 187096 263570
rect 187424 259412 187476 259418
rect 187424 259354 187476 259360
rect 187436 258194 187464 259354
rect 187424 258188 187476 258194
rect 187424 258130 187476 258136
rect 187056 251864 187108 251870
rect 187056 251806 187108 251812
rect 186228 249756 186280 249762
rect 186228 249698 186280 249704
rect 186228 241528 186280 241534
rect 186228 241470 186280 241476
rect 186134 214704 186190 214713
rect 186134 214639 186190 214648
rect 185582 208992 185638 209001
rect 185582 208927 185638 208936
rect 185584 196648 185636 196654
rect 185584 196590 185636 196596
rect 184848 182912 184900 182918
rect 184848 182854 184900 182860
rect 184386 182336 184442 182345
rect 184386 182271 184442 182280
rect 184400 164218 184428 182271
rect 184388 164212 184440 164218
rect 184388 164154 184440 164160
rect 184388 147688 184440 147694
rect 184388 147630 184440 147636
rect 184294 123448 184350 123457
rect 184294 123383 184350 123392
rect 184296 115252 184348 115258
rect 184296 115194 184348 115200
rect 184308 59362 184336 115194
rect 184400 96014 184428 147630
rect 184388 96008 184440 96014
rect 184388 95950 184440 95956
rect 184296 59356 184348 59362
rect 184296 59298 184348 59304
rect 185596 20641 185624 196590
rect 186240 185706 186268 241470
rect 187436 236706 187464 258130
rect 187424 236700 187476 236706
rect 187424 236642 187476 236648
rect 186964 234660 187016 234666
rect 186964 234602 187016 234608
rect 186320 222896 186372 222902
rect 186320 222838 186372 222844
rect 186332 220794 186360 222838
rect 186320 220788 186372 220794
rect 186320 220730 186372 220736
rect 186976 215286 187004 234602
rect 187056 233980 187108 233986
rect 187056 233922 187108 233928
rect 187068 226302 187096 233922
rect 187422 233200 187478 233209
rect 187422 233135 187478 233144
rect 187436 232558 187464 233135
rect 187424 232552 187476 232558
rect 187424 232494 187476 232500
rect 187056 226296 187108 226302
rect 187056 226238 187108 226244
rect 187528 222873 187556 281415
rect 188356 267102 188384 298794
rect 188448 273329 188476 302262
rect 188540 301510 188568 312530
rect 189092 302326 189120 360295
rect 189080 302320 189132 302326
rect 189080 302262 189132 302268
rect 188528 301504 188580 301510
rect 188528 301446 188580 301452
rect 188434 273320 188490 273329
rect 188434 273255 188490 273264
rect 188436 272536 188488 272542
rect 188436 272478 188488 272484
rect 188344 267096 188396 267102
rect 188344 267038 188396 267044
rect 187608 249076 187660 249082
rect 187608 249018 187660 249024
rect 187620 248470 187648 249018
rect 187608 248464 187660 248470
rect 187608 248406 187660 248412
rect 187514 222864 187570 222873
rect 187514 222799 187570 222808
rect 186964 215280 187016 215286
rect 186964 215222 187016 215228
rect 186228 185700 186280 185706
rect 186228 185642 186280 185648
rect 185768 185020 185820 185026
rect 185768 184962 185820 184968
rect 185674 179480 185730 179489
rect 185674 179415 185730 179424
rect 185688 155854 185716 179415
rect 185780 175982 185808 184962
rect 186976 180033 187004 215222
rect 186962 180024 187018 180033
rect 186962 179959 187018 179968
rect 185768 175976 185820 175982
rect 185768 175918 185820 175924
rect 185676 155848 185728 155854
rect 185676 155790 185728 155796
rect 186964 148368 187016 148374
rect 186964 148310 187016 148316
rect 185676 131164 185728 131170
rect 185676 131106 185728 131112
rect 185688 82657 185716 131106
rect 186976 94625 187004 148310
rect 187148 136672 187200 136678
rect 187148 136614 187200 136620
rect 187056 102264 187108 102270
rect 187056 102206 187108 102212
rect 186962 94616 187018 94625
rect 186962 94551 187018 94560
rect 186962 89040 187018 89049
rect 186962 88975 187018 88984
rect 185674 82648 185730 82657
rect 185674 82583 185730 82592
rect 185582 20632 185638 20641
rect 185582 20567 185638 20576
rect 186976 6225 187004 88975
rect 187068 67590 187096 102206
rect 187160 101425 187188 136614
rect 187146 101416 187202 101425
rect 187146 101351 187202 101360
rect 187620 93838 187648 248406
rect 188342 246528 188398 246537
rect 188342 246463 188398 246472
rect 187608 93832 187660 93838
rect 187608 93774 187660 93780
rect 187056 67584 187108 67590
rect 187056 67526 187108 67532
rect 188356 6769 188384 246463
rect 188448 234666 188476 272478
rect 188712 266484 188764 266490
rect 188712 266426 188764 266432
rect 188620 263696 188672 263702
rect 188620 263638 188672 263644
rect 188528 249756 188580 249762
rect 188528 249698 188580 249704
rect 188436 234660 188488 234666
rect 188436 234602 188488 234608
rect 188434 231840 188490 231849
rect 188434 231775 188490 231784
rect 188448 211857 188476 231775
rect 188434 211848 188490 211857
rect 188434 211783 188490 211792
rect 188434 202328 188490 202337
rect 188434 202263 188490 202272
rect 188448 44849 188476 202263
rect 188540 196722 188568 249698
rect 188632 231849 188660 263638
rect 188724 247722 188752 266426
rect 189078 257000 189134 257009
rect 189078 256935 189134 256944
rect 189092 256766 189120 256935
rect 189080 256760 189132 256766
rect 189080 256702 189132 256708
rect 188712 247716 188764 247722
rect 188712 247658 188764 247664
rect 188618 231840 188674 231849
rect 188618 231775 188674 231784
rect 189736 209710 189764 405690
rect 189814 382392 189870 382401
rect 189814 382327 189870 382336
rect 189828 327826 189856 382327
rect 191116 356289 191144 557534
rect 191654 552120 191710 552129
rect 191654 552055 191710 552064
rect 191196 471300 191248 471306
rect 191196 471242 191248 471248
rect 191208 367554 191236 471242
rect 191288 444032 191340 444038
rect 191288 443974 191340 443980
rect 191300 400450 191328 443974
rect 191288 400444 191340 400450
rect 191288 400386 191340 400392
rect 191288 397520 191340 397526
rect 191288 397462 191340 397468
rect 191300 369238 191328 397462
rect 191288 369232 191340 369238
rect 191288 369174 191340 369180
rect 191208 367526 191328 367554
rect 191300 364410 191328 367526
rect 191288 364404 191340 364410
rect 191288 364346 191340 364352
rect 191196 356856 191248 356862
rect 191196 356798 191248 356804
rect 191102 356280 191158 356289
rect 191102 356215 191158 356224
rect 189906 342544 189962 342553
rect 189906 342479 189962 342488
rect 189920 331945 189948 342479
rect 189906 331936 189962 331945
rect 189906 331871 189962 331880
rect 189816 327820 189868 327826
rect 189816 327762 189868 327768
rect 191116 312730 191144 356215
rect 191104 312724 191156 312730
rect 191104 312666 191156 312672
rect 189908 299600 189960 299606
rect 189908 299542 189960 299548
rect 189814 290592 189870 290601
rect 189814 290527 189870 290536
rect 189828 244934 189856 290527
rect 189920 287026 189948 299542
rect 191208 296070 191236 356798
rect 191300 322318 191328 364346
rect 191668 338745 191696 552055
rect 191760 444038 191788 702646
rect 218992 700330 219020 703520
rect 233884 702772 233936 702778
rect 233884 702714 233936 702720
rect 218980 700324 219032 700330
rect 218980 700266 219032 700272
rect 213920 568608 213972 568614
rect 213920 568550 213972 568556
rect 194600 563168 194652 563174
rect 194600 563110 194652 563116
rect 194508 560312 194560 560318
rect 194508 560254 194560 560260
rect 193956 549364 194008 549370
rect 193956 549306 194008 549312
rect 192484 548004 192536 548010
rect 192484 547946 192536 547952
rect 191748 444032 191800 444038
rect 191748 443974 191800 443980
rect 191748 398948 191800 398954
rect 191748 398890 191800 398896
rect 191760 397526 191788 398890
rect 191748 397520 191800 397526
rect 191748 397462 191800 397468
rect 192496 364334 192524 547946
rect 192574 545456 192630 545465
rect 192574 545391 192630 545400
rect 192588 518129 192616 545391
rect 193968 534818 193996 549306
rect 193956 534812 194008 534818
rect 193956 534754 194008 534760
rect 193864 534132 193916 534138
rect 193864 534074 193916 534080
rect 192574 518120 192630 518129
rect 192574 518055 192630 518064
rect 192576 398880 192628 398886
rect 192576 398822 192628 398828
rect 192588 376718 192616 398822
rect 192758 378176 192814 378185
rect 192758 378111 192814 378120
rect 192576 376712 192628 376718
rect 192576 376654 192628 376660
rect 192668 375420 192720 375426
rect 192668 375362 192720 375368
rect 192496 364306 192616 364334
rect 192588 353569 192616 364306
rect 192574 353560 192630 353569
rect 192574 353495 192630 353504
rect 192482 345944 192538 345953
rect 192482 345879 192538 345888
rect 191654 338736 191710 338745
rect 191654 338671 191710 338680
rect 191380 325712 191432 325718
rect 191380 325654 191432 325660
rect 191288 322312 191340 322318
rect 191288 322254 191340 322260
rect 191288 304360 191340 304366
rect 191288 304302 191340 304308
rect 191196 296064 191248 296070
rect 191196 296006 191248 296012
rect 191194 292632 191250 292641
rect 191194 292567 191250 292576
rect 190000 287156 190052 287162
rect 190000 287098 190052 287104
rect 189908 287020 189960 287026
rect 189908 286962 189960 286968
rect 189908 282260 189960 282266
rect 189908 282202 189960 282208
rect 189920 244934 189948 282202
rect 190012 259282 190040 287098
rect 191104 285796 191156 285802
rect 191104 285738 191156 285744
rect 190460 285048 190512 285054
rect 190460 284990 190512 284996
rect 190472 264897 190500 284990
rect 190458 264888 190514 264897
rect 190458 264823 190514 264832
rect 190000 259276 190052 259282
rect 190000 259218 190052 259224
rect 190274 257000 190330 257009
rect 190274 256935 190330 256944
rect 189816 244928 189868 244934
rect 189816 244870 189868 244876
rect 189908 244928 189960 244934
rect 189908 244870 189960 244876
rect 189816 244248 189868 244254
rect 189816 244190 189868 244196
rect 189828 221921 189856 244190
rect 190288 229945 190316 256935
rect 191116 254590 191144 285738
rect 191208 269822 191236 292567
rect 191300 276690 191328 304302
rect 191392 289134 191420 325654
rect 191380 289128 191432 289134
rect 191380 289070 191432 289076
rect 191748 285048 191800 285054
rect 191748 284990 191800 284996
rect 191760 284889 191788 284990
rect 191746 284880 191802 284889
rect 191746 284815 191802 284824
rect 191288 276684 191340 276690
rect 191288 276626 191340 276632
rect 191564 274780 191616 274786
rect 191564 274722 191616 274728
rect 191196 269816 191248 269822
rect 191196 269758 191248 269764
rect 191104 254584 191156 254590
rect 191104 254526 191156 254532
rect 191470 247072 191526 247081
rect 191470 247007 191526 247016
rect 190458 240952 190514 240961
rect 190458 240887 190514 240896
rect 190366 240816 190422 240825
rect 190366 240751 190422 240760
rect 190274 229936 190330 229945
rect 190274 229871 190330 229880
rect 189814 221912 189870 221921
rect 189814 221847 189870 221856
rect 189724 209704 189776 209710
rect 189724 209646 189776 209652
rect 188528 196716 188580 196722
rect 188528 196658 188580 196664
rect 189722 133920 189778 133929
rect 189722 133855 189778 133864
rect 188528 113280 188580 113286
rect 188528 113222 188580 113228
rect 188540 91050 188568 113222
rect 188528 91044 188580 91050
rect 188528 90986 188580 90992
rect 189736 51066 189764 133855
rect 189828 84182 189856 221847
rect 190380 175817 190408 240751
rect 190472 233170 190500 240887
rect 191484 234190 191512 247007
rect 191576 241505 191604 274722
rect 191748 268184 191800 268190
rect 191748 268126 191800 268132
rect 191760 267889 191788 268126
rect 191746 267880 191802 267889
rect 191746 267815 191802 267824
rect 191654 262984 191710 262993
rect 191654 262919 191710 262928
rect 191562 241496 191618 241505
rect 191562 241431 191618 241440
rect 191472 234184 191524 234190
rect 191472 234126 191524 234132
rect 190460 233164 190512 233170
rect 190460 233106 190512 233112
rect 191104 232552 191156 232558
rect 191104 232494 191156 232500
rect 190366 175808 190422 175817
rect 190366 175743 190422 175752
rect 189908 116000 189960 116006
rect 189908 115942 189960 115948
rect 189920 86970 189948 115942
rect 189908 86964 189960 86970
rect 189908 86906 189960 86912
rect 189816 84176 189868 84182
rect 189816 84118 189868 84124
rect 189724 51060 189776 51066
rect 189724 51002 189776 51008
rect 188434 44840 188490 44849
rect 188434 44775 188490 44784
rect 188342 6760 188398 6769
rect 188342 6695 188398 6704
rect 186962 6216 187018 6225
rect 186962 6151 187018 6160
rect 191116 4146 191144 232494
rect 191668 221513 191696 262919
rect 191654 221504 191710 221513
rect 191654 221439 191710 221448
rect 191760 185745 191788 267815
rect 191838 245712 191894 245721
rect 191838 245647 191840 245656
rect 191892 245647 191894 245656
rect 191840 245618 191892 245624
rect 191930 200832 191986 200841
rect 191930 200767 191986 200776
rect 191944 195974 191972 200767
rect 191932 195968 191984 195974
rect 191932 195910 191984 195916
rect 191746 185736 191802 185745
rect 191746 185671 191802 185680
rect 192496 178945 192524 345879
rect 192588 309126 192616 353495
rect 192680 349858 192708 375362
rect 192772 365022 192800 378111
rect 192760 365016 192812 365022
rect 192760 364958 192812 364964
rect 192668 349852 192720 349858
rect 192668 349794 192720 349800
rect 193036 309936 193088 309942
rect 193036 309878 193088 309884
rect 192576 309120 192628 309126
rect 192576 309062 192628 309068
rect 192944 252612 192996 252618
rect 192944 252554 192996 252560
rect 192668 243568 192720 243574
rect 192668 243510 192720 243516
rect 192680 241777 192708 243510
rect 192666 241768 192722 241777
rect 192666 241703 192722 241712
rect 192666 241632 192722 241641
rect 192666 241567 192722 241576
rect 192680 234569 192708 241567
rect 192666 234560 192722 234569
rect 192666 234495 192722 234504
rect 192576 234184 192628 234190
rect 192576 234126 192628 234132
rect 192482 178936 192538 178945
rect 192482 178871 192538 178880
rect 191194 131744 191250 131753
rect 191194 131679 191250 131688
rect 191208 33862 191236 131679
rect 192588 130422 192616 234126
rect 192956 233238 192984 252554
rect 193048 244254 193076 309878
rect 193876 292641 193904 534074
rect 193956 414044 194008 414050
rect 193956 413986 194008 413992
rect 193862 292632 193918 292641
rect 193862 292567 193918 292576
rect 193968 287881 193996 413986
rect 194520 383654 194548 560254
rect 194612 400926 194640 563110
rect 196624 563100 196676 563106
rect 196624 563042 196676 563048
rect 195888 556300 195940 556306
rect 195888 556242 195940 556248
rect 195334 545184 195390 545193
rect 195334 545119 195390 545128
rect 195242 542464 195298 542473
rect 195242 542399 195298 542408
rect 195256 538898 195284 542399
rect 195244 538892 195296 538898
rect 195244 538834 195296 538840
rect 195348 528554 195376 545119
rect 195796 538348 195848 538354
rect 195796 538290 195848 538296
rect 195256 528526 195376 528554
rect 195256 520946 195284 528526
rect 195244 520940 195296 520946
rect 195244 520882 195296 520888
rect 195244 455456 195296 455462
rect 195244 455398 195296 455404
rect 195256 441454 195284 455398
rect 195808 446457 195836 538290
rect 195794 446448 195850 446457
rect 195794 446383 195850 446392
rect 195336 445800 195388 445806
rect 195336 445742 195388 445748
rect 195348 445058 195376 445742
rect 195336 445052 195388 445058
rect 195336 444994 195388 445000
rect 195244 441448 195296 441454
rect 195244 441390 195296 441396
rect 195796 416832 195848 416838
rect 195796 416774 195848 416780
rect 194600 400920 194652 400926
rect 194600 400862 194652 400868
rect 194612 400246 194640 400862
rect 194600 400240 194652 400246
rect 194600 400182 194652 400188
rect 195244 400240 195296 400246
rect 195244 400182 195296 400188
rect 194428 383626 194548 383654
rect 194428 377534 194456 383626
rect 194508 380996 194560 381002
rect 194508 380938 194560 380944
rect 194416 377528 194468 377534
rect 194416 377470 194468 377476
rect 194140 377460 194192 377466
rect 194140 377402 194192 377408
rect 194152 356794 194180 377402
rect 194520 375329 194548 380938
rect 195256 376009 195284 400182
rect 195334 379536 195390 379545
rect 195334 379471 195390 379480
rect 195242 376000 195298 376009
rect 195242 375935 195298 375944
rect 194506 375320 194562 375329
rect 194506 375255 194562 375264
rect 195348 372609 195376 379471
rect 195428 375488 195480 375494
rect 195428 375430 195480 375436
rect 195334 372600 195390 372609
rect 195334 372535 195390 372544
rect 195440 371929 195468 375430
rect 195426 371920 195482 371929
rect 195426 371855 195482 371864
rect 195334 368520 195390 368529
rect 195334 368455 195390 368464
rect 194874 361856 194930 361865
rect 194874 361791 194930 361800
rect 194140 356788 194192 356794
rect 194140 356730 194192 356736
rect 194888 356697 194916 361791
rect 194046 356688 194102 356697
rect 194046 356623 194102 356632
rect 194874 356688 194930 356697
rect 194874 356623 194930 356632
rect 194060 329798 194088 356623
rect 195244 354000 195296 354006
rect 195244 353942 195296 353948
rect 195256 351218 195284 353942
rect 195348 351218 195376 368455
rect 195244 351212 195296 351218
rect 195244 351154 195296 351160
rect 195336 351212 195388 351218
rect 195336 351154 195388 351160
rect 194048 329792 194100 329798
rect 194048 329734 194100 329740
rect 195152 324964 195204 324970
rect 195152 324906 195204 324912
rect 195164 322250 195192 324906
rect 195152 322244 195204 322250
rect 195152 322186 195204 322192
rect 194048 305040 194100 305046
rect 194048 304982 194100 304988
rect 194060 296002 194088 304982
rect 194048 295996 194100 296002
rect 194048 295938 194100 295944
rect 194416 293276 194468 293282
rect 194416 293218 194468 293224
rect 194048 292664 194100 292670
rect 194048 292606 194100 292612
rect 193954 287872 194010 287881
rect 193954 287807 194010 287816
rect 193128 282192 193180 282198
rect 193128 282134 193180 282140
rect 193036 244248 193088 244254
rect 193036 244190 193088 244196
rect 192944 233232 192996 233238
rect 192944 233174 192996 233180
rect 192956 224942 192984 233174
rect 192944 224936 192996 224942
rect 192944 224878 192996 224884
rect 193140 200870 193168 282134
rect 193864 244316 193916 244322
rect 193864 244258 193916 244264
rect 193876 227497 193904 244258
rect 194060 240689 194088 292606
rect 194230 287464 194286 287473
rect 194230 287399 194286 287408
rect 194244 240825 194272 287399
rect 194428 256698 194456 293218
rect 194508 285864 194560 285870
rect 194508 285806 194560 285812
rect 194520 272377 194548 285806
rect 194506 272368 194562 272377
rect 194506 272303 194562 272312
rect 195150 265568 195206 265577
rect 195150 265503 195206 265512
rect 195164 265033 195192 265503
rect 195150 265024 195206 265033
rect 195150 264959 195206 264968
rect 194508 259820 194560 259826
rect 194508 259762 194560 259768
rect 194416 256692 194468 256698
rect 194416 256634 194468 256640
rect 194428 256018 194456 256634
rect 194416 256012 194468 256018
rect 194416 255954 194468 255960
rect 194416 253972 194468 253978
rect 194416 253914 194468 253920
rect 194428 253201 194456 253914
rect 194414 253192 194470 253201
rect 194414 253127 194470 253136
rect 194322 241496 194378 241505
rect 194322 241431 194378 241440
rect 194230 240816 194286 240825
rect 194230 240751 194286 240760
rect 194046 240680 194102 240689
rect 194046 240615 194102 240624
rect 194336 236774 194364 241431
rect 194324 236768 194376 236774
rect 194324 236710 194376 236716
rect 193954 236600 194010 236609
rect 193954 236535 194010 236544
rect 193862 227488 193918 227497
rect 193862 227423 193918 227432
rect 193968 224262 193996 236535
rect 194414 229800 194470 229809
rect 194414 229735 194470 229744
rect 194428 228449 194456 229735
rect 194414 228440 194470 228449
rect 194414 228375 194470 228384
rect 194324 227044 194376 227050
rect 194324 226986 194376 226992
rect 193956 224256 194008 224262
rect 193956 224198 194008 224204
rect 194336 222154 194364 226986
rect 194324 222148 194376 222154
rect 194324 222090 194376 222096
rect 194416 220108 194468 220114
rect 194416 220050 194468 220056
rect 194428 219366 194456 220050
rect 194416 219360 194468 219366
rect 194416 219302 194468 219308
rect 193862 212528 193918 212537
rect 193862 212463 193918 212472
rect 193128 200864 193180 200870
rect 193128 200806 193180 200812
rect 193126 199472 193182 199481
rect 193126 199407 193182 199416
rect 193140 195906 193168 199407
rect 193128 195900 193180 195906
rect 193128 195842 193180 195848
rect 193876 189786 193904 212463
rect 194324 199504 194376 199510
rect 194324 199446 194376 199452
rect 194336 195906 194364 199446
rect 194324 195900 194376 195906
rect 194324 195842 194376 195848
rect 193864 189780 193916 189786
rect 193864 189722 193916 189728
rect 193864 182912 193916 182918
rect 193864 182854 193916 182860
rect 192668 132524 192720 132530
rect 192668 132466 192720 132472
rect 192576 130416 192628 130422
rect 192576 130358 192628 130364
rect 192680 109721 192708 132466
rect 193876 118017 193904 182854
rect 194520 181393 194548 259762
rect 195256 245721 195284 351154
rect 195336 349172 195388 349178
rect 195336 349114 195388 349120
rect 195348 330546 195376 349114
rect 195518 348392 195574 348401
rect 195518 348327 195574 348336
rect 195532 331906 195560 348327
rect 195428 331900 195480 331906
rect 195428 331842 195480 331848
rect 195520 331900 195572 331906
rect 195520 331842 195572 331848
rect 195336 330540 195388 330546
rect 195336 330482 195388 330488
rect 195440 313954 195468 331842
rect 195428 313948 195480 313954
rect 195428 313890 195480 313896
rect 195336 306400 195388 306406
rect 195336 306342 195388 306348
rect 195348 279410 195376 306342
rect 195428 304292 195480 304298
rect 195428 304234 195480 304240
rect 195336 279404 195388 279410
rect 195336 279346 195388 279352
rect 195348 267734 195376 279346
rect 195440 278662 195468 304234
rect 195428 278656 195480 278662
rect 195428 278598 195480 278604
rect 195440 274786 195468 278598
rect 195428 274780 195480 274786
rect 195428 274722 195480 274728
rect 195348 267706 195744 267734
rect 195336 262268 195388 262274
rect 195336 262210 195388 262216
rect 195348 257689 195376 262210
rect 195428 262132 195480 262138
rect 195428 262074 195480 262080
rect 195440 260953 195468 262074
rect 195426 260944 195482 260953
rect 195426 260879 195482 260888
rect 195334 257680 195390 257689
rect 195334 257615 195390 257624
rect 195612 247172 195664 247178
rect 195612 247114 195664 247120
rect 195242 245712 195298 245721
rect 195242 245647 195298 245656
rect 195244 236700 195296 236706
rect 195244 236642 195296 236648
rect 195256 233986 195284 236642
rect 195244 233980 195296 233986
rect 195244 233922 195296 233928
rect 195242 231296 195298 231305
rect 195242 231231 195298 231240
rect 195256 230382 195284 231231
rect 195244 230376 195296 230382
rect 195244 230318 195296 230324
rect 195244 218068 195296 218074
rect 195244 218010 195296 218016
rect 194506 181384 194562 181393
rect 194506 181319 194562 181328
rect 193956 120216 194008 120222
rect 193956 120158 194008 120164
rect 193862 118008 193918 118017
rect 193862 117943 193918 117952
rect 193864 110560 193916 110566
rect 193864 110502 193916 110508
rect 192666 109712 192722 109721
rect 192666 109647 192722 109656
rect 192484 109132 192536 109138
rect 192484 109074 192536 109080
rect 192496 64870 192524 109074
rect 192574 103864 192630 103873
rect 192574 103799 192630 103808
rect 192588 81433 192616 103799
rect 192574 81424 192630 81433
rect 192574 81359 192630 81368
rect 192484 64864 192536 64870
rect 192484 64806 192536 64812
rect 193876 63510 193904 110502
rect 193968 85542 193996 120158
rect 193956 85536 194008 85542
rect 193956 85478 194008 85484
rect 193864 63504 193916 63510
rect 193864 63446 193916 63452
rect 191196 33856 191248 33862
rect 191196 33798 191248 33804
rect 191104 4140 191156 4146
rect 191104 4082 191156 4088
rect 195256 4049 195284 218010
rect 195624 188601 195652 247114
rect 195716 220726 195744 267706
rect 195808 252550 195836 416774
rect 195900 377641 195928 556242
rect 195980 382968 196032 382974
rect 195980 382910 196032 382916
rect 195886 377632 195942 377641
rect 195886 377567 195942 377576
rect 195992 375358 196020 382910
rect 195980 375352 196032 375358
rect 195980 375294 196032 375300
rect 196636 362982 196664 563042
rect 198464 559020 198516 559026
rect 198464 558962 198516 558968
rect 196716 558952 196768 558958
rect 196716 558894 196768 558900
rect 196728 387122 196756 558894
rect 198096 554804 198148 554810
rect 198096 554746 198148 554752
rect 196806 543960 196862 543969
rect 196806 543895 196862 543904
rect 196820 507142 196848 543895
rect 198004 535628 198056 535634
rect 198004 535570 198056 535576
rect 197358 534576 197414 534585
rect 197358 534511 197414 534520
rect 197372 534138 197400 534511
rect 197360 534132 197412 534138
rect 197360 534074 197412 534080
rect 197360 532704 197412 532710
rect 197360 532646 197412 532652
rect 197372 532273 197400 532646
rect 197358 532264 197414 532273
rect 197358 532199 197414 532208
rect 197360 529916 197412 529922
rect 197360 529858 197412 529864
rect 197372 529825 197400 529858
rect 197358 529816 197414 529825
rect 197358 529751 197414 529760
rect 197360 528556 197412 528562
rect 197360 528498 197412 528504
rect 197372 527377 197400 528498
rect 197358 527368 197414 527377
rect 197358 527303 197414 527312
rect 198016 525094 198044 535570
rect 198004 525088 198056 525094
rect 198004 525030 198056 525036
rect 197358 524784 197414 524793
rect 197358 524719 197414 524728
rect 197372 524482 197400 524719
rect 197360 524476 197412 524482
rect 197360 524418 197412 524424
rect 197358 522336 197414 522345
rect 197358 522271 197414 522280
rect 197372 521694 197400 522271
rect 197360 521688 197412 521694
rect 197360 521630 197412 521636
rect 197358 517440 197414 517449
rect 197358 517375 197414 517384
rect 197372 516186 197400 517375
rect 197360 516180 197412 516186
rect 197360 516122 197412 516128
rect 197358 514992 197414 515001
rect 197358 514927 197414 514936
rect 197372 514826 197400 514927
rect 197360 514820 197412 514826
rect 197360 514762 197412 514768
rect 198002 512544 198058 512553
rect 198002 512479 198058 512488
rect 197360 510604 197412 510610
rect 197360 510546 197412 510552
rect 197372 510241 197400 510546
rect 197358 510232 197414 510241
rect 197358 510167 197414 510176
rect 197358 507648 197414 507657
rect 197358 507583 197414 507592
rect 196808 507136 196860 507142
rect 196808 507078 196860 507084
rect 197372 504422 197400 507583
rect 197360 504416 197412 504422
rect 197360 504358 197412 504364
rect 197358 497856 197414 497865
rect 197358 497791 197414 497800
rect 197372 496874 197400 497791
rect 197360 496868 197412 496874
rect 197360 496810 197412 496816
rect 197358 495544 197414 495553
rect 197358 495479 197360 495488
rect 197412 495479 197414 495488
rect 197360 495450 197412 495456
rect 197358 492960 197414 492969
rect 197358 492895 197414 492904
rect 197372 492726 197400 492895
rect 197360 492720 197412 492726
rect 197360 492662 197412 492668
rect 197360 488504 197412 488510
rect 197360 488446 197412 488452
rect 197372 488209 197400 488446
rect 197358 488200 197414 488209
rect 197358 488135 197414 488144
rect 197358 485616 197414 485625
rect 197358 485551 197414 485560
rect 197372 483682 197400 485551
rect 197360 483676 197412 483682
rect 197360 483618 197412 483624
rect 197358 480720 197414 480729
rect 197358 480655 197414 480664
rect 197372 480282 197400 480655
rect 197360 480276 197412 480282
rect 197360 480218 197412 480224
rect 197358 478272 197414 478281
rect 197358 478207 197414 478216
rect 197372 477562 197400 478207
rect 197360 477556 197412 477562
rect 197360 477498 197412 477504
rect 197358 475824 197414 475833
rect 197358 475759 197414 475768
rect 197372 474774 197400 475759
rect 197360 474768 197412 474774
rect 197360 474710 197412 474716
rect 197360 473408 197412 473414
rect 197358 473376 197360 473385
rect 197412 473376 197414 473385
rect 197358 473311 197414 473320
rect 197266 470928 197322 470937
rect 197266 470863 197322 470872
rect 196716 387116 196768 387122
rect 196716 387058 196768 387064
rect 197174 382528 197230 382537
rect 197174 382463 197230 382472
rect 196808 371272 196860 371278
rect 196808 371214 196860 371220
rect 196624 362976 196676 362982
rect 196624 362918 196676 362924
rect 195980 333260 196032 333266
rect 195980 333202 196032 333208
rect 195992 327758 196020 333202
rect 195980 327752 196032 327758
rect 195980 327694 196032 327700
rect 196636 325038 196664 362918
rect 196714 353968 196770 353977
rect 196714 353903 196770 353912
rect 196624 325032 196676 325038
rect 196624 324974 196676 324980
rect 196624 320884 196676 320890
rect 196624 320826 196676 320832
rect 195980 284980 196032 284986
rect 195980 284922 196032 284928
rect 195992 278050 196020 284922
rect 195980 278044 196032 278050
rect 195980 277986 196032 277992
rect 195980 273964 196032 273970
rect 195980 273906 196032 273912
rect 195992 267734 196020 273906
rect 195992 267706 196112 267734
rect 195978 267200 196034 267209
rect 195978 267135 196034 267144
rect 195992 266490 196020 267135
rect 195980 266484 196032 266490
rect 195980 266426 196032 266432
rect 196084 259826 196112 267706
rect 196072 259820 196124 259826
rect 196072 259762 196124 259768
rect 195796 252544 195848 252550
rect 195796 252486 195848 252492
rect 195808 251666 195836 252486
rect 195796 251660 195848 251666
rect 195796 251602 195848 251608
rect 195704 220720 195756 220726
rect 195704 220662 195756 220668
rect 195808 196654 195836 251602
rect 196636 240553 196664 320826
rect 196728 309874 196756 353903
rect 196820 337414 196848 371214
rect 196808 337408 196860 337414
rect 196808 337350 196860 337356
rect 196716 309868 196768 309874
rect 196716 309810 196768 309816
rect 197188 287337 197216 382463
rect 197280 368490 197308 470863
rect 197358 468480 197414 468489
rect 197358 468415 197414 468424
rect 197372 467906 197400 468415
rect 197360 467900 197412 467906
rect 197360 467842 197412 467848
rect 197358 466032 197414 466041
rect 197358 465967 197414 465976
rect 197372 465118 197400 465967
rect 197360 465112 197412 465118
rect 197360 465054 197412 465060
rect 197358 463312 197414 463321
rect 197358 463247 197414 463256
rect 197372 462398 197400 463247
rect 197360 462392 197412 462398
rect 197360 462334 197412 462340
rect 197358 460864 197414 460873
rect 197358 460799 197414 460808
rect 197372 460222 197400 460799
rect 197360 460216 197412 460222
rect 197360 460158 197412 460164
rect 197358 458416 197414 458425
rect 197358 458351 197414 458360
rect 197372 458250 197400 458351
rect 197360 458244 197412 458250
rect 197360 458186 197412 458192
rect 197358 448624 197414 448633
rect 197358 448559 197360 448568
rect 197412 448559 197414 448568
rect 197360 448530 197412 448536
rect 197358 446176 197414 446185
rect 197358 446111 197414 446120
rect 197372 445806 197400 446111
rect 197360 445800 197412 445806
rect 197360 445742 197412 445748
rect 197360 444032 197412 444038
rect 197360 443974 197412 443980
rect 197372 443873 197400 443974
rect 197358 443864 197414 443873
rect 197358 443799 197414 443808
rect 197728 441448 197780 441454
rect 197726 441416 197728 441425
rect 197780 441416 197782 441425
rect 197726 441351 197782 441360
rect 197358 438968 197414 438977
rect 197358 438903 197360 438912
rect 197412 438903 197414 438912
rect 197360 438874 197412 438880
rect 197358 436384 197414 436393
rect 197358 436319 197414 436328
rect 197372 436150 197400 436319
rect 197360 436144 197412 436150
rect 197360 436086 197412 436092
rect 197358 431488 197414 431497
rect 197358 431423 197414 431432
rect 197372 430642 197400 431423
rect 197360 430636 197412 430642
rect 197360 430578 197412 430584
rect 197358 429040 197414 429049
rect 197358 428975 197414 428984
rect 197372 427854 197400 428975
rect 197360 427848 197412 427854
rect 197360 427790 197412 427796
rect 197358 426592 197414 426601
rect 197358 426527 197414 426536
rect 197372 426494 197400 426527
rect 197360 426488 197412 426494
rect 197360 426430 197412 426436
rect 197358 424144 197414 424153
rect 197358 424079 197414 424088
rect 197372 423706 197400 424079
rect 197360 423700 197412 423706
rect 197360 423642 197412 423648
rect 197358 419248 197414 419257
rect 197358 419183 197414 419192
rect 197372 418198 197400 419183
rect 197360 418192 197412 418198
rect 197360 418134 197412 418140
rect 197360 416832 197412 416838
rect 197358 416800 197360 416809
rect 197412 416800 197414 416809
rect 197358 416735 197414 416744
rect 197358 414352 197414 414361
rect 197358 414287 197414 414296
rect 197372 414050 197400 414287
rect 197360 414044 197412 414050
rect 197360 413986 197412 413992
rect 197358 411904 197414 411913
rect 197358 411839 197414 411848
rect 197372 411330 197400 411839
rect 197360 411324 197412 411330
rect 197360 411266 197412 411272
rect 197360 409828 197412 409834
rect 197360 409770 197412 409776
rect 197372 409601 197400 409770
rect 197358 409592 197414 409601
rect 197358 409527 197414 409536
rect 197358 407008 197414 407017
rect 197358 406943 197414 406952
rect 197372 405754 197400 406943
rect 197360 405748 197412 405754
rect 197360 405690 197412 405696
rect 197358 399664 197414 399673
rect 197358 399599 197414 399608
rect 197372 398954 197400 399599
rect 197360 398948 197412 398954
rect 197360 398890 197412 398896
rect 197358 397216 197414 397225
rect 197358 397151 197414 397160
rect 197372 396098 197400 397151
rect 197360 396092 197412 396098
rect 197360 396034 197412 396040
rect 197358 394768 197414 394777
rect 197358 394703 197360 394712
rect 197412 394703 197414 394712
rect 197360 394674 197412 394680
rect 197358 387424 197414 387433
rect 197358 387359 197414 387368
rect 197372 386442 197400 387359
rect 197360 386436 197412 386442
rect 197360 386378 197412 386384
rect 197358 380080 197414 380089
rect 197358 380015 197414 380024
rect 197372 379642 197400 380015
rect 197360 379636 197412 379642
rect 197360 379578 197412 379584
rect 197268 368484 197320 368490
rect 197268 368426 197320 368432
rect 198016 346633 198044 512479
rect 198108 471306 198136 554746
rect 198280 500948 198332 500954
rect 198280 500890 198332 500896
rect 198292 500449 198320 500890
rect 198278 500440 198334 500449
rect 198278 500375 198334 500384
rect 198096 471300 198148 471306
rect 198096 471242 198148 471248
rect 198476 419665 198504 558962
rect 198648 558204 198700 558210
rect 198648 558146 198700 558152
rect 198660 529825 198688 558146
rect 207662 556200 207718 556209
rect 207662 556135 207718 556144
rect 198830 554024 198886 554033
rect 198830 553959 198886 553968
rect 198740 537532 198792 537538
rect 198740 537474 198792 537480
rect 198752 534750 198780 537474
rect 198740 534744 198792 534750
rect 198740 534686 198792 534692
rect 198646 529816 198702 529825
rect 198646 529751 198702 529760
rect 198738 505200 198794 505209
rect 198738 505135 198794 505144
rect 198554 455968 198610 455977
rect 198554 455903 198610 455912
rect 198462 419656 198518 419665
rect 198462 419591 198518 419600
rect 198462 392320 198518 392329
rect 198462 392255 198518 392264
rect 198002 346624 198058 346633
rect 198002 346559 198058 346568
rect 197358 345128 197414 345137
rect 197358 345063 197360 345072
rect 197412 345063 197414 345072
rect 197360 345034 197412 345040
rect 197266 309768 197322 309777
rect 197266 309703 197322 309712
rect 197174 287328 197230 287337
rect 197174 287263 197230 287272
rect 196716 279472 196768 279478
rect 196716 279414 196768 279420
rect 196728 248742 196756 279414
rect 197280 275913 197308 309703
rect 198016 307834 198044 346559
rect 198004 307828 198056 307834
rect 198004 307770 198056 307776
rect 198016 306374 198044 307770
rect 198016 306346 198412 306374
rect 197358 282432 197414 282441
rect 197358 282367 197414 282376
rect 197372 282198 197400 282367
rect 197360 282192 197412 282198
rect 197360 282134 197412 282140
rect 197358 280256 197414 280265
rect 197358 280191 197360 280200
rect 197412 280191 197414 280200
rect 197360 280162 197412 280168
rect 197358 279440 197414 279449
rect 197358 279375 197360 279384
rect 197412 279375 197414 279384
rect 197360 279346 197412 279352
rect 197360 278656 197412 278662
rect 197358 278624 197360 278633
rect 197412 278624 197414 278633
rect 197358 278559 197414 278568
rect 198384 278089 198412 306346
rect 198370 278080 198426 278089
rect 198370 278015 198426 278024
rect 197360 277364 197412 277370
rect 197360 277306 197412 277312
rect 197372 276729 197400 277306
rect 197358 276720 197414 276729
rect 197358 276655 197414 276664
rect 197266 275904 197322 275913
rect 197266 275839 197322 275848
rect 197358 275088 197414 275097
rect 197358 275023 197414 275032
rect 197372 274718 197400 275023
rect 197360 274712 197412 274718
rect 197360 274654 197412 274660
rect 197450 274544 197506 274553
rect 197450 274479 197506 274488
rect 197464 273290 197492 274479
rect 197452 273284 197504 273290
rect 197452 273226 197504 273232
rect 197360 273216 197412 273222
rect 197360 273158 197412 273164
rect 197372 272921 197400 273158
rect 197358 272912 197414 272921
rect 197358 272847 197414 272856
rect 197358 271552 197414 271561
rect 197358 271487 197414 271496
rect 197372 270638 197400 271487
rect 197360 270632 197412 270638
rect 197360 270574 197412 270580
rect 196808 270564 196860 270570
rect 196808 270506 196860 270512
rect 196820 256766 196848 270506
rect 197358 269376 197414 269385
rect 197358 269311 197414 269320
rect 197372 269142 197400 269311
rect 197360 269136 197412 269142
rect 197360 269078 197412 269084
rect 197360 269000 197412 269006
rect 197360 268942 197412 268948
rect 197372 268025 197400 268942
rect 197450 268832 197506 268841
rect 197450 268767 197506 268776
rect 197464 268190 197492 268767
rect 197452 268184 197504 268190
rect 197452 268126 197504 268132
rect 197358 268016 197414 268025
rect 197358 267951 197414 267960
rect 197358 266656 197414 266665
rect 197358 266591 197414 266600
rect 197372 266422 197400 266591
rect 197360 266416 197412 266422
rect 197360 266358 197412 266364
rect 197450 264480 197506 264489
rect 197450 264415 197506 264424
rect 197464 263702 197492 264415
rect 197452 263696 197504 263702
rect 197358 263664 197414 263673
rect 197452 263638 197504 263644
rect 197358 263599 197360 263608
rect 197412 263599 197414 263608
rect 197360 263570 197412 263576
rect 198002 262304 198058 262313
rect 198002 262239 198004 262248
rect 198056 262239 198058 262248
rect 198004 262210 198056 262216
rect 197360 262200 197412 262206
rect 197360 262142 197412 262148
rect 197372 261497 197400 262142
rect 197358 261488 197414 261497
rect 197358 261423 197414 261432
rect 197358 260128 197414 260137
rect 197358 260063 197414 260072
rect 197268 259820 197320 259826
rect 197268 259762 197320 259768
rect 197280 259298 197308 259762
rect 197372 259486 197400 260063
rect 197360 259480 197412 259486
rect 197360 259422 197412 259428
rect 197358 259312 197414 259321
rect 197280 259270 197358 259298
rect 197358 259247 197414 259256
rect 197358 258768 197414 258777
rect 197358 258703 197414 258712
rect 197372 258194 197400 258703
rect 197360 258188 197412 258194
rect 197360 258130 197412 258136
rect 197358 257408 197414 257417
rect 197280 257366 197358 257394
rect 197280 256766 197308 257366
rect 197358 257343 197414 257352
rect 196808 256760 196860 256766
rect 196808 256702 196860 256708
rect 197268 256760 197320 256766
rect 197268 256702 197320 256708
rect 196808 254652 196860 254658
rect 196808 254594 196860 254600
rect 196716 248736 196768 248742
rect 196716 248678 196768 248684
rect 196728 247178 196756 248678
rect 196716 247172 196768 247178
rect 196716 247114 196768 247120
rect 196716 246356 196768 246362
rect 196716 246298 196768 246304
rect 196622 240544 196678 240553
rect 196622 240479 196678 240488
rect 196622 236736 196678 236745
rect 196622 236671 196678 236680
rect 195796 196648 195848 196654
rect 195796 196590 195848 196596
rect 195610 188592 195666 188601
rect 195610 188527 195666 188536
rect 195428 138032 195480 138038
rect 195428 137974 195480 137980
rect 195336 118720 195388 118726
rect 195336 118662 195388 118668
rect 195348 52426 195376 118662
rect 195440 71738 195468 137974
rect 195520 125656 195572 125662
rect 195520 125598 195572 125604
rect 195532 105602 195560 125598
rect 195520 105596 195572 105602
rect 195520 105538 195572 105544
rect 195428 71732 195480 71738
rect 195428 71674 195480 71680
rect 195336 52420 195388 52426
rect 195336 52362 195388 52368
rect 195242 4040 195298 4049
rect 195242 3975 195298 3984
rect 196636 3913 196664 236671
rect 196728 235958 196756 246298
rect 196820 237318 196848 254594
rect 197174 237960 197230 237969
rect 197174 237895 197230 237904
rect 197188 237425 197216 237895
rect 197174 237416 197230 237425
rect 197174 237351 197230 237360
rect 196808 237312 196860 237318
rect 196808 237254 196860 237260
rect 196716 235952 196768 235958
rect 196716 235894 196768 235900
rect 196714 211168 196770 211177
rect 196714 211103 196770 211112
rect 196728 191826 196756 211103
rect 197188 202162 197216 237351
rect 197176 202156 197228 202162
rect 197176 202098 197228 202104
rect 196808 196716 196860 196722
rect 196808 196658 196860 196664
rect 196716 191820 196768 191826
rect 196716 191762 196768 191768
rect 196820 178702 196848 196658
rect 197280 183025 197308 256702
rect 197360 256692 197412 256698
rect 197360 256634 197412 256640
rect 197372 256601 197400 256634
rect 197358 256592 197414 256601
rect 197358 256527 197414 256536
rect 197358 254416 197414 254425
rect 197358 254351 197414 254360
rect 197372 253978 197400 254351
rect 197360 253972 197412 253978
rect 197360 253914 197412 253920
rect 197358 253600 197414 253609
rect 197358 253535 197414 253544
rect 197372 253230 197400 253535
rect 197360 253224 197412 253230
rect 197360 253166 197412 253172
rect 197358 253056 197414 253065
rect 197358 252991 197414 253000
rect 197372 252618 197400 252991
rect 197360 252612 197412 252618
rect 197360 252554 197412 252560
rect 197358 251696 197414 251705
rect 197358 251631 197360 251640
rect 197412 251631 197414 251640
rect 197360 251602 197412 251608
rect 197450 250880 197506 250889
rect 197450 250815 197506 250824
rect 197358 250064 197414 250073
rect 197358 249999 197414 250008
rect 197372 249898 197400 249999
rect 197360 249892 197412 249898
rect 197360 249834 197412 249840
rect 197464 249830 197492 250815
rect 197452 249824 197504 249830
rect 197452 249766 197504 249772
rect 197358 249520 197414 249529
rect 197358 249455 197414 249464
rect 197372 248470 197400 249455
rect 197820 248736 197872 248742
rect 197818 248704 197820 248713
rect 197872 248704 197874 248713
rect 197818 248639 197874 248648
rect 197360 248464 197412 248470
rect 197360 248406 197412 248412
rect 198476 248414 198504 392255
rect 198568 305046 198596 455903
rect 198646 453520 198702 453529
rect 198646 453455 198702 453464
rect 198556 305040 198608 305046
rect 198556 304982 198608 304988
rect 198568 262857 198596 304982
rect 198660 299538 198688 453455
rect 198752 377330 198780 505135
rect 198844 463321 198872 553959
rect 204904 546576 204956 546582
rect 204904 546518 204956 546524
rect 199384 545216 199436 545222
rect 199384 545158 199436 545164
rect 198830 463312 198886 463321
rect 198830 463247 198886 463256
rect 198830 433936 198886 433945
rect 198830 433871 198886 433880
rect 198740 377324 198792 377330
rect 198740 377266 198792 377272
rect 198752 376786 198780 377266
rect 198740 376780 198792 376786
rect 198740 376722 198792 376728
rect 198844 376038 198872 433871
rect 198832 376032 198884 376038
rect 198832 375974 198884 375980
rect 199396 365838 199424 545158
rect 199476 543856 199528 543862
rect 199476 543798 199528 543804
rect 199488 530602 199516 543798
rect 201406 542736 201462 542745
rect 201406 542671 201462 542680
rect 201314 536072 201370 536081
rect 201314 536007 201370 536016
rect 199750 535936 199806 535945
rect 199750 535871 199806 535880
rect 199764 533361 199792 535871
rect 201328 535634 201356 536007
rect 201420 535945 201448 542671
rect 204074 538656 204130 538665
rect 204074 538591 204130 538600
rect 202786 538520 202842 538529
rect 202786 538455 202842 538464
rect 202800 538354 202828 538455
rect 202788 538348 202840 538354
rect 202788 538290 202840 538296
rect 201406 535936 201462 535945
rect 204088 535908 204116 538591
rect 204168 538280 204220 538286
rect 204166 538248 204168 538257
rect 204220 538248 204222 538257
rect 204166 538183 204222 538192
rect 201406 535871 201462 535880
rect 201316 535628 201368 535634
rect 201316 535570 201368 535576
rect 200394 535528 200450 535537
rect 202050 535528 202106 535537
rect 200450 535486 200790 535514
rect 201408 535492 201460 535498
rect 200394 535463 200450 535472
rect 202106 535486 202446 535514
rect 202050 535463 202106 535472
rect 201408 535434 201460 535440
rect 201420 535401 201448 535434
rect 201406 535392 201462 535401
rect 201406 535327 201462 535336
rect 204916 535294 204944 546518
rect 206282 545456 206338 545465
rect 206282 545391 206338 545400
rect 206296 536897 206324 545391
rect 207676 542337 207704 556135
rect 210424 553444 210476 553450
rect 210424 553386 210476 553392
rect 207018 542328 207074 542337
rect 207018 542263 207074 542272
rect 207662 542328 207718 542337
rect 207662 542263 207718 542272
rect 207032 541249 207060 542263
rect 207018 541240 207074 541249
rect 207018 541175 207074 541184
rect 206282 536888 206338 536897
rect 206282 536823 206338 536832
rect 206296 535922 206324 536823
rect 205758 535894 206324 535922
rect 207032 535922 207060 541175
rect 208400 538280 208452 538286
rect 208400 538222 208452 538228
rect 208412 537538 208440 538222
rect 208400 537532 208452 537538
rect 208400 537474 208452 537480
rect 208674 536072 208730 536081
rect 208674 536007 208730 536016
rect 208688 535922 208716 536007
rect 210436 535922 210464 553386
rect 212540 550656 212592 550662
rect 212540 550598 212592 550604
rect 207032 535894 207414 535922
rect 208688 535894 209070 535922
rect 210436 535894 210910 535922
rect 212552 535908 212580 550598
rect 213932 535922 213960 568550
rect 215300 560380 215352 560386
rect 215300 560322 215352 560328
rect 215312 557534 215340 560322
rect 216678 557560 216734 557569
rect 215312 557506 215432 557534
rect 215404 535922 215432 557506
rect 216734 557506 217088 557534
rect 216678 557495 216734 557504
rect 217060 535922 217088 557506
rect 226984 556232 227036 556238
rect 226984 556174 227036 556180
rect 223672 549364 223724 549370
rect 223672 549306 223724 549312
rect 220820 549296 220872 549302
rect 220820 549238 220872 549244
rect 218702 542736 218758 542745
rect 218702 542671 218758 542680
rect 218716 535922 218744 542671
rect 213932 535894 214222 535922
rect 215404 535894 215878 535922
rect 217060 535894 217534 535922
rect 218716 535894 219190 535922
rect 220832 535908 220860 549238
rect 222474 538520 222530 538529
rect 222474 538455 222530 538464
rect 221096 538348 221148 538354
rect 221096 538290 221148 538296
rect 221108 535401 221136 538290
rect 222488 535908 222516 538455
rect 223684 535922 223712 549306
rect 225326 546680 225382 546689
rect 225326 546615 225382 546624
rect 225340 535922 225368 546615
rect 226996 535922 227024 556174
rect 230478 545320 230534 545329
rect 230478 545255 230534 545264
rect 229100 543856 229152 543862
rect 229100 543798 229152 543804
rect 223684 535894 224158 535922
rect 225340 535894 225814 535922
rect 226996 535894 227470 535922
rect 229112 535908 229140 543798
rect 230492 535922 230520 545255
rect 232412 538348 232464 538354
rect 232412 538290 232464 538296
rect 230492 535894 230782 535922
rect 232424 535908 232452 538290
rect 233896 537169 233924 702714
rect 235184 702574 235212 703520
rect 267660 702982 267688 703520
rect 283852 702982 283880 703520
rect 267648 702976 267700 702982
rect 267648 702918 267700 702924
rect 283840 702976 283892 702982
rect 283840 702918 283892 702924
rect 273260 702908 273312 702914
rect 273260 702850 273312 702856
rect 276664 702908 276716 702914
rect 276664 702850 276716 702856
rect 235172 702568 235224 702574
rect 235172 702510 235224 702516
rect 264244 702568 264296 702574
rect 264244 702510 264296 702516
rect 255962 589384 256018 589393
rect 255962 589319 256018 589328
rect 241520 563168 241572 563174
rect 241520 563110 241572 563116
rect 241532 557534 241560 563110
rect 241532 557506 241928 557534
rect 237380 554872 237432 554878
rect 237380 554814 237432 554820
rect 235262 553480 235318 553489
rect 235262 553415 235318 553424
rect 233882 537160 233938 537169
rect 233882 537095 233938 537104
rect 233896 535922 233924 537095
rect 235276 535922 235304 553415
rect 233896 535894 234094 535922
rect 235276 535894 235750 535922
rect 237392 535908 237420 554814
rect 238760 552152 238812 552158
rect 238760 552094 238812 552100
rect 238772 535922 238800 552094
rect 240232 550724 240284 550730
rect 240232 550666 240284 550672
rect 240244 535922 240272 550666
rect 241900 535922 241928 557506
rect 247038 554840 247094 554849
rect 247038 554775 247094 554784
rect 245660 547936 245712 547942
rect 245660 547878 245712 547884
rect 243542 543960 243598 543969
rect 243542 543895 243598 543904
rect 243556 535922 243584 543895
rect 238772 535894 239062 535922
rect 240244 535894 240718 535922
rect 241900 535894 242374 535922
rect 243556 535894 244030 535922
rect 245672 535908 245700 547878
rect 247052 535922 247080 554775
rect 251824 546576 251876 546582
rect 251824 546518 251876 546524
rect 248510 545184 248566 545193
rect 248510 545119 248566 545128
rect 248524 535922 248552 545119
rect 250628 539640 250680 539646
rect 250628 539582 250680 539588
rect 247052 535894 247342 535922
rect 248524 535894 248998 535922
rect 250640 535908 250668 539582
rect 251836 535922 251864 546518
rect 253938 542600 253994 542609
rect 253938 542535 253994 542544
rect 251836 535894 252310 535922
rect 253952 535908 253980 542535
rect 255976 541249 256004 589319
rect 264256 560289 264284 702510
rect 268384 560312 268436 560318
rect 263598 560280 263654 560289
rect 263598 560215 263654 560224
rect 264242 560280 264298 560289
rect 268384 560254 268436 560260
rect 264242 560215 264298 560224
rect 263612 559065 263640 560215
rect 263598 559056 263654 559065
rect 263598 558991 263654 559000
rect 260104 553512 260156 553518
rect 260104 553454 260156 553460
rect 255962 541240 256018 541249
rect 255962 541175 256018 541184
rect 257342 541240 257398 541249
rect 257342 541175 257398 541184
rect 255594 538384 255650 538393
rect 255594 538319 255650 538328
rect 255608 535908 255636 538319
rect 257356 535922 257384 541175
rect 258448 541068 258500 541074
rect 258448 541010 258500 541016
rect 257278 535894 257384 535922
rect 258460 535922 258488 541010
rect 260116 535922 260144 553454
rect 262218 550760 262274 550769
rect 262218 550695 262274 550704
rect 258460 535894 258934 535922
rect 260116 535894 260590 535922
rect 262232 535908 262260 550695
rect 263612 535922 263640 558991
rect 268292 554804 268344 554810
rect 268292 554746 268344 554752
rect 266360 541000 266412 541006
rect 266360 540942 266412 540948
rect 266372 538801 266400 540942
rect 266358 538792 266414 538801
rect 266358 538727 266414 538736
rect 265530 538248 265586 538257
rect 265530 538183 265586 538192
rect 268304 538214 268332 554746
rect 268396 539578 268424 560254
rect 273272 559706 273300 702850
rect 276020 574796 276072 574802
rect 276020 574738 276072 574744
rect 276032 574462 276060 574738
rect 276676 574462 276704 702850
rect 281540 702840 281592 702846
rect 281540 702782 281592 702788
rect 276020 574456 276072 574462
rect 276020 574398 276072 574404
rect 276664 574456 276716 574462
rect 276664 574398 276716 574404
rect 273260 559700 273312 559706
rect 273260 559642 273312 559648
rect 273904 559700 273956 559706
rect 273904 559642 273956 559648
rect 273916 559026 273944 559642
rect 273904 559020 273956 559026
rect 273904 558962 273956 558968
rect 270500 557592 270552 557598
rect 270500 557534 270552 557540
rect 268384 539572 268436 539578
rect 268384 539514 268436 539520
rect 268304 538186 268608 538214
rect 263612 535894 263902 535922
rect 265544 535908 265572 538183
rect 267188 536852 267240 536858
rect 267188 536794 267240 536800
rect 267200 535908 267228 536794
rect 268580 535922 268608 538186
rect 270512 535922 270540 557534
rect 273916 539578 273944 558962
rect 276032 557534 276060 574398
rect 281552 557534 281580 702782
rect 300136 702642 300164 703520
rect 332520 703050 332548 703520
rect 331220 703044 331272 703050
rect 331220 702986 331272 702992
rect 332508 703044 332560 703050
rect 332508 702986 332560 702992
rect 300124 702636 300176 702642
rect 300124 702578 300176 702584
rect 300768 702636 300820 702642
rect 300768 702578 300820 702584
rect 300780 700330 300808 702578
rect 300768 700324 300820 700330
rect 300768 700266 300820 700272
rect 311900 565956 311952 565962
rect 311900 565898 311952 565904
rect 291200 565888 291252 565894
rect 291200 565830 291252 565836
rect 291212 557534 291240 565830
rect 303618 564496 303674 564505
rect 303618 564431 303674 564440
rect 309140 564460 309192 564466
rect 295984 563100 296036 563106
rect 295984 563042 296036 563048
rect 276032 557506 276888 557534
rect 281552 557506 281856 557534
rect 291212 557506 291792 557534
rect 272340 539572 272392 539578
rect 272340 539514 272392 539520
rect 273904 539572 273956 539578
rect 273904 539514 273956 539520
rect 275652 539572 275704 539578
rect 275652 539514 275704 539520
rect 268580 535894 269054 535922
rect 270512 535894 270710 535922
rect 272352 535908 272380 539514
rect 273994 538792 274050 538801
rect 273994 538727 274050 538736
rect 274008 535908 274036 538727
rect 275664 535908 275692 539514
rect 276860 535922 276888 557506
rect 278042 547904 278098 547913
rect 278042 547839 278098 547848
rect 278056 539578 278084 547839
rect 280160 542496 280212 542502
rect 280160 542438 280212 542444
rect 278044 539572 278096 539578
rect 278044 539514 278096 539520
rect 278964 539572 279016 539578
rect 278964 539514 279016 539520
rect 276860 535894 277334 535922
rect 278976 535908 279004 539514
rect 280172 535922 280200 542438
rect 281828 535922 281856 557506
rect 288440 556300 288492 556306
rect 288440 556242 288492 556248
rect 285126 552120 285182 552129
rect 285126 552055 285182 552064
rect 283932 539708 283984 539714
rect 283932 539650 283984 539656
rect 280172 535894 280646 535922
rect 281828 535894 282302 535922
rect 283944 535908 283972 539650
rect 285140 535922 285168 552055
rect 287060 548004 287112 548010
rect 287060 547946 287112 547952
rect 287072 535922 287100 547946
rect 288452 535922 288480 556242
rect 290094 549536 290150 549545
rect 290094 549471 290150 549480
rect 290108 535922 290136 549471
rect 291764 535922 291792 557506
rect 295340 547936 295392 547942
rect 295340 547878 295392 547884
rect 295352 535922 295380 547878
rect 295996 538354 296024 563042
rect 300030 546544 300086 546553
rect 300030 546479 300086 546488
rect 298376 545216 298428 545222
rect 298376 545158 298428 545164
rect 295984 538348 296036 538354
rect 295984 538290 296036 538296
rect 297180 538348 297232 538354
rect 297180 538290 297232 538296
rect 285140 535894 285614 535922
rect 287072 535894 287270 535922
rect 288452 535894 288926 535922
rect 290108 535894 290582 535922
rect 291764 535894 292238 535922
rect 295352 535894 295550 535922
rect 297192 535908 297220 538290
rect 298388 535922 298416 545158
rect 300044 535922 300072 546479
rect 303632 535922 303660 564431
rect 309140 564402 309192 564408
rect 309152 557534 309180 564402
rect 309152 557506 310008 557534
rect 305000 546508 305052 546514
rect 305000 546450 305052 546456
rect 305012 535922 305040 546450
rect 307114 539744 307170 539753
rect 307114 539679 307170 539688
rect 298388 535894 298862 535922
rect 300044 535894 300518 535922
rect 303632 535894 303830 535922
rect 305012 535894 305486 535922
rect 307128 535908 307156 539679
rect 309980 535922 310008 557506
rect 311912 535922 311940 565898
rect 331232 554033 331260 702986
rect 348804 700330 348832 703520
rect 351920 702976 351972 702982
rect 351920 702918 351972 702924
rect 349804 702840 349856 702846
rect 349804 702782 349856 702788
rect 341524 700324 341576 700330
rect 341524 700266 341576 700272
rect 342904 700324 342956 700330
rect 342904 700266 342956 700272
rect 348792 700324 348844 700330
rect 348792 700266 348844 700272
rect 332600 567248 332652 567254
rect 332600 567190 332652 567196
rect 332612 557534 332640 567190
rect 335360 561808 335412 561814
rect 335360 561750 335412 561756
rect 332612 557506 333376 557534
rect 331218 554024 331274 554033
rect 331218 553959 331274 553968
rect 316590 546544 316646 546553
rect 316590 546479 316646 546488
rect 327080 546508 327132 546514
rect 314936 545216 314988 545222
rect 314936 545158 314988 545164
rect 314948 535922 314976 545158
rect 316604 535922 316632 546479
rect 327080 546450 327132 546456
rect 324320 545148 324372 545154
rect 324320 545090 324372 545096
rect 318248 543856 318300 543862
rect 318248 543798 318300 543804
rect 318260 535922 318288 543798
rect 321560 543788 321612 543794
rect 321560 543730 321612 543736
rect 320178 541376 320234 541385
rect 320178 541311 320234 541320
rect 320192 535922 320220 541311
rect 321572 535922 321600 543730
rect 324332 540938 324360 545090
rect 324320 540932 324372 540938
rect 324320 540874 324372 540880
rect 324964 540932 325016 540938
rect 324964 540874 325016 540880
rect 323674 540152 323730 540161
rect 323674 540087 323730 540096
rect 323688 538354 323716 540087
rect 323676 538348 323728 538354
rect 323676 538290 323728 538296
rect 309980 535894 310454 535922
rect 311912 535894 312110 535922
rect 314948 535894 315422 535922
rect 316604 535894 317078 535922
rect 318260 535894 318734 535922
rect 320192 535894 320390 535922
rect 321572 535894 322046 535922
rect 323688 535908 323716 538290
rect 324976 535922 325004 540874
rect 327092 538214 327120 546450
rect 331680 545148 331732 545154
rect 331680 545090 331732 545096
rect 330024 543788 330076 543794
rect 330024 543730 330076 543736
rect 328828 539708 328880 539714
rect 328828 539650 328880 539656
rect 327092 538186 327212 538214
rect 324976 535894 325358 535922
rect 327184 535908 327212 538186
rect 328840 535908 328868 539650
rect 330036 535922 330064 543730
rect 331692 535922 331720 545090
rect 333348 535922 333376 557506
rect 335372 538214 335400 561750
rect 339958 549400 340014 549409
rect 339958 549335 340014 549344
rect 338304 542496 338356 542502
rect 338304 542438 338356 542444
rect 337106 538248 337162 538257
rect 335372 538186 335492 538214
rect 330036 535894 330510 535922
rect 331692 535894 332166 535922
rect 333348 535894 333822 535922
rect 335464 535908 335492 538186
rect 337106 538183 337162 538192
rect 337120 535908 337148 538183
rect 338316 535922 338344 542438
rect 339972 535922 340000 549335
rect 341536 540297 341564 700266
rect 342916 540938 342944 700266
rect 349816 596222 349844 702782
rect 349804 596216 349856 596222
rect 349804 596158 349856 596164
rect 343640 558952 343692 558958
rect 343640 558894 343692 558900
rect 342904 540932 342956 540938
rect 342904 540874 342956 540880
rect 341522 540288 341578 540297
rect 341522 540223 341578 540232
rect 340788 538348 340840 538354
rect 340788 538290 340840 538296
rect 340800 538218 340828 538290
rect 340788 538212 340840 538218
rect 343652 538214 343680 558894
rect 349816 557534 349844 596158
rect 349816 557506 350028 557534
rect 348238 541104 348294 541113
rect 348238 541039 348294 541048
rect 345386 539608 345442 539617
rect 345386 539543 345442 539552
rect 343652 538186 343772 538214
rect 340788 538154 340840 538160
rect 338316 535894 338790 535922
rect 339972 535894 340446 535922
rect 343744 535908 343772 538186
rect 345400 535908 345428 539543
rect 347044 538348 347096 538354
rect 347044 538290 347096 538296
rect 347056 535908 347084 538290
rect 348252 535922 348280 541039
rect 350000 539646 350028 557506
rect 351932 552090 351960 702918
rect 364996 702710 365024 703520
rect 397472 702794 397500 703520
rect 397380 702778 397500 702794
rect 397368 702772 397500 702778
rect 397420 702766 397500 702772
rect 397368 702714 397420 702720
rect 364984 702704 365036 702710
rect 364984 702646 365036 702652
rect 378784 702704 378836 702710
rect 378784 702646 378836 702652
rect 359464 702636 359516 702642
rect 359464 702578 359516 702584
rect 357532 561740 357584 561746
rect 357532 561682 357584 561688
rect 356242 560416 356298 560425
rect 356242 560351 356298 560360
rect 351920 552084 351972 552090
rect 351920 552026 351972 552032
rect 349988 539640 350040 539646
rect 349986 539608 349988 539617
rect 350040 539608 350042 539617
rect 349986 539543 350042 539552
rect 350354 538384 350410 538393
rect 350354 538319 350410 538328
rect 348252 535894 348726 535922
rect 350368 535908 350396 538319
rect 351932 538214 351960 552026
rect 353942 543824 353998 543833
rect 353942 543759 353998 543768
rect 351932 538186 352052 538214
rect 352024 535908 352052 538186
rect 353666 537024 353722 537033
rect 353666 536959 353722 536968
rect 353680 535908 353708 536959
rect 353956 536110 353984 543759
rect 356150 542464 356206 542473
rect 356150 542399 356206 542408
rect 353944 536104 353996 536110
rect 353944 536046 353996 536052
rect 354588 536104 354640 536110
rect 354588 536046 354640 536052
rect 313370 535800 313426 535809
rect 313426 535758 313766 535786
rect 313370 535735 313426 535744
rect 308402 535664 308458 535673
rect 342258 535664 342314 535673
rect 308458 535622 308798 535650
rect 342102 535622 342258 535650
rect 308402 535599 308458 535608
rect 342258 535599 342314 535608
rect 293500 535560 293552 535566
rect 302330 535528 302386 535537
rect 293552 535508 293894 535514
rect 293500 535502 293894 535508
rect 293512 535486 293894 535502
rect 302174 535486 302330 535514
rect 354600 535514 354628 536046
rect 354600 535486 354720 535514
rect 302330 535463 302386 535472
rect 354692 535401 354720 535486
rect 221094 535392 221150 535401
rect 221094 535327 221150 535336
rect 354678 535392 354734 535401
rect 355350 535350 355640 535378
rect 354678 535327 354734 535336
rect 355612 535294 355640 535350
rect 204904 535288 204956 535294
rect 204904 535230 204956 535236
rect 355600 535288 355652 535294
rect 355600 535230 355652 535236
rect 199844 534812 199896 534818
rect 199844 534754 199896 534760
rect 199750 533352 199806 533361
rect 199750 533287 199806 533296
rect 199476 530596 199528 530602
rect 199476 530538 199528 530544
rect 199658 378176 199714 378185
rect 199658 378111 199714 378120
rect 199672 377505 199700 378111
rect 199658 377496 199714 377505
rect 199658 377431 199714 377440
rect 199660 377324 199712 377330
rect 199660 377266 199712 377272
rect 199474 376544 199530 376553
rect 199474 376479 199530 376488
rect 199384 365832 199436 365838
rect 199384 365774 199436 365780
rect 199396 320929 199424 365774
rect 199382 320920 199438 320929
rect 199382 320855 199438 320864
rect 199488 314673 199516 376479
rect 199672 370530 199700 377266
rect 199856 376145 199884 534754
rect 356164 518894 356192 542399
rect 356256 523025 356284 560351
rect 357544 557534 357572 561682
rect 357544 557506 357940 557534
rect 357440 542428 357492 542434
rect 357440 542370 357492 542376
rect 356336 538280 356388 538286
rect 356336 538222 356388 538228
rect 356242 523016 356298 523025
rect 356242 522951 356298 522960
rect 356164 518866 356284 518894
rect 356256 496097 356284 518866
rect 356242 496088 356298 496097
rect 356242 496023 356298 496032
rect 356242 492688 356298 492697
rect 356242 492623 356298 492632
rect 356256 489914 356284 492623
rect 356348 490385 356376 538222
rect 357452 512689 357480 542370
rect 357622 540288 357678 540297
rect 357622 540223 357678 540232
rect 357636 519897 357664 540223
rect 357912 532137 357940 557506
rect 358818 538384 358874 538393
rect 358818 538319 358874 538328
rect 357898 532128 357954 532137
rect 357898 532063 357954 532072
rect 358726 532128 358782 532137
rect 358726 532063 358782 532072
rect 358740 532030 358768 532063
rect 358728 532024 358780 532030
rect 358728 531966 358780 531972
rect 358726 529680 358782 529689
rect 358726 529615 358782 529624
rect 358740 528630 358768 529615
rect 358728 528624 358780 528630
rect 358728 528566 358780 528572
rect 358726 527232 358782 527241
rect 358726 527167 358728 527176
rect 358780 527167 358782 527176
rect 358728 527138 358780 527144
rect 358726 524784 358782 524793
rect 358726 524719 358782 524728
rect 358740 524482 358768 524719
rect 358728 524476 358780 524482
rect 358728 524418 358780 524424
rect 358726 522336 358782 522345
rect 358726 522271 358782 522280
rect 358740 520946 358768 522271
rect 358728 520940 358780 520946
rect 358728 520882 358780 520888
rect 357622 519888 357678 519897
rect 357622 519823 357678 519832
rect 358726 519888 358782 519897
rect 358726 519823 358782 519832
rect 358740 519586 358768 519823
rect 358728 519580 358780 519586
rect 358728 519522 358780 519528
rect 358726 517440 358782 517449
rect 358726 517375 358782 517384
rect 358740 516186 358768 517375
rect 358728 516180 358780 516186
rect 358728 516122 358780 516128
rect 358082 514992 358138 515001
rect 358082 514927 358138 514936
rect 357438 512680 357494 512689
rect 357438 512615 357494 512624
rect 356702 507648 356758 507657
rect 356702 507583 356758 507592
rect 356334 490376 356390 490385
rect 356334 490311 356390 490320
rect 356164 489886 356284 489914
rect 202234 377632 202290 377641
rect 199842 376136 199898 376145
rect 199842 376071 199898 376080
rect 200040 374134 200068 377604
rect 201592 377528 201644 377534
rect 201406 377496 201462 377505
rect 201592 377470 201644 377476
rect 201406 377431 201462 377440
rect 200028 374128 200080 374134
rect 200028 374070 200080 374076
rect 199568 370524 199620 370530
rect 199568 370466 199620 370472
rect 199660 370524 199712 370530
rect 199660 370466 199712 370472
rect 199580 342990 199608 370466
rect 200212 368484 200264 368490
rect 200212 368426 200264 368432
rect 199568 342984 199620 342990
rect 199568 342926 199620 342932
rect 199660 336864 199712 336870
rect 199660 336806 199712 336812
rect 199568 330608 199620 330614
rect 199568 330550 199620 330556
rect 199474 314664 199530 314673
rect 199474 314599 199530 314608
rect 199580 307154 199608 330550
rect 199672 326466 199700 336806
rect 199660 326460 199712 326466
rect 199660 326402 199712 326408
rect 200118 314800 200174 314809
rect 200118 314735 200174 314744
rect 199658 314664 199714 314673
rect 199658 314599 199714 314608
rect 199672 313993 199700 314599
rect 199658 313984 199714 313993
rect 199658 313919 199714 313928
rect 199568 307148 199620 307154
rect 199568 307090 199620 307096
rect 200028 307080 200080 307086
rect 200028 307022 200080 307028
rect 198648 299532 198700 299538
rect 198648 299474 198700 299480
rect 198554 262848 198610 262857
rect 198554 262783 198610 262792
rect 198660 262313 198688 299474
rect 199934 293312 199990 293321
rect 199934 293247 199990 293256
rect 199290 287192 199346 287201
rect 199290 287127 199346 287136
rect 199304 282985 199332 287127
rect 199382 284472 199438 284481
rect 199382 284407 199438 284416
rect 199290 282976 199346 282985
rect 199290 282911 199346 282920
rect 198646 262304 198702 262313
rect 198646 262239 198702 262248
rect 199396 257378 199424 284407
rect 199476 284368 199528 284374
rect 199476 284310 199528 284316
rect 199488 272542 199516 284310
rect 199948 281625 199976 293247
rect 199934 281616 199990 281625
rect 199934 281551 199990 281560
rect 200040 280265 200068 307022
rect 200132 296714 200160 314735
rect 200224 301481 200252 368426
rect 201420 364993 201448 377431
rect 201406 364984 201462 364993
rect 201406 364919 201462 364928
rect 200764 362228 200816 362234
rect 200764 362170 200816 362176
rect 200776 314809 200804 362170
rect 201604 355230 201632 377470
rect 201696 375358 201724 377604
rect 355322 377632 355378 377641
rect 202234 377567 202290 377576
rect 202892 377590 203366 377618
rect 204272 377590 205022 377618
rect 201684 375352 201736 375358
rect 201684 375294 201736 375300
rect 201684 374128 201736 374134
rect 201684 374070 201736 374076
rect 201592 355224 201644 355230
rect 201592 355166 201644 355172
rect 201604 354754 201632 355166
rect 201592 354748 201644 354754
rect 201592 354690 201644 354696
rect 200856 331968 200908 331974
rect 200856 331910 200908 331916
rect 200762 314800 200818 314809
rect 200762 314735 200818 314744
rect 200210 301472 200266 301481
rect 200210 301407 200266 301416
rect 200868 300801 200896 331910
rect 201592 326392 201644 326398
rect 201592 326334 201644 326340
rect 201408 301504 201460 301510
rect 201406 301472 201408 301481
rect 201460 301472 201462 301481
rect 201406 301407 201462 301416
rect 200854 300792 200910 300801
rect 200854 300727 200910 300736
rect 200762 299432 200818 299441
rect 200762 299367 200818 299376
rect 200132 296686 200528 296714
rect 200394 286376 200450 286385
rect 200394 286311 200450 286320
rect 200408 284172 200436 286311
rect 200500 284186 200528 296686
rect 200776 285870 200804 299367
rect 201604 294545 201632 326334
rect 201696 298858 201724 374070
rect 202144 355224 202196 355230
rect 202144 355166 202196 355172
rect 202156 304881 202184 355166
rect 202248 343777 202276 377567
rect 202788 375352 202840 375358
rect 202788 375294 202840 375300
rect 202800 361865 202828 375294
rect 202892 369170 202920 377590
rect 202880 369164 202932 369170
rect 202880 369106 202932 369112
rect 203522 367432 203578 367441
rect 203522 367367 203578 367376
rect 202786 361856 202842 361865
rect 202786 361791 202842 361800
rect 202788 349852 202840 349858
rect 202788 349794 202840 349800
rect 202234 343768 202290 343777
rect 202234 343703 202290 343712
rect 202248 342922 202276 343703
rect 202236 342916 202288 342922
rect 202236 342858 202288 342864
rect 202800 317529 202828 349794
rect 203536 331809 203564 367367
rect 203522 331800 203578 331809
rect 203522 331735 203578 331744
rect 203522 329080 203578 329089
rect 203522 329015 203578 329024
rect 202786 317520 202842 317529
rect 202786 317455 202842 317464
rect 202142 304872 202198 304881
rect 202142 304807 202198 304816
rect 201684 298852 201736 298858
rect 201684 298794 201736 298800
rect 201590 294536 201646 294545
rect 201590 294471 201646 294480
rect 201604 293978 201632 294471
rect 201420 293950 201632 293978
rect 200764 285864 200816 285870
rect 200764 285806 200816 285812
rect 201224 285796 201276 285802
rect 201224 285738 201276 285744
rect 201130 285696 201186 285705
rect 201130 285631 201186 285640
rect 200500 284158 200790 284186
rect 201144 283966 201172 285631
rect 201236 283966 201264 285738
rect 201420 284186 201448 293950
rect 201682 291952 201738 291961
rect 201682 291887 201738 291896
rect 201498 289232 201554 289241
rect 201498 289167 201554 289176
rect 201512 284889 201540 289167
rect 201498 284880 201554 284889
rect 201498 284815 201554 284824
rect 201342 284158 201448 284186
rect 201696 284172 201724 291887
rect 202234 287328 202290 287337
rect 202234 287263 202290 287272
rect 202248 284172 202276 287263
rect 202800 284172 202828 317455
rect 202878 300792 202934 300801
rect 202878 300727 202934 300736
rect 202892 291961 202920 300727
rect 202878 291952 202934 291961
rect 202878 291887 202934 291896
rect 203536 291145 203564 329015
rect 204272 297430 204300 377590
rect 204352 376032 204404 376038
rect 204352 375974 204404 375980
rect 204260 297424 204312 297430
rect 204260 297366 204312 297372
rect 204364 293282 204392 375974
rect 206664 375358 206692 377604
rect 207032 377590 208334 377618
rect 209792 377590 209990 377618
rect 211172 377590 211646 377618
rect 212644 377590 213302 377618
rect 214576 377590 214958 377618
rect 205640 375352 205692 375358
rect 205640 375294 205692 375300
rect 206652 375352 206704 375358
rect 206652 375294 206704 375300
rect 205652 356833 205680 375294
rect 206376 371884 206428 371890
rect 206376 371826 206428 371832
rect 206284 369164 206336 369170
rect 206284 369106 206336 369112
rect 205638 356824 205694 356833
rect 205638 356759 205694 356768
rect 204444 347064 204496 347070
rect 204444 347006 204496 347012
rect 204456 299441 204484 347006
rect 205178 325136 205234 325145
rect 205178 325071 205234 325080
rect 204996 299464 205048 299470
rect 204442 299432 204498 299441
rect 204442 299367 204498 299376
rect 204994 299432 204996 299441
rect 205048 299432 205050 299441
rect 204994 299367 205050 299376
rect 204352 293276 204404 293282
rect 204352 293218 204404 293224
rect 204904 292664 204956 292670
rect 204904 292606 204956 292612
rect 204916 291242 204944 292606
rect 204904 291236 204956 291242
rect 204904 291178 204956 291184
rect 203522 291136 203578 291145
rect 203522 291071 203578 291080
rect 204166 291136 204222 291145
rect 204166 291071 204222 291080
rect 204180 289921 204208 291071
rect 204166 289912 204222 289921
rect 204166 289847 204222 289856
rect 203706 285832 203762 285841
rect 203706 285767 203762 285776
rect 203156 285728 203208 285734
rect 203156 285670 203208 285676
rect 203168 284172 203196 285670
rect 203720 284172 203748 285767
rect 204180 285734 204208 289847
rect 204718 288144 204774 288153
rect 204718 288079 204774 288088
rect 204258 287192 204314 287201
rect 204258 287127 204314 287136
rect 204168 285728 204220 285734
rect 204168 285670 204220 285676
rect 204272 284172 204300 287127
rect 204732 285977 204760 288079
rect 204718 285968 204774 285977
rect 204718 285903 204774 285912
rect 204628 285864 204680 285870
rect 204628 285806 204680 285812
rect 204640 284172 204668 285806
rect 204916 285734 204944 291178
rect 204904 285728 204956 285734
rect 204904 285670 204956 285676
rect 205192 284172 205220 325071
rect 206296 323785 206324 369106
rect 206388 341562 206416 371826
rect 207032 369918 207060 377590
rect 208490 376136 208546 376145
rect 208490 376071 208546 376080
rect 208400 372632 208452 372638
rect 208400 372574 208452 372580
rect 207020 369912 207072 369918
rect 207020 369854 207072 369860
rect 207664 369912 207716 369918
rect 207664 369854 207716 369860
rect 207676 358086 207704 369854
rect 207664 358080 207716 358086
rect 207664 358022 207716 358028
rect 206468 357468 206520 357474
rect 206468 357410 206520 357416
rect 206480 346390 206508 357410
rect 206468 346384 206520 346390
rect 206468 346326 206520 346332
rect 207662 344312 207718 344321
rect 207662 344247 207718 344256
rect 206376 341556 206428 341562
rect 206376 341498 206428 341504
rect 206466 340912 206522 340921
rect 206466 340847 206522 340856
rect 206374 337512 206430 337521
rect 206374 337447 206430 337456
rect 206282 323776 206338 323785
rect 206282 323711 206338 323720
rect 206284 319456 206336 319462
rect 206284 319398 206336 319404
rect 205916 317552 205968 317558
rect 205916 317494 205968 317500
rect 205928 312594 205956 317494
rect 205916 312588 205968 312594
rect 205916 312530 205968 312536
rect 206296 304298 206324 319398
rect 206388 311953 206416 337447
rect 206480 319433 206508 340847
rect 206560 325100 206612 325106
rect 206560 325042 206612 325048
rect 206466 319424 206522 319433
rect 206466 319359 206522 319368
rect 206374 311944 206430 311953
rect 206374 311879 206430 311888
rect 206572 310554 206600 325042
rect 206926 311944 206982 311953
rect 206926 311879 206982 311888
rect 206560 310548 206612 310554
rect 206560 310490 206612 310496
rect 206836 310548 206888 310554
rect 206836 310490 206888 310496
rect 206284 304292 206336 304298
rect 206284 304234 206336 304240
rect 206652 296064 206704 296070
rect 206652 296006 206704 296012
rect 206100 285728 206152 285734
rect 205546 285696 205602 285705
rect 206100 285670 206152 285676
rect 205546 285631 205602 285640
rect 205560 284172 205588 285631
rect 206112 284172 206140 285670
rect 206664 284172 206692 296006
rect 206848 285705 206876 310490
rect 206940 287054 206968 311879
rect 207676 311273 207704 344247
rect 207756 326392 207808 326398
rect 207756 326334 207808 326340
rect 207662 311264 207718 311273
rect 207662 311199 207718 311208
rect 207768 304366 207796 326334
rect 208412 306270 208440 372574
rect 208504 349110 208532 376071
rect 209688 374672 209740 374678
rect 209688 374614 209740 374620
rect 208492 349104 208544 349110
rect 208492 349046 208544 349052
rect 209044 349104 209096 349110
rect 209700 349081 209728 374614
rect 209044 349046 209096 349052
rect 209134 349072 209190 349081
rect 209056 347818 209084 349046
rect 209134 349007 209190 349016
rect 209686 349072 209742 349081
rect 209686 349007 209742 349016
rect 209148 348401 209176 349007
rect 209134 348392 209190 348401
rect 209134 348327 209190 348336
rect 209044 347812 209096 347818
rect 209044 347754 209096 347760
rect 209056 315314 209084 347754
rect 209136 319524 209188 319530
rect 209136 319466 209188 319472
rect 209044 315308 209096 315314
rect 209044 315250 209096 315256
rect 208490 311128 208546 311137
rect 208490 311063 208546 311072
rect 208504 307873 208532 311063
rect 208490 307864 208546 307873
rect 208490 307799 208546 307808
rect 208400 306264 208452 306270
rect 208400 306206 208452 306212
rect 208412 304994 208440 306206
rect 208320 304966 208440 304994
rect 207756 304360 207808 304366
rect 207756 304302 207808 304308
rect 208320 296714 208348 304966
rect 208136 296686 208348 296714
rect 206940 287026 207060 287054
rect 206834 285696 206890 285705
rect 206834 285631 206890 285640
rect 207032 284172 207060 287026
rect 207570 285696 207626 285705
rect 207570 285631 207626 285640
rect 207584 284172 207612 285631
rect 208136 284172 208164 296686
rect 208504 284172 208532 307799
rect 209148 298217 209176 319466
rect 209134 298208 209190 298217
rect 209134 298143 209190 298152
rect 209410 298208 209466 298217
rect 209410 298143 209466 298152
rect 209044 297424 209096 297430
rect 209044 297366 209096 297372
rect 209056 296750 209084 297366
rect 209044 296744 209096 296750
rect 209044 296686 209096 296692
rect 209056 284172 209084 296686
rect 209424 284172 209452 298143
rect 209792 297537 209820 377590
rect 211172 354006 211200 377590
rect 211802 376000 211858 376009
rect 211802 375935 211858 375944
rect 211160 354000 211212 354006
rect 211160 353942 211212 353948
rect 211068 316736 211120 316742
rect 211068 316678 211120 316684
rect 211080 316062 211108 316678
rect 209964 316056 210016 316062
rect 209964 315998 210016 316004
rect 211068 316056 211120 316062
rect 211068 315998 211120 316004
rect 209778 297528 209834 297537
rect 209778 297463 209834 297472
rect 209976 284172 210004 315998
rect 211816 302569 211844 375935
rect 211896 327820 211948 327826
rect 211896 327762 211948 327768
rect 211802 302560 211858 302569
rect 211802 302495 211858 302504
rect 211436 290488 211488 290494
rect 211436 290430 211488 290436
rect 211448 289950 211476 290430
rect 211436 289944 211488 289950
rect 211436 289886 211488 289892
rect 210976 289128 211028 289134
rect 210976 289070 211028 289076
rect 210988 288522 211016 289070
rect 210516 288516 210568 288522
rect 210516 288458 210568 288464
rect 210976 288516 211028 288522
rect 210976 288458 211028 288464
rect 210528 284172 210556 288458
rect 210884 284368 210936 284374
rect 210884 284310 210936 284316
rect 210896 284172 210924 284310
rect 211448 284172 211476 289886
rect 211816 288153 211844 302495
rect 211908 290465 211936 327762
rect 212644 326398 212672 377590
rect 214576 374105 214604 377590
rect 215208 376712 215260 376718
rect 215208 376654 215260 376660
rect 215220 375358 215248 376654
rect 215208 375352 215260 375358
rect 215208 375294 215260 375300
rect 214562 374096 214618 374105
rect 214562 374031 214618 374040
rect 213828 365016 213880 365022
rect 213828 364958 213880 364964
rect 212632 326392 212684 326398
rect 212632 326334 212684 326340
rect 212908 313948 212960 313954
rect 212908 313890 212960 313896
rect 212920 311914 212948 313890
rect 212908 311908 212960 311914
rect 212908 311850 212960 311856
rect 211894 290456 211950 290465
rect 211894 290391 211950 290400
rect 211802 288144 211858 288153
rect 211802 288079 211858 288088
rect 211908 287054 211936 290391
rect 211908 287026 212120 287054
rect 211986 285696 212042 285705
rect 211986 285631 212042 285640
rect 212000 284172 212028 285631
rect 212092 284186 212120 287026
rect 212092 284158 212382 284186
rect 212920 284172 212948 311850
rect 213460 285796 213512 285802
rect 213460 285738 213512 285744
rect 213472 284172 213500 285738
rect 213840 284172 213868 364958
rect 214576 324970 214604 374031
rect 214656 326392 214708 326398
rect 214656 326334 214708 326340
rect 214564 324964 214616 324970
rect 214564 324906 214616 324912
rect 214564 320884 214616 320890
rect 214564 320826 214616 320832
rect 214576 312497 214604 320826
rect 214668 316713 214696 326334
rect 214654 316704 214710 316713
rect 214654 316639 214710 316648
rect 215114 316704 215170 316713
rect 215114 316639 215170 316648
rect 214562 312488 214618 312497
rect 214562 312423 214618 312432
rect 215128 310457 215156 316639
rect 213918 310448 213974 310457
rect 213918 310383 213974 310392
rect 215114 310448 215170 310457
rect 215114 310383 215170 310392
rect 213932 285802 213960 310383
rect 214564 307148 214616 307154
rect 214564 307090 214616 307096
rect 214012 300892 214064 300898
rect 214012 300834 214064 300840
rect 213920 285796 213972 285802
rect 213920 285738 213972 285744
rect 214024 285705 214052 300834
rect 214576 286346 214604 307090
rect 215220 297430 215248 375294
rect 216600 374678 216628 377604
rect 218256 375358 218284 377604
rect 219452 377590 219926 377618
rect 221476 377590 221582 377618
rect 222212 377590 223238 377618
rect 223592 377590 224894 377618
rect 226352 377590 226550 377618
rect 227732 377590 228206 377618
rect 229112 377590 229862 377618
rect 230492 377590 231518 377618
rect 218244 375352 218296 375358
rect 218244 375294 218296 375300
rect 216588 374672 216640 374678
rect 216588 374614 216640 374620
rect 218702 369200 218758 369209
rect 218702 369135 218758 369144
rect 216126 363080 216182 363089
rect 216126 363015 216182 363024
rect 216034 358864 216090 358873
rect 216034 358799 216090 358808
rect 215944 342984 215996 342990
rect 215944 342926 215996 342932
rect 215852 315308 215904 315314
rect 215852 315250 215904 315256
rect 215864 306406 215892 315250
rect 215852 306400 215904 306406
rect 215852 306342 215904 306348
rect 215208 297424 215260 297430
rect 215208 297366 215260 297372
rect 214564 286340 214616 286346
rect 214564 286282 214616 286288
rect 215300 285796 215352 285802
rect 215300 285738 215352 285744
rect 214010 285696 214066 285705
rect 214010 285631 214066 285640
rect 214746 285696 214802 285705
rect 214746 285631 214802 285640
rect 214024 285025 214052 285631
rect 214010 285016 214066 285025
rect 214010 284951 214066 284960
rect 214760 284172 214788 285631
rect 215312 284172 215340 285738
rect 215864 284172 215892 306342
rect 215956 285841 215984 342926
rect 216048 327146 216076 358799
rect 216140 340105 216168 363015
rect 216680 340196 216732 340202
rect 216680 340138 216732 340144
rect 216126 340096 216182 340105
rect 216126 340031 216182 340040
rect 216128 338768 216180 338774
rect 216128 338710 216180 338716
rect 216036 327140 216088 327146
rect 216036 327082 216088 327088
rect 216048 325145 216076 327082
rect 216034 325136 216090 325145
rect 216034 325071 216090 325080
rect 216034 320784 216090 320793
rect 216034 320719 216090 320728
rect 216048 309806 216076 320719
rect 216140 309942 216168 338710
rect 216128 309936 216180 309942
rect 216128 309878 216180 309884
rect 216036 309800 216088 309806
rect 216036 309742 216088 309748
rect 216048 306374 216076 309742
rect 216048 306346 216260 306374
rect 216036 300892 216088 300898
rect 216036 300834 216088 300840
rect 216048 296070 216076 300834
rect 216036 296064 216088 296070
rect 216036 296006 216088 296012
rect 215942 285832 215998 285841
rect 215942 285767 215998 285776
rect 216232 285705 216260 306346
rect 216692 287745 216720 340138
rect 217324 333328 217376 333334
rect 217324 333270 217376 333276
rect 217336 313954 217364 333270
rect 217324 313948 217376 313954
rect 217324 313890 217376 313896
rect 218058 304872 218114 304881
rect 218058 304807 218114 304816
rect 218072 304502 218100 304807
rect 218060 304496 218112 304502
rect 218060 304438 218112 304444
rect 218716 301073 218744 369135
rect 219346 321600 219402 321609
rect 219346 321535 219402 321544
rect 219360 304502 219388 321535
rect 219452 314129 219480 377590
rect 221476 374105 221504 377590
rect 221462 374096 221518 374105
rect 221462 374031 221518 374040
rect 221476 355337 221504 374031
rect 221462 355328 221518 355337
rect 221462 355263 221518 355272
rect 222212 349761 222240 377590
rect 222842 365800 222898 365809
rect 222842 365735 222898 365744
rect 222198 349752 222254 349761
rect 222198 349687 222254 349696
rect 221556 343732 221608 343738
rect 221556 343674 221608 343680
rect 221464 326460 221516 326466
rect 221464 326402 221516 326408
rect 220084 323604 220136 323610
rect 220084 323546 220136 323552
rect 219438 314120 219494 314129
rect 219438 314055 219494 314064
rect 219348 304496 219400 304502
rect 219348 304438 219400 304444
rect 218242 301064 218298 301073
rect 218242 300999 218298 301008
rect 218702 301064 218758 301073
rect 218702 300999 218758 301008
rect 218058 297120 218114 297129
rect 218058 297055 218114 297064
rect 218072 295089 218100 297055
rect 218058 295080 218114 295089
rect 218058 295015 218114 295024
rect 218060 289944 218112 289950
rect 218060 289886 218112 289892
rect 218072 289377 218100 289886
rect 218058 289368 218114 289377
rect 218058 289303 218114 289312
rect 216678 287736 216734 287745
rect 216678 287671 216734 287680
rect 216692 287054 216720 287671
rect 217690 287328 217746 287337
rect 217690 287263 217746 287272
rect 216772 287156 216824 287162
rect 216772 287098 216824 287104
rect 216600 287026 216720 287054
rect 216600 285802 216628 287026
rect 216588 285796 216640 285802
rect 216588 285738 216640 285744
rect 216218 285696 216274 285705
rect 216218 285631 216274 285640
rect 216784 284172 216812 287098
rect 217322 284472 217378 284481
rect 217322 284407 217378 284416
rect 217336 284172 217364 284407
rect 217704 284172 217732 287263
rect 218058 285832 218114 285841
rect 218058 285767 218114 285776
rect 218072 285666 218100 285767
rect 218060 285660 218112 285666
rect 218060 285602 218112 285608
rect 218256 284172 218284 300999
rect 219714 300792 219770 300801
rect 219714 300727 219770 300736
rect 218702 300112 218758 300121
rect 218702 300047 218758 300056
rect 218716 295225 218744 300047
rect 219728 299713 219756 300727
rect 219714 299704 219770 299713
rect 219714 299639 219770 299648
rect 218702 295216 218758 295225
rect 218702 295151 218758 295160
rect 218612 285660 218664 285666
rect 218612 285602 218664 285608
rect 218624 284172 218652 285602
rect 219728 284172 219756 299639
rect 220096 291174 220124 323546
rect 220176 322312 220228 322318
rect 220176 322254 220228 322260
rect 220188 300801 220216 322254
rect 221188 304496 221240 304502
rect 221188 304438 221240 304444
rect 220174 300792 220230 300801
rect 220174 300727 220230 300736
rect 220726 292632 220782 292641
rect 220636 292596 220688 292602
rect 220726 292567 220782 292576
rect 220636 292538 220688 292544
rect 220084 291168 220136 291174
rect 220084 291110 220136 291116
rect 220648 287162 220676 292538
rect 220740 290601 220768 292567
rect 220726 290592 220782 290601
rect 220726 290527 220782 290536
rect 220636 287156 220688 287162
rect 220636 287098 220688 287104
rect 220082 285832 220138 285841
rect 220082 285767 220138 285776
rect 220096 284172 220124 285767
rect 220648 284172 220676 287098
rect 221200 284172 221228 304438
rect 221476 285705 221504 326402
rect 221568 312594 221596 343674
rect 221648 312724 221700 312730
rect 221648 312666 221700 312672
rect 221556 312588 221608 312594
rect 221556 312530 221608 312536
rect 221660 289921 221688 312666
rect 222856 304366 222884 365735
rect 223592 352646 223620 377590
rect 223580 352640 223632 352646
rect 223580 352582 223632 352588
rect 223592 351966 223620 352582
rect 223580 351960 223632 351966
rect 223580 351902 223632 351908
rect 224316 351960 224368 351966
rect 224316 351902 224368 351908
rect 224224 351212 224276 351218
rect 224224 351154 224276 351160
rect 222934 338192 222990 338201
rect 222934 338127 222990 338136
rect 222844 304360 222896 304366
rect 222844 304302 222896 304308
rect 222948 294098 222976 338127
rect 223028 316056 223080 316062
rect 223028 315998 223080 316004
rect 223040 306338 223068 315998
rect 223028 306332 223080 306338
rect 223028 306274 223080 306280
rect 223212 305108 223264 305114
rect 223212 305050 223264 305056
rect 223026 304192 223082 304201
rect 223026 304127 223082 304136
rect 223040 295361 223068 304127
rect 223224 299470 223252 305050
rect 223212 299464 223264 299470
rect 223212 299406 223264 299412
rect 223026 295352 223082 295361
rect 223026 295287 223082 295296
rect 222476 294092 222528 294098
rect 222476 294034 222528 294040
rect 222936 294092 222988 294098
rect 222936 294034 222988 294040
rect 222108 291168 222160 291174
rect 222108 291110 222160 291116
rect 222120 289950 222148 291110
rect 222108 289944 222160 289950
rect 221646 289912 221702 289921
rect 222108 289886 222160 289892
rect 221646 289847 221702 289856
rect 221462 285696 221518 285705
rect 221462 285631 221518 285640
rect 221660 284186 221688 289847
rect 221582 284158 221688 284186
rect 222120 284172 222148 289886
rect 222488 284172 222516 294034
rect 222842 288552 222898 288561
rect 222842 288487 222898 288496
rect 222856 286385 222884 288487
rect 222842 286376 222898 286385
rect 222842 286311 222898 286320
rect 223040 284172 223068 295287
rect 224236 290018 224264 351154
rect 224328 344321 224356 351902
rect 224314 344312 224370 344321
rect 224314 344247 224370 344256
rect 225602 343768 225658 343777
rect 225602 343703 225658 343712
rect 224316 336048 224368 336054
rect 224316 335990 224368 335996
rect 224224 290012 224276 290018
rect 224224 289954 224276 289960
rect 223580 287088 223632 287094
rect 223580 287030 223632 287036
rect 201132 283960 201184 283966
rect 201132 283902 201184 283908
rect 201224 283960 201276 283966
rect 214470 283928 214526 283937
rect 201224 283902 201276 283908
rect 214406 283886 214470 283914
rect 216402 283928 216458 283937
rect 216246 283886 216402 283914
rect 214470 283863 214526 283872
rect 216402 283863 216458 283872
rect 218794 283928 218850 283937
rect 223592 283914 223620 287030
rect 224236 284186 224264 289954
rect 224328 284481 224356 335990
rect 224408 289876 224460 289882
rect 224408 289818 224460 289824
rect 224420 287094 224448 289818
rect 224408 287088 224460 287094
rect 224408 287030 224460 287036
rect 224314 284472 224370 284481
rect 224314 284407 224370 284416
rect 223974 284158 224264 284186
rect 224420 284186 224448 287030
rect 225052 286340 225104 286346
rect 225052 286282 225104 286288
rect 225064 285977 225092 286282
rect 225050 285968 225106 285977
rect 225050 285903 225106 285912
rect 224420 284158 224526 284186
rect 225064 284172 225092 285903
rect 225420 285728 225472 285734
rect 225616 285705 225644 343703
rect 225694 322144 225750 322153
rect 225694 322079 225750 322088
rect 225708 299577 225736 322079
rect 226248 313336 226300 313342
rect 226248 313278 226300 313284
rect 226260 309126 226288 313278
rect 226248 309120 226300 309126
rect 226248 309062 226300 309068
rect 225694 299568 225750 299577
rect 225694 299503 225750 299512
rect 225970 298752 226026 298761
rect 225970 298687 226026 298696
rect 225420 285670 225472 285676
rect 225602 285696 225658 285705
rect 225432 284172 225460 285670
rect 225602 285631 225658 285640
rect 225984 284172 226012 298687
rect 226352 297401 226380 377590
rect 227076 356788 227128 356794
rect 227076 356730 227128 356736
rect 226984 354000 227036 354006
rect 226984 353942 227036 353948
rect 226996 340785 227024 353942
rect 227088 344486 227116 356730
rect 227732 348537 227760 377590
rect 228364 374672 228416 374678
rect 228364 374614 228416 374620
rect 227718 348528 227774 348537
rect 227718 348463 227774 348472
rect 227628 345024 227680 345030
rect 227628 344966 227680 344972
rect 227640 344486 227668 344966
rect 227076 344480 227128 344486
rect 227076 344422 227128 344428
rect 227628 344480 227680 344486
rect 227628 344422 227680 344428
rect 226982 340776 227038 340785
rect 226982 340711 227038 340720
rect 226892 309120 226944 309126
rect 226892 309062 226944 309068
rect 226338 297392 226394 297401
rect 226338 297327 226394 297336
rect 226522 285696 226578 285705
rect 226522 285631 226578 285640
rect 226536 284172 226564 285631
rect 226904 284172 226932 309062
rect 227442 299568 227498 299577
rect 227442 299503 227498 299512
rect 226984 295384 227036 295390
rect 226984 295326 227036 295332
rect 226996 285734 227024 295326
rect 226984 285728 227036 285734
rect 226984 285670 227036 285676
rect 227456 284172 227484 299503
rect 227640 295390 227668 344422
rect 228376 343670 228404 374614
rect 229112 357406 229140 377590
rect 229100 357400 229152 357406
rect 229100 357342 229152 357348
rect 228454 353424 228510 353433
rect 228454 353359 228510 353368
rect 228364 343664 228416 343670
rect 228364 343606 228416 343612
rect 228376 308446 228404 343606
rect 228468 336054 228496 353359
rect 229192 338156 229244 338162
rect 229192 338098 229244 338104
rect 228456 336048 228508 336054
rect 228456 335990 228508 335996
rect 228456 325032 228508 325038
rect 228456 324974 228508 324980
rect 228364 308440 228416 308446
rect 228364 308382 228416 308388
rect 228364 298240 228416 298246
rect 228364 298182 228416 298188
rect 227628 295384 227680 295390
rect 227628 295326 227680 295332
rect 228376 295225 228404 298182
rect 228468 296714 228496 324974
rect 228914 296984 228970 296993
rect 228914 296919 228970 296928
rect 228928 296714 228956 296919
rect 228468 296686 228956 296714
rect 228362 295216 228418 295225
rect 228362 295151 228418 295160
rect 228376 284172 228404 295151
rect 228928 284172 228956 296686
rect 223762 283928 223818 283937
rect 218850 283886 219190 283914
rect 223592 283900 223762 283914
rect 223606 283886 223762 283900
rect 218794 283863 218850 283872
rect 227994 283928 228050 283937
rect 227838 283886 227994 283914
rect 223762 283863 223818 283872
rect 229204 283914 229232 338098
rect 229742 332616 229798 332625
rect 229742 332551 229798 332560
rect 229756 287201 229784 332551
rect 230492 331129 230520 377590
rect 233160 374678 233188 377604
rect 234632 377590 234830 377618
rect 236012 377590 236486 377618
rect 233882 376000 233938 376009
rect 233882 375935 233938 375944
rect 233896 375193 233924 375935
rect 233882 375184 233938 375193
rect 233882 375119 233938 375128
rect 233884 375080 233936 375086
rect 233884 375022 233936 375028
rect 233148 374672 233200 374678
rect 233148 374614 233200 374620
rect 232504 369164 232556 369170
rect 232504 369106 232556 369112
rect 232516 358154 232544 369106
rect 232596 361616 232648 361622
rect 232596 361558 232648 361564
rect 232504 358148 232556 358154
rect 232504 358090 232556 358096
rect 232502 356688 232558 356697
rect 232502 356623 232558 356632
rect 231122 341456 231178 341465
rect 231122 341391 231178 341400
rect 230478 331120 230534 331129
rect 230478 331055 230534 331064
rect 231136 309777 231164 341391
rect 231214 331120 231270 331129
rect 231214 331055 231270 331064
rect 231122 309768 231178 309777
rect 231122 309703 231178 309712
rect 231228 306649 231256 331055
rect 231674 311264 231730 311273
rect 231674 311199 231730 311208
rect 231688 309233 231716 311199
rect 231674 309224 231730 309233
rect 231674 309159 231730 309168
rect 231214 306640 231270 306649
rect 231214 306575 231270 306584
rect 231228 296714 231256 306575
rect 231136 296686 231256 296714
rect 231136 293321 231164 296686
rect 231122 293312 231178 293321
rect 231122 293247 231178 293256
rect 230386 292088 230442 292097
rect 230386 292023 230442 292032
rect 229742 287192 229798 287201
rect 229742 287127 229798 287136
rect 229756 284186 229784 287127
rect 229756 284158 229862 284186
rect 230400 284172 230428 292023
rect 231308 288448 231360 288454
rect 231308 288390 231360 288396
rect 230756 285864 230808 285870
rect 230756 285806 230808 285812
rect 230768 284172 230796 285806
rect 229466 283928 229522 283937
rect 229204 283886 229466 283914
rect 227994 283863 228050 283872
rect 231320 283914 231348 288390
rect 231688 284172 231716 309159
rect 232226 307728 232282 307737
rect 232226 307663 232282 307672
rect 232240 306513 232268 307663
rect 232226 306504 232282 306513
rect 232226 306439 232282 306448
rect 232240 284172 232268 306439
rect 232516 289785 232544 356623
rect 232608 342922 232636 361558
rect 232596 342916 232648 342922
rect 232596 342858 232648 342864
rect 232596 320952 232648 320958
rect 232596 320894 232648 320900
rect 232608 307737 232636 320894
rect 233896 319569 233924 375022
rect 234632 374134 234660 377590
rect 234620 374128 234672 374134
rect 234620 374070 234672 374076
rect 234632 373998 234660 374070
rect 234620 373992 234672 373998
rect 234620 373934 234672 373940
rect 235264 371748 235316 371754
rect 235264 371690 235316 371696
rect 234528 353320 234580 353326
rect 234528 353262 234580 353268
rect 234068 322244 234120 322250
rect 234068 322186 234120 322192
rect 233976 321632 234028 321638
rect 233976 321574 234028 321580
rect 233882 319560 233938 319569
rect 233882 319495 233938 319504
rect 232594 307728 232650 307737
rect 232594 307663 232650 307672
rect 233148 305040 233200 305046
rect 233148 304982 233200 304988
rect 233700 305040 233752 305046
rect 233700 304982 233752 304988
rect 233160 297498 233188 304982
rect 233148 297492 233200 297498
rect 233148 297434 233200 297440
rect 232594 296848 232650 296857
rect 232594 296783 232650 296792
rect 232502 289776 232558 289785
rect 232502 289711 232558 289720
rect 232608 287881 232636 296783
rect 232594 287872 232650 287881
rect 232594 287807 232650 287816
rect 232778 285968 232834 285977
rect 232778 285903 232834 285912
rect 232792 284172 232820 285903
rect 233148 285728 233200 285734
rect 233148 285670 233200 285676
rect 233160 284172 233188 285670
rect 233712 284172 233740 304982
rect 233988 285734 234016 321574
rect 234080 306374 234108 322186
rect 234080 306346 234292 306374
rect 234264 292602 234292 306346
rect 234540 305046 234568 353262
rect 235276 337521 235304 371690
rect 236012 338774 236040 377590
rect 238128 375086 238156 377604
rect 238772 377590 239798 377618
rect 240152 377590 241454 377618
rect 242912 377590 243110 377618
rect 244292 377590 244766 377618
rect 245672 377590 246422 377618
rect 238116 375080 238168 375086
rect 238116 375022 238168 375028
rect 238024 374128 238076 374134
rect 238024 374070 238076 374076
rect 236642 348392 236698 348401
rect 236642 348327 236698 348336
rect 236656 338774 236684 348327
rect 236000 338768 236052 338774
rect 236000 338710 236052 338716
rect 236644 338768 236696 338774
rect 236644 338710 236696 338716
rect 235262 337512 235318 337521
rect 235262 337447 235318 337456
rect 236642 330032 236698 330041
rect 236642 329967 236698 329976
rect 235264 329112 235316 329118
rect 235264 329054 235316 329060
rect 235276 311137 235304 329054
rect 236656 322998 236684 329967
rect 236644 322992 236696 322998
rect 236644 322934 236696 322940
rect 237288 322992 237340 322998
rect 237288 322934 237340 322940
rect 236000 313948 236052 313954
rect 236000 313890 236052 313896
rect 235262 311128 235318 311137
rect 235262 311063 235318 311072
rect 235538 311128 235594 311137
rect 235538 311063 235594 311072
rect 234528 305040 234580 305046
rect 234528 304982 234580 304988
rect 234620 304360 234672 304366
rect 234620 304302 234672 304308
rect 234632 303686 234660 304302
rect 234620 303680 234672 303686
rect 234620 303622 234672 303628
rect 234252 292596 234304 292602
rect 234252 292538 234304 292544
rect 233976 285728 234028 285734
rect 233976 285670 234028 285676
rect 234264 284172 234292 292538
rect 234632 284172 234660 303622
rect 235172 288924 235224 288930
rect 235172 288866 235224 288872
rect 234710 286376 234766 286385
rect 234710 286311 234766 286320
rect 234724 285054 234752 286311
rect 234712 285048 234764 285054
rect 234712 284990 234764 284996
rect 235184 284172 235212 288866
rect 235448 285796 235500 285802
rect 235448 285738 235500 285744
rect 235460 284986 235488 285738
rect 235448 284980 235500 284986
rect 235448 284922 235500 284928
rect 235552 284172 235580 311063
rect 236012 289105 236040 313890
rect 236092 295996 236144 296002
rect 236092 295938 236144 295944
rect 235998 289096 236054 289105
rect 235998 289031 236054 289040
rect 236012 288930 236040 289031
rect 236000 288924 236052 288930
rect 236000 288866 236052 288872
rect 236104 287054 236132 295938
rect 236642 289776 236698 289785
rect 236642 289711 236698 289720
rect 236104 287026 236408 287054
rect 236092 285728 236144 285734
rect 236092 285670 236144 285676
rect 236104 284172 236132 285670
rect 236380 283937 236408 287026
rect 236656 285705 236684 289711
rect 237300 285734 237328 322934
rect 238036 313954 238064 374070
rect 238772 371754 238800 377590
rect 238760 371748 238812 371754
rect 238760 371690 238812 371696
rect 238116 357400 238168 357406
rect 238116 357342 238168 357348
rect 238128 325009 238156 357342
rect 240152 353326 240180 377590
rect 242912 371385 242940 377590
rect 242898 371376 242954 371385
rect 242898 371311 242954 371320
rect 243634 371376 243690 371385
rect 243634 371311 243690 371320
rect 242164 370524 242216 370530
rect 242164 370466 242216 370472
rect 240140 353320 240192 353326
rect 240140 353262 240192 353268
rect 241428 348492 241480 348498
rect 241428 348434 241480 348440
rect 240876 347064 240928 347070
rect 240876 347006 240928 347012
rect 240140 346384 240192 346390
rect 240140 346326 240192 346332
rect 238942 334248 238998 334257
rect 238942 334183 238998 334192
rect 238666 327312 238722 327321
rect 238666 327247 238722 327256
rect 238680 325718 238708 327247
rect 238668 325712 238720 325718
rect 238668 325654 238720 325660
rect 238114 325000 238170 325009
rect 238114 324935 238170 324944
rect 238024 313948 238076 313954
rect 238024 313890 238076 313896
rect 237378 287328 237434 287337
rect 237378 287263 237434 287272
rect 237288 285728 237340 285734
rect 236642 285696 236698 285705
rect 237288 285670 237340 285676
rect 237392 285666 237420 287263
rect 238680 285870 238708 325654
rect 237564 285864 237616 285870
rect 237564 285806 237616 285812
rect 238668 285864 238720 285870
rect 238668 285806 238720 285812
rect 236642 285631 236698 285640
rect 237380 285660 237432 285666
rect 236656 284172 236684 285631
rect 237380 285602 237432 285608
rect 237576 284172 237604 285806
rect 238484 285728 238536 285734
rect 238484 285670 238536 285676
rect 238114 284472 238170 284481
rect 238114 284407 238170 284416
rect 238128 284172 238156 284407
rect 238496 284172 238524 285670
rect 238956 285666 238984 334183
rect 239126 331936 239182 331945
rect 239126 331871 239182 331880
rect 239140 327758 239168 331871
rect 239128 327752 239180 327758
rect 239128 327694 239180 327700
rect 239036 309868 239088 309874
rect 239036 309810 239088 309816
rect 240048 309868 240100 309874
rect 240048 309810 240100 309816
rect 238944 285660 238996 285666
rect 238944 285602 238996 285608
rect 239048 284172 239076 309810
rect 240060 309194 240088 309810
rect 240048 309188 240100 309194
rect 240048 309130 240100 309136
rect 240152 306374 240180 346326
rect 240784 343664 240836 343670
rect 240784 343606 240836 343612
rect 240796 307086 240824 343606
rect 240888 316742 240916 347006
rect 241440 346390 241468 348434
rect 241428 346384 241480 346390
rect 241428 346326 241480 346332
rect 241978 326496 242034 326505
rect 241978 326431 242034 326440
rect 241992 320210 242020 326431
rect 241980 320204 242032 320210
rect 241980 320146 242032 320152
rect 240968 317484 241020 317490
rect 240968 317426 241020 317432
rect 240876 316736 240928 316742
rect 240876 316678 240928 316684
rect 240784 307080 240836 307086
rect 240784 307022 240836 307028
rect 240152 306346 240640 306374
rect 239954 292632 240010 292641
rect 239954 292567 240010 292576
rect 239218 289368 239274 289377
rect 239218 289303 239274 289312
rect 239232 287745 239260 289303
rect 239218 287736 239274 287745
rect 239218 287671 239274 287680
rect 239588 285660 239640 285666
rect 239588 285602 239640 285608
rect 239600 284172 239628 285602
rect 239968 284172 239996 292567
rect 240508 289128 240560 289134
rect 240508 289070 240560 289076
rect 240520 284172 240548 289070
rect 240612 284186 240640 306346
rect 240980 289785 241008 317426
rect 241426 293992 241482 294001
rect 241426 293927 241482 293936
rect 241440 291242 241468 293927
rect 241428 291236 241480 291242
rect 241428 291178 241480 291184
rect 240966 289776 241022 289785
rect 240966 289711 241022 289720
rect 240612 284158 240902 284186
rect 241440 284172 241468 291178
rect 241992 284172 242020 320146
rect 242176 295361 242204 370466
rect 243542 344312 243598 344321
rect 243542 344247 243598 344256
rect 242254 323640 242310 323649
rect 242254 323575 242310 323584
rect 242268 295934 242296 323575
rect 242256 295928 242308 295934
rect 242256 295870 242308 295876
rect 243452 295928 243504 295934
rect 243452 295870 243504 295876
rect 243464 295458 243492 295870
rect 243452 295452 243504 295458
rect 243452 295394 243504 295400
rect 242162 295352 242218 295361
rect 242162 295287 242218 295296
rect 242176 284186 242204 295287
rect 242806 293992 242862 294001
rect 242806 293927 242862 293936
rect 242820 289649 242848 293927
rect 242806 289640 242862 289649
rect 242806 289575 242862 289584
rect 242820 289241 242848 289575
rect 242806 289232 242862 289241
rect 242806 289167 242862 289176
rect 242898 288416 242954 288425
rect 242898 288351 242954 288360
rect 242912 287201 242940 288351
rect 242898 287192 242954 287201
rect 242898 287127 242954 287136
rect 242176 284158 242374 284186
rect 242912 284172 242940 287127
rect 243464 284172 243492 295394
rect 243556 288425 243584 344247
rect 243648 341601 243676 371311
rect 244292 347750 244320 377590
rect 245014 363624 245070 363633
rect 245014 363559 245070 363568
rect 244280 347744 244332 347750
rect 244280 347686 244332 347692
rect 244924 347744 244976 347750
rect 244924 347686 244976 347692
rect 243634 341592 243690 341601
rect 243634 341527 243690 341536
rect 244738 326360 244794 326369
rect 244738 326295 244794 326304
rect 243636 323060 243688 323066
rect 243636 323002 243688 323008
rect 243648 308553 243676 323002
rect 244752 322833 244780 326295
rect 244738 322824 244794 322833
rect 244738 322759 244794 322768
rect 244752 321745 244780 322759
rect 244738 321736 244794 321745
rect 244738 321671 244794 321680
rect 243634 308544 243690 308553
rect 243634 308479 243690 308488
rect 244280 308440 244332 308446
rect 244280 308382 244332 308388
rect 243818 289640 243874 289649
rect 243818 289575 243874 289584
rect 243542 288416 243598 288425
rect 243542 288351 243598 288360
rect 243832 284172 243860 289575
rect 244002 287328 244058 287337
rect 244002 287263 244058 287272
rect 244016 284889 244044 287263
rect 244188 285796 244240 285802
rect 244188 285738 244240 285744
rect 244094 285016 244150 285025
rect 244094 284951 244150 284960
rect 244002 284880 244058 284889
rect 244002 284815 244058 284824
rect 244002 284336 244058 284345
rect 244002 284271 244058 284280
rect 231490 283928 231546 283937
rect 231320 283900 231490 283914
rect 231334 283886 231490 283900
rect 229466 283863 229522 283872
rect 231490 283863 231546 283872
rect 236366 283928 236422 283937
rect 236366 283863 236422 283872
rect 236734 283928 236790 283937
rect 236790 283886 237038 283914
rect 236734 283863 236790 283872
rect 200026 280256 200082 280265
rect 200026 280191 200082 280200
rect 244016 277394 244044 284271
rect 244108 284073 244136 284951
rect 244094 284064 244150 284073
rect 244094 283999 244150 284008
rect 244200 283626 244228 285738
rect 244188 283620 244240 283626
rect 244188 283562 244240 283568
rect 244292 278089 244320 308382
rect 244936 300830 244964 347686
rect 245028 330614 245056 363559
rect 245672 355434 245700 377590
rect 248064 376038 248092 377604
rect 247040 376032 247092 376038
rect 247040 375974 247092 375980
rect 248052 376032 248104 376038
rect 248052 375974 248104 375980
rect 247052 375329 247080 375974
rect 247038 375320 247094 375329
rect 247038 375255 247094 375264
rect 246396 374128 246448 374134
rect 246396 374070 246448 374076
rect 245660 355428 245712 355434
rect 245660 355370 245712 355376
rect 246302 351928 246358 351937
rect 246302 351863 246358 351872
rect 245108 341556 245160 341562
rect 245108 341498 245160 341504
rect 245016 330608 245068 330614
rect 245016 330550 245068 330556
rect 245120 319530 245148 341498
rect 245108 319524 245160 319530
rect 245108 319466 245160 319472
rect 245660 316124 245712 316130
rect 245660 316066 245712 316072
rect 245672 311846 245700 316066
rect 245660 311840 245712 311846
rect 245660 311782 245712 311788
rect 244924 300824 244976 300830
rect 244924 300766 244976 300772
rect 244372 299600 244424 299606
rect 244372 299542 244424 299548
rect 244384 298790 244412 299542
rect 244372 298784 244424 298790
rect 244372 298726 244424 298732
rect 244464 298716 244516 298722
rect 244464 298658 244516 298664
rect 244370 282432 244426 282441
rect 244370 282367 244426 282376
rect 244278 278080 244334 278089
rect 244278 278015 244334 278024
rect 244016 277366 244136 277394
rect 199934 276720 199990 276729
rect 199934 276655 199990 276664
rect 199476 272536 199528 272542
rect 199476 272478 199528 272484
rect 199842 270192 199898 270201
rect 199842 270127 199898 270136
rect 199384 257372 199436 257378
rect 199384 257314 199436 257320
rect 198476 248386 198596 248414
rect 197358 247888 197414 247897
rect 197358 247823 197414 247832
rect 197372 247110 197400 247823
rect 197360 247104 197412 247110
rect 197360 247046 197412 247052
rect 197726 245168 197782 245177
rect 197726 245103 197782 245112
rect 197740 244934 197768 245103
rect 197728 244928 197780 244934
rect 197728 244870 197780 244876
rect 198568 244361 198596 248386
rect 198832 245676 198884 245682
rect 198832 245618 198884 245624
rect 198646 245168 198702 245177
rect 198646 245103 198702 245112
rect 198554 244352 198610 244361
rect 198554 244287 198610 244296
rect 197360 244248 197412 244254
rect 197360 244190 197412 244196
rect 197372 243817 197400 244190
rect 197358 243808 197414 243817
rect 197358 243743 197414 243752
rect 197358 242176 197414 242185
rect 197358 242111 197414 242120
rect 197372 241534 197400 242111
rect 197360 241528 197412 241534
rect 197360 241470 197412 241476
rect 198568 238754 198596 244287
rect 198660 243114 198688 245103
rect 198660 243086 198780 243114
rect 198752 240417 198780 243086
rect 198844 241641 198872 245618
rect 199750 241904 199806 241913
rect 199750 241839 199806 241848
rect 198830 241632 198886 241641
rect 198830 241567 198886 241576
rect 199566 240680 199622 240689
rect 199566 240615 199622 240624
rect 198738 240408 198794 240417
rect 199580 240378 199608 240615
rect 199658 240544 199714 240553
rect 199658 240479 199714 240488
rect 199672 240446 199700 240479
rect 199660 240440 199712 240446
rect 199660 240382 199712 240388
rect 198738 240343 198794 240352
rect 199568 240372 199620 240378
rect 199568 240314 199620 240320
rect 199764 240145 199792 241839
rect 199750 240136 199806 240145
rect 199750 240071 199806 240080
rect 198568 238726 198688 238754
rect 198002 214704 198058 214713
rect 198002 214639 198058 214648
rect 198016 191146 198044 214639
rect 198004 191140 198056 191146
rect 198004 191082 198056 191088
rect 197266 183016 197322 183025
rect 197266 182951 197322 182960
rect 196808 178696 196860 178702
rect 196808 178638 196860 178644
rect 198096 178084 198148 178090
rect 198096 178026 198148 178032
rect 196714 177168 196770 177177
rect 196714 177103 196770 177112
rect 196728 160002 196756 177103
rect 198004 173188 198056 173194
rect 198004 173130 198056 173136
rect 198016 163538 198044 173130
rect 198108 169658 198136 178026
rect 198660 177342 198688 238726
rect 199384 236768 199436 236774
rect 199384 236710 199436 236716
rect 198740 231736 198792 231742
rect 198740 231678 198792 231684
rect 198752 231198 198780 231678
rect 198740 231192 198792 231198
rect 198740 231134 198792 231140
rect 198738 225040 198794 225049
rect 198738 224975 198794 224984
rect 198752 193118 198780 224975
rect 198830 204368 198886 204377
rect 198830 204303 198886 204312
rect 198844 204105 198872 204303
rect 198830 204096 198886 204105
rect 198830 204031 198886 204040
rect 198740 193112 198792 193118
rect 198740 193054 198792 193060
rect 198752 192574 198780 193054
rect 198740 192568 198792 192574
rect 198740 192510 198792 192516
rect 199396 182918 199424 236710
rect 199856 231198 199884 270127
rect 199948 236706 199976 276655
rect 200026 273728 200082 273737
rect 200026 273663 200082 273672
rect 199936 236700 199988 236706
rect 199936 236642 199988 236648
rect 199844 231192 199896 231198
rect 199844 231134 199896 231140
rect 199476 220720 199528 220726
rect 199476 220662 199528 220668
rect 199488 191214 199516 220662
rect 200040 219502 200068 273663
rect 244108 263430 244136 277366
rect 244280 270224 244332 270230
rect 244278 270192 244280 270201
rect 244332 270192 244334 270201
rect 244278 270127 244334 270136
rect 244096 263424 244148 263430
rect 244096 263366 244148 263372
rect 244002 254688 244058 254697
rect 244002 254623 244058 254632
rect 200120 240848 200172 240854
rect 200120 240790 200172 240796
rect 200132 237386 200160 240790
rect 200224 240145 200252 240244
rect 200210 240136 200266 240145
rect 200210 240071 200266 240080
rect 200224 237425 200252 240071
rect 200592 240009 200620 240244
rect 201038 240136 201094 240145
rect 201144 240122 201172 240244
rect 201224 240168 201276 240174
rect 201144 240116 201224 240122
rect 201144 240110 201276 240116
rect 201144 240094 201264 240110
rect 201038 240071 201094 240080
rect 200578 240000 200634 240009
rect 200578 239935 200634 239944
rect 200210 237416 200266 237425
rect 200120 237380 200172 237386
rect 200210 237351 200266 237360
rect 200120 237322 200172 237328
rect 200764 236700 200816 236706
rect 200764 236642 200816 236648
rect 200028 219496 200080 219502
rect 200028 219438 200080 219444
rect 200776 194546 200804 236642
rect 201052 229094 201080 240071
rect 201236 238754 201264 240094
rect 201406 240000 201462 240009
rect 201406 239935 201462 239944
rect 201236 238726 201356 238754
rect 201052 229066 201172 229094
rect 201144 214674 201172 229066
rect 201132 214668 201184 214674
rect 201132 214610 201184 214616
rect 201328 196722 201356 238726
rect 201420 237402 201448 239935
rect 201512 238754 201540 240244
rect 201512 238726 201632 238754
rect 201420 237374 201540 237402
rect 201406 237280 201462 237289
rect 201406 237215 201462 237224
rect 201316 196716 201368 196722
rect 201316 196658 201368 196664
rect 200764 194540 200816 194546
rect 200764 194482 200816 194488
rect 199476 191208 199528 191214
rect 199476 191150 199528 191156
rect 201420 187241 201448 237215
rect 201512 233889 201540 237374
rect 201604 234297 201632 238726
rect 202064 237969 202092 240244
rect 202328 240168 202380 240174
rect 202616 240145 202644 240244
rect 202328 240110 202380 240116
rect 202602 240136 202658 240145
rect 202050 237960 202106 237969
rect 202050 237895 202106 237904
rect 202144 237448 202196 237454
rect 202144 237390 202196 237396
rect 201590 234288 201646 234297
rect 201590 234223 201646 234232
rect 201498 233880 201554 233889
rect 201498 233815 201554 233824
rect 201498 229936 201554 229945
rect 201498 229871 201554 229880
rect 201512 222902 201540 229871
rect 201500 222896 201552 222902
rect 201500 222838 201552 222844
rect 201500 219496 201552 219502
rect 201500 219438 201552 219444
rect 201512 198694 201540 219438
rect 201590 210352 201646 210361
rect 201590 210287 201646 210296
rect 201604 206417 201632 210287
rect 201590 206408 201646 206417
rect 201590 206343 201646 206352
rect 201500 198688 201552 198694
rect 201500 198630 201552 198636
rect 202156 198014 202184 237390
rect 202234 233880 202290 233889
rect 202234 233815 202290 233824
rect 202248 213926 202276 233815
rect 202340 230382 202368 240110
rect 202602 240071 202658 240080
rect 202616 238746 202644 240071
rect 202984 238754 203012 240244
rect 202604 238740 202656 238746
rect 202984 238726 203104 238754
rect 202604 238682 202656 238688
rect 202616 237454 202644 238682
rect 202604 237448 202656 237454
rect 202604 237390 202656 237396
rect 202880 237448 202932 237454
rect 202880 237390 202932 237396
rect 202788 237312 202840 237318
rect 202786 237280 202788 237289
rect 202840 237280 202842 237289
rect 202786 237215 202842 237224
rect 202418 234288 202474 234297
rect 202418 234223 202474 234232
rect 202328 230376 202380 230382
rect 202328 230318 202380 230324
rect 202236 213920 202288 213926
rect 202236 213862 202288 213868
rect 202144 198008 202196 198014
rect 202144 197950 202196 197956
rect 202248 196761 202276 213862
rect 202432 213246 202460 234223
rect 202892 231169 202920 237390
rect 202878 231160 202934 231169
rect 202878 231095 202934 231104
rect 203076 221882 203104 238726
rect 203536 237017 203564 240244
rect 203984 240168 204036 240174
rect 204088 240122 204116 240244
rect 204036 240116 204116 240122
rect 203984 240110 204116 240116
rect 203996 240094 204116 240110
rect 203522 237008 203578 237017
rect 203522 236943 203578 236952
rect 203064 221876 203116 221882
rect 203064 221818 203116 221824
rect 203076 221474 203104 221818
rect 203064 221468 203116 221474
rect 203064 221410 203116 221416
rect 202420 213240 202472 213246
rect 202420 213182 202472 213188
rect 202418 196888 202474 196897
rect 202418 196823 202474 196832
rect 202234 196752 202290 196761
rect 202234 196687 202290 196696
rect 202144 189848 202196 189854
rect 202432 189825 202460 196823
rect 202144 189790 202196 189796
rect 202418 189816 202474 189825
rect 201406 187232 201462 187241
rect 201406 187167 201462 187176
rect 199384 182912 199436 182918
rect 199384 182854 199436 182860
rect 200764 182844 200816 182850
rect 200764 182786 200816 182792
rect 198648 177336 198700 177342
rect 198648 177278 198700 177284
rect 198096 169652 198148 169658
rect 198096 169594 198148 169600
rect 198004 163532 198056 163538
rect 198004 163474 198056 163480
rect 196716 159996 196768 160002
rect 196716 159938 196768 159944
rect 198096 150476 198148 150482
rect 198096 150418 198148 150424
rect 196716 135992 196768 135998
rect 196716 135934 196768 135940
rect 196728 101522 196756 135934
rect 198004 127016 198056 127022
rect 198004 126958 198056 126964
rect 196808 121576 196860 121582
rect 196808 121518 196860 121524
rect 196716 101516 196768 101522
rect 196716 101458 196768 101464
rect 196820 93673 196848 121518
rect 196900 100768 196952 100774
rect 196900 100710 196952 100716
rect 196806 93664 196862 93673
rect 196806 93599 196862 93608
rect 196912 87718 196940 100710
rect 196900 87712 196952 87718
rect 196900 87654 196952 87660
rect 196808 87644 196860 87650
rect 196808 87586 196860 87592
rect 196622 3904 196678 3913
rect 196622 3839 196678 3848
rect 196820 3369 196848 87586
rect 198016 60722 198044 126958
rect 198108 116618 198136 150418
rect 199474 127256 199530 127265
rect 199474 127191 199530 127200
rect 199382 124808 199438 124817
rect 199382 124743 199438 124752
rect 198280 117428 198332 117434
rect 198280 117370 198332 117376
rect 198096 116612 198148 116618
rect 198096 116554 198148 116560
rect 198096 114572 198148 114578
rect 198096 114514 198148 114520
rect 198108 85377 198136 114514
rect 198188 104916 198240 104922
rect 198188 104858 198240 104864
rect 198094 85368 198150 85377
rect 198094 85303 198150 85312
rect 198096 82204 198148 82210
rect 198096 82146 198148 82152
rect 198004 60716 198056 60722
rect 198004 60658 198056 60664
rect 198108 18630 198136 82146
rect 198200 77217 198228 104858
rect 198292 104242 198320 117370
rect 198646 104816 198702 104825
rect 198646 104751 198702 104760
rect 198280 104236 198332 104242
rect 198280 104178 198332 104184
rect 198660 96014 198688 104751
rect 198648 96008 198700 96014
rect 198648 95950 198700 95956
rect 198186 77208 198242 77217
rect 198186 77143 198242 77152
rect 199396 68950 199424 124743
rect 199488 80073 199516 127191
rect 199474 80064 199530 80073
rect 200776 80034 200804 182786
rect 200856 129804 200908 129810
rect 200856 129746 200908 129752
rect 200868 115258 200896 129746
rect 200948 116068 201000 116074
rect 200948 116010 201000 116016
rect 200856 115252 200908 115258
rect 200856 115194 200908 115200
rect 200856 93152 200908 93158
rect 200856 93094 200908 93100
rect 199474 79999 199530 80008
rect 200764 80028 200816 80034
rect 200764 79970 200816 79976
rect 199384 68944 199436 68950
rect 199384 68886 199436 68892
rect 200868 62082 200896 93094
rect 200960 89729 200988 116010
rect 200946 89720 201002 89729
rect 200946 89655 201002 89664
rect 200856 62076 200908 62082
rect 200856 62018 200908 62024
rect 202156 18630 202184 189790
rect 202418 189751 202474 189760
rect 202236 151088 202288 151094
rect 202236 151030 202288 151036
rect 202248 90409 202276 151030
rect 202420 128376 202472 128382
rect 202420 128318 202472 128324
rect 202328 94512 202380 94518
rect 202328 94454 202380 94460
rect 202234 90400 202290 90409
rect 202234 90335 202290 90344
rect 202340 57934 202368 94454
rect 202432 93945 202460 128318
rect 202418 93936 202474 93945
rect 202418 93871 202474 93880
rect 203536 85542 203564 236943
rect 204088 231130 204116 240094
rect 204076 231124 204128 231130
rect 204076 231066 204128 231072
rect 204166 228440 204222 228449
rect 204166 228375 204222 228384
rect 204180 226001 204208 228375
rect 204456 227361 204484 240244
rect 205008 237454 205036 240244
rect 204996 237448 205048 237454
rect 204996 237390 205048 237396
rect 205376 233170 205404 240244
rect 205928 238754 205956 240244
rect 205836 238726 205956 238754
rect 205836 238649 205864 238726
rect 205822 238640 205878 238649
rect 205822 238575 205878 238584
rect 205640 235272 205692 235278
rect 205638 235240 205640 235249
rect 205692 235240 205694 235249
rect 205638 235175 205694 235184
rect 205364 233164 205416 233170
rect 205364 233106 205416 233112
rect 204442 227352 204498 227361
rect 204442 227287 204498 227296
rect 204456 226409 204484 227287
rect 204442 226400 204498 226409
rect 204442 226335 204498 226344
rect 204904 226364 204956 226370
rect 204904 226306 204956 226312
rect 204166 225992 204222 226001
rect 204166 225927 204222 225936
rect 203616 221876 203668 221882
rect 203616 221818 203668 221824
rect 203628 210361 203656 221818
rect 203614 210352 203670 210361
rect 203614 210287 203670 210296
rect 204720 209092 204772 209098
rect 204720 209034 204772 209040
rect 204732 206961 204760 209034
rect 204718 206952 204774 206961
rect 204718 206887 204774 206896
rect 203616 200864 203668 200870
rect 203616 200806 203668 200812
rect 203628 175137 203656 200806
rect 204260 194540 204312 194546
rect 204260 194482 204312 194488
rect 204272 192506 204300 194482
rect 204916 193225 204944 226306
rect 205376 219434 205404 233106
rect 205640 231600 205692 231606
rect 205640 231542 205692 231548
rect 205008 219406 205404 219434
rect 204902 193216 204958 193225
rect 204902 193151 204958 193160
rect 204260 192500 204312 192506
rect 204260 192442 204312 192448
rect 204904 188352 204956 188358
rect 204904 188294 204956 188300
rect 204916 184278 204944 188294
rect 204168 184272 204220 184278
rect 204168 184214 204220 184220
rect 204904 184272 204956 184278
rect 204904 184214 204956 184220
rect 204180 183530 204208 184214
rect 204168 183524 204220 183530
rect 204168 183466 204220 183472
rect 204904 181552 204956 181558
rect 204904 181494 204956 181500
rect 203614 175128 203670 175137
rect 203614 175063 203670 175072
rect 203708 118788 203760 118794
rect 203708 118730 203760 118736
rect 203616 114640 203668 114646
rect 203616 114582 203668 114588
rect 203524 85536 203576 85542
rect 203524 85478 203576 85484
rect 202328 57928 202380 57934
rect 202328 57870 202380 57876
rect 203628 55214 203656 114582
rect 203720 84114 203748 118730
rect 203708 84108 203760 84114
rect 203708 84050 203760 84056
rect 203616 55208 203668 55214
rect 203616 55150 203668 55156
rect 204916 22681 204944 181494
rect 205008 81394 205036 219406
rect 205652 213874 205680 231542
rect 205836 229094 205864 238575
rect 206376 234660 206428 234666
rect 206376 234602 206428 234608
rect 205836 229066 206324 229094
rect 205560 213846 205680 213874
rect 205086 200968 205142 200977
rect 205086 200903 205142 200912
rect 205100 186969 205128 200903
rect 205560 200190 205588 213846
rect 205638 213752 205694 213761
rect 205638 213687 205694 213696
rect 205652 213314 205680 213687
rect 205640 213308 205692 213314
rect 205640 213250 205692 213256
rect 206296 209545 206324 229066
rect 206282 209536 206338 209545
rect 206282 209471 206338 209480
rect 205548 200184 205600 200190
rect 205548 200126 205600 200132
rect 206296 193934 206324 209471
rect 206284 193928 206336 193934
rect 206284 193870 206336 193876
rect 205640 187740 205692 187746
rect 205640 187682 205692 187688
rect 205086 186960 205142 186969
rect 205086 186895 205142 186904
rect 205652 186289 205680 187682
rect 206284 187060 206336 187066
rect 206284 187002 206336 187008
rect 205638 186280 205694 186289
rect 205638 186215 205694 186224
rect 205272 140820 205324 140826
rect 205272 140762 205324 140768
rect 205180 128444 205232 128450
rect 205180 128386 205232 128392
rect 205088 106412 205140 106418
rect 205088 106354 205140 106360
rect 204996 81388 205048 81394
rect 204996 81330 205048 81336
rect 205100 67522 205128 106354
rect 205192 93809 205220 128386
rect 205284 106962 205312 140762
rect 205272 106956 205324 106962
rect 205272 106898 205324 106904
rect 205178 93800 205234 93809
rect 205178 93735 205234 93744
rect 205088 67516 205140 67522
rect 205088 67458 205140 67464
rect 206296 55185 206324 187002
rect 206388 181558 206416 234602
rect 206480 231606 206508 240244
rect 206848 235890 206876 240244
rect 207400 238754 207428 240244
rect 207952 240145 207980 240244
rect 208320 240145 208348 240244
rect 208400 240168 208452 240174
rect 207938 240136 207994 240145
rect 207938 240071 207994 240080
rect 208306 240136 208362 240145
rect 208400 240110 208452 240116
rect 208306 240071 208362 240080
rect 207400 238726 207704 238754
rect 207112 237448 207164 237454
rect 207112 237390 207164 237396
rect 206836 235884 206888 235890
rect 206836 235826 206888 235832
rect 206848 234666 206876 235826
rect 206836 234660 206888 234666
rect 206836 234602 206888 234608
rect 206468 231600 206520 231606
rect 206468 231542 206520 231548
rect 206468 214668 206520 214674
rect 206468 214610 206520 214616
rect 206480 200122 206508 214610
rect 207124 206825 207152 237390
rect 207676 237153 207704 238726
rect 207952 237454 207980 240071
rect 208320 238241 208348 240071
rect 208306 238232 208362 238241
rect 208306 238167 208362 238176
rect 207940 237448 207992 237454
rect 207940 237390 207992 237396
rect 207662 237144 207718 237153
rect 207662 237079 207718 237088
rect 207572 230376 207624 230382
rect 207572 230318 207624 230324
rect 207584 228449 207612 230318
rect 207570 228440 207626 228449
rect 207570 228375 207626 228384
rect 207676 218754 207704 237079
rect 208320 236706 208348 238167
rect 208412 237289 208440 240110
rect 208872 238754 208900 240244
rect 208872 238726 209084 238754
rect 208398 237280 208454 237289
rect 208398 237215 208454 237224
rect 208308 236700 208360 236706
rect 208308 236642 208360 236648
rect 208400 230988 208452 230994
rect 208400 230930 208452 230936
rect 208412 229094 208440 230930
rect 208412 229066 208532 229094
rect 208400 221468 208452 221474
rect 208400 221410 208452 221416
rect 207664 218748 207716 218754
rect 207664 218690 207716 218696
rect 208412 218006 208440 221410
rect 208504 219065 208532 229066
rect 209056 228993 209084 238726
rect 209240 230994 209268 240244
rect 209688 237448 209740 237454
rect 209688 237390 209740 237396
rect 209228 230988 209280 230994
rect 209228 230930 209280 230936
rect 209700 229129 209728 237390
rect 209686 229120 209742 229129
rect 209686 229055 209742 229064
rect 209042 228984 209098 228993
rect 209042 228919 209098 228928
rect 208490 219056 208546 219065
rect 208490 218991 208546 219000
rect 208400 218000 208452 218006
rect 208400 217942 208452 217948
rect 208504 214985 208532 218991
rect 208490 214976 208546 214985
rect 208490 214911 208546 214920
rect 207110 206816 207166 206825
rect 207110 206751 207166 206760
rect 207124 205737 207152 206751
rect 207110 205728 207166 205737
rect 207110 205663 207166 205672
rect 207662 205728 207718 205737
rect 207662 205663 207718 205672
rect 206468 200116 206520 200122
rect 206468 200058 206520 200064
rect 207676 185638 207704 205663
rect 209056 200841 209084 228919
rect 209700 226370 209728 229055
rect 209688 226364 209740 226370
rect 209688 226306 209740 226312
rect 209792 220697 209820 240244
rect 210344 237454 210372 240244
rect 210712 240145 210740 240244
rect 210698 240136 210754 240145
rect 210698 240071 210754 240080
rect 210332 237448 210384 237454
rect 210712 237425 210740 240071
rect 210332 237390 210384 237396
rect 210698 237416 210754 237425
rect 210698 237351 210754 237360
rect 211264 235521 211292 240244
rect 211250 235512 211306 235521
rect 211250 235447 211306 235456
rect 210608 233980 210660 233986
rect 210608 233922 210660 233928
rect 209778 220688 209834 220697
rect 209778 220623 209834 220632
rect 210422 220688 210478 220697
rect 210422 220623 210478 220632
rect 209686 215112 209742 215121
rect 209686 215047 209742 215056
rect 209042 200832 209098 200841
rect 209042 200767 209098 200776
rect 209228 193860 209280 193866
rect 209228 193802 209280 193808
rect 207664 185632 207716 185638
rect 207664 185574 207716 185580
rect 206376 181552 206428 181558
rect 206376 181494 206428 181500
rect 209042 178936 209098 178945
rect 209042 178871 209098 178880
rect 206374 135552 206430 135561
rect 206374 135487 206430 135496
rect 206388 94489 206416 135487
rect 206468 130416 206520 130422
rect 206468 130358 206520 130364
rect 206374 94480 206430 94489
rect 206374 94415 206430 94424
rect 206480 93809 206508 130358
rect 207756 124296 207808 124302
rect 207756 124238 207808 124244
rect 207664 107772 207716 107778
rect 207664 107714 207716 107720
rect 206466 93800 206522 93809
rect 206466 93735 206522 93744
rect 206376 90364 206428 90370
rect 206376 90306 206428 90312
rect 206282 55176 206338 55185
rect 206282 55111 206338 55120
rect 206388 36650 206416 90306
rect 207676 66230 207704 107714
rect 207768 90982 207796 124238
rect 207756 90976 207808 90982
rect 207756 90918 207808 90924
rect 207664 66224 207716 66230
rect 207664 66166 207716 66172
rect 209056 37262 209084 178871
rect 209240 178809 209268 193802
rect 209226 178800 209282 178809
rect 209226 178735 209282 178744
rect 209228 142248 209280 142254
rect 209228 142190 209280 142196
rect 209136 132592 209188 132598
rect 209136 132534 209188 132540
rect 209148 92313 209176 132534
rect 209240 124817 209268 142190
rect 209226 124808 209282 124817
rect 209226 124743 209282 124752
rect 209318 118008 209374 118017
rect 209318 117943 209374 117952
rect 209332 92449 209360 117943
rect 209700 92478 209728 215047
rect 210436 206281 210464 220623
rect 210620 220153 210648 233922
rect 211816 233170 211844 240244
rect 211894 236056 211950 236065
rect 211894 235991 211950 236000
rect 211804 233164 211856 233170
rect 211804 233106 211856 233112
rect 211908 223582 211936 235991
rect 211896 223576 211948 223582
rect 211896 223518 211948 223524
rect 210606 220144 210662 220153
rect 210606 220079 210662 220088
rect 210422 206272 210478 206281
rect 210422 206207 210478 206216
rect 211804 202836 211856 202842
rect 211804 202778 211856 202784
rect 210422 201104 210478 201113
rect 210422 201039 210478 201048
rect 210436 177449 210464 201039
rect 210422 177440 210478 177449
rect 210422 177375 210478 177384
rect 210424 133952 210476 133958
rect 210424 133894 210476 133900
rect 210436 93158 210464 133894
rect 210516 129872 210568 129878
rect 210516 129814 210568 129820
rect 210424 93152 210476 93158
rect 210424 93094 210476 93100
rect 209688 92472 209740 92478
rect 209318 92440 209374 92449
rect 209688 92414 209740 92420
rect 209318 92375 209374 92384
rect 209134 92304 209190 92313
rect 209134 92239 209190 92248
rect 210528 91633 210556 129814
rect 210606 98696 210662 98705
rect 210606 98631 210662 98640
rect 210514 91624 210570 91633
rect 210514 91559 210570 91568
rect 209136 89004 209188 89010
rect 209136 88946 209188 88952
rect 209044 37256 209096 37262
rect 209044 37198 209096 37204
rect 206376 36644 206428 36650
rect 206376 36586 206428 36592
rect 209148 22846 209176 88946
rect 210424 84856 210476 84862
rect 210424 84798 210476 84804
rect 209136 22840 209188 22846
rect 209136 22782 209188 22788
rect 204902 22672 204958 22681
rect 204902 22607 204958 22616
rect 210436 18698 210464 84798
rect 210620 74526 210648 98631
rect 211816 95878 211844 202778
rect 211908 180169 211936 223518
rect 212184 202842 212212 240244
rect 212446 235512 212502 235521
rect 212446 235447 212502 235456
rect 212460 204270 212488 235447
rect 212736 207913 212764 240244
rect 212816 233164 212868 233170
rect 212816 233106 212868 233112
rect 212722 207904 212778 207913
rect 212722 207839 212778 207848
rect 212736 207097 212764 207839
rect 212722 207088 212778 207097
rect 212722 207023 212778 207032
rect 212448 204264 212500 204270
rect 212448 204206 212500 204212
rect 212460 203590 212488 204206
rect 212828 204202 212856 233106
rect 213104 229094 213132 240244
rect 213104 229066 213316 229094
rect 213184 225480 213236 225486
rect 213184 225422 213236 225428
rect 212816 204196 212868 204202
rect 212816 204138 212868 204144
rect 212448 203584 212500 203590
rect 212448 203526 212500 203532
rect 212172 202836 212224 202842
rect 212172 202778 212224 202784
rect 213196 202230 213224 225422
rect 213288 222154 213316 229066
rect 213656 226302 213684 240244
rect 214208 239426 214236 240244
rect 214196 239420 214248 239426
rect 214196 239362 214248 239368
rect 214208 231849 214236 239362
rect 214194 231840 214250 231849
rect 214194 231775 214250 231784
rect 213644 226296 213696 226302
rect 213644 226238 213696 226244
rect 213656 225486 213684 226238
rect 213644 225480 213696 225486
rect 213644 225422 213696 225428
rect 213276 222148 213328 222154
rect 213276 222090 213328 222096
rect 213288 212537 213316 222090
rect 214576 213761 214604 240244
rect 215128 240009 215156 240244
rect 215114 240000 215170 240009
rect 215114 239935 215170 239944
rect 215128 238754 215156 239935
rect 215128 238726 215248 238754
rect 214562 213752 214618 213761
rect 214562 213687 214618 213696
rect 213274 212528 213330 212537
rect 213274 212463 213330 212472
rect 215116 212424 215168 212430
rect 215116 212366 215168 212372
rect 215128 211818 215156 212366
rect 215116 211812 215168 211818
rect 215116 211754 215168 211760
rect 213274 207088 213330 207097
rect 213274 207023 213330 207032
rect 213184 202224 213236 202230
rect 213184 202166 213236 202172
rect 213288 198082 213316 207023
rect 214472 205624 214524 205630
rect 214470 205592 214472 205601
rect 214524 205592 214526 205601
rect 214470 205527 214526 205536
rect 214484 204338 214512 205527
rect 214472 204332 214524 204338
rect 214472 204274 214524 204280
rect 213828 204196 213880 204202
rect 213828 204138 213880 204144
rect 213840 203658 213868 204138
rect 213828 203652 213880 203658
rect 213828 203594 213880 203600
rect 215128 198082 215156 211754
rect 213276 198076 213328 198082
rect 213276 198018 213328 198024
rect 215116 198076 215168 198082
rect 215116 198018 215168 198024
rect 215220 180794 215248 238726
rect 215298 235784 215354 235793
rect 215298 235719 215354 235728
rect 215312 235249 215340 235719
rect 215298 235240 215354 235249
rect 215298 235175 215354 235184
rect 215300 233980 215352 233986
rect 215300 233922 215352 233928
rect 215312 231305 215340 233922
rect 215298 231296 215354 231305
rect 215298 231231 215354 231240
rect 215298 213888 215354 213897
rect 215298 213823 215354 213832
rect 215312 213314 215340 213823
rect 215300 213308 215352 213314
rect 215300 213250 215352 213256
rect 215298 212664 215354 212673
rect 215298 212599 215354 212608
rect 215312 211138 215340 212599
rect 215680 212430 215708 240244
rect 216048 232558 216076 240244
rect 216600 235249 216628 240244
rect 216678 237416 216734 237425
rect 216678 237351 216734 237360
rect 216586 235240 216642 235249
rect 216586 235175 216642 235184
rect 216036 232552 216088 232558
rect 216036 232494 216088 232500
rect 216048 229094 216076 232494
rect 215956 229066 216076 229094
rect 215956 214033 215984 229066
rect 216034 219464 216090 219473
rect 216034 219399 216090 219408
rect 215942 214024 215998 214033
rect 215942 213959 215998 213968
rect 215668 212424 215720 212430
rect 215668 212366 215720 212372
rect 215300 211132 215352 211138
rect 215300 211074 215352 211080
rect 215852 200184 215904 200190
rect 215852 200126 215904 200132
rect 215864 193905 215892 200126
rect 215850 193896 215906 193905
rect 215850 193831 215906 193840
rect 215128 180766 215248 180794
rect 214562 180704 214618 180713
rect 214562 180639 214618 180648
rect 211894 180160 211950 180169
rect 214576 180130 214604 180639
rect 211894 180095 211950 180104
rect 214564 180124 214616 180130
rect 214564 180066 214616 180072
rect 214104 179444 214156 179450
rect 214104 179386 214156 179392
rect 212448 176724 212500 176730
rect 212448 176666 212500 176672
rect 212460 173806 212488 176666
rect 213920 176656 213972 176662
rect 213920 176598 213972 176604
rect 213932 175681 213960 176598
rect 213918 175672 213974 175681
rect 213918 175607 213974 175616
rect 213920 175228 213972 175234
rect 213920 175170 213972 175176
rect 213932 175001 213960 175170
rect 214012 175160 214064 175166
rect 214012 175102 214064 175108
rect 213918 174992 213974 175001
rect 213918 174927 213974 174936
rect 214024 174321 214052 175102
rect 214010 174312 214066 174321
rect 214010 174247 214066 174256
rect 213920 173868 213972 173874
rect 213920 173810 213972 173816
rect 212448 173800 212500 173806
rect 212448 173742 212500 173748
rect 213932 173641 213960 173810
rect 214012 173800 214064 173806
rect 214012 173742 214064 173748
rect 213918 173632 213974 173641
rect 213918 173567 213974 173576
rect 214024 172961 214052 173742
rect 214010 172952 214066 172961
rect 214010 172887 214066 172896
rect 213920 172508 213972 172514
rect 213920 172450 213972 172456
rect 213932 172281 213960 172450
rect 213918 172272 213974 172281
rect 213918 172207 213974 172216
rect 214116 171601 214144 179386
rect 215128 178770 215156 180766
rect 215116 178764 215168 178770
rect 215116 178706 215168 178712
rect 215392 177404 215444 177410
rect 215392 177346 215444 177352
rect 214838 177304 214894 177313
rect 214838 177239 214894 177248
rect 214472 175976 214524 175982
rect 214472 175918 214524 175924
rect 214102 171592 214158 171601
rect 214102 171527 214158 171536
rect 214012 171080 214064 171086
rect 213918 171048 213974 171057
rect 214012 171022 214064 171028
rect 213918 170983 213920 170992
rect 213972 170983 213974 170992
rect 213920 170954 213972 170960
rect 214024 170377 214052 171022
rect 214010 170368 214066 170377
rect 214010 170303 214066 170312
rect 214012 169720 214064 169726
rect 213918 169688 213974 169697
rect 214012 169662 214064 169668
rect 213918 169623 213920 169632
rect 213972 169623 213974 169632
rect 213920 169594 213972 169600
rect 214024 169017 214052 169662
rect 214010 169008 214066 169017
rect 214010 168943 214066 168952
rect 213920 168360 213972 168366
rect 213918 168328 213920 168337
rect 213972 168328 213974 168337
rect 213918 168263 213974 168272
rect 214012 168292 214064 168298
rect 214012 168234 214064 168240
rect 214024 167657 214052 168234
rect 214010 167648 214066 167657
rect 214010 167583 214066 167592
rect 213920 167000 213972 167006
rect 213918 166968 213920 166977
rect 213972 166968 213974 166977
rect 213918 166903 213974 166912
rect 214012 166932 214064 166938
rect 214012 166874 214064 166880
rect 214024 166433 214052 166874
rect 214010 166424 214066 166433
rect 214010 166359 214066 166368
rect 213920 165572 213972 165578
rect 213920 165514 213972 165520
rect 213932 165073 213960 165514
rect 214012 165504 214064 165510
rect 214012 165446 214064 165452
rect 213918 165064 213974 165073
rect 213918 164999 213974 165008
rect 214024 164393 214052 165446
rect 214010 164384 214066 164393
rect 214010 164319 214066 164328
rect 213920 164212 213972 164218
rect 213920 164154 213972 164160
rect 213932 163033 213960 164154
rect 214484 163713 214512 175918
rect 214562 175264 214618 175273
rect 214562 175199 214564 175208
rect 214616 175199 214618 175208
rect 214564 175170 214616 175176
rect 214562 175128 214618 175137
rect 214562 175063 214618 175072
rect 214576 173942 214604 175063
rect 214564 173936 214616 173942
rect 214564 173878 214616 173884
rect 214852 165753 214880 177239
rect 215300 175296 215352 175302
rect 215300 175238 215352 175244
rect 215312 172446 215340 175238
rect 215404 173913 215432 177346
rect 215956 177313 215984 213959
rect 216048 213625 216076 219399
rect 216034 213616 216090 213625
rect 216034 213551 216090 213560
rect 216692 208049 216720 237351
rect 217152 227050 217180 240244
rect 217520 240145 217548 240244
rect 217506 240136 217562 240145
rect 217506 240071 217562 240080
rect 217520 237425 217548 240071
rect 218072 238754 218100 240244
rect 218440 240145 218468 240244
rect 218426 240136 218482 240145
rect 218426 240071 218482 240080
rect 218072 238726 218284 238754
rect 217506 237416 217562 237425
rect 217506 237351 217562 237360
rect 218150 237416 218206 237425
rect 218150 237351 218206 237360
rect 217140 227044 217192 227050
rect 217140 226986 217192 226992
rect 217324 219496 217376 219502
rect 217324 219438 217376 219444
rect 217336 210497 217364 219438
rect 217322 210488 217378 210497
rect 217322 210423 217378 210432
rect 216678 208040 216734 208049
rect 216678 207975 216734 207984
rect 216692 207097 216720 207975
rect 216678 207088 216734 207097
rect 216678 207023 216734 207032
rect 217322 207088 217378 207097
rect 217322 207023 217378 207032
rect 217336 199442 217364 207023
rect 217324 199436 217376 199442
rect 217324 199378 217376 199384
rect 217232 186992 217284 186998
rect 217232 186934 217284 186940
rect 217244 186454 217272 186934
rect 218164 186454 218192 237351
rect 218256 216481 218284 238726
rect 218440 237425 218468 240071
rect 218992 239873 219020 240244
rect 218978 239864 219034 239873
rect 218978 239799 219034 239808
rect 219346 239864 219402 239873
rect 219346 239799 219402 239808
rect 218426 237416 218482 237425
rect 218426 237351 218482 237360
rect 218242 216472 218298 216481
rect 218242 216407 218298 216416
rect 219360 215286 219388 239799
rect 219440 238808 219492 238814
rect 219440 238750 219492 238756
rect 219452 237153 219480 238750
rect 219544 237289 219572 240244
rect 219530 237280 219586 237289
rect 219530 237215 219586 237224
rect 219438 237144 219494 237153
rect 219438 237079 219494 237088
rect 219912 225622 219940 240244
rect 220464 238754 220492 240244
rect 220820 239488 220872 239494
rect 220820 239430 220872 239436
rect 220280 238726 220492 238754
rect 220280 235958 220308 238726
rect 220832 238377 220860 239430
rect 221016 238513 221044 240244
rect 221002 238504 221058 238513
rect 221002 238439 221058 238448
rect 220818 238368 220874 238377
rect 220818 238303 220874 238312
rect 221016 237425 221044 238439
rect 221002 237416 221058 237425
rect 221002 237351 221058 237360
rect 220358 236600 220414 236609
rect 220358 236535 220414 236544
rect 220268 235952 220320 235958
rect 220268 235894 220320 235900
rect 220082 234696 220138 234705
rect 220082 234631 220138 234640
rect 219900 225616 219952 225622
rect 219900 225558 219952 225564
rect 220096 220794 220124 234631
rect 220174 226400 220230 226409
rect 220174 226335 220230 226344
rect 220084 220788 220136 220794
rect 220084 220730 220136 220736
rect 219348 215280 219400 215286
rect 219348 215222 219400 215228
rect 217232 186448 217284 186454
rect 217232 186390 217284 186396
rect 218152 186448 218204 186454
rect 218152 186390 218204 186396
rect 215942 177304 215998 177313
rect 215942 177239 215998 177248
rect 215390 173904 215446 173913
rect 215390 173839 215446 173848
rect 215300 172440 215352 172446
rect 215300 172382 215352 172388
rect 214838 165744 214894 165753
rect 214838 165679 214894 165688
rect 214470 163704 214526 163713
rect 214470 163639 214526 163648
rect 214840 163532 214892 163538
rect 214840 163474 214892 163480
rect 213918 163024 213974 163033
rect 213918 162959 213974 162968
rect 213920 162852 213972 162858
rect 213920 162794 213972 162800
rect 213932 162353 213960 162794
rect 214012 162784 214064 162790
rect 214012 162726 214064 162732
rect 213918 162344 213974 162353
rect 213918 162279 213974 162288
rect 214024 161809 214052 162726
rect 214010 161800 214066 161809
rect 214010 161735 214066 161744
rect 213920 161424 213972 161430
rect 213920 161366 213972 161372
rect 213932 161129 213960 161366
rect 214012 161356 214064 161362
rect 214012 161298 214064 161304
rect 213918 161120 213974 161129
rect 213918 161055 213974 161064
rect 214024 160449 214052 161298
rect 214010 160440 214066 160449
rect 214010 160375 214066 160384
rect 213920 160064 213972 160070
rect 213920 160006 213972 160012
rect 213932 159769 213960 160006
rect 214012 159996 214064 160002
rect 214012 159938 214064 159944
rect 213918 159760 213974 159769
rect 213918 159695 213974 159704
rect 214024 159089 214052 159938
rect 214010 159080 214066 159089
rect 214010 159015 214066 159024
rect 213920 158704 213972 158710
rect 213920 158646 213972 158652
rect 213932 158409 213960 158646
rect 213918 158400 213974 158409
rect 213918 158335 213974 158344
rect 214564 158024 214616 158030
rect 214564 157966 214616 157972
rect 213920 157344 213972 157350
rect 213920 157286 213972 157292
rect 213932 157185 213960 157286
rect 214012 157276 214064 157282
rect 214012 157218 214064 157224
rect 213918 157176 213974 157185
rect 213918 157111 213974 157120
rect 214024 156505 214052 157218
rect 214010 156496 214066 156505
rect 214010 156431 214066 156440
rect 213920 155916 213972 155922
rect 213920 155858 213972 155864
rect 213932 155825 213960 155858
rect 214012 155848 214064 155854
rect 213918 155816 213974 155825
rect 214012 155790 214064 155796
rect 213918 155751 213974 155760
rect 214024 155145 214052 155790
rect 214010 155136 214066 155145
rect 214010 155071 214066 155080
rect 214010 154456 214066 154465
rect 214010 154391 214066 154400
rect 213918 153776 213974 153785
rect 213918 153711 213974 153720
rect 211896 153332 211948 153338
rect 211896 153274 211948 153280
rect 211908 131782 211936 153274
rect 213932 153270 213960 153711
rect 214024 153338 214052 154391
rect 214012 153332 214064 153338
rect 214012 153274 214064 153280
rect 213920 153264 213972 153270
rect 213920 153206 213972 153212
rect 213918 153096 213974 153105
rect 213918 153031 213974 153040
rect 213366 151872 213422 151881
rect 213932 151842 213960 153031
rect 214470 152552 214526 152561
rect 214470 152487 214526 152496
rect 213366 151807 213422 151816
rect 213920 151836 213972 151842
rect 213274 147248 213330 147257
rect 213274 147183 213330 147192
rect 213182 139904 213238 139913
rect 213182 139839 213238 139848
rect 211986 136640 212042 136649
rect 211986 136575 212042 136584
rect 211896 131776 211948 131782
rect 211896 131718 211948 131724
rect 212000 119377 212028 136575
rect 211986 119368 212042 119377
rect 211986 119303 212042 119312
rect 211896 103556 211948 103562
rect 211896 103498 211948 103504
rect 211804 95872 211856 95878
rect 211804 95814 211856 95820
rect 211908 90545 211936 103498
rect 211988 99476 212040 99482
rect 211988 99418 212040 99424
rect 211894 90536 211950 90545
rect 211894 90471 211950 90480
rect 212000 88097 212028 99418
rect 213196 95946 213224 139839
rect 213288 126274 213316 147183
rect 213380 135930 213408 151807
rect 213920 151778 213972 151784
rect 213918 150512 213974 150521
rect 213918 150447 213920 150456
rect 213972 150447 213974 150456
rect 213920 150418 213972 150424
rect 214012 150408 214064 150414
rect 214012 150350 214064 150356
rect 213920 150340 213972 150346
rect 213920 150282 213972 150288
rect 213932 149161 213960 150282
rect 214024 149841 214052 150350
rect 214010 149832 214066 149841
rect 214010 149767 214066 149776
rect 213918 149152 213974 149161
rect 213918 149087 213974 149096
rect 213918 147928 213974 147937
rect 213918 147863 213974 147872
rect 213932 147694 213960 147863
rect 213920 147688 213972 147694
rect 213920 147630 213972 147636
rect 213918 146568 213974 146577
rect 213918 146503 213974 146512
rect 213932 146334 213960 146503
rect 213920 146328 213972 146334
rect 213920 146270 213972 146276
rect 214010 145888 214066 145897
rect 214010 145823 214066 145832
rect 213918 145208 213974 145217
rect 213918 145143 213974 145152
rect 213932 144974 213960 145143
rect 214024 145042 214052 145823
rect 214012 145036 214064 145042
rect 214012 144978 214064 144984
rect 213920 144968 213972 144974
rect 213920 144910 213972 144916
rect 213918 143848 213974 143857
rect 213918 143783 213974 143792
rect 213932 143614 213960 143783
rect 213920 143608 213972 143614
rect 213920 143550 213972 143556
rect 214010 143304 214066 143313
rect 214010 143239 214066 143248
rect 213918 142624 213974 142633
rect 213918 142559 213974 142568
rect 213932 142254 213960 142559
rect 213920 142248 213972 142254
rect 213920 142190 213972 142196
rect 214024 142186 214052 143239
rect 214012 142180 214064 142186
rect 214484 142154 214512 152487
rect 214576 148481 214604 157966
rect 214852 157729 214880 163474
rect 214838 157720 214894 157729
rect 214838 157655 214894 157664
rect 214654 151192 214710 151201
rect 214654 151127 214710 151136
rect 214562 148472 214618 148481
rect 214562 148407 214618 148416
rect 214012 142122 214064 142128
rect 214392 142126 214512 142154
rect 213918 141944 213974 141953
rect 213918 141879 213974 141888
rect 213932 140826 213960 141879
rect 213920 140820 213972 140826
rect 213920 140762 213972 140768
rect 213918 140584 213974 140593
rect 213918 140519 213974 140528
rect 213932 139466 213960 140519
rect 213920 139460 213972 139466
rect 213920 139402 213972 139408
rect 214010 139224 214066 139233
rect 214010 139159 214066 139168
rect 213918 138680 213974 138689
rect 213918 138615 213974 138624
rect 213932 138038 213960 138615
rect 213920 138032 213972 138038
rect 213920 137974 213972 137980
rect 213918 137320 213974 137329
rect 213918 137255 213974 137264
rect 213932 136678 213960 137255
rect 213920 136672 213972 136678
rect 213920 136614 213972 136620
rect 214024 135998 214052 139159
rect 214392 138718 214420 142126
rect 214668 141438 214696 151127
rect 215942 144528 215998 144537
rect 215942 144463 215998 144472
rect 214656 141432 214708 141438
rect 214656 141374 214708 141380
rect 214562 141264 214618 141273
rect 214562 141199 214618 141208
rect 214380 138712 214432 138718
rect 214380 138654 214432 138660
rect 214102 138000 214158 138009
rect 214102 137935 214158 137944
rect 214012 135992 214064 135998
rect 214012 135934 214064 135940
rect 213368 135924 213420 135930
rect 213368 135866 213420 135872
rect 213918 134600 213974 134609
rect 214116 134570 214144 137935
rect 213918 134535 213974 134544
rect 214104 134564 214156 134570
rect 213932 133958 213960 134535
rect 214104 134506 214156 134512
rect 213920 133952 213972 133958
rect 213920 133894 213972 133900
rect 214010 133376 214066 133385
rect 214010 133311 214066 133320
rect 213918 132696 213974 132705
rect 213918 132631 213974 132640
rect 213932 132598 213960 132631
rect 213920 132592 213972 132598
rect 213920 132534 213972 132540
rect 214024 132530 214052 133311
rect 214012 132524 214064 132530
rect 214012 132466 214064 132472
rect 213918 132016 213974 132025
rect 213918 131951 213974 131960
rect 213932 131170 213960 131951
rect 213920 131164 213972 131170
rect 213920 131106 213972 131112
rect 213918 130656 213974 130665
rect 213918 130591 213974 130600
rect 213932 129810 213960 130591
rect 214010 129976 214066 129985
rect 214010 129911 214066 129920
rect 214024 129878 214052 129911
rect 214012 129872 214064 129878
rect 214012 129814 214064 129820
rect 213920 129804 213972 129810
rect 213920 129746 213972 129752
rect 214010 129296 214066 129305
rect 214010 129231 214066 129240
rect 213918 128752 213974 128761
rect 213918 128687 213974 128696
rect 213932 128450 213960 128687
rect 213920 128444 213972 128450
rect 213920 128386 213972 128392
rect 214024 128382 214052 129231
rect 214012 128376 214064 128382
rect 214012 128318 214064 128324
rect 213918 128072 213974 128081
rect 213918 128007 213974 128016
rect 213932 127022 213960 128007
rect 213920 127016 213972 127022
rect 213920 126958 213972 126964
rect 213918 126712 213974 126721
rect 213918 126647 213974 126656
rect 213276 126268 213328 126274
rect 213276 126210 213328 126216
rect 213932 125662 213960 126647
rect 213920 125656 213972 125662
rect 213920 125598 213972 125604
rect 214010 125352 214066 125361
rect 214010 125287 214066 125296
rect 213918 124672 213974 124681
rect 213918 124607 213974 124616
rect 213932 124234 213960 124607
rect 214024 124302 214052 125287
rect 214012 124296 214064 124302
rect 214012 124238 214064 124244
rect 213920 124228 213972 124234
rect 213920 124170 213972 124176
rect 213918 124128 213974 124137
rect 213918 124063 213974 124072
rect 213458 123448 213514 123457
rect 213458 123383 213514 123392
rect 213274 118824 213330 118833
rect 213274 118759 213330 118768
rect 213288 97306 213316 118759
rect 213366 106176 213422 106185
rect 213366 106111 213422 106120
rect 213276 97300 213328 97306
rect 213276 97242 213328 97248
rect 213184 95940 213236 95946
rect 213184 95882 213236 95888
rect 213184 93220 213236 93226
rect 213184 93162 213236 93168
rect 211986 88088 212042 88097
rect 211986 88023 212042 88032
rect 211802 87680 211858 87689
rect 211802 87615 211858 87624
rect 210608 74520 210660 74526
rect 210608 74462 210660 74468
rect 211816 44946 211844 87615
rect 211804 44940 211856 44946
rect 211804 44882 211856 44888
rect 210424 18692 210476 18698
rect 210424 18634 210476 18640
rect 198096 18624 198148 18630
rect 198096 18566 198148 18572
rect 202144 18624 202196 18630
rect 202144 18566 202196 18572
rect 213196 10402 213224 93162
rect 213276 83496 213328 83502
rect 213276 83438 213328 83444
rect 213288 35290 213316 83438
rect 213380 82142 213408 106111
rect 213472 101454 213500 123383
rect 213932 122874 213960 124063
rect 213920 122868 213972 122874
rect 213920 122810 213972 122816
rect 214010 122768 214066 122777
rect 214010 122703 214066 122712
rect 213918 122088 213974 122097
rect 213918 122023 213974 122032
rect 213932 121582 213960 122023
rect 213920 121576 213972 121582
rect 213920 121518 213972 121524
rect 214024 121514 214052 122703
rect 214012 121508 214064 121514
rect 214012 121450 214064 121456
rect 214010 121408 214066 121417
rect 214010 121343 214066 121352
rect 213918 120728 213974 120737
rect 213918 120663 213974 120672
rect 213932 120222 213960 120663
rect 213920 120216 213972 120222
rect 213920 120158 213972 120164
rect 214024 120154 214052 121343
rect 214012 120148 214064 120154
rect 214012 120090 214064 120096
rect 214010 120048 214066 120057
rect 214010 119983 214066 119992
rect 213918 119504 213974 119513
rect 213918 119439 213974 119448
rect 213932 118794 213960 119439
rect 213920 118788 213972 118794
rect 213920 118730 213972 118736
rect 214024 118726 214052 119983
rect 214012 118720 214064 118726
rect 214012 118662 214064 118668
rect 214010 118144 214066 118153
rect 214010 118079 214066 118088
rect 213918 117464 213974 117473
rect 214024 117434 214052 118079
rect 213918 117399 213974 117408
rect 214012 117428 214064 117434
rect 213932 117366 213960 117399
rect 214012 117370 214064 117376
rect 213920 117360 213972 117366
rect 213920 117302 213972 117308
rect 214010 116784 214066 116793
rect 214010 116719 214066 116728
rect 213918 116104 213974 116113
rect 214024 116074 214052 116719
rect 213918 116039 213974 116048
rect 214012 116068 214064 116074
rect 213932 116006 213960 116039
rect 214012 116010 214064 116016
rect 213920 116000 213972 116006
rect 213920 115942 213972 115948
rect 214010 115424 214066 115433
rect 214010 115359 214066 115368
rect 213918 114880 213974 114889
rect 213918 114815 213974 114824
rect 213932 114578 213960 114815
rect 214024 114646 214052 115359
rect 214012 114640 214064 114646
rect 214012 114582 214064 114588
rect 213920 114572 213972 114578
rect 213920 114514 213972 114520
rect 214010 114200 214066 114209
rect 214010 114135 214066 114144
rect 213918 113520 213974 113529
rect 213918 113455 213974 113464
rect 213932 113286 213960 113455
rect 213920 113280 213972 113286
rect 213920 113222 213972 113228
rect 214024 113218 214052 114135
rect 214012 113212 214064 113218
rect 214012 113154 214064 113160
rect 214010 112840 214066 112849
rect 214010 112775 214066 112784
rect 213918 112160 213974 112169
rect 213918 112095 213974 112104
rect 213932 111858 213960 112095
rect 214024 111926 214052 112775
rect 214012 111920 214064 111926
rect 214012 111862 214064 111868
rect 213920 111852 213972 111858
rect 213920 111794 213972 111800
rect 214010 111480 214066 111489
rect 214010 111415 214066 111424
rect 213918 110800 213974 110809
rect 213918 110735 213974 110744
rect 213932 110498 213960 110735
rect 214024 110566 214052 111415
rect 214012 110560 214064 110566
rect 214012 110502 214064 110508
rect 213920 110492 213972 110498
rect 213920 110434 213972 110440
rect 214010 110256 214066 110265
rect 214010 110191 214066 110200
rect 213918 109576 213974 109585
rect 213918 109511 213974 109520
rect 213932 109070 213960 109511
rect 214024 109138 214052 110191
rect 214012 109132 214064 109138
rect 214012 109074 214064 109080
rect 213920 109064 213972 109070
rect 213920 109006 213972 109012
rect 214010 108896 214066 108905
rect 214010 108831 214066 108840
rect 213918 108216 213974 108225
rect 213918 108151 213974 108160
rect 213932 107710 213960 108151
rect 214024 107778 214052 108831
rect 214012 107772 214064 107778
rect 214012 107714 214064 107720
rect 213920 107704 213972 107710
rect 213920 107646 213972 107652
rect 214010 107536 214066 107545
rect 214010 107471 214066 107480
rect 213918 106856 213974 106865
rect 213918 106791 213974 106800
rect 213932 106350 213960 106791
rect 214024 106418 214052 107471
rect 214012 106412 214064 106418
rect 214012 106354 214064 106360
rect 213920 106344 213972 106350
rect 213920 106286 213972 106292
rect 213918 104952 213974 104961
rect 213918 104887 213920 104896
rect 213972 104887 213974 104896
rect 213920 104858 213972 104864
rect 214576 104174 214604 141199
rect 214838 135280 214894 135289
rect 214838 135215 214894 135224
rect 214654 131336 214710 131345
rect 214654 131271 214710 131280
rect 214564 104168 214616 104174
rect 214564 104110 214616 104116
rect 213918 103592 213974 103601
rect 213918 103527 213920 103536
rect 213972 103527 213974 103536
rect 213920 103498 213972 103504
rect 214010 102912 214066 102921
rect 214010 102847 214066 102856
rect 214024 102270 214052 102847
rect 214012 102264 214064 102270
rect 213918 102232 213974 102241
rect 214012 102206 214064 102212
rect 213918 102167 213920 102176
rect 213972 102167 213974 102176
rect 213920 102138 213972 102144
rect 213918 101552 213974 101561
rect 213918 101487 213974 101496
rect 213460 101448 213512 101454
rect 213460 101390 213512 101396
rect 213932 100774 213960 101487
rect 214562 101008 214618 101017
rect 214562 100943 214618 100952
rect 213920 100768 213972 100774
rect 213920 100710 213972 100716
rect 213918 100328 213974 100337
rect 213918 100263 213974 100272
rect 213932 99414 213960 100263
rect 214470 99648 214526 99657
rect 214470 99583 214526 99592
rect 214484 99482 214512 99583
rect 214472 99476 214524 99482
rect 214472 99418 214524 99424
rect 213920 99408 213972 99414
rect 213920 99350 213972 99356
rect 214010 98968 214066 98977
rect 214010 98903 214066 98912
rect 213918 98288 213974 98297
rect 213918 98223 213974 98232
rect 213932 98054 213960 98223
rect 214024 98122 214052 98903
rect 214012 98116 214064 98122
rect 214012 98058 214064 98064
rect 213920 98048 213972 98054
rect 213920 97990 213972 97996
rect 213918 97608 213974 97617
rect 213918 97543 213974 97552
rect 213932 96694 213960 97543
rect 213920 96688 213972 96694
rect 213920 96630 213972 96636
rect 214576 89185 214604 100943
rect 214668 94518 214696 131271
rect 214852 127634 214880 135215
rect 214840 127628 214892 127634
rect 214840 127570 214892 127576
rect 215298 100056 215354 100065
rect 215298 99991 215354 100000
rect 215312 97986 215340 99991
rect 215956 98705 215984 144463
rect 216034 126032 216090 126041
rect 216034 125967 216090 125976
rect 215942 98696 215998 98705
rect 215942 98631 215998 98640
rect 215300 97980 215352 97986
rect 215300 97922 215352 97928
rect 214746 96928 214802 96937
rect 214746 96863 214802 96872
rect 214656 94512 214708 94518
rect 214656 94454 214708 94460
rect 214562 89176 214618 89185
rect 214562 89111 214618 89120
rect 214564 86352 214616 86358
rect 214564 86294 214616 86300
rect 213368 82136 213420 82142
rect 213368 82078 213420 82084
rect 213276 35284 213328 35290
rect 213276 35226 213328 35232
rect 213184 10396 213236 10402
rect 213184 10338 213236 10344
rect 214576 7682 214604 86294
rect 214760 73166 214788 96863
rect 214838 96384 214894 96393
rect 214838 96319 214894 96328
rect 214852 86873 214880 96319
rect 215944 91792 215996 91798
rect 215944 91734 215996 91740
rect 214838 86864 214894 86873
rect 214838 86799 214894 86808
rect 214748 73160 214800 73166
rect 214748 73102 214800 73108
rect 214564 7676 214616 7682
rect 214564 7618 214616 7624
rect 215956 6186 215984 91734
rect 216048 53786 216076 125967
rect 216126 106720 216182 106729
rect 216126 106655 216182 106664
rect 216140 95130 216168 106655
rect 216128 95124 216180 95130
rect 216128 95066 216180 95072
rect 217244 89690 217272 186390
rect 218060 186380 218112 186386
rect 218060 186322 218112 186328
rect 218072 183530 218100 186322
rect 218060 183524 218112 183530
rect 218060 183466 218112 183472
rect 220096 182850 220124 220730
rect 220188 190369 220216 226335
rect 220280 216034 220308 235894
rect 220372 227633 220400 236535
rect 220358 227624 220414 227633
rect 220358 227559 220414 227568
rect 220360 225616 220412 225622
rect 220360 225558 220412 225564
rect 220372 216646 220400 225558
rect 221384 219434 221412 240244
rect 221462 237416 221518 237425
rect 221462 237351 221518 237360
rect 221476 224942 221504 237351
rect 221464 224936 221516 224942
rect 221464 224878 221516 224884
rect 221372 219428 221424 219434
rect 221372 219370 221424 219376
rect 220360 216640 220412 216646
rect 220360 216582 220412 216588
rect 220268 216028 220320 216034
rect 220268 215970 220320 215976
rect 221462 212664 221518 212673
rect 221462 212599 221518 212608
rect 220174 190360 220230 190369
rect 220174 190295 220230 190304
rect 220084 182844 220136 182850
rect 220084 182786 220136 182792
rect 221476 178945 221504 212599
rect 221936 209545 221964 240244
rect 222304 238678 222332 240244
rect 222292 238672 222344 238678
rect 222292 238614 222344 238620
rect 222304 230382 222332 238614
rect 222292 230376 222344 230382
rect 222292 230318 222344 230324
rect 222856 227730 222884 240244
rect 223408 238649 223436 240244
rect 223394 238640 223450 238649
rect 223394 238575 223450 238584
rect 223408 237862 223436 238575
rect 223396 237856 223448 237862
rect 223396 237798 223448 237804
rect 223776 237386 223804 240244
rect 223764 237380 223816 237386
rect 223764 237322 223816 237328
rect 223776 236065 223804 237322
rect 223762 236056 223818 236065
rect 223762 235991 223818 236000
rect 222936 235340 222988 235346
rect 222936 235282 222988 235288
rect 222844 227724 222896 227730
rect 222844 227666 222896 227672
rect 222108 218748 222160 218754
rect 222108 218690 222160 218696
rect 222120 214577 222148 218690
rect 222106 214568 222162 214577
rect 222106 214503 222162 214512
rect 221922 209536 221978 209545
rect 221922 209471 221978 209480
rect 222856 187678 222884 227666
rect 222948 226234 222976 235282
rect 224224 235272 224276 235278
rect 224224 235214 224276 235220
rect 224236 234705 224264 235214
rect 224222 234696 224278 234705
rect 224222 234631 224278 234640
rect 224224 231124 224276 231130
rect 224224 231066 224276 231072
rect 222936 226228 222988 226234
rect 222936 226170 222988 226176
rect 223488 224256 223540 224262
rect 223488 224198 223540 224204
rect 223500 222154 223528 224198
rect 223488 222148 223540 222154
rect 223488 222090 223540 222096
rect 223488 214600 223540 214606
rect 223488 214542 223540 214548
rect 223500 213926 223528 214542
rect 223488 213920 223540 213926
rect 223488 213862 223540 213868
rect 223488 192568 223540 192574
rect 223488 192510 223540 192516
rect 223500 189961 223528 192510
rect 223486 189952 223542 189961
rect 223486 189887 223542 189896
rect 224236 189854 224264 231066
rect 224328 229090 224356 240244
rect 224880 238134 224908 240244
rect 225052 240168 225104 240174
rect 225052 240110 225104 240116
rect 225064 238513 225092 240110
rect 225050 238504 225106 238513
rect 225050 238439 225106 238448
rect 224868 238128 224920 238134
rect 224868 238070 224920 238076
rect 225142 237416 225198 237425
rect 225142 237351 225198 237360
rect 224316 229084 224368 229090
rect 224316 229026 224368 229032
rect 224328 227118 224356 229026
rect 224316 227112 224368 227118
rect 224316 227054 224368 227060
rect 225156 212498 225184 237351
rect 225248 217938 225276 240244
rect 225800 240145 225828 240244
rect 225786 240136 225842 240145
rect 225786 240071 225842 240080
rect 225800 237425 225828 240071
rect 225786 237416 225842 237425
rect 225786 237351 225842 237360
rect 226168 234433 226196 240244
rect 226720 240122 226748 240244
rect 226800 240168 226852 240174
rect 226720 240116 226800 240122
rect 226720 240110 226852 240116
rect 226720 240094 226840 240110
rect 226812 238754 226840 240094
rect 226812 238726 227024 238754
rect 226996 238377 227024 238726
rect 226982 238368 227038 238377
rect 226982 238303 227038 238312
rect 226154 234424 226210 234433
rect 226154 234359 226210 234368
rect 226168 219434 226196 234359
rect 226340 227044 226392 227050
rect 226340 226986 226392 226992
rect 225708 219406 226196 219434
rect 225236 217932 225288 217938
rect 225236 217874 225288 217880
rect 225248 213217 225276 217874
rect 225234 213208 225290 213217
rect 225234 213143 225290 213152
rect 225144 212492 225196 212498
rect 225144 212434 225196 212440
rect 225604 212492 225656 212498
rect 225604 212434 225656 212440
rect 224316 204332 224368 204338
rect 224316 204274 224368 204280
rect 224328 192574 224356 204274
rect 224316 192568 224368 192574
rect 224316 192510 224368 192516
rect 224224 189848 224276 189854
rect 224224 189790 224276 189796
rect 222844 187672 222896 187678
rect 222844 187614 222896 187620
rect 224958 183560 225014 183569
rect 224958 183495 225014 183504
rect 224972 182986 225000 183495
rect 224960 182980 225012 182986
rect 224960 182922 225012 182928
rect 225616 182889 225644 212434
rect 225708 204950 225736 219406
rect 226352 209778 226380 226986
rect 226340 209772 226392 209778
rect 226340 209714 226392 209720
rect 226352 208418 226380 209714
rect 226340 208412 226392 208418
rect 226340 208354 226392 208360
rect 225696 204944 225748 204950
rect 225696 204886 225748 204892
rect 225878 183696 225934 183705
rect 225878 183631 225934 183640
rect 225696 182912 225748 182918
rect 225602 182880 225658 182889
rect 225696 182854 225748 182860
rect 225602 182815 225658 182824
rect 221462 178936 221518 178945
rect 221462 178871 221518 178880
rect 225708 178022 225736 182854
rect 225892 180810 225920 183631
rect 226246 182336 226302 182345
rect 226246 182271 226302 182280
rect 225880 180804 225932 180810
rect 225880 180746 225932 180752
rect 225696 178016 225748 178022
rect 225696 177958 225748 177964
rect 226260 177410 226288 182271
rect 226996 181529 227024 238303
rect 227074 233336 227130 233345
rect 227074 233271 227130 233280
rect 227088 226409 227116 233271
rect 227074 226400 227130 226409
rect 227074 226335 227130 226344
rect 227272 220794 227300 240244
rect 227536 238128 227588 238134
rect 227536 238070 227588 238076
rect 227548 237425 227576 238070
rect 227534 237416 227590 237425
rect 227534 237351 227590 237360
rect 227260 220788 227312 220794
rect 227260 220730 227312 220736
rect 227272 219366 227300 220730
rect 227260 219360 227312 219366
rect 227260 219302 227312 219308
rect 227076 208412 227128 208418
rect 227076 208354 227128 208360
rect 226982 181520 227038 181529
rect 226982 181455 227038 181464
rect 227088 178945 227116 208354
rect 226338 178936 226394 178945
rect 226338 178871 226394 178880
rect 227074 178936 227130 178945
rect 227074 178871 227130 178880
rect 226248 177404 226300 177410
rect 226248 177346 226300 177352
rect 226352 176905 226380 178871
rect 226338 176896 226394 176905
rect 226338 176831 226394 176840
rect 227548 176050 227576 237351
rect 227640 233345 227668 240244
rect 227626 233336 227682 233345
rect 227626 233271 227682 233280
rect 227718 233200 227774 233209
rect 227718 233135 227774 233144
rect 227732 232558 227760 233135
rect 228192 232937 228220 240244
rect 228364 240168 228416 240174
rect 228364 240110 228416 240116
rect 228178 232928 228234 232937
rect 228178 232863 228234 232872
rect 227720 232552 227772 232558
rect 227720 232494 227772 232500
rect 228192 231130 228220 232863
rect 228180 231124 228232 231130
rect 228180 231066 228232 231072
rect 228376 207058 228404 240110
rect 228744 240106 228772 240244
rect 228732 240100 228784 240106
rect 228732 240042 228784 240048
rect 228744 221474 228772 240042
rect 229112 236774 229140 240244
rect 229376 237856 229428 237862
rect 229376 237798 229428 237804
rect 229100 236768 229152 236774
rect 229100 236710 229152 236716
rect 228732 221468 228784 221474
rect 228732 221410 228784 221416
rect 228364 207052 228416 207058
rect 228364 206994 228416 207000
rect 227720 206916 227772 206922
rect 227720 206858 227772 206864
rect 227732 205737 227760 206858
rect 227718 205728 227774 205737
rect 227718 205663 227774 205672
rect 227720 182980 227772 182986
rect 227720 182922 227772 182928
rect 227732 182209 227760 182922
rect 227718 182200 227774 182209
rect 227718 182135 227774 182144
rect 227812 181484 227864 181490
rect 227812 181426 227864 181432
rect 227718 178664 227774 178673
rect 227718 178599 227774 178608
rect 227536 176044 227588 176050
rect 227536 175986 227588 175992
rect 227732 175982 227760 178599
rect 227824 176633 227852 181426
rect 228376 179081 228404 206994
rect 229388 190454 229416 237798
rect 229664 236065 229692 240244
rect 229836 237720 229888 237726
rect 229836 237662 229888 237668
rect 229848 236609 229876 237662
rect 230216 237454 230244 240244
rect 230584 240145 230612 240244
rect 231032 240168 231084 240174
rect 230570 240136 230626 240145
rect 231136 240122 231164 240244
rect 231084 240116 231164 240122
rect 231032 240110 231164 240116
rect 231044 240094 231164 240110
rect 230570 240071 230626 240080
rect 230204 237448 230256 237454
rect 230204 237390 230256 237396
rect 229834 236600 229890 236609
rect 229834 236535 229890 236544
rect 229650 236056 229706 236065
rect 229650 235991 229706 236000
rect 229664 232801 229692 235991
rect 229650 232792 229706 232801
rect 229650 232727 229706 232736
rect 230584 231713 230612 240071
rect 230570 231704 230626 231713
rect 230570 231639 230626 231648
rect 230480 231192 230532 231198
rect 230480 231134 230532 231140
rect 229744 213240 229796 213246
rect 229744 213182 229796 213188
rect 229756 207670 229784 213182
rect 229744 207664 229796 207670
rect 229744 207606 229796 207612
rect 229388 190426 229600 190454
rect 228638 183560 228694 183569
rect 228638 183495 228694 183504
rect 228652 180810 228680 183495
rect 228640 180804 228692 180810
rect 228640 180746 228692 180752
rect 229374 180160 229430 180169
rect 229374 180095 229430 180104
rect 228362 179072 228418 179081
rect 228362 179007 228418 179016
rect 229284 178764 229336 178770
rect 229284 178706 229336 178712
rect 229100 178016 229152 178022
rect 229100 177958 229152 177964
rect 227810 176624 227866 176633
rect 227810 176559 227866 176568
rect 227810 176080 227866 176089
rect 227810 176015 227866 176024
rect 227720 175976 227772 175982
rect 221186 175944 221242 175953
rect 221186 175879 221242 175888
rect 224222 175944 224278 175953
rect 227720 175918 227772 175924
rect 227824 175914 227852 176015
rect 224222 175879 224278 175888
rect 227812 175908 227864 175914
rect 221200 175846 221228 175879
rect 224236 175846 224264 175879
rect 227812 175850 227864 175856
rect 221188 175840 221240 175846
rect 221188 175782 221240 175788
rect 224224 175840 224276 175846
rect 224224 175782 224276 175788
rect 229008 175160 229060 175166
rect 229008 175102 229060 175108
rect 229020 174078 229048 175102
rect 229008 174072 229060 174078
rect 229008 174014 229060 174020
rect 229112 173777 229140 177958
rect 229192 174072 229244 174078
rect 229190 174040 229192 174049
rect 229244 174040 229246 174049
rect 229190 173975 229246 173984
rect 229296 173890 229324 178706
rect 229204 173862 229324 173890
rect 229098 173768 229154 173777
rect 229098 173703 229154 173712
rect 229204 164393 229232 173862
rect 229388 173754 229416 180095
rect 229296 173726 229416 173754
rect 229296 170921 229324 173726
rect 229572 173618 229600 190426
rect 229744 187672 229796 187678
rect 229744 187614 229796 187620
rect 229756 176769 229784 187614
rect 230388 180124 230440 180130
rect 230388 180066 230440 180072
rect 230400 179761 230428 180066
rect 230386 179752 230442 179761
rect 230386 179687 230442 179696
rect 229742 176760 229798 176769
rect 229742 176695 229798 176704
rect 229388 173590 229600 173618
rect 229282 170912 229338 170921
rect 229282 170847 229338 170856
rect 229190 164384 229246 164393
rect 229190 164319 229246 164328
rect 229388 155825 229416 173590
rect 229742 170368 229798 170377
rect 229742 170303 229798 170312
rect 229374 155816 229430 155825
rect 229374 155751 229430 155760
rect 229756 146305 229784 170303
rect 230492 166326 230520 231134
rect 231504 229094 231532 240244
rect 231858 239456 231914 239465
rect 231858 239391 231914 239400
rect 231584 234660 231636 234666
rect 231584 234602 231636 234608
rect 231596 230450 231624 234602
rect 231584 230444 231636 230450
rect 231584 230386 231636 230392
rect 231136 229066 231532 229094
rect 231136 217977 231164 229066
rect 231504 228993 231532 229066
rect 231490 228984 231546 228993
rect 231490 228919 231546 228928
rect 231122 217968 231178 217977
rect 231122 217903 231178 217912
rect 231124 189780 231176 189786
rect 231124 189722 231176 189728
rect 231136 179382 231164 189722
rect 231124 179376 231176 179382
rect 231124 179318 231176 179324
rect 230570 178664 230626 178673
rect 230570 178599 230626 178608
rect 230584 174729 230612 178599
rect 230662 176624 230718 176633
rect 230662 176559 230718 176568
rect 230570 174720 230626 174729
rect 230570 174655 230626 174664
rect 230570 174448 230626 174457
rect 230570 174383 230626 174392
rect 230584 168298 230612 174383
rect 230572 168292 230624 168298
rect 230572 168234 230624 168240
rect 230480 166320 230532 166326
rect 230480 166262 230532 166268
rect 229834 162072 229890 162081
rect 229834 162007 229890 162016
rect 229848 152561 229876 162007
rect 230676 160993 230704 176559
rect 231124 175228 231176 175234
rect 231124 175170 231176 175176
rect 230756 173392 230808 173398
rect 230754 173360 230756 173369
rect 230808 173360 230810 173369
rect 230754 173295 230810 173304
rect 230756 171012 230808 171018
rect 230756 170954 230808 170960
rect 230768 170513 230796 170954
rect 230754 170504 230810 170513
rect 230754 170439 230810 170448
rect 230848 168292 230900 168298
rect 230848 168234 230900 168240
rect 230756 166320 230808 166326
rect 230756 166262 230808 166268
rect 230662 160984 230718 160993
rect 230662 160919 230718 160928
rect 230572 159384 230624 159390
rect 230572 159326 230624 159332
rect 230584 158137 230612 159326
rect 230768 158681 230796 166262
rect 230754 158672 230810 158681
rect 230754 158607 230810 158616
rect 230570 158128 230626 158137
rect 230570 158063 230626 158072
rect 230860 157729 230888 168234
rect 231136 166161 231164 175170
rect 231584 172508 231636 172514
rect 231584 172450 231636 172456
rect 231596 171465 231624 172450
rect 231768 172168 231820 172174
rect 231768 172110 231820 172116
rect 231780 171873 231808 172110
rect 231766 171864 231822 171873
rect 231766 171799 231822 171808
rect 231582 171456 231638 171465
rect 231582 171391 231638 171400
rect 231768 171080 231820 171086
rect 231768 171022 231820 171028
rect 231780 169969 231808 171022
rect 231766 169960 231822 169969
rect 231766 169895 231822 169904
rect 231768 169720 231820 169726
rect 231768 169662 231820 169668
rect 231216 169244 231268 169250
rect 231216 169186 231268 169192
rect 231228 169017 231256 169186
rect 231214 169008 231270 169017
rect 231214 168943 231270 168952
rect 231780 168609 231808 169662
rect 231766 168600 231822 168609
rect 231766 168535 231822 168544
rect 231400 168224 231452 168230
rect 231400 168166 231452 168172
rect 231412 168065 231440 168166
rect 231398 168056 231454 168065
rect 231398 167991 231454 168000
rect 231766 167648 231822 167657
rect 231872 167634 231900 239391
rect 232056 235958 232084 240244
rect 232608 240145 232636 240244
rect 232594 240136 232650 240145
rect 232594 240071 232650 240080
rect 232976 238754 233004 240244
rect 232792 238726 233004 238754
rect 232792 238377 232820 238726
rect 232778 238368 232834 238377
rect 232778 238303 232834 238312
rect 232504 237448 232556 237454
rect 232504 237390 232556 237396
rect 232044 235952 232096 235958
rect 232044 235894 232096 235900
rect 232056 235346 232084 235894
rect 232044 235340 232096 235346
rect 232044 235282 232096 235288
rect 232516 225049 232544 237390
rect 232594 228440 232650 228449
rect 232594 228375 232650 228384
rect 232502 225040 232558 225049
rect 232502 224975 232558 224984
rect 231950 216064 232006 216073
rect 231950 215999 232006 216008
rect 231822 167606 231900 167634
rect 231766 167583 231822 167592
rect 231768 166728 231820 166734
rect 231766 166696 231768 166705
rect 231820 166696 231822 166705
rect 231766 166631 231822 166640
rect 231122 166152 231178 166161
rect 231122 166087 231178 166096
rect 231492 165504 231544 165510
rect 231492 165446 231544 165452
rect 231504 164801 231532 165446
rect 231490 164792 231546 164801
rect 231490 164727 231546 164736
rect 231768 164212 231820 164218
rect 231768 164154 231820 164160
rect 231676 164144 231728 164150
rect 231676 164086 231728 164092
rect 231688 162897 231716 164086
rect 231780 163849 231808 164154
rect 231766 163840 231822 163849
rect 231766 163775 231822 163784
rect 231674 162888 231730 162897
rect 231674 162823 231730 162832
rect 230940 162716 230992 162722
rect 230940 162658 230992 162664
rect 230952 161945 230980 162658
rect 230938 161936 230994 161945
rect 230938 161871 230994 161880
rect 231768 160744 231820 160750
rect 231768 160686 231820 160692
rect 231780 159633 231808 160686
rect 231766 159624 231822 159633
rect 231766 159559 231822 159568
rect 231124 159316 231176 159322
rect 231124 159258 231176 159264
rect 231136 159089 231164 159258
rect 231122 159080 231178 159089
rect 231122 159015 231178 159024
rect 231308 158024 231360 158030
rect 231308 157966 231360 157972
rect 231674 157992 231730 158001
rect 230846 157720 230902 157729
rect 230846 157655 230902 157664
rect 231124 156664 231176 156670
rect 231124 156606 231176 156612
rect 230020 155236 230072 155242
rect 230020 155178 230072 155184
rect 229834 152552 229890 152561
rect 229834 152487 229890 152496
rect 229742 146296 229798 146305
rect 229742 146231 229798 146240
rect 229650 144120 229706 144129
rect 229650 144055 229706 144064
rect 229664 141681 229692 144055
rect 229650 141672 229706 141681
rect 229650 141607 229706 141616
rect 229098 140720 229154 140729
rect 229098 140655 229154 140664
rect 229112 113174 229140 140655
rect 229836 138032 229888 138038
rect 229836 137974 229888 137980
rect 229742 136912 229798 136921
rect 229742 136847 229798 136856
rect 229756 133657 229784 136847
rect 229742 133648 229798 133657
rect 229742 133583 229798 133592
rect 229742 123312 229798 123321
rect 229742 123247 229798 123256
rect 229112 113146 229232 113174
rect 229098 96792 229154 96801
rect 229020 96750 229098 96778
rect 225052 96076 225104 96082
rect 225052 96018 225104 96024
rect 226432 96076 226484 96082
rect 226432 96018 226484 96024
rect 222476 96008 222528 96014
rect 225064 95985 225092 96018
rect 226444 95985 226472 96018
rect 229020 95985 229048 96750
rect 229098 96727 229154 96736
rect 222476 95950 222528 95956
rect 225050 95976 225106 95985
rect 222488 95198 222516 95950
rect 225050 95911 225106 95920
rect 226430 95976 226486 95985
rect 226430 95911 226486 95920
rect 229006 95976 229062 95985
rect 229006 95911 229062 95920
rect 229008 95872 229060 95878
rect 229008 95814 229060 95820
rect 229020 95577 229048 95814
rect 229006 95568 229062 95577
rect 229006 95503 229062 95512
rect 228546 95296 228602 95305
rect 226432 95260 226484 95266
rect 228546 95231 228602 95240
rect 226432 95202 226484 95208
rect 222476 95192 222528 95198
rect 222476 95134 222528 95140
rect 220818 94752 220874 94761
rect 220818 94687 220874 94696
rect 220832 93838 220860 94687
rect 224222 94616 224278 94625
rect 224222 94551 224278 94560
rect 225602 94616 225658 94625
rect 225602 94551 225658 94560
rect 220820 93832 220872 93838
rect 220820 93774 220872 93780
rect 222844 93152 222896 93158
rect 218794 93120 218850 93129
rect 222844 93094 222896 93100
rect 218794 93055 218850 93064
rect 217232 89684 217284 89690
rect 217232 89626 217284 89632
rect 217322 89176 217378 89185
rect 217322 89111 217378 89120
rect 216128 82136 216180 82142
rect 216128 82078 216180 82084
rect 216036 53780 216088 53786
rect 216036 53722 216088 53728
rect 216140 20058 216168 82078
rect 216128 20052 216180 20058
rect 216128 19994 216180 20000
rect 217336 11830 217364 89111
rect 218704 73908 218756 73914
rect 218704 73850 218756 73856
rect 218716 33794 218744 73850
rect 218808 73846 218836 93055
rect 221462 91760 221518 91769
rect 221462 91695 221518 91704
rect 220084 90432 220136 90438
rect 220084 90374 220136 90380
rect 218796 73840 218848 73846
rect 218796 73782 218848 73788
rect 218704 33788 218756 33794
rect 218704 33730 218756 33736
rect 217324 11824 217376 11830
rect 217324 11766 217376 11772
rect 220096 9042 220124 90374
rect 220174 83464 220230 83473
rect 220174 83399 220230 83408
rect 220188 15978 220216 83399
rect 221476 53145 221504 91695
rect 221462 53136 221518 53145
rect 221462 53071 221518 53080
rect 220176 15972 220228 15978
rect 220176 15914 220228 15920
rect 220084 9036 220136 9042
rect 220084 8978 220136 8984
rect 215944 6180 215996 6186
rect 215944 6122 215996 6128
rect 196806 3360 196862 3369
rect 196806 3295 196862 3304
rect 184202 2680 184258 2689
rect 184202 2615 184258 2624
rect 222856 2174 222884 93094
rect 222934 84960 222990 84969
rect 222934 84895 222990 84904
rect 222948 10334 222976 84895
rect 224236 20670 224264 94551
rect 224316 87712 224368 87718
rect 224316 87654 224368 87660
rect 224224 20664 224276 20670
rect 224224 20606 224276 20612
rect 224328 19990 224356 87654
rect 225616 44878 225644 94551
rect 226444 87553 226472 95202
rect 226430 87544 226486 87553
rect 226430 87479 226486 87488
rect 228362 79656 228418 79665
rect 228362 79591 228418 79600
rect 225604 44872 225656 44878
rect 225604 44814 225656 44820
rect 228376 22778 228404 79591
rect 228560 79529 228588 95231
rect 229204 95130 229232 113146
rect 229192 95124 229244 95130
rect 229192 95066 229244 95072
rect 228546 79520 228602 79529
rect 228546 79455 228602 79464
rect 229756 28354 229784 123247
rect 229848 86358 229876 137974
rect 229926 131472 229982 131481
rect 229926 131407 229982 131416
rect 229940 93129 229968 131407
rect 230032 123593 230060 155178
rect 230664 153944 230716 153950
rect 230664 153886 230716 153892
rect 230570 153776 230626 153785
rect 230570 153711 230626 153720
rect 230584 152017 230612 153711
rect 230570 152008 230626 152017
rect 230570 151943 230626 151952
rect 230388 151088 230440 151094
rect 230676 151065 230704 153886
rect 230756 152516 230808 152522
rect 230756 152458 230808 152464
rect 230388 151030 230440 151036
rect 230662 151056 230718 151065
rect 230400 143041 230428 151030
rect 230662 150991 230718 151000
rect 230572 150408 230624 150414
rect 230572 150350 230624 150356
rect 230584 149161 230612 150350
rect 230570 149152 230626 149161
rect 230570 149087 230626 149096
rect 230572 149048 230624 149054
rect 230572 148990 230624 148996
rect 230584 147801 230612 148990
rect 230768 148209 230796 152458
rect 231136 149705 231164 156606
rect 231320 155281 231348 157966
rect 231674 157927 231730 157936
rect 231306 155272 231362 155281
rect 231306 155207 231362 155216
rect 231584 154556 231636 154562
rect 231584 154498 231636 154504
rect 231596 153377 231624 154498
rect 231688 154329 231716 157927
rect 231964 156670 231992 215999
rect 232516 199481 232544 224975
rect 232608 215966 232636 228375
rect 232792 226273 232820 238303
rect 232778 226264 232834 226273
rect 232778 226199 232834 226208
rect 233332 216028 233384 216034
rect 233332 215970 233384 215976
rect 232596 215960 232648 215966
rect 232596 215902 232648 215908
rect 232596 200184 232648 200190
rect 232596 200126 232648 200132
rect 232502 199472 232558 199481
rect 232502 199407 232558 199416
rect 232044 184272 232096 184278
rect 232044 184214 232096 184220
rect 232056 175234 232084 184214
rect 232608 184210 232636 200126
rect 232504 184204 232556 184210
rect 232504 184146 232556 184152
rect 232596 184204 232648 184210
rect 232596 184146 232648 184152
rect 232044 175228 232096 175234
rect 232044 175170 232096 175176
rect 232042 174040 232098 174049
rect 232042 173975 232098 173984
rect 231952 156664 232004 156670
rect 231952 156606 232004 156612
rect 231768 156596 231820 156602
rect 231768 156538 231820 156544
rect 231674 154320 231730 154329
rect 231674 154255 231730 154264
rect 231780 153921 231808 156538
rect 231766 153912 231822 153921
rect 231766 153847 231822 153856
rect 231582 153368 231638 153377
rect 231582 153303 231638 153312
rect 232056 151814 232084 173975
rect 232516 171018 232544 184146
rect 233238 178120 233294 178129
rect 233238 178055 233294 178064
rect 233252 173398 233280 178055
rect 233240 173392 233292 173398
rect 233240 173334 233292 173340
rect 232504 171012 232556 171018
rect 232504 170954 232556 170960
rect 233344 169250 233372 215970
rect 233528 215257 233556 240244
rect 234080 238785 234108 240244
rect 234066 238776 234122 238785
rect 234066 238711 234122 238720
rect 234080 234666 234108 238711
rect 234068 234660 234120 234666
rect 234068 234602 234120 234608
rect 233514 215248 233570 215257
rect 233514 215183 233570 215192
rect 233528 211818 233556 215183
rect 233516 211812 233568 211818
rect 233516 211754 233568 211760
rect 234448 209098 234476 240244
rect 235000 216714 235028 240244
rect 235368 227633 235396 240244
rect 235354 227624 235410 227633
rect 235354 227559 235410 227568
rect 234988 216708 235040 216714
rect 234988 216650 235040 216656
rect 235000 216617 235028 216650
rect 235920 216617 235948 240244
rect 236000 233912 236052 233918
rect 236000 233854 236052 233860
rect 236012 233170 236040 233854
rect 236000 233164 236052 233170
rect 236000 233106 236052 233112
rect 236472 219366 236500 240244
rect 236840 240009 236868 240244
rect 237392 240038 237420 240244
rect 237944 240145 237972 240244
rect 237930 240136 237986 240145
rect 237930 240071 237986 240080
rect 237380 240032 237432 240038
rect 236826 240000 236882 240009
rect 237380 239974 237432 239980
rect 238116 240032 238168 240038
rect 238116 239974 238168 239980
rect 236826 239935 236882 239944
rect 236840 237726 236868 239935
rect 238024 238808 238076 238814
rect 238024 238750 238076 238756
rect 236828 237720 236880 237726
rect 236828 237662 236880 237668
rect 236644 233164 236696 233170
rect 236644 233106 236696 233112
rect 236460 219360 236512 219366
rect 236460 219302 236512 219308
rect 234986 216608 235042 216617
rect 234986 216543 235042 216552
rect 235906 216608 235962 216617
rect 235906 216543 235962 216552
rect 235262 214704 235318 214713
rect 235262 214639 235318 214648
rect 234436 209092 234488 209098
rect 234436 209034 234488 209040
rect 234448 208457 234476 209034
rect 234434 208448 234490 208457
rect 234434 208383 234490 208392
rect 234620 200796 234672 200802
rect 234620 200738 234672 200744
rect 233516 182844 233568 182850
rect 233516 182786 233568 182792
rect 233424 173936 233476 173942
rect 233424 173878 233476 173884
rect 233332 169244 233384 169250
rect 233332 169186 233384 169192
rect 232780 165640 232832 165646
rect 232780 165582 232832 165588
rect 232686 157856 232742 157865
rect 232686 157791 232742 157800
rect 231872 151786 232084 151814
rect 232596 151836 232648 151842
rect 231216 149728 231268 149734
rect 231122 149696 231178 149705
rect 231216 149670 231268 149676
rect 231122 149631 231178 149640
rect 230754 148200 230810 148209
rect 230754 148135 230810 148144
rect 230570 147792 230626 147801
rect 230570 147727 230626 147736
rect 230756 147620 230808 147626
rect 230756 147562 230808 147568
rect 230768 147257 230796 147562
rect 230754 147248 230810 147257
rect 230754 147183 230810 147192
rect 231124 146940 231176 146946
rect 231124 146882 231176 146888
rect 230664 146260 230716 146266
rect 230664 146202 230716 146208
rect 230676 144945 230704 146202
rect 230662 144936 230718 144945
rect 230662 144871 230718 144880
rect 230386 143032 230442 143041
rect 230386 142967 230442 142976
rect 230572 136604 230624 136610
rect 230572 136546 230624 136552
rect 230584 136377 230612 136546
rect 230570 136368 230626 136377
rect 230570 136303 230626 136312
rect 230664 133204 230716 133210
rect 230664 133146 230716 133152
rect 230676 127945 230704 133146
rect 231136 132494 231164 146882
rect 231228 135969 231256 149670
rect 231306 149152 231362 149161
rect 231306 149087 231362 149096
rect 231320 145353 231348 149087
rect 231872 147778 231900 151786
rect 232596 151778 232648 151784
rect 231780 147750 231900 147778
rect 231780 146849 231808 147750
rect 231766 146840 231822 146849
rect 231766 146775 231822 146784
rect 231674 145752 231730 145761
rect 231674 145687 231730 145696
rect 231400 145580 231452 145586
rect 231400 145522 231452 145528
rect 231306 145344 231362 145353
rect 231306 145279 231362 145288
rect 231308 136196 231360 136202
rect 231308 136138 231360 136144
rect 231214 135960 231270 135969
rect 231214 135895 231270 135904
rect 231320 135425 231348 136138
rect 231306 135416 231362 135425
rect 231306 135351 231362 135360
rect 231308 135312 231360 135318
rect 231308 135254 231360 135260
rect 231044 132466 231164 132494
rect 231044 129849 231072 132466
rect 231124 131028 231176 131034
rect 231124 130970 231176 130976
rect 231136 130665 231164 130970
rect 231122 130656 231178 130665
rect 231122 130591 231178 130600
rect 231030 129840 231086 129849
rect 231030 129775 231086 129784
rect 230756 129736 230808 129742
rect 230756 129678 230808 129684
rect 230768 128897 230796 129678
rect 231320 129305 231348 135254
rect 231412 132569 231440 145522
rect 231688 144401 231716 145687
rect 231768 144900 231820 144906
rect 231768 144842 231820 144848
rect 231674 144392 231730 144401
rect 231674 144327 231730 144336
rect 231780 143993 231808 144842
rect 231766 143984 231822 143993
rect 231766 143919 231822 143928
rect 231768 143472 231820 143478
rect 231766 143440 231768 143449
rect 231820 143440 231822 143449
rect 231766 143375 231822 143384
rect 232504 142180 232556 142186
rect 232504 142122 232556 142128
rect 231584 141432 231636 141438
rect 231584 141374 231636 141380
rect 231596 135318 231624 141374
rect 231768 139392 231820 139398
rect 231768 139334 231820 139340
rect 231780 138281 231808 139334
rect 231766 138272 231822 138281
rect 231766 138207 231822 138216
rect 231768 137964 231820 137970
rect 231768 137906 231820 137912
rect 231780 137873 231808 137906
rect 231766 137864 231822 137873
rect 231766 137799 231822 137808
rect 231584 135312 231636 135318
rect 231584 135254 231636 135260
rect 231492 135244 231544 135250
rect 231492 135186 231544 135192
rect 231504 134065 231532 135186
rect 231768 135176 231820 135182
rect 231768 135118 231820 135124
rect 231780 135017 231808 135118
rect 231766 135008 231822 135017
rect 231766 134943 231822 134952
rect 231490 134056 231546 134065
rect 231490 133991 231546 134000
rect 231492 133884 231544 133890
rect 231492 133826 231544 133832
rect 231504 133113 231532 133826
rect 231490 133104 231546 133113
rect 231490 133039 231546 133048
rect 231398 132560 231454 132569
rect 231398 132495 231454 132504
rect 231768 132456 231820 132462
rect 231768 132398 231820 132404
rect 231400 131708 231452 131714
rect 231400 131650 231452 131656
rect 231412 131209 231440 131650
rect 231780 131617 231808 132398
rect 231766 131608 231822 131617
rect 231766 131543 231822 131552
rect 231398 131200 231454 131209
rect 231398 131135 231454 131144
rect 231768 131096 231820 131102
rect 231768 131038 231820 131044
rect 231780 130257 231808 131038
rect 231766 130248 231822 130257
rect 231766 130183 231822 130192
rect 231306 129296 231362 129305
rect 231306 129231 231362 129240
rect 230754 128888 230810 128897
rect 230754 128823 230810 128832
rect 231674 128344 231730 128353
rect 231674 128279 231730 128288
rect 231768 128308 231820 128314
rect 231688 128246 231716 128279
rect 231768 128250 231820 128256
rect 231676 128240 231728 128246
rect 231676 128182 231728 128188
rect 231674 128072 231730 128081
rect 231674 128007 231730 128016
rect 230662 127936 230718 127945
rect 230662 127871 230718 127880
rect 231308 126948 231360 126954
rect 231308 126890 231360 126896
rect 231214 126848 231270 126857
rect 231214 126783 231270 126792
rect 230572 126744 230624 126750
rect 230572 126686 230624 126692
rect 230584 126041 230612 126686
rect 230570 126032 230626 126041
rect 230570 125967 230626 125976
rect 230756 125588 230808 125594
rect 230756 125530 230808 125536
rect 230768 124545 230796 125530
rect 230754 124536 230810 124545
rect 230754 124471 230810 124480
rect 231124 123956 231176 123962
rect 231124 123898 231176 123904
rect 230018 123584 230074 123593
rect 230018 123519 230074 123528
rect 230664 123480 230716 123486
rect 230664 123422 230716 123428
rect 230676 118969 230704 123422
rect 231032 122732 231084 122738
rect 231032 122674 231084 122680
rect 231044 122233 231072 122674
rect 231030 122224 231086 122233
rect 231030 122159 231086 122168
rect 230662 118960 230718 118969
rect 230662 118895 230718 118904
rect 230572 118652 230624 118658
rect 230572 118594 230624 118600
rect 230584 117473 230612 118594
rect 230570 117464 230626 117473
rect 230570 117399 230626 117408
rect 230848 117156 230900 117162
rect 230848 117098 230900 117104
rect 230860 117065 230888 117098
rect 230846 117056 230902 117065
rect 230846 116991 230902 117000
rect 230664 115252 230716 115258
rect 230664 115194 230716 115200
rect 230676 113665 230704 115194
rect 231136 114617 231164 123898
rect 231228 121689 231256 126783
rect 231320 126449 231348 126890
rect 231306 126440 231362 126449
rect 231306 126375 231362 126384
rect 231492 125180 231544 125186
rect 231492 125122 231544 125128
rect 231504 125089 231532 125122
rect 231490 125080 231546 125089
rect 231490 125015 231546 125024
rect 231306 124808 231362 124817
rect 231306 124743 231362 124752
rect 231214 121680 231270 121689
rect 231214 121615 231270 121624
rect 231214 120592 231270 120601
rect 231214 120527 231270 120536
rect 231122 114608 231178 114617
rect 231122 114543 231178 114552
rect 230662 113656 230718 113665
rect 230662 113591 230718 113600
rect 231032 113076 231084 113082
rect 231032 113018 231084 113024
rect 231044 112713 231072 113018
rect 231030 112704 231086 112713
rect 231030 112639 231086 112648
rect 231122 112160 231178 112169
rect 231122 112095 231178 112104
rect 230572 111784 230624 111790
rect 230572 111726 230624 111732
rect 230584 111353 230612 111726
rect 230570 111344 230626 111353
rect 230570 111279 230626 111288
rect 230940 107568 230992 107574
rect 230940 107510 230992 107516
rect 230952 107137 230980 107510
rect 230938 107128 230994 107137
rect 230938 107063 230994 107072
rect 230754 104680 230810 104689
rect 230754 104615 230810 104624
rect 230480 101516 230532 101522
rect 230480 101458 230532 101464
rect 230492 100881 230520 101458
rect 230478 100872 230534 100881
rect 230478 100807 230534 100816
rect 230572 99748 230624 99754
rect 230572 99690 230624 99696
rect 230584 99521 230612 99690
rect 230570 99512 230626 99521
rect 230570 99447 230626 99456
rect 230768 98977 230796 104615
rect 231032 99340 231084 99346
rect 231032 99282 231084 99288
rect 230754 98968 230810 98977
rect 230754 98903 230810 98912
rect 230756 98864 230808 98870
rect 230756 98806 230808 98812
rect 230768 98569 230796 98806
rect 230754 98560 230810 98569
rect 230754 98495 230810 98504
rect 231044 98025 231072 99282
rect 231030 98016 231086 98025
rect 231030 97951 231086 97960
rect 230478 96248 230534 96257
rect 230478 96183 230534 96192
rect 230492 95538 230520 96183
rect 230480 95532 230532 95538
rect 230480 95474 230532 95480
rect 229926 93120 229982 93129
rect 229926 93055 229982 93064
rect 229836 86352 229888 86358
rect 229836 86294 229888 86300
rect 229744 28348 229796 28354
rect 229744 28290 229796 28296
rect 228364 22772 228416 22778
rect 228364 22714 228416 22720
rect 224316 19984 224368 19990
rect 224316 19926 224368 19932
rect 231136 15910 231164 112095
rect 231228 103329 231256 120527
rect 231320 111761 231348 124743
rect 231688 124137 231716 128007
rect 231780 127401 231808 128250
rect 231766 127392 231822 127401
rect 231766 127327 231822 127336
rect 231674 124128 231730 124137
rect 231674 124063 231730 124072
rect 231768 122800 231820 122806
rect 231768 122742 231820 122748
rect 231780 122641 231808 122742
rect 231766 122632 231822 122641
rect 231766 122567 231822 122576
rect 231768 121440 231820 121446
rect 231768 121382 231820 121388
rect 231780 120737 231808 121382
rect 231766 120728 231822 120737
rect 231492 120692 231544 120698
rect 231766 120663 231822 120672
rect 231492 120634 231544 120640
rect 231504 120329 231532 120634
rect 231490 120320 231546 120329
rect 231490 120255 231546 120264
rect 231768 120080 231820 120086
rect 231674 120048 231730 120057
rect 231768 120022 231820 120028
rect 231674 119983 231730 119992
rect 231688 119377 231716 119983
rect 231780 119785 231808 120022
rect 231766 119776 231822 119785
rect 231766 119711 231822 119720
rect 231674 119368 231730 119377
rect 231674 119303 231730 119312
rect 231676 118040 231728 118046
rect 231676 117982 231728 117988
rect 231398 116376 231454 116385
rect 231398 116311 231454 116320
rect 231306 111752 231362 111761
rect 231306 111687 231362 111696
rect 231412 105641 231440 116311
rect 231688 116113 231716 117982
rect 231768 117224 231820 117230
rect 231768 117166 231820 117172
rect 231780 116521 231808 117166
rect 231766 116512 231822 116521
rect 231766 116447 231822 116456
rect 231674 116104 231730 116113
rect 231674 116039 231730 116048
rect 231492 115932 231544 115938
rect 231492 115874 231544 115880
rect 231504 115161 231532 115874
rect 231490 115152 231546 115161
rect 231490 115087 231546 115096
rect 231676 114504 231728 114510
rect 231676 114446 231728 114452
rect 231492 114232 231544 114238
rect 231490 114200 231492 114209
rect 231544 114200 231546 114209
rect 231490 114135 231546 114144
rect 231688 113257 231716 114446
rect 231674 113248 231730 113257
rect 231674 113183 231730 113192
rect 231768 113144 231820 113150
rect 231768 113086 231820 113092
rect 231780 112305 231808 113086
rect 231766 112296 231822 112305
rect 231766 112231 231822 112240
rect 231768 111716 231820 111722
rect 231768 111658 231820 111664
rect 231674 111072 231730 111081
rect 231674 111007 231730 111016
rect 231688 109857 231716 111007
rect 231780 110809 231808 111658
rect 231766 110800 231822 110809
rect 231766 110735 231822 110744
rect 231768 110424 231820 110430
rect 231768 110366 231820 110372
rect 231674 109848 231730 109857
rect 231674 109783 231730 109792
rect 231676 109744 231728 109750
rect 231676 109686 231728 109692
rect 231492 108996 231544 109002
rect 231492 108938 231544 108944
rect 231504 107953 231532 108938
rect 231490 107944 231546 107953
rect 231490 107879 231546 107888
rect 231584 107636 231636 107642
rect 231584 107578 231636 107584
rect 231596 106593 231624 107578
rect 231582 106584 231638 106593
rect 231582 106519 231638 106528
rect 231584 106276 231636 106282
rect 231584 106218 231636 106224
rect 231398 105632 231454 105641
rect 231398 105567 231454 105576
rect 231596 105233 231624 106218
rect 231582 105224 231638 105233
rect 231582 105159 231638 105168
rect 231492 104780 231544 104786
rect 231492 104722 231544 104728
rect 231504 103737 231532 104722
rect 231490 103728 231546 103737
rect 231490 103663 231546 103672
rect 231688 103514 231716 109686
rect 231780 109449 231808 110366
rect 231766 109440 231822 109449
rect 231766 109375 231822 109384
rect 231768 108928 231820 108934
rect 231768 108870 231820 108876
rect 231780 108497 231808 108870
rect 231766 108488 231822 108497
rect 231766 108423 231822 108432
rect 231768 104848 231820 104854
rect 231768 104790 231820 104796
rect 231780 104281 231808 104790
rect 231766 104272 231822 104281
rect 231766 104207 231822 104216
rect 231504 103486 231716 103514
rect 231768 103488 231820 103494
rect 231400 103420 231452 103426
rect 231400 103362 231452 103368
rect 231214 103320 231270 103329
rect 231214 103255 231270 103264
rect 231412 102785 231440 103362
rect 231398 102776 231454 102785
rect 231398 102711 231454 102720
rect 231504 101833 231532 103486
rect 231768 103430 231820 103436
rect 231674 102776 231730 102785
rect 231674 102711 231730 102720
rect 231490 101824 231546 101833
rect 231490 101759 231546 101768
rect 231214 101280 231270 101289
rect 231214 101215 231270 101224
rect 231228 29714 231256 101215
rect 231688 99929 231716 102711
rect 231780 102377 231808 103430
rect 231766 102368 231822 102377
rect 231766 102303 231822 102312
rect 231768 102128 231820 102134
rect 231768 102070 231820 102076
rect 231780 101425 231808 102070
rect 231766 101416 231822 101425
rect 231766 101351 231822 101360
rect 231768 100632 231820 100638
rect 231768 100574 231820 100580
rect 231780 100473 231808 100574
rect 231766 100464 231822 100473
rect 231766 100399 231822 100408
rect 231674 99920 231730 99929
rect 231674 99855 231730 99864
rect 232516 99754 232544 142122
rect 232608 111790 232636 151778
rect 232700 117162 232728 157791
rect 232792 126750 232820 165582
rect 233436 162722 233464 173878
rect 233424 162716 233476 162722
rect 233424 162658 233476 162664
rect 233528 147626 233556 182786
rect 234632 172174 234660 200738
rect 234712 176044 234764 176050
rect 234712 175986 234764 175992
rect 234620 172168 234672 172174
rect 234620 172110 234672 172116
rect 234724 169561 234752 175986
rect 234710 169552 234766 169561
rect 234710 169487 234766 169496
rect 234618 168600 234674 168609
rect 234618 168535 234674 168544
rect 234632 165209 234660 168535
rect 235276 166734 235304 214639
rect 236000 191208 236052 191214
rect 236000 191150 236052 191156
rect 235356 175296 235408 175302
rect 235356 175238 235408 175244
rect 235264 166728 235316 166734
rect 235264 166670 235316 166676
rect 234618 165200 234674 165209
rect 234618 165135 234674 165144
rect 234068 164280 234120 164286
rect 234068 164222 234120 164228
rect 233976 157412 234028 157418
rect 233976 157354 234028 157360
rect 233882 155272 233938 155281
rect 233882 155207 233938 155216
rect 233516 147620 233568 147626
rect 233516 147562 233568 147568
rect 233792 147008 233844 147014
rect 233792 146950 233844 146956
rect 233804 145897 233832 146950
rect 233790 145888 233846 145897
rect 233790 145823 233846 145832
rect 232780 126744 232832 126750
rect 232780 126686 232832 126692
rect 232688 117156 232740 117162
rect 232688 117098 232740 117104
rect 232778 116648 232834 116657
rect 232778 116583 232834 116592
rect 232596 111784 232648 111790
rect 232596 111726 232648 111732
rect 232594 105496 232650 105505
rect 232594 105431 232650 105440
rect 232504 99748 232556 99754
rect 232504 99690 232556 99696
rect 231398 98696 231454 98705
rect 231398 98631 231454 98640
rect 231412 97617 231440 98631
rect 231398 97608 231454 97617
rect 231398 97543 231454 97552
rect 231306 96656 231362 96665
rect 231306 96591 231362 96600
rect 231320 82793 231348 96591
rect 232504 95532 232556 95538
rect 232504 95474 232556 95480
rect 231306 82784 231362 82793
rect 231306 82719 231362 82728
rect 231320 31074 231348 82719
rect 231308 31068 231360 31074
rect 231308 31010 231360 31016
rect 231216 29708 231268 29714
rect 231216 29650 231268 29656
rect 231124 15904 231176 15910
rect 231124 15846 231176 15852
rect 222936 10328 222988 10334
rect 222936 10270 222988 10276
rect 232516 4214 232544 95474
rect 232608 93226 232636 105431
rect 232596 93220 232648 93226
rect 232596 93162 232648 93168
rect 232792 82210 232820 116583
rect 233896 114238 233924 155207
rect 233988 118658 234016 157354
rect 234080 125186 234108 164222
rect 234160 140140 234212 140146
rect 234160 140082 234212 140088
rect 234172 131714 234200 140082
rect 235262 135824 235318 135833
rect 235262 135759 235318 135768
rect 234160 131708 234212 131714
rect 234160 131650 234212 131656
rect 234068 125180 234120 125186
rect 234068 125122 234120 125128
rect 234158 123448 234214 123457
rect 234158 123383 234214 123392
rect 234066 122088 234122 122097
rect 234066 122023 234122 122032
rect 233976 118652 234028 118658
rect 233976 118594 234028 118600
rect 233884 114232 233936 114238
rect 233884 114174 233936 114180
rect 233882 105632 233938 105641
rect 233882 105567 233938 105576
rect 232780 82204 232832 82210
rect 232780 82146 232832 82152
rect 232504 4208 232556 4214
rect 232504 4150 232556 4156
rect 222844 2168 222896 2174
rect 222844 2110 222896 2116
rect 233896 2106 233924 105567
rect 233976 99408 234028 99414
rect 233976 99350 234028 99356
rect 233988 11762 234016 99350
rect 234080 89010 234108 122023
rect 234172 98870 234200 123383
rect 234160 98864 234212 98870
rect 234160 98806 234212 98812
rect 234068 89004 234120 89010
rect 234068 88946 234120 88952
rect 235276 13190 235304 135759
rect 235368 104689 235396 175238
rect 235538 166288 235594 166297
rect 235538 166223 235594 166232
rect 235448 161492 235500 161498
rect 235448 161434 235500 161440
rect 235460 126857 235488 161434
rect 235552 158001 235580 166223
rect 236012 165510 236040 191150
rect 236092 185700 236144 185706
rect 236092 185642 236144 185648
rect 236104 168473 236132 185642
rect 236090 168464 236146 168473
rect 236090 168399 236146 168408
rect 236000 165504 236052 165510
rect 236000 165446 236052 165452
rect 235538 157992 235594 158001
rect 235538 157927 235594 157936
rect 235540 154624 235592 154630
rect 235540 154566 235592 154572
rect 235446 126848 235502 126857
rect 235446 126783 235502 126792
rect 235552 123962 235580 154566
rect 236656 143478 236684 233106
rect 237380 202224 237432 202230
rect 237380 202166 237432 202172
rect 236826 168464 236882 168473
rect 236826 168399 236882 168408
rect 236736 166320 236788 166326
rect 236736 166262 236788 166268
rect 236644 143472 236696 143478
rect 236644 143414 236696 143420
rect 236748 136202 236776 166262
rect 236736 136196 236788 136202
rect 236736 136138 236788 136144
rect 236840 128246 236868 168399
rect 237392 166297 237420 202166
rect 237472 178696 237524 178702
rect 237472 178638 237524 178644
rect 237484 168230 237512 178638
rect 238036 174593 238064 238750
rect 238128 223553 238156 239974
rect 238312 231305 238340 240244
rect 238864 232937 238892 240244
rect 239232 237454 239260 240244
rect 239220 237448 239272 237454
rect 239220 237390 239272 237396
rect 239496 236700 239548 236706
rect 239496 236642 239548 236648
rect 238850 232928 238906 232937
rect 238850 232863 238906 232872
rect 239402 232928 239458 232937
rect 239402 232863 239458 232872
rect 239416 231985 239444 232863
rect 239402 231976 239458 231985
rect 239402 231911 239458 231920
rect 238298 231296 238354 231305
rect 238298 231231 238354 231240
rect 238114 223544 238170 223553
rect 238114 223479 238170 223488
rect 239416 220833 239444 231911
rect 239508 227050 239536 236642
rect 239496 227044 239548 227050
rect 239496 226986 239548 226992
rect 239402 220824 239458 220833
rect 239402 220759 239458 220768
rect 238758 210352 238814 210361
rect 238758 210287 238814 210296
rect 238772 207777 238800 210287
rect 239784 209846 239812 240244
rect 240336 238746 240364 240244
rect 240324 238740 240376 238746
rect 240324 238682 240376 238688
rect 240048 237516 240100 237522
rect 240048 237458 240100 237464
rect 240060 223417 240088 237458
rect 240336 235657 240364 238682
rect 240322 235648 240378 235657
rect 240322 235583 240378 235592
rect 240704 235385 240732 240244
rect 240968 237448 241020 237454
rect 240968 237390 241020 237396
rect 240784 236020 240836 236026
rect 240784 235962 240836 235968
rect 240690 235376 240746 235385
rect 240690 235311 240746 235320
rect 240704 230489 240732 235311
rect 240690 230480 240746 230489
rect 240690 230415 240746 230424
rect 240796 227497 240824 235962
rect 240876 234660 240928 234666
rect 240876 234602 240928 234608
rect 240782 227488 240838 227497
rect 240782 227423 240838 227432
rect 240692 227112 240744 227118
rect 240692 227054 240744 227060
rect 240704 225690 240732 227054
rect 240692 225684 240744 225690
rect 240692 225626 240744 225632
rect 240046 223408 240102 223417
rect 240046 223343 240102 223352
rect 238852 209840 238904 209846
rect 238852 209782 238904 209788
rect 239772 209840 239824 209846
rect 239772 209782 239824 209788
rect 238864 208321 238892 209782
rect 240232 208344 240284 208350
rect 238850 208312 238906 208321
rect 240232 208286 240284 208292
rect 238850 208247 238906 208256
rect 238758 207768 238814 207777
rect 238758 207703 238814 207712
rect 238760 203652 238812 203658
rect 238760 203594 238812 203600
rect 238116 192500 238168 192506
rect 238116 192442 238168 192448
rect 238128 177410 238156 192442
rect 238116 177404 238168 177410
rect 238116 177346 238168 177352
rect 238022 174584 238078 174593
rect 238022 174519 238078 174528
rect 238116 173188 238168 173194
rect 238116 173130 238168 173136
rect 237472 168224 237524 168230
rect 237472 168166 237524 168172
rect 237378 166288 237434 166297
rect 237378 166223 237434 166232
rect 238022 164520 238078 164529
rect 238022 164455 238078 164464
rect 236920 160132 236972 160138
rect 236920 160074 236972 160080
rect 236828 128240 236880 128246
rect 236828 128182 236880 128188
rect 236736 127016 236788 127022
rect 236736 126958 236788 126964
rect 236644 124228 236696 124234
rect 236644 124170 236696 124176
rect 235540 123956 235592 123962
rect 235540 123898 235592 123904
rect 235448 122868 235500 122874
rect 235448 122810 235500 122816
rect 235354 104680 235410 104689
rect 235354 104615 235410 104624
rect 235356 96688 235408 96694
rect 235356 96630 235408 96636
rect 235368 36582 235396 96630
rect 235460 82113 235488 122810
rect 235446 82104 235502 82113
rect 235446 82039 235502 82048
rect 236656 76673 236684 124170
rect 236748 84969 236776 126958
rect 236932 120698 236960 160074
rect 237012 142860 237064 142866
rect 237012 142802 237064 142808
rect 237024 125497 237052 142802
rect 238036 128081 238064 164455
rect 238128 154873 238156 173130
rect 238390 167648 238446 167657
rect 238390 167583 238446 167592
rect 238300 164348 238352 164354
rect 238300 164290 238352 164296
rect 238208 158772 238260 158778
rect 238208 158714 238260 158720
rect 238114 154864 238170 154873
rect 238114 154799 238170 154808
rect 238116 147688 238168 147694
rect 238116 147630 238168 147636
rect 238022 128072 238078 128081
rect 238022 128007 238078 128016
rect 237010 125488 237066 125497
rect 237010 125423 237066 125432
rect 238024 124296 238076 124302
rect 238024 124238 238076 124244
rect 236920 120692 236972 120698
rect 236920 120634 236972 120640
rect 236734 84960 236790 84969
rect 236734 84895 236790 84904
rect 236642 76664 236698 76673
rect 236642 76599 236698 76608
rect 235356 36576 235408 36582
rect 235356 36518 235408 36524
rect 235264 13184 235316 13190
rect 235264 13126 235316 13132
rect 233976 11756 234028 11762
rect 233976 11698 234028 11704
rect 238036 4826 238064 124238
rect 238128 107574 238156 147630
rect 238220 118017 238248 158714
rect 238312 125594 238340 164290
rect 238404 159322 238432 167583
rect 238392 159316 238444 159322
rect 238392 159258 238444 159264
rect 238772 158030 238800 203594
rect 240140 196716 240192 196722
rect 240140 196658 240192 196664
rect 238944 186380 238996 186386
rect 238944 186322 238996 186328
rect 238852 181552 238904 181558
rect 238852 181494 238904 181500
rect 238760 158024 238812 158030
rect 238760 157966 238812 157972
rect 238864 146266 238892 181494
rect 238956 170377 238984 186322
rect 239034 176080 239090 176089
rect 239034 176015 239090 176024
rect 238942 170368 238998 170377
rect 238942 170303 238998 170312
rect 239048 163441 239076 176015
rect 239034 163432 239090 163441
rect 239034 163367 239090 163376
rect 239864 155984 239916 155990
rect 239864 155926 239916 155932
rect 238852 146260 238904 146266
rect 238852 146202 238904 146208
rect 239588 144968 239640 144974
rect 239588 144910 239640 144916
rect 239402 139496 239458 139505
rect 239402 139431 239458 139440
rect 238392 126268 238444 126274
rect 238392 126210 238444 126216
rect 238300 125588 238352 125594
rect 238300 125530 238352 125536
rect 238206 118008 238262 118017
rect 238206 117943 238262 117952
rect 238300 117972 238352 117978
rect 238300 117914 238352 117920
rect 238116 107568 238168 107574
rect 238116 107510 238168 107516
rect 238114 104000 238170 104009
rect 238114 103935 238170 103944
rect 238128 13122 238156 103935
rect 238312 101522 238340 117914
rect 238300 101516 238352 101522
rect 238300 101458 238352 101464
rect 238404 90438 238432 126210
rect 238392 90432 238444 90438
rect 238392 90374 238444 90380
rect 238116 13116 238168 13122
rect 238116 13058 238168 13064
rect 239416 6254 239444 139431
rect 239494 118824 239550 118833
rect 239494 118759 239550 118768
rect 239508 35222 239536 118759
rect 239600 103426 239628 144910
rect 239876 115569 239904 155926
rect 240152 154562 240180 196658
rect 240244 172514 240272 208286
rect 240796 182918 240824 227423
rect 240888 208350 240916 234602
rect 240980 211041 241008 237390
rect 241256 237386 241284 240244
rect 241808 240122 241836 240244
rect 241888 240168 241940 240174
rect 241808 240116 241888 240122
rect 241808 240110 241940 240116
rect 241808 240094 241928 240110
rect 241702 237552 241758 237561
rect 241702 237487 241758 237496
rect 241244 237380 241296 237386
rect 241244 237322 241296 237328
rect 241256 236026 241284 237322
rect 241244 236020 241296 236026
rect 241244 235962 241296 235968
rect 240966 211032 241022 211041
rect 240966 210967 241022 210976
rect 240876 208344 240928 208350
rect 240876 208286 240928 208292
rect 241612 198076 241664 198082
rect 241612 198018 241664 198024
rect 240784 182912 240836 182918
rect 240784 182854 240836 182860
rect 241058 179616 241114 179625
rect 241058 179551 241114 179560
rect 240876 173936 240928 173942
rect 240876 173878 240928 173884
rect 240232 172508 240284 172514
rect 240232 172450 240284 172456
rect 240784 168428 240836 168434
rect 240784 168370 240836 168376
rect 240140 154556 240192 154562
rect 240140 154498 240192 154504
rect 240796 129742 240824 168370
rect 240888 146985 240916 173878
rect 240968 171148 241020 171154
rect 240968 171090 241020 171096
rect 240874 146976 240930 146985
rect 240874 146911 240930 146920
rect 240980 145586 241008 171090
rect 241072 168450 241100 179551
rect 241520 177404 241572 177410
rect 241520 177346 241572 177352
rect 241532 171086 241560 177346
rect 241520 171080 241572 171086
rect 241520 171022 241572 171028
rect 241072 168422 241560 168450
rect 241532 160750 241560 168422
rect 241520 160744 241572 160750
rect 241520 160686 241572 160692
rect 241624 153950 241652 198018
rect 241716 174321 241744 237487
rect 241808 237425 241836 240094
rect 242176 239442 242204 240244
rect 242084 239414 242204 239442
rect 242084 238678 242112 239414
rect 242162 239320 242218 239329
rect 242162 239255 242218 239264
rect 242072 238672 242124 238678
rect 242072 238614 242124 238620
rect 241794 237416 241850 237425
rect 241794 237351 241850 237360
rect 242084 229094 242112 238614
rect 242176 238513 242204 239255
rect 242162 238504 242218 238513
rect 242162 238439 242218 238448
rect 242728 237522 242756 240244
rect 242716 237516 242768 237522
rect 242716 237458 242768 237464
rect 242256 236768 242308 236774
rect 242256 236710 242308 236716
rect 242268 234054 242296 236710
rect 243280 234666 243308 240244
rect 243648 238649 243676 240244
rect 243912 240236 243964 240242
rect 243912 240178 243964 240184
rect 243924 240106 243952 240178
rect 243912 240100 243964 240106
rect 243912 240042 243964 240048
rect 244016 238754 244044 254623
rect 244094 241360 244150 241369
rect 244094 241295 244150 241304
rect 244108 240310 244136 241295
rect 244096 240304 244148 240310
rect 244096 240246 244148 240252
rect 243924 238726 244044 238754
rect 243634 238640 243690 238649
rect 243634 238575 243690 238584
rect 243268 234660 243320 234666
rect 243268 234602 243320 234608
rect 242256 234048 242308 234054
rect 242256 233990 242308 233996
rect 242084 229066 242204 229094
rect 241702 174312 241758 174321
rect 241702 174247 241758 174256
rect 241612 153944 241664 153950
rect 241612 153886 241664 153892
rect 241060 153876 241112 153882
rect 241060 153818 241112 153824
rect 240968 145580 241020 145586
rect 240968 145522 241020 145528
rect 240968 143608 241020 143614
rect 240968 143550 241020 143556
rect 240784 129736 240836 129742
rect 240784 129678 240836 129684
rect 240874 128752 240930 128761
rect 240874 128687 240930 128696
rect 240784 116000 240836 116006
rect 240784 115942 240836 115948
rect 239862 115560 239918 115569
rect 239862 115495 239918 115504
rect 239678 115152 239734 115161
rect 239678 115087 239734 115096
rect 239588 103420 239640 103426
rect 239588 103362 239640 103368
rect 239692 73914 239720 115087
rect 239680 73908 239732 73914
rect 239680 73850 239732 73856
rect 239496 35216 239548 35222
rect 239496 35158 239548 35164
rect 240796 28286 240824 115942
rect 240888 47666 240916 128687
rect 240980 103494 241008 143550
rect 241072 114510 241100 153818
rect 242176 144906 242204 229066
rect 242268 219201 242296 233990
rect 243648 233073 243676 238575
rect 243634 233064 243690 233073
rect 243634 232999 243690 233008
rect 243544 229152 243596 229158
rect 243544 229094 243596 229100
rect 242900 229016 242952 229022
rect 242900 228958 242952 228964
rect 242912 228614 242940 228958
rect 242900 228608 242952 228614
rect 242900 228550 242952 228556
rect 242808 227792 242860 227798
rect 242808 227734 242860 227740
rect 242820 226001 242848 227734
rect 242806 225992 242862 226001
rect 242806 225927 242862 225936
rect 242254 219192 242310 219201
rect 242254 219127 242310 219136
rect 242254 172952 242310 172961
rect 242254 172887 242310 172896
rect 242164 144900 242216 144906
rect 242164 144842 242216 144848
rect 242268 133521 242296 172887
rect 242912 164150 242940 228550
rect 242992 189848 243044 189854
rect 242992 189790 243044 189796
rect 242900 164144 242952 164150
rect 242900 164086 242952 164092
rect 242438 150104 242494 150113
rect 242438 150039 242494 150048
rect 242346 146704 242402 146713
rect 242346 146639 242402 146648
rect 242254 133512 242310 133521
rect 242254 133447 242310 133456
rect 242162 117600 242218 117609
rect 242162 117535 242218 117544
rect 241060 114504 241112 114510
rect 241060 114446 241112 114452
rect 241152 113824 241204 113830
rect 241152 113766 241204 113772
rect 240968 103488 241020 103494
rect 240968 103430 241020 103436
rect 241060 100768 241112 100774
rect 241060 100710 241112 100716
rect 240968 78056 241020 78062
rect 240968 77998 241020 78004
rect 240876 47660 240928 47666
rect 240876 47602 240928 47608
rect 240784 28280 240836 28286
rect 240784 28222 240836 28228
rect 239404 6248 239456 6254
rect 239404 6190 239456 6196
rect 238024 4820 238076 4826
rect 238024 4762 238076 4768
rect 235816 4208 235868 4214
rect 235816 4150 235868 4156
rect 233884 2100 233936 2106
rect 233884 2042 233936 2048
rect 235828 480 235856 4150
rect 240508 3528 240560 3534
rect 240508 3470 240560 3476
rect 239312 2984 239364 2990
rect 239312 2926 239364 2932
rect 239324 480 239352 2926
rect 240520 480 240548 3470
rect 240980 2990 241008 77998
rect 241072 77994 241100 100710
rect 241164 83473 241192 113766
rect 241518 95704 241574 95713
rect 241518 95639 241574 95648
rect 241532 95266 241560 95639
rect 241520 95260 241572 95266
rect 241520 95202 241572 95208
rect 241150 83464 241206 83473
rect 241150 83399 241206 83408
rect 241060 77988 241112 77994
rect 241060 77930 241112 77936
rect 241520 51060 241572 51066
rect 241520 51002 241572 51008
rect 241532 16574 241560 51002
rect 242176 17270 242204 117535
rect 242254 110800 242310 110809
rect 242254 110735 242310 110744
rect 242268 50386 242296 110735
rect 242360 104825 242388 146639
rect 242452 108934 242480 150039
rect 243004 148753 243032 189790
rect 243556 169726 243584 229094
rect 243924 228614 243952 238726
rect 243912 228608 243964 228614
rect 243912 228550 243964 228556
rect 244292 172825 244320 270127
rect 244384 226137 244412 282367
rect 244476 271017 244504 298658
rect 245476 287088 245528 287094
rect 245476 287030 245528 287036
rect 244556 285048 244608 285054
rect 244556 284990 244608 284996
rect 244462 271008 244518 271017
rect 244462 270943 244518 270952
rect 244568 258233 244596 284990
rect 245488 284986 245516 287030
rect 245476 284980 245528 284986
rect 245476 284922 245528 284928
rect 245672 276729 245700 311782
rect 246316 311166 246344 351863
rect 246408 348430 246436 374070
rect 246396 348424 246448 348430
rect 246396 348366 246448 348372
rect 249616 346384 249668 346390
rect 249616 346326 249668 346332
rect 249628 345710 249656 346326
rect 248512 345704 248564 345710
rect 248512 345646 248564 345652
rect 249616 345704 249668 345710
rect 249616 345646 249668 345652
rect 248524 345545 248552 345646
rect 248510 345536 248566 345545
rect 248510 345471 248566 345480
rect 248420 339516 248472 339522
rect 248420 339458 248472 339464
rect 247682 335608 247738 335617
rect 247682 335543 247738 335552
rect 247222 334112 247278 334121
rect 247222 334047 247278 334056
rect 246304 311160 246356 311166
rect 246304 311102 246356 311108
rect 247132 304292 247184 304298
rect 247132 304234 247184 304240
rect 247040 300824 247092 300830
rect 247040 300766 247092 300772
rect 245750 289776 245806 289785
rect 245750 289711 245806 289720
rect 245764 288561 245792 289711
rect 245750 288552 245806 288561
rect 245750 288487 245806 288496
rect 245658 276720 245714 276729
rect 245658 276655 245714 276664
rect 245764 276162 245792 288487
rect 247052 287706 247080 300766
rect 247040 287700 247092 287706
rect 247040 287642 247092 287648
rect 247052 287054 247080 287642
rect 246960 287026 247080 287054
rect 246960 283801 246988 287026
rect 246946 283792 247002 283801
rect 246946 283727 247002 283736
rect 246854 283248 246910 283257
rect 246854 283183 246856 283192
rect 246908 283183 246910 283192
rect 246856 283154 246908 283160
rect 245936 282872 245988 282878
rect 245936 282814 245988 282820
rect 245948 281625 245976 282814
rect 245934 281616 245990 281625
rect 245934 281551 245990 281560
rect 245934 281072 245990 281081
rect 245934 281007 245990 281016
rect 245948 280838 245976 281007
rect 245936 280832 245988 280838
rect 245936 280774 245988 280780
rect 245936 280152 245988 280158
rect 245936 280094 245988 280100
rect 245948 278905 245976 280094
rect 245934 278896 245990 278905
rect 245934 278831 245990 278840
rect 246302 278080 246358 278089
rect 246302 278015 246358 278024
rect 245934 277536 245990 277545
rect 245934 277471 245990 277480
rect 245948 277438 245976 277471
rect 245936 277432 245988 277438
rect 245936 277374 245988 277380
rect 245672 276134 245792 276162
rect 245672 274553 245700 276134
rect 245752 276004 245804 276010
rect 245752 275946 245804 275952
rect 245764 275369 245792 275946
rect 245936 275936 245988 275942
rect 245934 275904 245936 275913
rect 245988 275904 245990 275913
rect 245934 275839 245990 275848
rect 245750 275360 245806 275369
rect 245750 275295 245806 275304
rect 245658 274544 245714 274553
rect 245658 274479 245714 274488
rect 245842 273728 245898 273737
rect 245842 273663 245898 273672
rect 245856 273290 245884 273663
rect 245844 273284 245896 273290
rect 245844 273226 245896 273232
rect 245936 273216 245988 273222
rect 245750 273184 245806 273193
rect 245936 273158 245988 273164
rect 245750 273119 245806 273128
rect 245764 272542 245792 273119
rect 245752 272536 245804 272542
rect 245752 272478 245804 272484
rect 245948 272377 245976 273158
rect 245934 272368 245990 272377
rect 245934 272303 245990 272312
rect 245934 271552 245990 271561
rect 245934 271487 245990 271496
rect 245948 271454 245976 271487
rect 245936 271448 245988 271454
rect 245936 271390 245988 271396
rect 245844 270496 245896 270502
rect 245844 270438 245896 270444
rect 245856 269657 245884 270438
rect 245842 269648 245898 269657
rect 245842 269583 245898 269592
rect 246316 268394 246344 278015
rect 246304 268388 246356 268394
rect 246304 268330 246356 268336
rect 245752 267708 245804 267714
rect 245752 267650 245804 267656
rect 245764 266665 245792 267650
rect 245750 266656 245806 266665
rect 245750 266591 245806 266600
rect 245660 265872 245712 265878
rect 245658 265840 245660 265849
rect 245712 265840 245714 265849
rect 245658 265775 245714 265784
rect 245844 264920 245896 264926
rect 245844 264862 245896 264868
rect 245856 263945 245884 264862
rect 246026 264480 246082 264489
rect 246026 264415 246082 264424
rect 245842 263936 245898 263945
rect 245842 263871 245898 263880
rect 245660 263424 245712 263430
rect 245660 263366 245712 263372
rect 244554 258224 244610 258233
rect 244554 258159 244610 258168
rect 244568 258126 244596 258159
rect 244556 258120 244608 258126
rect 244556 258062 244608 258068
rect 245672 256601 245700 263366
rect 245934 262304 245990 262313
rect 245934 262239 245936 262248
rect 245988 262239 245990 262248
rect 245936 262210 245988 262216
rect 245750 261760 245806 261769
rect 245750 261695 245806 261704
rect 245764 259894 245792 261695
rect 246040 261497 246068 264415
rect 246026 261488 246082 261497
rect 246026 261423 246082 261432
rect 245844 260976 245896 260982
rect 245842 260944 245844 260953
rect 245896 260944 245898 260953
rect 245842 260879 245898 260888
rect 245752 259888 245804 259894
rect 245752 259830 245804 259836
rect 246394 259584 246450 259593
rect 246394 259519 246450 259528
rect 246408 259486 246436 259519
rect 246396 259480 246448 259486
rect 246396 259422 246448 259428
rect 245752 259412 245804 259418
rect 245752 259354 245804 259360
rect 245764 258777 245792 259354
rect 245750 258768 245806 258777
rect 245750 258703 245806 258712
rect 245752 258052 245804 258058
rect 245752 257994 245804 258000
rect 245764 257417 245792 257994
rect 245750 257408 245806 257417
rect 245750 257343 245806 257352
rect 245658 256592 245714 256601
rect 245658 256527 245714 256536
rect 245672 256018 245700 256527
rect 245750 256048 245806 256057
rect 245660 256012 245712 256018
rect 245750 255983 245806 255992
rect 245660 255954 245712 255960
rect 245764 255406 245792 255983
rect 245752 255400 245804 255406
rect 245752 255342 245804 255348
rect 245844 255264 245896 255270
rect 245844 255206 245896 255212
rect 245856 254425 245884 255206
rect 245842 254416 245898 254425
rect 245842 254351 245898 254360
rect 246028 253904 246080 253910
rect 245934 253872 245990 253881
rect 246028 253846 246080 253852
rect 245934 253807 245936 253816
rect 245988 253807 245990 253816
rect 245936 253778 245988 253784
rect 246040 253065 246068 253846
rect 246026 253056 246082 253065
rect 246026 252991 246082 253000
rect 245936 252544 245988 252550
rect 245936 252486 245988 252492
rect 245948 252249 245976 252486
rect 245934 252240 245990 252249
rect 245934 252175 245990 252184
rect 245936 251864 245988 251870
rect 245936 251806 245988 251812
rect 245948 251705 245976 251806
rect 245934 251696 245990 251705
rect 245934 251631 245990 251640
rect 245844 251184 245896 251190
rect 245844 251126 245896 251132
rect 245856 250345 245884 251126
rect 245934 250880 245990 250889
rect 245934 250815 245990 250824
rect 245842 250336 245898 250345
rect 245842 250271 245898 250280
rect 245948 249762 245976 250815
rect 245936 249756 245988 249762
rect 245936 249698 245988 249704
rect 244462 248704 244518 248713
rect 244462 248639 244518 248648
rect 244476 233170 244504 248639
rect 245658 248160 245714 248169
rect 245658 248095 245714 248104
rect 245672 247722 245700 248095
rect 245660 247716 245712 247722
rect 245660 247658 245712 247664
rect 245934 247344 245990 247353
rect 245934 247279 245990 247288
rect 245948 247110 245976 247279
rect 245936 247104 245988 247110
rect 245936 247046 245988 247052
rect 245842 246528 245898 246537
rect 245842 246463 245898 246472
rect 244556 245744 244608 245750
rect 244556 245686 244608 245692
rect 244568 240038 244596 245686
rect 245856 245682 245884 246463
rect 245934 245984 245990 245993
rect 245934 245919 245990 245928
rect 245844 245676 245896 245682
rect 245844 245618 245896 245624
rect 245658 245168 245714 245177
rect 245658 245103 245714 245112
rect 244556 240032 244608 240038
rect 244556 239974 244608 239980
rect 244464 233164 244516 233170
rect 244464 233106 244516 233112
rect 244370 226128 244426 226137
rect 244370 226063 244426 226072
rect 244384 225321 244412 226063
rect 244370 225312 244426 225321
rect 244370 225247 244426 225256
rect 244370 225176 244426 225185
rect 244370 225111 244426 225120
rect 244384 219337 244412 225111
rect 244370 219328 244426 219337
rect 244370 219263 244426 219272
rect 245672 213926 245700 245103
rect 245948 244322 245976 245919
rect 246302 244624 246358 244633
rect 246302 244559 246358 244568
rect 245936 244316 245988 244322
rect 245936 244258 245988 244264
rect 245842 243808 245898 243817
rect 245842 243743 245898 243752
rect 245856 242962 245884 243743
rect 245844 242956 245896 242962
rect 245844 242898 245896 242904
rect 245750 241632 245806 241641
rect 245750 241567 245806 241576
rect 245764 241534 245792 241567
rect 245752 241528 245804 241534
rect 245752 241470 245804 241476
rect 245948 239329 245976 244258
rect 245934 239320 245990 239329
rect 245934 239255 245990 239264
rect 246316 224670 246344 244559
rect 246394 242448 246450 242457
rect 246394 242383 246450 242392
rect 246408 241602 246436 242383
rect 246396 241596 246448 241602
rect 246396 241538 246448 241544
rect 246946 240816 247002 240825
rect 247002 240774 247080 240802
rect 246946 240751 247002 240760
rect 247052 238754 247080 240774
rect 247144 240174 247172 304234
rect 247236 283218 247264 334047
rect 247696 302938 247724 335543
rect 247684 302932 247736 302938
rect 247684 302874 247736 302880
rect 247408 288516 247460 288522
rect 247408 288458 247460 288464
rect 247314 287872 247370 287881
rect 247314 287807 247370 287816
rect 247224 283212 247276 283218
rect 247224 283154 247276 283160
rect 247328 260137 247356 287807
rect 247314 260128 247370 260137
rect 247314 260063 247370 260072
rect 247224 241596 247276 241602
rect 247224 241538 247276 241544
rect 247132 240168 247184 240174
rect 247132 240110 247184 240116
rect 247052 238726 247172 238754
rect 246304 224664 246356 224670
rect 246304 224606 246356 224612
rect 246302 223408 246358 223417
rect 246302 223343 246358 223352
rect 245660 213920 245712 213926
rect 245660 213862 245712 213868
rect 244464 187740 244516 187746
rect 244464 187682 244516 187688
rect 244370 180024 244426 180033
rect 244370 179959 244426 179968
rect 244278 172816 244334 172825
rect 244278 172751 244334 172760
rect 243820 169788 243872 169794
rect 243820 169730 243872 169736
rect 243544 169720 243596 169726
rect 243544 169662 243596 169668
rect 243728 160200 243780 160206
rect 243728 160142 243780 160148
rect 242990 148744 243046 148753
rect 242990 148679 243046 148688
rect 243636 145036 243688 145042
rect 243636 144978 243688 144984
rect 242532 140072 242584 140078
rect 242532 140014 242584 140020
rect 242544 111722 242572 140014
rect 243542 138136 243598 138145
rect 243542 138071 243598 138080
rect 242532 111716 242584 111722
rect 242532 111658 242584 111664
rect 242440 108928 242492 108934
rect 242440 108870 242492 108876
rect 242346 104816 242402 104825
rect 242346 104751 242402 104760
rect 242530 104136 242586 104145
rect 242530 104071 242586 104080
rect 242346 100056 242402 100065
rect 242346 99991 242402 100000
rect 242360 75313 242388 99991
rect 242544 91798 242572 104071
rect 242532 91792 242584 91798
rect 242532 91734 242584 91740
rect 242346 75304 242402 75313
rect 242346 75239 242402 75248
rect 242256 50380 242308 50386
rect 242256 50322 242308 50328
rect 243556 49026 243584 138071
rect 243648 104786 243676 144978
rect 243740 120086 243768 160142
rect 243832 140146 243860 169730
rect 243910 153232 243966 153241
rect 243910 153167 243966 153176
rect 243820 140140 243872 140146
rect 243820 140082 243872 140088
rect 243924 124817 243952 153167
rect 244384 137970 244412 179959
rect 244476 156602 244504 187682
rect 244924 174548 244976 174554
rect 244924 174490 244976 174496
rect 244936 159390 244964 174490
rect 245016 162920 245068 162926
rect 245016 162862 245068 162868
rect 244924 159384 244976 159390
rect 244924 159326 244976 159332
rect 244924 157480 244976 157486
rect 244924 157422 244976 157428
rect 244464 156596 244516 156602
rect 244464 156538 244516 156544
rect 244372 137964 244424 137970
rect 244372 137906 244424 137912
rect 243910 124808 243966 124817
rect 243910 124743 243966 124752
rect 243728 120080 243780 120086
rect 243728 120022 243780 120028
rect 244936 117230 244964 157422
rect 245028 122738 245056 162862
rect 245672 150482 245700 213862
rect 245752 192568 245804 192574
rect 245752 192510 245804 192516
rect 245660 150476 245712 150482
rect 245660 150418 245712 150424
rect 245198 145616 245254 145625
rect 245198 145551 245254 145560
rect 245108 125656 245160 125662
rect 245108 125598 245160 125604
rect 245016 122732 245068 122738
rect 245016 122674 245068 122680
rect 244924 117224 244976 117230
rect 244924 117166 244976 117172
rect 244922 113384 244978 113393
rect 244922 113319 244978 113328
rect 243728 110492 243780 110498
rect 243728 110434 243780 110440
rect 243636 104780 243688 104786
rect 243636 104722 243688 104728
rect 243740 93158 243768 110434
rect 243728 93152 243780 93158
rect 243728 93094 243780 93100
rect 244280 54596 244332 54602
rect 244280 54538 244332 54544
rect 243544 49020 243596 49026
rect 243544 48962 243596 48968
rect 242898 26888 242954 26897
rect 242898 26823 242954 26832
rect 242164 17264 242216 17270
rect 242164 17206 242216 17212
rect 241532 16546 241744 16574
rect 240968 2984 241020 2990
rect 240968 2926 241020 2932
rect 241716 480 241744 16546
rect 242912 11762 242940 26823
rect 244292 16574 244320 54538
rect 244936 39370 244964 113319
rect 245016 104916 245068 104922
rect 245016 104858 245068 104864
rect 245028 60042 245056 104858
rect 245120 84862 245148 125598
rect 245212 107545 245240 145551
rect 245764 140185 245792 192510
rect 246316 182850 246344 223343
rect 247144 206922 247172 238726
rect 247236 233986 247264 241538
rect 247224 233980 247276 233986
rect 247224 233922 247276 233928
rect 247224 224664 247276 224670
rect 247224 224606 247276 224612
rect 247236 206990 247264 224606
rect 247224 206984 247276 206990
rect 247224 206926 247276 206932
rect 247132 206916 247184 206922
rect 247132 206858 247184 206864
rect 247236 200114 247264 206926
rect 247052 200086 247264 200114
rect 246304 182844 246356 182850
rect 246304 182786 246356 182792
rect 245842 181384 245898 181393
rect 245842 181319 245898 181328
rect 245750 140176 245806 140185
rect 245750 140111 245806 140120
rect 245856 136610 245884 181319
rect 245934 174584 245990 174593
rect 245934 174519 245990 174528
rect 245948 144129 245976 174519
rect 247052 167113 247080 200086
rect 247224 175976 247276 175982
rect 247224 175918 247276 175924
rect 247038 167104 247094 167113
rect 247038 167039 247094 167048
rect 246488 151156 246540 151162
rect 246488 151098 246540 151104
rect 245934 144120 245990 144129
rect 245934 144055 245990 144064
rect 246396 143676 246448 143682
rect 246396 143618 246448 143624
rect 245844 136604 245896 136610
rect 245844 136546 245896 136552
rect 245290 135960 245346 135969
rect 245290 135895 245346 135904
rect 245304 126274 245332 135895
rect 245292 126268 245344 126274
rect 245292 126210 245344 126216
rect 246302 121680 246358 121689
rect 246302 121615 246358 121624
rect 245198 107536 245254 107545
rect 245198 107471 245254 107480
rect 245108 84856 245160 84862
rect 245108 84798 245160 84804
rect 245016 60036 245068 60042
rect 245016 59978 245068 59984
rect 244924 39364 244976 39370
rect 244924 39306 244976 39312
rect 246316 32502 246344 121615
rect 246408 109750 246436 143618
rect 246500 118046 246528 151098
rect 247236 147014 247264 175918
rect 247420 164218 247448 288458
rect 248432 270230 248460 339458
rect 248696 291304 248748 291310
rect 248696 291246 248748 291252
rect 248512 287156 248564 287162
rect 248512 287098 248564 287104
rect 248420 270224 248472 270230
rect 248420 270166 248472 270172
rect 248420 260976 248472 260982
rect 248420 260918 248472 260924
rect 247960 171216 248012 171222
rect 247960 171158 248012 171164
rect 247408 164212 247460 164218
rect 247408 164154 247460 164160
rect 247776 161560 247828 161566
rect 247776 161502 247828 161508
rect 247224 147008 247276 147014
rect 247224 146950 247276 146956
rect 246670 132832 246726 132841
rect 246670 132767 246726 132776
rect 246488 118040 246540 118046
rect 246488 117982 246540 117988
rect 246396 109744 246448 109750
rect 246396 109686 246448 109692
rect 246578 108080 246634 108089
rect 246578 108015 246634 108024
rect 246488 106344 246540 106350
rect 246488 106286 246540 106292
rect 246396 76560 246448 76566
rect 246396 76502 246448 76508
rect 246304 32496 246356 32502
rect 246304 32438 246356 32444
rect 244292 16546 245240 16574
rect 242900 11756 242952 11762
rect 242900 11698 242952 11704
rect 244096 11756 244148 11762
rect 244096 11698 244148 11704
rect 242898 7576 242954 7585
rect 242898 7511 242954 7520
rect 242912 2786 242940 7511
rect 242900 2780 242952 2786
rect 242900 2722 242952 2728
rect 242912 480 242940 2722
rect 244108 480 244136 11698
rect 245212 480 245240 16546
rect 246212 4820 246264 4826
rect 246212 4762 246264 4768
rect 246224 3913 246252 4762
rect 246210 3904 246266 3913
rect 246266 3862 246344 3890
rect 246210 3839 246266 3848
rect 246316 2938 246344 3862
rect 246408 3534 246436 76502
rect 246500 64297 246528 106286
rect 246592 76537 246620 108015
rect 246684 105641 246712 132767
rect 247684 131164 247736 131170
rect 247684 131106 247736 131112
rect 246670 105632 246726 105641
rect 246670 105567 246726 105576
rect 246578 76528 246634 76537
rect 246578 76463 246634 76472
rect 246486 64288 246542 64297
rect 246486 64223 246542 64232
rect 247696 57225 247724 131106
rect 247788 121446 247816 161502
rect 247866 141400 247922 141409
rect 247866 141335 247922 141344
rect 247776 121440 247828 121446
rect 247776 121382 247828 121388
rect 247880 102134 247908 141335
rect 247972 132462 248000 171158
rect 248052 158840 248104 158846
rect 248052 158782 248104 158788
rect 247960 132456 248012 132462
rect 247960 132398 248012 132404
rect 248064 123486 248092 158782
rect 248432 145761 248460 260918
rect 248524 229158 248552 287098
rect 248604 271448 248656 271454
rect 248604 271390 248656 271396
rect 248512 229152 248564 229158
rect 248512 229094 248564 229100
rect 248616 222154 248644 271390
rect 248708 260982 248736 291246
rect 249720 282266 249748 377604
rect 251376 374746 251404 377604
rect 252572 377590 253046 377618
rect 250444 374740 250496 374746
rect 250444 374682 250496 374688
rect 251364 374740 251416 374746
rect 251364 374682 251416 374688
rect 249892 340944 249944 340950
rect 249892 340886 249944 340892
rect 249800 283212 249852 283218
rect 249800 283154 249852 283160
rect 249708 282260 249760 282266
rect 249708 282202 249760 282208
rect 249706 279440 249762 279449
rect 249706 279375 249762 279384
rect 249720 278798 249748 279375
rect 249708 278792 249760 278798
rect 249708 278734 249760 278740
rect 248696 260976 248748 260982
rect 248696 260918 248748 260924
rect 248696 249756 248748 249762
rect 248696 249698 248748 249704
rect 248604 222148 248656 222154
rect 248604 222090 248656 222096
rect 248616 222057 248644 222090
rect 248602 222048 248658 222057
rect 248602 221983 248658 221992
rect 248708 211070 248736 249698
rect 249706 213752 249762 213761
rect 249706 213687 249762 213696
rect 249720 212566 249748 213687
rect 249708 212560 249760 212566
rect 249708 212502 249760 212508
rect 248696 211064 248748 211070
rect 248696 211006 248748 211012
rect 248708 200114 248736 211006
rect 248524 200086 248736 200114
rect 248524 156777 248552 200086
rect 249246 174312 249302 174321
rect 249246 174247 249302 174256
rect 249062 159080 249118 159089
rect 249062 159015 249118 159024
rect 248510 156768 248566 156777
rect 248510 156703 248566 156712
rect 248418 145752 248474 145761
rect 248418 145687 248474 145696
rect 248052 123480 248104 123486
rect 248052 123422 248104 123428
rect 247960 119400 248012 119406
rect 247960 119342 248012 119348
rect 247868 102128 247920 102134
rect 247868 102070 247920 102076
rect 247774 100872 247830 100881
rect 247774 100807 247830 100816
rect 247682 57216 247738 57225
rect 247682 57151 247738 57160
rect 247684 49020 247736 49026
rect 247684 48962 247736 48968
rect 247696 6914 247724 48962
rect 247788 48929 247816 100807
rect 247972 87650 248000 119342
rect 249076 118697 249104 159015
rect 249156 146328 249208 146334
rect 249156 146270 249208 146276
rect 249062 118688 249118 118697
rect 249062 118623 249118 118632
rect 249064 110560 249116 110566
rect 249064 110502 249116 110508
rect 247960 87644 248012 87650
rect 247960 87586 248012 87592
rect 247774 48920 247830 48929
rect 247774 48855 247830 48864
rect 249076 40798 249104 110502
rect 249168 106282 249196 146270
rect 249260 135182 249288 174247
rect 249812 151094 249840 283154
rect 249904 265878 249932 340886
rect 249982 297120 250038 297129
rect 249982 297055 250038 297064
rect 249892 265872 249944 265878
rect 249892 265814 249944 265820
rect 249892 259888 249944 259894
rect 249892 259830 249944 259836
rect 249904 205562 249932 259830
rect 249996 255406 250024 297055
rect 249984 255400 250036 255406
rect 249984 255342 250036 255348
rect 249892 205556 249944 205562
rect 249892 205498 249944 205504
rect 249904 162489 249932 205498
rect 250456 202473 250484 374682
rect 252572 356794 252600 377590
rect 254688 374814 254716 377604
rect 255976 377590 256358 377618
rect 256804 377590 258014 377618
rect 259472 377590 259854 377618
rect 254676 374808 254728 374814
rect 254676 374750 254728 374756
rect 255412 374808 255464 374814
rect 255412 374750 255464 374756
rect 253202 364984 253258 364993
rect 253202 364919 253258 364928
rect 252560 356788 252612 356794
rect 252560 356730 252612 356736
rect 252650 332888 252706 332897
rect 252650 332823 252706 332832
rect 252468 318096 252520 318102
rect 252468 318038 252520 318044
rect 251272 313948 251324 313954
rect 251272 313890 251324 313896
rect 251180 302932 251232 302938
rect 251180 302874 251232 302880
rect 251192 272542 251220 302874
rect 251180 272536 251232 272542
rect 251180 272478 251232 272484
rect 251088 255400 251140 255406
rect 251088 255342 251140 255348
rect 251100 254590 251128 255342
rect 251088 254584 251140 254590
rect 251088 254526 251140 254532
rect 250442 202464 250498 202473
rect 250442 202399 250498 202408
rect 250720 168496 250772 168502
rect 250720 168438 250772 168444
rect 250442 166016 250498 166025
rect 250442 165951 250498 165960
rect 249890 162480 249946 162489
rect 249890 162415 249946 162424
rect 249800 151088 249852 151094
rect 249800 151030 249852 151036
rect 249340 141500 249392 141506
rect 249340 141442 249392 141448
rect 249248 135176 249300 135182
rect 249248 135118 249300 135124
rect 249248 120760 249300 120766
rect 249248 120702 249300 120708
rect 249156 106276 249208 106282
rect 249156 106218 249208 106224
rect 249156 102196 249208 102202
rect 249156 102138 249208 102144
rect 249168 65521 249196 102138
rect 249260 82142 249288 120702
rect 249352 113082 249380 141442
rect 250456 126954 250484 165951
rect 250534 150920 250590 150929
rect 250534 150855 250590 150864
rect 250444 126948 250496 126954
rect 250444 126890 250496 126896
rect 250444 117360 250496 117366
rect 250444 117302 250496 117308
rect 249340 113076 249392 113082
rect 249340 113018 249392 113024
rect 249248 82136 249300 82142
rect 249248 82078 249300 82084
rect 249154 65512 249210 65521
rect 249154 65447 249210 65456
rect 249800 51060 249852 51066
rect 249800 51002 249852 51008
rect 249812 50969 249840 51002
rect 249798 50960 249854 50969
rect 249798 50895 249854 50904
rect 249154 46200 249210 46209
rect 249154 46135 249210 46144
rect 249064 40792 249116 40798
rect 249064 40734 249116 40740
rect 249168 16590 249196 46135
rect 249156 16584 249208 16590
rect 249156 16526 249208 16532
rect 249708 16584 249760 16590
rect 249708 16526 249760 16532
rect 247604 6886 247724 6914
rect 247604 4146 247632 6886
rect 247592 4140 247644 4146
rect 247592 4082 247644 4088
rect 246396 3528 246448 3534
rect 246396 3470 246448 3476
rect 246316 2910 246436 2938
rect 246408 480 246436 2910
rect 247604 480 247632 4082
rect 249720 3534 249748 16526
rect 249982 13832 250038 13841
rect 249982 13767 250038 13776
rect 248788 3528 248840 3534
rect 248788 3470 248840 3476
rect 249708 3528 249760 3534
rect 249708 3470 249760 3476
rect 248800 480 248828 3470
rect 249996 480 250024 13767
rect 250456 8974 250484 117302
rect 250548 111081 250576 150855
rect 250732 146946 250760 168438
rect 251192 160041 251220 272478
rect 251284 249801 251312 313890
rect 251824 285728 251876 285734
rect 251824 285670 251876 285676
rect 251836 272610 251864 285670
rect 251824 272604 251876 272610
rect 251824 272546 251876 272552
rect 251362 252512 251418 252521
rect 251362 252447 251418 252456
rect 251376 251870 251404 252447
rect 251364 251864 251416 251870
rect 251364 251806 251416 251812
rect 252376 251864 252428 251870
rect 252376 251806 252428 251812
rect 252388 251258 252416 251806
rect 252376 251252 252428 251258
rect 252376 251194 252428 251200
rect 251270 249792 251326 249801
rect 251270 249727 251326 249736
rect 252374 249792 252430 249801
rect 252374 249727 252430 249736
rect 251284 248985 251312 249727
rect 251270 248976 251326 248985
rect 251270 248911 251326 248920
rect 251272 247104 251324 247110
rect 251272 247046 251324 247052
rect 251284 210769 251312 247046
rect 252388 244934 252416 249727
rect 252376 244928 252428 244934
rect 252376 244870 252428 244876
rect 252480 238746 252508 318038
rect 252560 294092 252612 294098
rect 252560 294034 252612 294040
rect 252468 238740 252520 238746
rect 252468 238682 252520 238688
rect 252480 238134 252508 238682
rect 252468 238128 252520 238134
rect 252468 238070 252520 238076
rect 251914 215928 251970 215937
rect 251914 215863 251970 215872
rect 251928 215257 251956 215863
rect 251914 215248 251970 215257
rect 251914 215183 251970 215192
rect 251270 210760 251326 210769
rect 251270 210695 251326 210704
rect 252572 173194 252600 294034
rect 252664 238678 252692 332823
rect 253216 319462 253244 364919
rect 254582 338736 254638 338745
rect 254582 338671 254638 338680
rect 254596 323610 254624 338671
rect 255424 326398 255452 374750
rect 255976 374134 256004 377590
rect 255964 374128 256016 374134
rect 255964 374070 256016 374076
rect 255412 326392 255464 326398
rect 255412 326334 255464 326340
rect 254584 323604 254636 323610
rect 254584 323546 254636 323552
rect 255320 319524 255372 319530
rect 255320 319466 255372 319472
rect 253204 319456 253256 319462
rect 253204 319398 253256 319404
rect 253938 318880 253994 318889
rect 253938 318815 253994 318824
rect 252836 312588 252888 312594
rect 252836 312530 252888 312536
rect 252742 261488 252798 261497
rect 252742 261423 252798 261432
rect 252652 238672 252704 238678
rect 252652 238614 252704 238620
rect 252756 195906 252784 261423
rect 252848 255270 252876 312530
rect 253952 275942 253980 318815
rect 254214 308544 254270 308553
rect 254214 308479 254270 308488
rect 254124 282260 254176 282266
rect 254124 282202 254176 282208
rect 254032 278044 254084 278050
rect 254032 277986 254084 277992
rect 254044 277438 254072 277986
rect 254032 277432 254084 277438
rect 254032 277374 254084 277380
rect 253940 275936 253992 275942
rect 253940 275878 253992 275884
rect 253952 275330 253980 275878
rect 253940 275324 253992 275330
rect 253940 275266 253992 275272
rect 253940 273284 253992 273290
rect 253940 273226 253992 273232
rect 253202 269240 253258 269249
rect 253202 269175 253258 269184
rect 253216 268462 253244 269175
rect 253204 268456 253256 268462
rect 253204 268398 253256 268404
rect 252836 255264 252888 255270
rect 252836 255206 252888 255212
rect 252848 254658 252876 255206
rect 252836 254652 252888 254658
rect 252836 254594 252888 254600
rect 253202 211848 253258 211857
rect 253202 211783 253258 211792
rect 252744 195900 252796 195906
rect 252744 195842 252796 195848
rect 252650 183696 252706 183705
rect 252650 183631 252706 183640
rect 252560 173188 252612 173194
rect 252560 173130 252612 173136
rect 251822 168600 251878 168609
rect 251822 168535 251878 168544
rect 251178 160032 251234 160041
rect 251178 159967 251234 159976
rect 250720 146940 250772 146946
rect 250720 146882 250772 146888
rect 250628 146396 250680 146402
rect 250628 146338 250680 146344
rect 250534 111072 250590 111081
rect 250534 111007 250590 111016
rect 250536 109064 250588 109070
rect 250536 109006 250588 109012
rect 250548 54534 250576 109006
rect 250640 104854 250668 146338
rect 251836 141438 251864 168535
rect 252100 167068 252152 167074
rect 252100 167010 252152 167016
rect 251914 154864 251970 154873
rect 251914 154799 251970 154808
rect 251824 141432 251876 141438
rect 251824 141374 251876 141380
rect 251824 131232 251876 131238
rect 251824 131174 251876 131180
rect 250718 105632 250774 105641
rect 250718 105567 250774 105576
rect 250628 104848 250680 104854
rect 250628 104790 250680 104796
rect 250732 87689 250760 105567
rect 250718 87680 250774 87689
rect 250718 87615 250774 87624
rect 250536 54528 250588 54534
rect 250536 54470 250588 54476
rect 251836 51785 251864 131174
rect 251928 115258 251956 154799
rect 252008 150476 252060 150482
rect 252008 150418 252060 150424
rect 251916 115252 251968 115258
rect 251916 115194 251968 115200
rect 251916 111852 251968 111858
rect 251916 111794 251968 111800
rect 251928 69698 251956 111794
rect 252020 110430 252048 150418
rect 252112 128314 252140 167010
rect 252664 149054 252692 183631
rect 252756 172417 252784 195842
rect 253216 192506 253244 211783
rect 253204 192500 253256 192506
rect 253204 192442 253256 192448
rect 253952 178673 253980 273226
rect 254044 217841 254072 277374
rect 254136 231849 254164 282202
rect 254228 273222 254256 308479
rect 254584 289944 254636 289950
rect 254584 289886 254636 289892
rect 254596 282198 254624 289886
rect 254584 282192 254636 282198
rect 254584 282134 254636 282140
rect 254216 273216 254268 273222
rect 254216 273158 254268 273164
rect 254228 272542 254256 273158
rect 254216 272536 254268 272542
rect 254216 272478 254268 272484
rect 255332 267889 255360 319466
rect 255976 310321 256004 374070
rect 256700 311160 256752 311166
rect 256700 311102 256752 311108
rect 256146 310448 256202 310457
rect 256146 310383 256202 310392
rect 255962 310312 256018 310321
rect 255962 310247 256018 310256
rect 255962 298208 256018 298217
rect 255962 298143 256018 298152
rect 255410 291816 255466 291825
rect 255410 291751 255466 291760
rect 255318 267880 255374 267889
rect 255318 267815 255374 267824
rect 255332 265674 255360 267815
rect 255424 266257 255452 291751
rect 255504 286340 255556 286346
rect 255504 286282 255556 286288
rect 255516 280158 255544 286282
rect 255504 280152 255556 280158
rect 255504 280094 255556 280100
rect 255410 266248 255466 266257
rect 255410 266183 255466 266192
rect 255320 265668 255372 265674
rect 255320 265610 255372 265616
rect 255424 265577 255452 266183
rect 255410 265568 255466 265577
rect 255410 265503 255466 265512
rect 255320 262268 255372 262274
rect 255320 262210 255372 262216
rect 254122 231840 254178 231849
rect 254122 231775 254178 231784
rect 254136 231169 254164 231775
rect 254122 231160 254178 231169
rect 254122 231095 254178 231104
rect 254030 217832 254086 217841
rect 254030 217767 254086 217776
rect 255332 200802 255360 262210
rect 255410 245712 255466 245721
rect 255410 245647 255412 245656
rect 255464 245647 255466 245656
rect 255412 245618 255464 245624
rect 255320 200796 255372 200802
rect 255320 200738 255372 200744
rect 255424 195974 255452 245618
rect 255976 196722 256004 298143
rect 256160 291825 256188 310383
rect 256146 291816 256202 291825
rect 256146 291751 256202 291760
rect 256712 240281 256740 311102
rect 256804 310457 256832 377590
rect 258724 375352 258776 375358
rect 258724 375294 258776 375300
rect 258078 367704 258134 367713
rect 258078 367639 258134 367648
rect 256790 310448 256846 310457
rect 256790 310383 256846 310392
rect 257342 310312 257398 310321
rect 257342 310247 257398 310256
rect 256790 303784 256846 303793
rect 256790 303719 256846 303728
rect 256804 258058 256832 303719
rect 256792 258052 256844 258058
rect 256792 257994 256844 258000
rect 256804 257378 256832 257994
rect 256792 257372 256844 257378
rect 256792 257314 256844 257320
rect 256698 240272 256754 240281
rect 256698 240207 256754 240216
rect 256712 233918 256740 240207
rect 256700 233912 256752 233918
rect 256700 233854 256752 233860
rect 255964 196716 256016 196722
rect 255964 196658 256016 196664
rect 255412 195968 255464 195974
rect 255412 195910 255464 195916
rect 254032 184204 254084 184210
rect 254032 184146 254084 184152
rect 253938 178664 253994 178673
rect 253938 178599 253994 178608
rect 252742 172408 252798 172417
rect 252742 172343 252798 172352
rect 253478 171592 253534 171601
rect 253478 171527 253534 171536
rect 253296 156052 253348 156058
rect 253296 155994 253348 156000
rect 252652 149048 252704 149054
rect 252652 148990 252704 148996
rect 253202 132968 253258 132977
rect 253202 132903 253258 132912
rect 252100 128308 252152 128314
rect 252100 128250 252152 128256
rect 252100 122120 252152 122126
rect 252100 122062 252152 122068
rect 252008 110424 252060 110430
rect 252008 110366 252060 110372
rect 252112 83502 252140 122062
rect 252100 83496 252152 83502
rect 252100 83438 252152 83444
rect 251916 69692 251968 69698
rect 251916 69634 251968 69640
rect 253216 62830 253244 132903
rect 253308 115938 253336 155994
rect 253388 149116 253440 149122
rect 253388 149058 253440 149064
rect 253296 115932 253348 115938
rect 253296 115874 253348 115880
rect 253400 109002 253428 149058
rect 253492 132433 253520 171527
rect 254044 139398 254072 184146
rect 254584 180124 254636 180130
rect 254584 180066 254636 180072
rect 254596 152969 254624 180066
rect 254676 172576 254728 172582
rect 254676 172518 254728 172524
rect 254582 152960 254638 152969
rect 254582 152895 254638 152904
rect 254584 139460 254636 139466
rect 254584 139402 254636 139408
rect 254032 139392 254084 139398
rect 254032 139334 254084 139340
rect 253478 132424 253534 132433
rect 253478 132359 253534 132368
rect 253480 113212 253532 113218
rect 253480 113154 253532 113160
rect 253388 108996 253440 109002
rect 253388 108938 253440 108944
rect 253294 107808 253350 107817
rect 253294 107743 253350 107752
rect 253204 62824 253256 62830
rect 253204 62766 253256 62772
rect 251822 51776 251878 51785
rect 251822 51711 251878 51720
rect 253308 43518 253336 107743
rect 253492 75177 253520 113154
rect 253478 75168 253534 75177
rect 253478 75103 253534 75112
rect 254596 68377 254624 139402
rect 254688 133890 254716 172518
rect 256056 167136 256108 167142
rect 256056 167078 256108 167084
rect 255964 162988 256016 162994
rect 255964 162930 256016 162936
rect 254766 151872 254822 151881
rect 254766 151807 254822 151816
rect 254676 133884 254728 133890
rect 254676 133826 254728 133832
rect 254674 114608 254730 114617
rect 254674 114543 254730 114552
rect 254582 68368 254638 68377
rect 254582 68303 254638 68312
rect 254688 50289 254716 114543
rect 254780 110401 254808 151807
rect 255976 142769 256004 162930
rect 255962 142760 256018 142769
rect 255962 142695 256018 142704
rect 256068 133210 256096 167078
rect 256240 147756 256292 147762
rect 256240 147698 256292 147704
rect 256146 142760 256202 142769
rect 256146 142695 256202 142704
rect 256056 133204 256108 133210
rect 256056 133146 256108 133152
rect 255964 132524 256016 132530
rect 255964 132466 256016 132472
rect 254860 128376 254912 128382
rect 254860 128318 254912 128324
rect 254872 113830 254900 128318
rect 254860 113824 254912 113830
rect 254860 113766 254912 113772
rect 254766 110392 254822 110401
rect 254766 110327 254822 110336
rect 254768 103556 254820 103562
rect 254768 103498 254820 103504
rect 254780 91769 254808 103498
rect 254766 91760 254822 91769
rect 254766 91695 254822 91704
rect 255976 65657 256004 132466
rect 256056 109132 256108 109138
rect 256056 109074 256108 109080
rect 255962 65648 256018 65657
rect 255962 65583 256018 65592
rect 256068 55894 256096 109074
rect 256160 100638 256188 142695
rect 256252 116521 256280 147698
rect 256238 116512 256294 116521
rect 256238 116447 256294 116456
rect 256240 114572 256292 114578
rect 256240 114514 256292 114520
rect 256148 100632 256200 100638
rect 256148 100574 256200 100580
rect 256252 87718 256280 114514
rect 256240 87712 256292 87718
rect 256240 87654 256292 87660
rect 257356 86970 257384 310247
rect 258092 219434 258120 367639
rect 258736 360874 258764 375294
rect 258172 360868 258224 360874
rect 258172 360810 258224 360816
rect 258724 360868 258776 360874
rect 258724 360810 258776 360816
rect 258184 289134 258212 360810
rect 259472 359514 259500 377590
rect 261496 375358 261524 377604
rect 262232 377590 263166 377618
rect 263704 377590 264822 377618
rect 266372 377590 266478 377618
rect 267752 377590 268134 377618
rect 269132 377590 269790 377618
rect 270512 377590 271446 377618
rect 272720 377590 273102 377618
rect 261484 375352 261536 375358
rect 261484 375294 261536 375300
rect 261484 374740 261536 374746
rect 261484 374682 261536 374688
rect 259460 359508 259512 359514
rect 259460 359450 259512 359456
rect 259368 327752 259420 327758
rect 259368 327694 259420 327700
rect 259380 327078 259408 327694
rect 259368 327072 259420 327078
rect 259368 327014 259420 327020
rect 258264 302252 258316 302258
rect 258264 302194 258316 302200
rect 258172 289128 258224 289134
rect 258172 289070 258224 289076
rect 258172 284980 258224 284986
rect 258172 284922 258224 284928
rect 258080 219428 258132 219434
rect 258080 219370 258132 219376
rect 258184 174554 258212 284922
rect 258276 253842 258304 302194
rect 258264 253836 258316 253842
rect 258264 253778 258316 253784
rect 259276 253836 259328 253842
rect 259276 253778 259328 253784
rect 259288 253298 259316 253778
rect 259276 253292 259328 253298
rect 259276 253234 259328 253240
rect 259276 243568 259328 243574
rect 259276 243510 259328 243516
rect 259288 242962 259316 243510
rect 258264 242956 258316 242962
rect 258264 242898 258316 242904
rect 259276 242956 259328 242962
rect 259276 242898 259328 242904
rect 258276 227798 258304 242898
rect 258264 227792 258316 227798
rect 258264 227734 258316 227740
rect 258724 227792 258776 227798
rect 258724 227734 258776 227740
rect 258736 185706 258764 227734
rect 259276 219428 259328 219434
rect 259276 219370 259328 219376
rect 259288 218754 259316 219370
rect 259276 218748 259328 218754
rect 259276 218690 259328 218696
rect 259380 211041 259408 327014
rect 259472 321638 259500 359450
rect 261496 346390 261524 374682
rect 261484 346384 261536 346390
rect 261484 346326 261536 346332
rect 260104 342916 260156 342922
rect 260104 342858 260156 342864
rect 260116 332586 260144 342858
rect 260932 337408 260984 337414
rect 260932 337350 260984 337356
rect 260104 332580 260156 332586
rect 260104 332522 260156 332528
rect 260116 331294 260144 332522
rect 260104 331288 260156 331294
rect 260104 331230 260156 331236
rect 260748 331288 260800 331294
rect 260748 331230 260800 331236
rect 259552 329792 259604 329798
rect 259552 329734 259604 329740
rect 259564 328545 259592 329734
rect 259550 328536 259606 328545
rect 259550 328471 259606 328480
rect 259460 321632 259512 321638
rect 259460 321574 259512 321580
rect 260104 321632 260156 321638
rect 260104 321574 260156 321580
rect 259460 317552 259512 317558
rect 259460 317494 259512 317500
rect 259472 251190 259500 317494
rect 260116 312594 260144 321574
rect 260104 312588 260156 312594
rect 260104 312530 260156 312536
rect 260104 287700 260156 287706
rect 260104 287642 260156 287648
rect 259550 285968 259606 285977
rect 259550 285903 259606 285912
rect 259460 251184 259512 251190
rect 259460 251126 259512 251132
rect 259564 222193 259592 285903
rect 260116 248414 260144 287642
rect 260760 282946 260788 331230
rect 260840 283620 260892 283626
rect 260840 283562 260892 283568
rect 260748 282940 260800 282946
rect 260748 282882 260800 282888
rect 260748 251184 260800 251190
rect 260748 251126 260800 251132
rect 260760 250510 260788 251126
rect 260748 250504 260800 250510
rect 260748 250446 260800 250452
rect 260116 248386 260236 248414
rect 260104 245676 260156 245682
rect 260104 245618 260156 245624
rect 260116 240009 260144 245618
rect 260208 240786 260236 248386
rect 260746 242992 260802 243001
rect 260746 242927 260748 242936
rect 260800 242927 260802 242936
rect 260748 242898 260800 242904
rect 260196 240780 260248 240786
rect 260196 240722 260248 240728
rect 260102 240000 260158 240009
rect 260102 239935 260158 239944
rect 260748 239420 260800 239426
rect 260748 239362 260800 239368
rect 260104 238060 260156 238066
rect 260104 238002 260156 238008
rect 259550 222184 259606 222193
rect 259550 222119 259606 222128
rect 259366 211032 259422 211041
rect 259366 210967 259422 210976
rect 260116 209681 260144 238002
rect 260760 229094 260788 239362
rect 260668 229066 260788 229094
rect 260668 221354 260696 229066
rect 260746 222184 260802 222193
rect 260746 222119 260802 222128
rect 260760 221474 260788 222119
rect 260748 221468 260800 221474
rect 260748 221410 260800 221416
rect 260668 221326 260788 221354
rect 260760 220794 260788 221326
rect 260748 220788 260800 220794
rect 260748 220730 260800 220736
rect 260760 220114 260788 220730
rect 260748 220108 260800 220114
rect 260748 220050 260800 220056
rect 260102 209672 260158 209681
rect 260102 209607 260158 209616
rect 258724 185700 258776 185706
rect 258724 185642 258776 185648
rect 260748 181484 260800 181490
rect 260748 181426 260800 181432
rect 258172 174548 258224 174554
rect 258172 174490 258224 174496
rect 258724 174004 258776 174010
rect 258724 173946 258776 173952
rect 257434 163160 257490 163169
rect 257434 163095 257490 163104
rect 257448 122806 257476 163095
rect 258736 149734 258764 173946
rect 259000 172644 259052 172650
rect 259000 172586 259052 172592
rect 258906 161936 258962 161945
rect 258906 161871 258962 161880
rect 258724 149728 258776 149734
rect 257526 149696 257582 149705
rect 258724 149670 258776 149676
rect 257526 149631 257582 149640
rect 257436 122800 257488 122806
rect 257436 122742 257488 122748
rect 257436 116068 257488 116074
rect 257436 116010 257488 116016
rect 257344 86964 257396 86970
rect 257344 86906 257396 86912
rect 257448 64161 257476 116010
rect 257540 109041 257568 149631
rect 258724 136672 258776 136678
rect 258724 136614 258776 136620
rect 257526 109032 257582 109041
rect 257526 108967 257582 108976
rect 257620 108316 257672 108322
rect 257620 108258 257672 108264
rect 257632 101425 257660 108258
rect 257618 101416 257674 101425
rect 257618 101351 257674 101360
rect 257528 99476 257580 99482
rect 257528 99418 257580 99424
rect 257540 77897 257568 99418
rect 257988 86964 258040 86970
rect 257988 86906 258040 86912
rect 257526 77888 257582 77897
rect 257526 77823 257582 77832
rect 257434 64152 257490 64161
rect 257434 64087 257490 64096
rect 256056 55888 256108 55894
rect 256056 55830 256108 55836
rect 254674 50280 254730 50289
rect 254674 50215 254730 50224
rect 253296 43512 253348 43518
rect 253296 43454 253348 43460
rect 251822 33824 251878 33833
rect 251822 33759 251878 33768
rect 250536 22772 250588 22778
rect 250536 22714 250588 22720
rect 250548 15201 250576 22714
rect 250534 15192 250590 15201
rect 250534 15127 250590 15136
rect 250548 13841 250576 15127
rect 250534 13832 250590 13841
rect 250534 13767 250590 13776
rect 251836 12442 251864 33759
rect 255962 25664 256018 25673
rect 255962 25599 256018 25608
rect 254582 24168 254638 24177
rect 254582 24103 254638 24112
rect 253478 15872 253534 15881
rect 253478 15807 253534 15816
rect 253492 15337 253520 15807
rect 254596 15337 254624 24103
rect 253478 15328 253534 15337
rect 253478 15263 253534 15272
rect 254582 15328 254638 15337
rect 254582 15263 254638 15272
rect 251824 12436 251876 12442
rect 251824 12378 251876 12384
rect 251836 11966 251864 12378
rect 251180 11960 251232 11966
rect 251180 11902 251232 11908
rect 251824 11960 251876 11966
rect 251824 11902 251876 11908
rect 250444 8968 250496 8974
rect 250444 8910 250496 8916
rect 251192 480 251220 11902
rect 253202 11792 253258 11801
rect 253202 11727 253258 11736
rect 253216 3534 253244 11727
rect 252376 3528 252428 3534
rect 252376 3470 252428 3476
rect 253204 3528 253256 3534
rect 253204 3470 253256 3476
rect 252388 480 252416 3470
rect 253492 480 253520 15263
rect 255976 15162 256004 25599
rect 257344 25560 257396 25566
rect 257344 25502 257396 25508
rect 255964 15156 256016 15162
rect 255964 15098 256016 15104
rect 256608 15156 256660 15162
rect 256608 15098 256660 15104
rect 254676 4140 254728 4146
rect 254676 4082 254728 4088
rect 254688 480 254716 4082
rect 256620 3505 256648 15098
rect 257356 4049 257384 25502
rect 257066 4040 257122 4049
rect 257066 3975 257122 3984
rect 257342 4040 257398 4049
rect 258000 4026 258028 86906
rect 258080 37256 258132 37262
rect 258080 37198 258132 37204
rect 258092 4146 258120 37198
rect 258736 14482 258764 136614
rect 258816 135380 258868 135386
rect 258816 135322 258868 135328
rect 258828 53106 258856 135322
rect 258920 121417 258948 161871
rect 259012 135250 259040 172586
rect 260102 170232 260158 170241
rect 260102 170167 260158 170176
rect 259000 135244 259052 135250
rect 259000 135186 259052 135192
rect 260116 131034 260144 170167
rect 260288 153264 260340 153270
rect 260288 153206 260340 153212
rect 260196 135312 260248 135318
rect 260196 135254 260248 135260
rect 260104 131028 260156 131034
rect 260104 130970 260156 130976
rect 258906 121408 258962 121417
rect 258906 121343 258962 121352
rect 259000 120148 259052 120154
rect 259000 120090 259052 120096
rect 258908 114640 258960 114646
rect 258908 114582 258960 114588
rect 258920 73817 258948 114582
rect 259012 105505 259040 120090
rect 259276 118720 259328 118726
rect 259276 118662 259328 118668
rect 259288 115161 259316 118662
rect 260102 117872 260158 117881
rect 260102 117807 260158 117816
rect 259274 115152 259330 115161
rect 259274 115087 259330 115096
rect 258998 105496 259054 105505
rect 258998 105431 259054 105440
rect 258906 73808 258962 73817
rect 258906 73743 258962 73752
rect 259458 53952 259514 53961
rect 259458 53887 259514 53896
rect 258816 53100 258868 53106
rect 258816 53042 258868 53048
rect 259368 40792 259420 40798
rect 259368 40734 259420 40740
rect 259380 37262 259408 40734
rect 259368 37256 259420 37262
rect 259368 37198 259420 37204
rect 258724 14476 258776 14482
rect 258724 14418 258776 14424
rect 258080 4140 258132 4146
rect 258080 4082 258132 4088
rect 258000 3998 258304 4026
rect 257342 3975 257398 3984
rect 255870 3496 255926 3505
rect 255870 3431 255926 3440
rect 256606 3496 256662 3505
rect 256606 3431 256662 3440
rect 255884 480 255912 3431
rect 257080 480 257108 3975
rect 258276 480 258304 3998
rect 259472 480 259500 53887
rect 260116 29646 260144 117807
rect 260208 69737 260236 135254
rect 260300 113150 260328 153206
rect 260288 113144 260340 113150
rect 260288 113086 260340 113092
rect 260288 104984 260340 104990
rect 260288 104926 260340 104932
rect 260194 69728 260250 69737
rect 260194 69663 260250 69672
rect 260300 58682 260328 104926
rect 260760 93770 260788 181426
rect 260852 152522 260880 283562
rect 260944 237289 260972 337350
rect 261024 331900 261076 331906
rect 261024 331842 261076 331848
rect 261036 252550 261064 331842
rect 262232 293185 262260 377590
rect 262864 374672 262916 374678
rect 262864 374614 262916 374620
rect 262312 314696 262364 314702
rect 262312 314638 262364 314644
rect 262218 293176 262274 293185
rect 262218 293111 262274 293120
rect 262220 272604 262272 272610
rect 262220 272546 262272 272552
rect 261024 252544 261076 252550
rect 261024 252486 261076 252492
rect 262128 252544 262180 252550
rect 262128 252486 262180 252492
rect 262140 251870 262168 252486
rect 262128 251864 262180 251870
rect 262128 251806 262180 251812
rect 260930 237280 260986 237289
rect 260930 237215 260986 237224
rect 260944 236706 260972 237215
rect 260932 236700 260984 236706
rect 260932 236642 260984 236648
rect 262232 180130 262260 272546
rect 262324 270502 262352 314638
rect 262404 294024 262456 294030
rect 262404 293966 262456 293972
rect 262312 270496 262364 270502
rect 262312 270438 262364 270444
rect 262310 266384 262366 266393
rect 262310 266319 262366 266328
rect 262324 226953 262352 266319
rect 262416 253910 262444 293966
rect 262680 270496 262732 270502
rect 262680 270438 262732 270444
rect 262692 269822 262720 270438
rect 262680 269816 262732 269822
rect 262680 269758 262732 269764
rect 262770 266248 262826 266257
rect 262770 266183 262826 266192
rect 262784 262886 262812 266183
rect 262772 262880 262824 262886
rect 262772 262822 262824 262828
rect 262404 253904 262456 253910
rect 262404 253846 262456 253852
rect 262680 253904 262732 253910
rect 262680 253846 262732 253852
rect 262692 253230 262720 253846
rect 262680 253224 262732 253230
rect 262680 253166 262732 253172
rect 262876 241369 262904 374614
rect 263600 355428 263652 355434
rect 263600 355370 263652 355376
rect 262956 292664 263008 292670
rect 262956 292606 263008 292612
rect 262968 273970 262996 292606
rect 262956 273964 263008 273970
rect 262956 273906 263008 273912
rect 262862 241360 262918 241369
rect 262862 241295 262918 241304
rect 262864 238128 262916 238134
rect 262864 238070 262916 238076
rect 262310 226944 262366 226953
rect 262310 226879 262366 226888
rect 262876 207738 262904 238070
rect 263612 212537 263640 355370
rect 263704 347721 263732 377590
rect 265070 349208 265126 349217
rect 265070 349143 265126 349152
rect 263690 347712 263746 347721
rect 263690 347647 263746 347656
rect 264242 347712 264298 347721
rect 264242 347647 264298 347656
rect 264256 346497 264284 347647
rect 264242 346488 264298 346497
rect 264242 346423 264298 346432
rect 263784 338768 263836 338774
rect 263784 338710 263836 338716
rect 263690 301064 263746 301073
rect 263690 300999 263746 301008
rect 263598 212528 263654 212537
rect 263598 212463 263654 212472
rect 263612 211886 263640 212463
rect 263600 211880 263652 211886
rect 263600 211822 263652 211828
rect 263704 209774 263732 300999
rect 263796 276010 263824 338710
rect 263784 276004 263836 276010
rect 263784 275946 263836 275952
rect 263796 275398 263824 275946
rect 263784 275392 263836 275398
rect 263784 275334 263836 275340
rect 264256 249150 264284 346423
rect 264980 319456 265032 319462
rect 264980 319398 265032 319404
rect 264334 269784 264390 269793
rect 264334 269719 264390 269728
rect 264348 268462 264376 269719
rect 264336 268456 264388 268462
rect 264336 268398 264388 268404
rect 264244 249144 264296 249150
rect 264244 249086 264296 249092
rect 263612 209746 263732 209774
rect 262864 207732 262916 207738
rect 262864 207674 262916 207680
rect 263612 204241 263640 209746
rect 263598 204232 263654 204241
rect 263598 204167 263654 204176
rect 263612 203561 263640 204167
rect 263598 203552 263654 203561
rect 263598 203487 263654 203496
rect 262220 180124 262272 180130
rect 262220 180066 262272 180072
rect 264348 180033 264376 268398
rect 264992 192545 265020 319398
rect 265084 267714 265112 349143
rect 265164 298784 265216 298790
rect 265164 298726 265216 298732
rect 265072 267708 265124 267714
rect 265072 267650 265124 267656
rect 265084 267034 265112 267650
rect 265072 267028 265124 267034
rect 265072 266970 265124 266976
rect 265176 262018 265204 298726
rect 266372 296177 266400 377590
rect 266452 330540 266504 330546
rect 266452 330482 266504 330488
rect 266464 328438 266492 330482
rect 266452 328432 266504 328438
rect 266452 328374 266504 328380
rect 267648 328432 267700 328438
rect 267648 328374 267700 328380
rect 267096 298172 267148 298178
rect 267096 298114 267148 298120
rect 266358 296168 266414 296177
rect 266358 296103 266414 296112
rect 267004 294160 267056 294166
rect 267004 294102 267056 294108
rect 266360 264920 266412 264926
rect 266360 264862 266412 264868
rect 266372 264246 266400 264862
rect 266360 264240 266412 264246
rect 266360 264182 266412 264188
rect 265084 261990 265204 262018
rect 265084 259418 265112 261990
rect 265624 261588 265676 261594
rect 265624 261530 265676 261536
rect 265072 259412 265124 259418
rect 265072 259354 265124 259360
rect 265084 258806 265112 259354
rect 265072 258800 265124 258806
rect 265072 258742 265124 258748
rect 265636 234054 265664 261530
rect 265624 234048 265676 234054
rect 265624 233990 265676 233996
rect 264978 192536 265034 192545
rect 264978 192471 265034 192480
rect 264334 180024 264390 180033
rect 264334 179959 264390 179968
rect 265636 178702 265664 233990
rect 267016 225622 267044 294102
rect 267108 285666 267136 298114
rect 267096 285660 267148 285666
rect 267096 285602 267148 285608
rect 267660 264246 267688 328374
rect 267648 264240 267700 264246
rect 267648 264182 267700 264188
rect 267004 225616 267056 225622
rect 267004 225558 267056 225564
rect 267016 193866 267044 225558
rect 267752 215286 267780 377590
rect 267832 369232 267884 369238
rect 267832 369174 267884 369180
rect 267740 215280 267792 215286
rect 267740 215222 267792 215228
rect 267844 209545 267872 369174
rect 269132 294166 269160 377590
rect 269762 351248 269818 351257
rect 269762 351183 269818 351192
rect 269212 313336 269264 313342
rect 269212 313278 269264 313284
rect 269120 294160 269172 294166
rect 269120 294102 269172 294108
rect 268384 292596 268436 292602
rect 268384 292538 268436 292544
rect 268396 276690 268424 292538
rect 268384 276684 268436 276690
rect 268384 276626 268436 276632
rect 268384 264308 268436 264314
rect 268384 264250 268436 264256
rect 268396 235958 268424 264250
rect 268384 235952 268436 235958
rect 268384 235894 268436 235900
rect 267830 209536 267886 209545
rect 267830 209471 267886 209480
rect 267844 209098 267872 209471
rect 267832 209092 267884 209098
rect 267832 209034 267884 209040
rect 267004 193860 267056 193866
rect 267004 193802 267056 193808
rect 268396 188358 268424 235894
rect 269028 215280 269080 215286
rect 269028 215222 269080 215228
rect 269040 214606 269068 215222
rect 269028 214600 269080 214606
rect 269028 214542 269080 214548
rect 268384 188352 268436 188358
rect 268384 188294 268436 188300
rect 269224 181490 269252 313278
rect 269776 219366 269804 351183
rect 270408 293276 270460 293282
rect 270408 293218 270460 293224
rect 269854 231296 269910 231305
rect 269854 231231 269910 231240
rect 269764 219360 269816 219366
rect 269764 219302 269816 219308
rect 269776 218822 269804 219302
rect 269764 218816 269816 218822
rect 269764 218758 269816 218764
rect 269212 181484 269264 181490
rect 269212 181426 269264 181432
rect 265624 178696 265676 178702
rect 265624 178638 265676 178644
rect 269868 176662 269896 231231
rect 270420 230518 270448 293218
rect 270512 233238 270540 377590
rect 272720 376825 272748 377590
rect 272706 376816 272762 376825
rect 272706 376751 272762 376760
rect 274744 374746 274772 377604
rect 276032 377590 276414 377618
rect 277412 377590 278070 377618
rect 274732 374740 274784 374746
rect 274732 374682 274784 374688
rect 271880 367124 271932 367130
rect 271880 367066 271932 367072
rect 270590 331800 270646 331809
rect 270590 331735 270646 331744
rect 270500 233232 270552 233238
rect 270500 233174 270552 233180
rect 270408 230512 270460 230518
rect 270408 230454 270460 230460
rect 270604 216617 270632 331735
rect 271142 284064 271198 284073
rect 271142 283999 271198 284008
rect 270590 216608 270646 216617
rect 270590 216543 270646 216552
rect 271156 183025 271184 283999
rect 271892 227633 271920 367066
rect 273904 354068 273956 354074
rect 273904 354010 273956 354016
rect 273258 313984 273314 313993
rect 273258 313919 273314 313928
rect 272522 302424 272578 302433
rect 272522 302359 272578 302368
rect 272536 256902 272564 302359
rect 273272 286385 273300 313919
rect 273258 286376 273314 286385
rect 273258 286311 273260 286320
rect 273312 286311 273314 286320
rect 273260 286282 273312 286288
rect 273272 286251 273300 286282
rect 272524 256896 272576 256902
rect 272524 256838 272576 256844
rect 273916 239426 273944 354010
rect 275284 327140 275336 327146
rect 275284 327082 275336 327088
rect 274086 309224 274142 309233
rect 274086 309159 274142 309168
rect 273994 285832 274050 285841
rect 273994 285767 274050 285776
rect 273904 239420 273956 239426
rect 273904 239362 273956 239368
rect 271878 227624 271934 227633
rect 271878 227559 271934 227568
rect 271892 226953 271920 227559
rect 271878 226944 271934 226953
rect 271878 226879 271934 226888
rect 271786 216608 271842 216617
rect 271786 216543 271842 216552
rect 271800 215937 271828 216543
rect 271786 215928 271842 215937
rect 271786 215863 271842 215872
rect 272616 207664 272668 207670
rect 272616 207606 272668 207612
rect 272524 203584 272576 203590
rect 272524 203526 272576 203532
rect 271142 183016 271198 183025
rect 271142 182951 271198 182960
rect 272062 182200 272118 182209
rect 272062 182135 272118 182144
rect 272076 181393 272104 182135
rect 272062 181384 272118 181393
rect 272062 181319 272118 181328
rect 272536 180130 272564 203526
rect 272628 195294 272656 207606
rect 272616 195288 272668 195294
rect 272616 195230 272668 195236
rect 272524 180124 272576 180130
rect 272524 180066 272576 180072
rect 274008 178673 274036 285767
rect 274100 225593 274128 309159
rect 274180 301504 274232 301510
rect 274180 301446 274232 301452
rect 274192 271182 274220 301446
rect 274180 271176 274232 271182
rect 274180 271118 274232 271124
rect 274086 225584 274142 225593
rect 274086 225519 274142 225528
rect 275296 186998 275324 327082
rect 275374 296984 275430 296993
rect 275374 296919 275430 296928
rect 275284 186992 275336 186998
rect 275284 186934 275336 186940
rect 275284 180872 275336 180878
rect 275284 180814 275336 180820
rect 275296 179382 275324 180814
rect 275284 179376 275336 179382
rect 275284 179318 275336 179324
rect 275388 178809 275416 296919
rect 276032 224942 276060 377590
rect 277412 320890 277440 377590
rect 279712 375358 279740 377604
rect 281382 377590 281488 377618
rect 283038 377590 283604 377618
rect 281460 376689 281488 377590
rect 281446 376680 281502 376689
rect 281446 376615 281502 376624
rect 278136 375352 278188 375358
rect 278136 375294 278188 375300
rect 279700 375352 279752 375358
rect 281460 375329 281488 376615
rect 279700 375294 279752 375300
rect 281446 375320 281502 375329
rect 277400 320884 277452 320890
rect 277400 320826 277452 320832
rect 276756 310548 276808 310554
rect 276756 310490 276808 310496
rect 276664 307828 276716 307834
rect 276664 307770 276716 307776
rect 276020 224936 276072 224942
rect 276020 224878 276072 224884
rect 276032 224262 276060 224878
rect 276020 224256 276072 224262
rect 276020 224198 276072 224204
rect 275374 178800 275430 178809
rect 275374 178735 275430 178744
rect 273994 178664 274050 178673
rect 273994 178599 274050 178608
rect 276676 178022 276704 307770
rect 276768 207641 276796 310490
rect 278042 305008 278098 305017
rect 278042 304943 278098 304952
rect 277398 280800 277454 280809
rect 277398 280735 277454 280744
rect 277412 273222 277440 280735
rect 276848 273216 276900 273222
rect 276848 273158 276900 273164
rect 277400 273216 277452 273222
rect 277400 273158 277452 273164
rect 276860 219473 276888 273158
rect 276940 220108 276992 220114
rect 276940 220050 276992 220056
rect 276846 219464 276902 219473
rect 276846 219399 276902 219408
rect 276754 207632 276810 207641
rect 276754 207567 276810 207576
rect 276756 193860 276808 193866
rect 276756 193802 276808 193808
rect 276768 178770 276796 193802
rect 276756 178764 276808 178770
rect 276756 178706 276808 178712
rect 276664 178016 276716 178022
rect 276664 177958 276716 177964
rect 269856 176656 269908 176662
rect 269856 176598 269908 176604
rect 276860 176594 276888 219399
rect 276952 192574 276980 220050
rect 276940 192568 276992 192574
rect 276940 192510 276992 192516
rect 278056 176769 278084 304943
rect 278148 293282 278176 375294
rect 281446 375255 281502 375264
rect 281460 374105 281488 375255
rect 279422 374096 279478 374105
rect 279422 374031 279478 374040
rect 281446 374096 281502 374105
rect 281446 374031 281502 374040
rect 278226 314800 278282 314809
rect 278226 314735 278282 314744
rect 278136 293276 278188 293282
rect 278136 293218 278188 293224
rect 278134 287736 278190 287745
rect 278134 287671 278190 287680
rect 278148 220114 278176 287671
rect 278240 250578 278268 314735
rect 279436 304201 279464 374031
rect 281460 363730 281488 374031
rect 283576 367169 283604 377590
rect 284312 377590 284694 377618
rect 285692 377590 286350 377618
rect 287072 377590 288006 377618
rect 288452 377590 289662 377618
rect 291212 377590 291318 377618
rect 292592 377590 292974 377618
rect 283378 367160 283434 367169
rect 283378 367095 283434 367104
rect 283562 367160 283618 367169
rect 283562 367095 283618 367104
rect 283392 366353 283420 367095
rect 283378 366344 283434 366353
rect 283378 366279 283434 366288
rect 281448 363724 281500 363730
rect 281448 363666 281500 363672
rect 282184 356720 282236 356726
rect 282184 356662 282236 356668
rect 280804 338768 280856 338774
rect 280804 338710 280856 338716
rect 279422 304192 279478 304201
rect 279422 304127 279478 304136
rect 279516 298240 279568 298246
rect 279516 298182 279568 298188
rect 278778 289096 278834 289105
rect 278778 289031 278834 289040
rect 278792 282878 278820 289031
rect 278780 282872 278832 282878
rect 278780 282814 278832 282820
rect 279424 282192 279476 282198
rect 279424 282134 279476 282140
rect 278228 250572 278280 250578
rect 278228 250514 278280 250520
rect 278136 220108 278188 220114
rect 278136 220050 278188 220056
rect 278136 207732 278188 207738
rect 278136 207674 278188 207680
rect 278148 180674 278176 207674
rect 279436 193905 279464 282134
rect 279528 274650 279556 298182
rect 280344 280832 280396 280838
rect 280344 280774 280396 280780
rect 280356 280265 280384 280774
rect 280342 280256 280398 280265
rect 280342 280191 280398 280200
rect 279516 274644 279568 274650
rect 279516 274586 279568 274592
rect 279516 256896 279568 256902
rect 279516 256838 279568 256844
rect 279422 193896 279478 193905
rect 279422 193831 279478 193840
rect 279424 185632 279476 185638
rect 279424 185574 279476 185580
rect 278688 180804 278740 180810
rect 278688 180746 278740 180752
rect 278700 180690 278728 180746
rect 278136 180668 278188 180674
rect 278700 180662 278820 180690
rect 278136 180610 278188 180616
rect 278792 177177 278820 180662
rect 279240 178764 279292 178770
rect 279240 178706 279292 178712
rect 278778 177168 278834 177177
rect 278778 177103 278834 177112
rect 278042 176760 278098 176769
rect 278042 176695 278098 176704
rect 276848 176588 276900 176594
rect 276848 176530 276900 176536
rect 264978 175672 265034 175681
rect 264978 175607 265034 175616
rect 264992 175302 265020 175607
rect 264980 175296 265032 175302
rect 264980 175238 265032 175244
rect 265070 175264 265126 175273
rect 265070 175199 265126 175208
rect 264978 174040 265034 174049
rect 265084 174010 265112 175199
rect 265714 174856 265770 174865
rect 265714 174791 265770 174800
rect 264978 173975 265034 173984
rect 265072 174004 265124 174010
rect 264992 173942 265020 173975
rect 265072 173946 265124 173952
rect 264980 173936 265032 173942
rect 264980 173878 265032 173884
rect 265070 173632 265126 173641
rect 265070 173567 265126 173576
rect 264978 172680 265034 172689
rect 265084 172650 265112 173567
rect 264978 172615 265034 172624
rect 265072 172644 265124 172650
rect 264992 172582 265020 172615
rect 265072 172586 265124 172592
rect 264980 172576 265032 172582
rect 264980 172518 265032 172524
rect 265070 172272 265126 172281
rect 265070 172207 265126 172216
rect 264978 171456 265034 171465
rect 264978 171391 265034 171400
rect 264992 171222 265020 171391
rect 264980 171216 265032 171222
rect 264980 171158 265032 171164
rect 265084 171154 265112 172207
rect 265072 171148 265124 171154
rect 265072 171090 265124 171096
rect 264978 171048 265034 171057
rect 264978 170983 265034 170992
rect 264242 170096 264298 170105
rect 264242 170031 264298 170040
rect 262862 166968 262918 166977
rect 262862 166903 262918 166912
rect 260840 152516 260892 152522
rect 260840 152458 260892 152464
rect 261668 140820 261720 140826
rect 261668 140762 261720 140768
rect 261576 127084 261628 127090
rect 261576 127026 261628 127032
rect 261482 119368 261538 119377
rect 261482 119303 261538 119312
rect 260748 93764 260800 93770
rect 260748 93706 260800 93712
rect 260760 93673 260788 93706
rect 260746 93664 260802 93673
rect 260746 93599 260802 93608
rect 260288 58676 260340 58682
rect 260288 58618 260340 58624
rect 260380 55888 260432 55894
rect 260380 55830 260432 55836
rect 260392 55185 260420 55830
rect 260378 55176 260434 55185
rect 260378 55111 260434 55120
rect 260392 53961 260420 55111
rect 260378 53952 260434 53961
rect 260378 53887 260434 53896
rect 260104 29640 260156 29646
rect 260104 29582 260156 29588
rect 260102 10296 260158 10305
rect 260102 10231 260158 10240
rect 260116 3641 260144 10231
rect 261496 7614 261524 119303
rect 261588 69601 261616 127026
rect 261680 98705 261708 140762
rect 262770 137592 262826 137601
rect 262770 137527 262826 137536
rect 262784 137193 262812 137527
rect 262770 137184 262826 137193
rect 262770 137119 262826 137128
rect 262678 136368 262734 136377
rect 262678 136303 262734 136312
rect 262692 135833 262720 136303
rect 262678 135824 262734 135833
rect 262678 135759 262734 135768
rect 262770 133240 262826 133249
rect 262770 133175 262826 133184
rect 262784 132841 262812 133175
rect 262770 132832 262826 132841
rect 262770 132767 262826 132776
rect 262876 126993 262904 166903
rect 263138 145616 263194 145625
rect 263138 145551 263194 145560
rect 262862 126984 262918 126993
rect 262862 126919 262918 126928
rect 263048 126948 263100 126954
rect 263048 126890 263100 126896
rect 262862 120728 262918 120737
rect 262862 120663 262918 120672
rect 262876 119406 262904 120663
rect 262954 120320 263010 120329
rect 262954 120255 263010 120264
rect 262864 119400 262916 119406
rect 262864 119342 262916 119348
rect 262968 113174 262996 120255
rect 262876 113146 262996 113174
rect 261760 100836 261812 100842
rect 261760 100778 261812 100784
rect 261666 98696 261722 98705
rect 261666 98631 261722 98640
rect 261772 86290 261800 100778
rect 261852 98048 261904 98054
rect 261852 97990 261904 97996
rect 261864 89049 261892 97990
rect 261850 89040 261906 89049
rect 261850 88975 261906 88984
rect 261760 86284 261812 86290
rect 261760 86226 261812 86232
rect 261574 69592 261630 69601
rect 261574 69527 261630 69536
rect 262876 46238 262904 113146
rect 262954 106448 263010 106457
rect 262954 106383 263010 106392
rect 262968 61402 262996 106383
rect 263060 99346 263088 126890
rect 263152 120873 263180 145551
rect 264256 131102 264284 170031
rect 264992 169794 265020 170983
rect 264980 169788 265032 169794
rect 264980 169730 265032 169736
rect 264978 169688 265034 169697
rect 264978 169623 265034 169632
rect 264992 168502 265020 169623
rect 265070 168872 265126 168881
rect 265070 168807 265126 168816
rect 264980 168496 265032 168502
rect 264980 168438 265032 168444
rect 265084 168434 265112 168807
rect 265072 168428 265124 168434
rect 265072 168370 265124 168376
rect 264978 167920 265034 167929
rect 264978 167855 265034 167864
rect 264992 167142 265020 167855
rect 265070 167512 265126 167521
rect 265070 167447 265126 167456
rect 264980 167136 265032 167142
rect 264980 167078 265032 167084
rect 265084 167074 265112 167447
rect 265072 167068 265124 167074
rect 265072 167010 265124 167016
rect 265728 166326 265756 174791
rect 279252 172258 279280 178706
rect 279332 178016 279384 178022
rect 279332 177958 279384 177964
rect 279344 173777 279372 177958
rect 279330 173768 279386 173777
rect 279330 173703 279386 173712
rect 279330 172272 279386 172281
rect 279252 172230 279330 172258
rect 279330 172207 279386 172216
rect 279436 169153 279464 185574
rect 279528 181490 279556 256838
rect 280816 238066 280844 338710
rect 282196 316713 282224 356662
rect 282276 323604 282328 323610
rect 282276 323546 282328 323552
rect 282182 316704 282238 316713
rect 282182 316639 282238 316648
rect 282182 291952 282238 291961
rect 282182 291887 282238 291896
rect 280896 289128 280948 289134
rect 280896 289070 280948 289076
rect 280908 262954 280936 289070
rect 281448 281512 281500 281518
rect 281448 281454 281500 281460
rect 281460 280838 281488 281454
rect 281448 280832 281500 280838
rect 281448 280774 281500 280780
rect 281448 276752 281500 276758
rect 281448 276694 281500 276700
rect 280896 262948 280948 262954
rect 280896 262890 280948 262896
rect 280804 238060 280856 238066
rect 280804 238002 280856 238008
rect 280804 233300 280856 233306
rect 280804 233242 280856 233248
rect 279608 196648 279660 196654
rect 279608 196590 279660 196596
rect 279516 181484 279568 181490
rect 279516 181426 279568 181432
rect 279516 177336 279568 177342
rect 279516 177278 279568 177284
rect 279422 169144 279478 169153
rect 279422 169079 279478 169088
rect 279528 166841 279556 177278
rect 279620 175982 279648 196590
rect 280250 187232 280306 187241
rect 280250 187167 280306 187176
rect 279884 176656 279936 176662
rect 279884 176598 279936 176604
rect 279896 176089 279924 176598
rect 280068 176588 280120 176594
rect 280068 176530 280120 176536
rect 280080 176497 280108 176530
rect 280066 176488 280122 176497
rect 280066 176423 280122 176432
rect 279882 176080 279938 176089
rect 279882 176015 279938 176024
rect 279608 175976 279660 175982
rect 279608 175918 279660 175924
rect 280160 175976 280212 175982
rect 280160 175918 280212 175924
rect 279606 175808 279662 175817
rect 279606 175743 279662 175752
rect 279620 174321 279648 175743
rect 279606 174312 279662 174321
rect 279606 174247 279662 174256
rect 280172 171134 280200 175918
rect 279712 171106 280200 171134
rect 279514 166832 279570 166841
rect 279514 166767 279570 166776
rect 265716 166320 265768 166326
rect 264978 166288 265034 166297
rect 265716 166262 265768 166268
rect 264978 166223 265034 166232
rect 264992 165646 265020 166223
rect 265622 165880 265678 165889
rect 265622 165815 265678 165824
rect 264980 165640 265032 165646
rect 264980 165582 265032 165588
rect 265070 165336 265126 165345
rect 265070 165271 265126 165280
rect 264978 164928 265034 164937
rect 264978 164863 265034 164872
rect 264992 164354 265020 164863
rect 264980 164348 265032 164354
rect 264980 164290 265032 164296
rect 265084 164286 265112 165271
rect 265072 164280 265124 164286
rect 265072 164222 265124 164228
rect 265254 164112 265310 164121
rect 265254 164047 265310 164056
rect 265070 163704 265126 163713
rect 265070 163639 265126 163648
rect 265084 162994 265112 163639
rect 265072 162988 265124 162994
rect 265072 162930 265124 162936
rect 264980 162920 265032 162926
rect 264978 162888 264980 162897
rect 265032 162888 265034 162897
rect 264978 162823 265034 162832
rect 265070 162344 265126 162353
rect 265070 162279 265126 162288
rect 264980 161560 265032 161566
rect 264978 161528 264980 161537
rect 265032 161528 265034 161537
rect 265084 161498 265112 162279
rect 264978 161463 265034 161472
rect 265072 161492 265124 161498
rect 265072 161434 265124 161440
rect 265070 161120 265126 161129
rect 265070 161055 265126 161064
rect 264978 160712 265034 160721
rect 264978 160647 265034 160656
rect 264992 160206 265020 160647
rect 264980 160200 265032 160206
rect 264980 160142 265032 160148
rect 265084 160138 265112 161055
rect 265072 160132 265124 160138
rect 265072 160074 265124 160080
rect 265070 159760 265126 159769
rect 265070 159695 265126 159704
rect 264978 158944 265034 158953
rect 264978 158879 265034 158888
rect 264992 158778 265020 158879
rect 265084 158846 265112 159695
rect 265072 158840 265124 158846
rect 265072 158782 265124 158788
rect 264980 158772 265032 158778
rect 264980 158714 265032 158720
rect 265070 158536 265126 158545
rect 265070 158471 265126 158480
rect 264978 157720 265034 157729
rect 264978 157655 265034 157664
rect 264992 157486 265020 157655
rect 264980 157480 265032 157486
rect 264980 157422 265032 157428
rect 265084 157418 265112 158471
rect 265072 157412 265124 157418
rect 265072 157354 265124 157360
rect 265070 156768 265126 156777
rect 265070 156703 265126 156712
rect 264978 156360 265034 156369
rect 264978 156295 265034 156304
rect 264992 156058 265020 156295
rect 264980 156052 265032 156058
rect 264980 155994 265032 156000
rect 265084 155990 265112 156703
rect 265072 155984 265124 155990
rect 265072 155926 265124 155932
rect 265162 155952 265218 155961
rect 265162 155887 265218 155896
rect 265176 154630 265204 155887
rect 265268 155242 265296 164047
rect 265256 155236 265308 155242
rect 265256 155178 265308 155184
rect 265164 154624 265216 154630
rect 264978 154592 265034 154601
rect 265164 154566 265216 154572
rect 264978 154527 265034 154536
rect 264992 153882 265020 154527
rect 264980 153876 265032 153882
rect 264980 153818 265032 153824
rect 264978 153776 265034 153785
rect 264978 153711 265034 153720
rect 264992 153270 265020 153711
rect 264980 153264 265032 153270
rect 264980 153206 265032 153212
rect 264978 152960 265034 152969
rect 264978 152895 265034 152904
rect 264334 152552 264390 152561
rect 264334 152487 264390 152496
rect 264348 140078 264376 152487
rect 264992 151842 265020 152895
rect 264980 151836 265032 151842
rect 264980 151778 265032 151784
rect 264978 151192 265034 151201
rect 264978 151127 265034 151136
rect 264992 150482 265020 151127
rect 265070 150784 265126 150793
rect 265070 150719 265126 150728
rect 264980 150476 265032 150482
rect 264980 150418 265032 150424
rect 264978 149968 265034 149977
rect 264978 149903 265034 149912
rect 264992 149122 265020 149903
rect 265084 149705 265112 150719
rect 265070 149696 265126 149705
rect 265070 149631 265126 149640
rect 265162 149560 265218 149569
rect 265162 149495 265218 149504
rect 264980 149116 265032 149122
rect 264980 149058 265032 149064
rect 265070 149016 265126 149025
rect 265070 148951 265126 148960
rect 264978 147792 265034 147801
rect 264978 147727 264980 147736
rect 265032 147727 265034 147736
rect 264980 147698 265032 147704
rect 265084 147694 265112 148951
rect 265072 147688 265124 147694
rect 265072 147630 265124 147636
rect 265070 147384 265126 147393
rect 265070 147319 265126 147328
rect 264978 146432 265034 146441
rect 264978 146367 264980 146376
rect 265032 146367 265034 146376
rect 264980 146338 265032 146344
rect 265084 146334 265112 147319
rect 265072 146328 265124 146334
rect 265072 146270 265124 146276
rect 265070 146024 265126 146033
rect 265070 145959 265126 145968
rect 264978 145208 265034 145217
rect 264978 145143 265034 145152
rect 264992 144974 265020 145143
rect 265084 145042 265112 145959
rect 265176 145761 265204 149495
rect 265162 145752 265218 145761
rect 265162 145687 265218 145696
rect 265072 145036 265124 145042
rect 265072 144978 265124 144984
rect 264980 144968 265032 144974
rect 264980 144910 265032 144916
rect 265070 144800 265126 144809
rect 265070 144735 265126 144744
rect 264978 144392 265034 144401
rect 264978 144327 265034 144336
rect 264992 143682 265020 144327
rect 264980 143676 265032 143682
rect 264980 143618 265032 143624
rect 265084 143614 265112 144735
rect 265162 143848 265218 143857
rect 265162 143783 265218 143792
rect 265072 143608 265124 143614
rect 265072 143550 265124 143556
rect 264610 142624 264666 142633
rect 264610 142559 264666 142568
rect 264336 140072 264388 140078
rect 264336 140014 264388 140020
rect 264334 139224 264390 139233
rect 264334 139159 264390 139168
rect 264244 131096 264296 131102
rect 264244 131038 264296 131044
rect 263138 120864 263194 120873
rect 263138 120799 263194 120808
rect 263140 111920 263192 111926
rect 263140 111862 263192 111868
rect 263048 99340 263100 99346
rect 263048 99282 263100 99288
rect 263152 90370 263180 111862
rect 264242 108760 264298 108769
rect 264242 108695 264298 108704
rect 263140 90364 263192 90370
rect 263140 90306 263192 90312
rect 262956 61396 263008 61402
rect 262956 61338 263008 61344
rect 262954 57216 263010 57225
rect 262954 57151 263010 57160
rect 262864 46232 262916 46238
rect 262864 46174 262916 46180
rect 262968 27606 262996 57151
rect 262220 27600 262272 27606
rect 262220 27542 262272 27548
rect 262956 27600 263008 27606
rect 262956 27542 263008 27548
rect 262232 16574 262260 27542
rect 263600 26920 263652 26926
rect 263600 26862 263652 26868
rect 263612 16574 263640 26862
rect 264256 21418 264284 108695
rect 264348 108322 264376 139159
rect 264624 132494 264652 142559
rect 264978 142216 265034 142225
rect 264978 142151 264980 142160
rect 265032 142151 265034 142160
rect 264980 142122 265032 142128
rect 265176 141409 265204 143783
rect 265636 142866 265664 165815
rect 279712 161474 279740 171106
rect 280264 164937 280292 187167
rect 280816 184210 280844 233242
rect 280804 184204 280856 184210
rect 280804 184146 280856 184152
rect 280436 182912 280488 182918
rect 280436 182854 280488 182860
rect 280344 180668 280396 180674
rect 280344 180610 280396 180616
rect 280250 164928 280306 164937
rect 280250 164863 280306 164872
rect 279068 161446 279740 161474
rect 265806 157176 265862 157185
rect 265806 157111 265862 157120
rect 265820 151162 265848 157111
rect 265990 154184 266046 154193
rect 265990 154119 266046 154128
rect 265808 151156 265860 151162
rect 265808 151098 265860 151104
rect 265714 148608 265770 148617
rect 265714 148543 265770 148552
rect 265624 142860 265676 142866
rect 265624 142802 265676 142808
rect 265162 141400 265218 141409
rect 265162 141335 265218 141344
rect 264978 140856 265034 140865
rect 264978 140791 264980 140800
rect 265032 140791 265034 140800
rect 264980 140762 265032 140768
rect 264978 140040 265034 140049
rect 264978 139975 265034 139984
rect 264992 139466 265020 139975
rect 264980 139460 265032 139466
rect 264980 139402 265032 139408
rect 264978 138680 265034 138689
rect 264978 138615 265034 138624
rect 264992 138038 265020 138615
rect 264980 138032 265032 138038
rect 264980 137974 265032 137980
rect 264978 137048 265034 137057
rect 264978 136983 265034 136992
rect 264992 136678 265020 136983
rect 264980 136672 265032 136678
rect 264980 136614 265032 136620
rect 264978 136232 265034 136241
rect 264978 136167 265034 136176
rect 264992 135318 265020 136167
rect 265070 135688 265126 135697
rect 265070 135623 265126 135632
rect 265084 135386 265112 135623
rect 265072 135380 265124 135386
rect 265072 135322 265124 135328
rect 264980 135312 265032 135318
rect 264980 135254 265032 135260
rect 264978 132696 265034 132705
rect 264978 132631 265034 132640
rect 264992 132530 265020 132631
rect 264532 132466 264652 132494
rect 264980 132524 265032 132530
rect 264980 132466 265032 132472
rect 264426 108624 264482 108633
rect 264426 108559 264482 108568
rect 264336 108316 264388 108322
rect 264336 108258 264388 108264
rect 264334 105224 264390 105233
rect 264334 105159 264390 105168
rect 264348 42090 264376 105159
rect 264440 57254 264468 108559
rect 264532 102785 264560 132466
rect 265070 131880 265126 131889
rect 265070 131815 265126 131824
rect 264978 131472 265034 131481
rect 264978 131407 265034 131416
rect 264992 131238 265020 131407
rect 264980 131232 265032 131238
rect 264980 131174 265032 131180
rect 265084 131170 265112 131815
rect 265072 131164 265124 131170
rect 265072 131106 265124 131112
rect 264978 129704 265034 129713
rect 264978 129639 265034 129648
rect 264992 128450 265020 129639
rect 265622 128480 265678 128489
rect 264980 128444 265032 128450
rect 265622 128415 265678 128424
rect 264980 128386 265032 128392
rect 264612 128376 264664 128382
rect 264612 128318 264664 128324
rect 264624 107642 264652 128318
rect 264978 127936 265034 127945
rect 264978 127871 265034 127880
rect 264992 127022 265020 127871
rect 265070 127120 265126 127129
rect 265070 127055 265072 127064
rect 265124 127055 265126 127064
rect 265072 127026 265124 127032
rect 264980 127016 265032 127022
rect 264980 126958 265032 126964
rect 264978 126304 265034 126313
rect 264978 126239 265034 126248
rect 264992 125662 265020 126239
rect 264980 125656 265032 125662
rect 264980 125598 265032 125604
rect 265070 125352 265126 125361
rect 265070 125287 265126 125296
rect 264978 124536 265034 124545
rect 264978 124471 265034 124480
rect 264992 124302 265020 124471
rect 264980 124296 265032 124302
rect 264980 124238 265032 124244
rect 265084 124234 265112 125287
rect 265072 124228 265124 124234
rect 265072 124170 265124 124176
rect 264978 124128 265034 124137
rect 264978 124063 265034 124072
rect 264992 122874 265020 124063
rect 265070 123720 265126 123729
rect 265070 123655 265126 123664
rect 264980 122868 265032 122874
rect 264980 122810 265032 122816
rect 265084 122126 265112 123655
rect 265072 122120 265124 122126
rect 265072 122062 265124 122068
rect 264978 121952 265034 121961
rect 264978 121887 265034 121896
rect 264992 120766 265020 121887
rect 265070 121136 265126 121145
rect 265070 121071 265126 121080
rect 264980 120760 265032 120766
rect 264980 120702 265032 120708
rect 265084 120154 265112 121071
rect 265072 120148 265124 120154
rect 265072 120090 265124 120096
rect 264978 119776 265034 119785
rect 264978 119711 265034 119720
rect 264992 118726 265020 119711
rect 264980 118720 265032 118726
rect 264980 118662 265032 118668
rect 264978 118552 265034 118561
rect 264978 118487 265034 118496
rect 264992 117366 265020 118487
rect 264980 117360 265032 117366
rect 264980 117302 265032 117308
rect 265070 117192 265126 117201
rect 265070 117127 265126 117136
rect 264978 116376 265034 116385
rect 264978 116311 265034 116320
rect 264992 116074 265020 116311
rect 264980 116068 265032 116074
rect 264980 116010 265032 116016
rect 265084 116006 265112 117127
rect 265072 116000 265124 116006
rect 265072 115942 265124 115948
rect 265070 115560 265126 115569
rect 265070 115495 265126 115504
rect 264978 115152 265034 115161
rect 264978 115087 265034 115096
rect 264992 114578 265020 115087
rect 265084 114646 265112 115495
rect 265072 114640 265124 114646
rect 265072 114582 265124 114588
rect 264980 114572 265032 114578
rect 264980 114514 265032 114520
rect 264978 113792 265034 113801
rect 264978 113727 265034 113736
rect 264992 113218 265020 113727
rect 264980 113212 265032 113218
rect 264980 113154 265032 113160
rect 265254 112568 265310 112577
rect 265254 112503 265310 112512
rect 264978 112024 265034 112033
rect 264978 111959 265034 111968
rect 264992 111858 265020 111959
rect 265268 111926 265296 112503
rect 265256 111920 265308 111926
rect 265256 111862 265308 111868
rect 264980 111852 265032 111858
rect 264980 111794 265032 111800
rect 265070 111616 265126 111625
rect 265070 111551 265126 111560
rect 264978 111208 265034 111217
rect 264978 111143 265034 111152
rect 264992 110498 265020 111143
rect 265084 110566 265112 111551
rect 265072 110560 265124 110566
rect 265072 110502 265124 110508
rect 264980 110492 265032 110498
rect 264980 110434 265032 110440
rect 265070 109984 265126 109993
rect 265070 109919 265126 109928
rect 264978 109576 265034 109585
rect 264978 109511 265034 109520
rect 264992 109138 265020 109511
rect 264980 109132 265032 109138
rect 264980 109074 265032 109080
rect 265084 109070 265112 109919
rect 265072 109064 265124 109070
rect 265072 109006 265124 109012
rect 264612 107636 264664 107642
rect 264612 107578 264664 107584
rect 264978 106992 265034 107001
rect 264978 106927 265034 106936
rect 264992 106350 265020 106927
rect 264980 106344 265032 106350
rect 264980 106286 265032 106292
rect 264978 106040 265034 106049
rect 264978 105975 265034 105984
rect 264992 104922 265020 105975
rect 265070 105632 265126 105641
rect 265070 105567 265126 105576
rect 265084 104990 265112 105567
rect 265072 104984 265124 104990
rect 265072 104926 265124 104932
rect 264980 104916 265032 104922
rect 264980 104858 265032 104864
rect 264978 103864 265034 103873
rect 264978 103799 265034 103808
rect 264992 103562 265020 103799
rect 264980 103556 265032 103562
rect 264980 103498 265032 103504
rect 264978 103456 265034 103465
rect 264978 103391 265034 103400
rect 264518 102776 264574 102785
rect 264518 102711 264574 102720
rect 264886 102640 264942 102649
rect 264886 102575 264942 102584
rect 264900 94625 264928 102575
rect 264992 102202 265020 103391
rect 264980 102196 265032 102202
rect 264980 102138 265032 102144
rect 264978 101824 265034 101833
rect 264978 101759 265034 101768
rect 264992 100774 265020 101759
rect 265070 101280 265126 101289
rect 265070 101215 265126 101224
rect 265084 100842 265112 101215
rect 265072 100836 265124 100842
rect 265072 100778 265124 100784
rect 264980 100768 265032 100774
rect 264980 100710 265032 100716
rect 265070 100056 265126 100065
rect 265070 99991 265126 100000
rect 264978 99648 265034 99657
rect 264978 99583 265034 99592
rect 264992 99414 265020 99583
rect 265084 99482 265112 99991
rect 265072 99476 265124 99482
rect 265072 99418 265124 99424
rect 264980 99408 265032 99414
rect 264980 99350 265032 99356
rect 264978 98696 265034 98705
rect 264978 98631 265034 98640
rect 264992 98054 265020 98631
rect 264980 98048 265032 98054
rect 264980 97990 265032 97996
rect 265070 97880 265126 97889
rect 265070 97815 265126 97824
rect 264980 97300 265032 97306
rect 264980 97242 265032 97248
rect 264992 97073 265020 97242
rect 264978 97064 265034 97073
rect 264978 96999 265034 97008
rect 265084 96694 265112 97815
rect 265072 96688 265124 96694
rect 265072 96630 265124 96636
rect 264886 94616 264942 94625
rect 264886 94551 264942 94560
rect 264428 57248 264480 57254
rect 264428 57190 264480 57196
rect 265636 43450 265664 128415
rect 265728 128382 265756 148543
rect 265806 143440 265862 143449
rect 265806 143375 265862 143384
rect 265716 128376 265768 128382
rect 265716 128318 265768 128324
rect 265714 125896 265770 125905
rect 265714 125831 265770 125840
rect 265728 66881 265756 125831
rect 265820 117978 265848 143375
rect 265898 141808 265954 141817
rect 265898 141743 265954 141752
rect 265912 123457 265940 141743
rect 266004 141506 266032 154119
rect 279068 151814 279096 161446
rect 280356 161129 280384 180610
rect 280342 161120 280398 161129
rect 280342 161055 280398 161064
rect 280068 157412 280120 157418
rect 280068 157354 280120 157360
rect 279068 151786 279372 151814
rect 279344 144809 279372 151786
rect 279330 144800 279386 144809
rect 279330 144735 279386 144744
rect 280080 142154 280108 157354
rect 279160 142126 280108 142154
rect 265992 141500 266044 141506
rect 265992 141442 266044 141448
rect 266082 141264 266138 141273
rect 266082 141199 266138 141208
rect 266096 126954 266124 141199
rect 267002 134464 267058 134473
rect 267002 134399 267058 134408
rect 266084 126948 266136 126954
rect 266084 126890 266136 126896
rect 265898 123448 265954 123457
rect 265898 123383 265954 123392
rect 265808 117972 265860 117978
rect 265808 117914 265860 117920
rect 266266 109032 266322 109041
rect 266266 108967 266322 108976
rect 265806 98288 265862 98297
rect 265806 98223 265862 98232
rect 265820 79393 265848 98223
rect 266280 93838 266308 108967
rect 266268 93832 266320 93838
rect 266268 93774 266320 93780
rect 265806 79384 265862 79393
rect 265806 79319 265862 79328
rect 265714 66872 265770 66881
rect 265714 66807 265770 66816
rect 267016 58585 267044 134399
rect 279160 133362 279188 142126
rect 279330 133376 279386 133385
rect 279160 133334 279330 133362
rect 279330 133311 279386 133320
rect 267094 122904 267150 122913
rect 267094 122839 267150 122848
rect 267108 68241 267136 122839
rect 280158 121408 280214 121417
rect 280158 121343 280214 121352
rect 279330 120184 279386 120193
rect 279330 120119 279386 120128
rect 267646 115968 267702 115977
rect 267646 115903 267702 115912
rect 267186 100464 267242 100473
rect 267186 100399 267242 100408
rect 267200 72593 267228 100399
rect 267660 95470 267688 115903
rect 279344 113174 279372 120119
rect 279068 113146 279372 113174
rect 267738 110392 267794 110401
rect 267738 110327 267794 110336
rect 267648 95464 267700 95470
rect 267648 95406 267700 95412
rect 267186 72584 267242 72593
rect 267186 72519 267242 72528
rect 267094 68232 267150 68241
rect 267094 68167 267150 68176
rect 267002 58576 267058 58585
rect 267002 58511 267058 58520
rect 267752 51746 267780 110327
rect 267830 95568 267886 95577
rect 267830 95503 267886 95512
rect 267844 88330 267872 95503
rect 269212 95464 269264 95470
rect 269212 95406 269264 95412
rect 267832 88324 267884 88330
rect 267832 88266 267884 88272
rect 269120 60308 269172 60314
rect 269120 60250 269172 60256
rect 267740 51740 267792 51746
rect 267740 51682 267792 51688
rect 265624 43444 265676 43450
rect 265624 43386 265676 43392
rect 264336 42084 264388 42090
rect 264336 42026 264388 42032
rect 268384 42084 268436 42090
rect 268384 42026 268436 42032
rect 264244 21412 264296 21418
rect 264244 21354 264296 21360
rect 268396 19281 268424 42026
rect 267738 19272 267794 19281
rect 267738 19207 267794 19216
rect 268382 19272 268438 19281
rect 268382 19207 268438 19216
rect 262232 16546 262536 16574
rect 263612 16546 264192 16574
rect 261758 11656 261814 11665
rect 261758 11591 261814 11600
rect 261772 9654 261800 11591
rect 261760 9648 261812 9654
rect 261760 9590 261812 9596
rect 261484 7608 261536 7614
rect 261484 7550 261536 7556
rect 260102 3632 260158 3641
rect 260102 3567 260158 3576
rect 260654 3632 260710 3641
rect 260654 3567 260710 3576
rect 260668 480 260696 3567
rect 261772 480 261800 9590
rect 262508 490 262536 16546
rect 262784 598 262996 626
rect 262784 490 262812 598
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262508 462 262812 490
rect 262968 480 262996 598
rect 264164 480 264192 16546
rect 264980 12504 265032 12510
rect 264980 12446 265032 12452
rect 264992 490 265020 12446
rect 266360 3528 266412 3534
rect 266360 3470 266412 3476
rect 266544 3528 266596 3534
rect 266544 3470 266596 3476
rect 266372 3369 266400 3470
rect 266358 3360 266414 3369
rect 266358 3295 266414 3304
rect 265176 598 265388 626
rect 265176 490 265204 598
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 264992 462 265204 490
rect 265360 480 265388 598
rect 266556 480 266584 3470
rect 267752 3466 267780 19207
rect 269132 16574 269160 60250
rect 269224 40730 269252 95406
rect 270498 94616 270554 94625
rect 270498 94551 270554 94560
rect 270512 78674 270540 94551
rect 271878 94480 271934 94489
rect 271878 94415 271934 94424
rect 270500 78668 270552 78674
rect 270500 78610 270552 78616
rect 271052 78668 271104 78674
rect 271052 78610 271104 78616
rect 271064 78062 271092 78610
rect 271052 78056 271104 78062
rect 271052 77998 271104 78004
rect 271892 60722 271920 94415
rect 274008 93770 274036 96084
rect 275928 94512 275980 94518
rect 275928 94454 275980 94460
rect 273996 93764 274048 93770
rect 273996 93706 274048 93712
rect 273904 93152 273956 93158
rect 273904 93094 273956 93100
rect 271880 60716 271932 60722
rect 271880 60658 271932 60664
rect 271892 60314 271920 60658
rect 271880 60308 271932 60314
rect 271880 60250 271932 60256
rect 271144 58676 271196 58682
rect 271144 58618 271196 58624
rect 269212 40724 269264 40730
rect 269212 40666 269264 40672
rect 270500 20664 270552 20670
rect 270500 20606 270552 20612
rect 270512 16574 270540 20606
rect 269132 16546 270080 16574
rect 270512 16546 270816 16574
rect 267740 3460 267792 3466
rect 267740 3402 267792 3408
rect 268844 3460 268896 3466
rect 268844 3402 268896 3408
rect 267740 3324 267792 3330
rect 267740 3266 267792 3272
rect 267752 480 267780 3266
rect 268856 480 268884 3402
rect 270052 480 270080 16546
rect 270788 490 270816 16546
rect 271156 3534 271184 58618
rect 273916 30297 273944 93094
rect 275940 92313 275968 94454
rect 275926 92304 275982 92313
rect 275926 92239 275982 92248
rect 275940 91202 275968 92239
rect 275940 91174 276060 91202
rect 273994 62792 274050 62801
rect 273994 62727 274050 62736
rect 273258 30288 273314 30297
rect 273258 30223 273314 30232
rect 273902 30288 273958 30297
rect 273902 30223 273958 30232
rect 271788 28280 271840 28286
rect 271788 28222 271840 28228
rect 271800 20670 271828 28222
rect 271788 20664 271840 20670
rect 271788 20606 271840 20612
rect 271144 3528 271196 3534
rect 271144 3470 271196 3476
rect 272432 2984 272484 2990
rect 272432 2926 272484 2932
rect 271064 598 271276 626
rect 271064 490 271092 598
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 270788 462 271092 490
rect 271248 480 271276 598
rect 272444 480 272472 2926
rect 273272 490 273300 30223
rect 274008 2990 274036 62727
rect 275284 32428 275336 32434
rect 275284 32370 275336 32376
rect 275296 31822 275324 32370
rect 275284 31816 275336 31822
rect 275284 31758 275336 31764
rect 275296 3534 275324 31758
rect 276032 3602 276060 91174
rect 279068 89690 279096 113146
rect 279330 104272 279386 104281
rect 279330 104207 279386 104216
rect 279344 93838 279372 104207
rect 279332 93832 279384 93838
rect 279332 93774 279384 93780
rect 279056 89684 279108 89690
rect 279056 89626 279108 89632
rect 278042 86184 278098 86193
rect 278042 86119 278098 86128
rect 276664 36576 276716 36582
rect 276664 36518 276716 36524
rect 276676 31822 276704 36518
rect 276664 31816 276716 31822
rect 276664 31758 276716 31764
rect 278056 31074 278084 86119
rect 280172 85542 280200 121343
rect 280448 119241 280476 182854
rect 281460 172961 281488 276694
rect 281540 245744 281592 245750
rect 281540 245686 281592 245692
rect 281446 172952 281502 172961
rect 281446 172887 281502 172896
rect 281552 157418 281580 245686
rect 282196 232558 282224 291887
rect 282288 276690 282316 323546
rect 282366 306640 282422 306649
rect 282366 306575 282422 306584
rect 282380 283626 282408 306575
rect 283194 299704 283250 299713
rect 283194 299639 283250 299648
rect 282368 283620 282420 283626
rect 282368 283562 282420 283568
rect 282276 276684 282328 276690
rect 282276 276626 282328 276632
rect 282276 271856 282328 271862
rect 282276 271798 282328 271804
rect 282288 270609 282316 271798
rect 282274 270600 282330 270609
rect 282274 270535 282330 270544
rect 282184 232552 282236 232558
rect 282184 232494 282236 232500
rect 282184 230512 282236 230518
rect 282184 230454 282236 230460
rect 281632 193928 281684 193934
rect 281632 193870 281684 193876
rect 281540 157412 281592 157418
rect 281540 157354 281592 157360
rect 281644 129033 281672 193870
rect 281724 185700 281776 185706
rect 281724 185642 281776 185648
rect 281736 151881 281764 185642
rect 282196 179790 282224 230454
rect 282184 179784 282236 179790
rect 282184 179726 282236 179732
rect 282918 179480 282974 179489
rect 282918 179415 282974 179424
rect 281814 175536 281870 175545
rect 281814 175471 281870 175480
rect 281828 175302 281856 175471
rect 281816 175296 281868 175302
rect 281816 175238 281868 175244
rect 282828 175160 282880 175166
rect 282828 175102 282880 175108
rect 282840 174729 282868 175102
rect 282826 174720 282882 174729
rect 282826 174655 282882 174664
rect 282734 174312 282790 174321
rect 282734 174247 282790 174256
rect 282748 173890 282776 174247
rect 282826 174040 282882 174049
rect 282932 174026 282960 179415
rect 283012 178696 283064 178702
rect 283012 178638 283064 178644
rect 282882 173998 282960 174026
rect 282826 173975 282882 173984
rect 282748 173862 282960 173890
rect 281816 171012 281868 171018
rect 281816 170954 281868 170960
rect 281828 170921 281856 170954
rect 281814 170912 281870 170921
rect 281814 170847 281870 170856
rect 282828 169720 282880 169726
rect 282828 169662 282880 169668
rect 282840 169425 282868 169662
rect 282826 169416 282882 169425
rect 282826 169351 282882 169360
rect 282736 168360 282788 168366
rect 282736 168302 282788 168308
rect 282748 167113 282776 168302
rect 282828 168020 282880 168026
rect 282828 167962 282880 167968
rect 282840 167929 282868 167962
rect 282826 167920 282882 167929
rect 282826 167855 282882 167864
rect 282734 167104 282790 167113
rect 282734 167039 282790 167048
rect 282826 165608 282882 165617
rect 282826 165543 282882 165552
rect 282840 165238 282868 165543
rect 282828 165232 282880 165238
rect 282828 165174 282880 165180
rect 282184 164212 282236 164218
rect 282184 164154 282236 164160
rect 281816 164144 281868 164150
rect 281814 164112 281816 164121
rect 281868 164112 281870 164121
rect 281814 164047 281870 164056
rect 282196 163305 282224 164154
rect 282182 163296 282238 163305
rect 282182 163231 282238 163240
rect 282276 162784 282328 162790
rect 282276 162726 282328 162732
rect 282288 161809 282316 162726
rect 282826 162616 282882 162625
rect 282932 162602 282960 173862
rect 282882 162574 282960 162602
rect 282826 162551 282882 162560
rect 282274 161800 282330 161809
rect 282274 161735 282330 161744
rect 282644 161424 282696 161430
rect 282644 161366 282696 161372
rect 282656 160313 282684 161366
rect 282642 160304 282698 160313
rect 282642 160239 282698 160248
rect 282828 160064 282880 160070
rect 282828 160006 282880 160012
rect 282736 159996 282788 160002
rect 282736 159938 282788 159944
rect 282748 158817 282776 159938
rect 282840 159497 282868 160006
rect 282826 159488 282882 159497
rect 282826 159423 282882 159432
rect 282734 158808 282790 158817
rect 282734 158743 282790 158752
rect 282092 158704 282144 158710
rect 282092 158646 282144 158652
rect 282104 158001 282132 158646
rect 282184 158024 282236 158030
rect 282090 157992 282146 158001
rect 282184 157966 282236 157972
rect 282090 157927 282146 157936
rect 281722 151872 281778 151881
rect 281722 151807 281778 151816
rect 281908 150408 281960 150414
rect 281908 150350 281960 150356
rect 281920 149705 281948 150350
rect 281906 149696 281962 149705
rect 281906 149631 281962 149640
rect 281724 138984 281776 138990
rect 281722 138952 281724 138961
rect 281776 138952 281778 138961
rect 281722 138887 281778 138896
rect 282196 136649 282224 157966
rect 282828 156664 282880 156670
rect 282828 156606 282880 156612
rect 282552 155712 282604 155718
rect 282550 155680 282552 155689
rect 282604 155680 282606 155689
rect 282550 155615 282606 155624
rect 282368 154556 282420 154562
rect 282368 154498 282420 154504
rect 282380 153513 282408 154498
rect 282840 154193 282868 156606
rect 282826 154184 282882 154193
rect 282826 154119 282882 154128
rect 282736 153876 282788 153882
rect 282736 153818 282788 153824
rect 282366 153504 282422 153513
rect 282366 153439 282422 153448
rect 282748 151201 282776 153818
rect 282828 153196 282880 153202
rect 282828 153138 282880 153144
rect 282840 152697 282868 153138
rect 282826 152688 282882 152697
rect 282826 152623 282882 152632
rect 282734 151192 282790 151201
rect 282734 151127 282790 151136
rect 282736 151088 282788 151094
rect 282736 151030 282788 151036
rect 282748 148889 282776 151030
rect 282826 150376 282882 150385
rect 282826 150311 282828 150320
rect 282880 150311 282882 150320
rect 282828 150282 282880 150288
rect 282828 149048 282880 149054
rect 282828 148990 282880 148996
rect 282734 148880 282790 148889
rect 282734 148815 282790 148824
rect 282840 148073 282868 148990
rect 282826 148064 282882 148073
rect 282826 147999 282882 148008
rect 282736 147620 282788 147626
rect 282736 147562 282788 147568
rect 282748 146577 282776 147562
rect 282828 147552 282880 147558
rect 282828 147494 282880 147500
rect 282840 147393 282868 147494
rect 282826 147384 282882 147393
rect 282826 147319 282882 147328
rect 282734 146568 282790 146577
rect 282734 146503 282790 146512
rect 282552 146260 282604 146266
rect 282552 146202 282604 146208
rect 282564 145081 282592 146202
rect 282828 146192 282880 146198
rect 282828 146134 282880 146140
rect 282840 145897 282868 146134
rect 282826 145888 282882 145897
rect 282826 145823 282882 145832
rect 282550 145072 282606 145081
rect 282550 145007 282606 145016
rect 282460 144900 282512 144906
rect 282460 144842 282512 144848
rect 282472 143585 282500 144842
rect 282458 143576 282514 143585
rect 282458 143511 282514 143520
rect 282826 142760 282882 142769
rect 282826 142695 282882 142704
rect 282840 142458 282868 142695
rect 282828 142452 282880 142458
rect 282828 142394 282880 142400
rect 282828 142112 282880 142118
rect 282826 142080 282828 142089
rect 282880 142080 282882 142089
rect 282736 142044 282788 142050
rect 282826 142015 282882 142024
rect 282736 141986 282788 141992
rect 282748 141273 282776 141986
rect 282734 141264 282790 141273
rect 282734 141199 282790 141208
rect 282828 140752 282880 140758
rect 282828 140694 282880 140700
rect 282840 140457 282868 140694
rect 282826 140448 282882 140457
rect 282826 140383 282882 140392
rect 282644 139392 282696 139398
rect 282644 139334 282696 139340
rect 282656 138281 282684 139334
rect 282642 138272 282698 138281
rect 282642 138207 282698 138216
rect 282828 137964 282880 137970
rect 282828 137906 282880 137912
rect 282840 137465 282868 137906
rect 282826 137456 282882 137465
rect 282826 137391 282882 137400
rect 282182 136640 282238 136649
rect 282182 136575 282238 136584
rect 282828 136604 282880 136610
rect 282828 136546 282880 136552
rect 282840 135969 282868 136546
rect 282826 135960 282882 135969
rect 282276 135924 282328 135930
rect 282826 135895 282882 135904
rect 282276 135866 282328 135872
rect 282288 132494 282316 135866
rect 282828 135244 282880 135250
rect 282828 135186 282880 135192
rect 282840 135153 282868 135186
rect 282826 135144 282882 135153
rect 282826 135079 282882 135088
rect 282460 134972 282512 134978
rect 282460 134914 282512 134920
rect 282472 134473 282500 134914
rect 282458 134464 282514 134473
rect 282458 134399 282514 134408
rect 283024 132494 283052 178638
rect 283208 171018 283236 299639
rect 283564 291848 283616 291854
rect 283564 291790 283616 291796
rect 283576 245750 283604 291790
rect 283564 245744 283616 245750
rect 283564 245686 283616 245692
rect 283564 211880 283616 211886
rect 283564 211822 283616 211828
rect 283576 180033 283604 211822
rect 284312 200025 284340 377590
rect 285586 367160 285642 367169
rect 285586 367095 285642 367104
rect 284944 299532 284996 299538
rect 284944 299474 284996 299480
rect 284484 225684 284536 225690
rect 284484 225626 284536 225632
rect 284496 225010 284524 225626
rect 284484 225004 284536 225010
rect 284484 224946 284536 224952
rect 284392 204944 284444 204950
rect 284392 204886 284444 204892
rect 284298 200016 284354 200025
rect 284298 199951 284354 199960
rect 284312 199481 284340 199951
rect 284298 199472 284354 199481
rect 284298 199407 284354 199416
rect 283562 180024 283618 180033
rect 283562 179959 283618 179968
rect 283196 171012 283248 171018
rect 283196 170954 283248 170960
rect 283564 156732 283616 156738
rect 283564 156674 283616 156680
rect 282196 132466 282316 132494
rect 282932 132466 283052 132494
rect 281630 129024 281686 129033
rect 281630 128959 281686 128968
rect 281538 126848 281594 126857
rect 281538 126783 281594 126792
rect 280434 119232 280490 119241
rect 280434 119167 280490 119176
rect 280160 85536 280212 85542
rect 280160 85478 280212 85484
rect 281552 81394 281580 126783
rect 282092 126268 282144 126274
rect 282092 126210 282144 126216
rect 281632 125588 281684 125594
rect 281632 125530 281684 125536
rect 281644 124545 281672 125530
rect 281630 124536 281686 124545
rect 281630 124471 281686 124480
rect 282104 123729 282132 126210
rect 282196 125225 282224 132466
rect 282828 132456 282880 132462
rect 282828 132398 282880 132404
rect 282840 131345 282868 132398
rect 282826 131336 282882 131345
rect 282826 131271 282882 131280
rect 282276 131096 282328 131102
rect 282276 131038 282328 131044
rect 282288 130665 282316 131038
rect 282644 131028 282696 131034
rect 282644 130970 282696 130976
rect 282274 130656 282330 130665
rect 282274 130591 282330 130600
rect 282656 129849 282684 130970
rect 282642 129840 282698 129849
rect 282642 129775 282698 129784
rect 282826 128344 282882 128353
rect 282826 128279 282882 128288
rect 282840 128246 282868 128279
rect 282828 128240 282880 128246
rect 282828 128182 282880 128188
rect 282826 127528 282882 127537
rect 282932 127514 282960 132466
rect 282882 127486 282960 127514
rect 282826 127463 282882 127472
rect 282828 126948 282880 126954
rect 282828 126890 282880 126896
rect 282840 126041 282868 126890
rect 282826 126032 282882 126041
rect 282826 125967 282882 125976
rect 282182 125216 282238 125225
rect 282182 125151 282238 125160
rect 282644 124160 282696 124166
rect 282644 124102 282696 124108
rect 282090 123720 282146 123729
rect 282090 123655 282146 123664
rect 282656 123049 282684 124102
rect 282642 123040 282698 123049
rect 282642 122975 282698 122984
rect 282826 122224 282882 122233
rect 282826 122159 282882 122168
rect 282840 121650 282868 122159
rect 282828 121644 282880 121650
rect 282828 121586 282880 121592
rect 282828 120080 282880 120086
rect 282828 120022 282880 120028
rect 282840 119921 282868 120022
rect 282826 119912 282882 119921
rect 282826 119847 282882 119856
rect 282184 119400 282236 119406
rect 282184 119342 282236 119348
rect 281724 115932 281776 115938
rect 281724 115874 281776 115880
rect 281736 115433 281764 115874
rect 281722 115424 281778 115433
rect 281722 115359 281778 115368
rect 282196 108497 282224 119342
rect 282828 118652 282880 118658
rect 282828 118594 282880 118600
rect 282840 118425 282868 118594
rect 282826 118416 282882 118425
rect 282826 118351 282882 118360
rect 282828 118108 282880 118114
rect 282828 118050 282880 118056
rect 282840 117609 282868 118050
rect 282826 117600 282882 117609
rect 282826 117535 282882 117544
rect 282828 117292 282880 117298
rect 282828 117234 282880 117240
rect 282840 116929 282868 117234
rect 282826 116920 282882 116929
rect 282826 116855 282882 116864
rect 282276 116748 282328 116754
rect 282276 116690 282328 116696
rect 282288 116113 282316 116690
rect 282274 116104 282330 116113
rect 282274 116039 282330 116048
rect 282460 115864 282512 115870
rect 282460 115806 282512 115812
rect 282472 114617 282500 115806
rect 282458 114608 282514 114617
rect 282458 114543 282514 114552
rect 282276 114164 282328 114170
rect 282276 114106 282328 114112
rect 282288 113801 282316 114106
rect 282274 113792 282330 113801
rect 282274 113727 282330 113736
rect 282828 113144 282880 113150
rect 282826 113112 282828 113121
rect 282880 113112 282882 113121
rect 282826 113047 282882 113056
rect 282828 112668 282880 112674
rect 282828 112610 282880 112616
rect 282840 112305 282868 112610
rect 282826 112296 282882 112305
rect 282826 112231 282882 112240
rect 282276 111784 282328 111790
rect 282276 111726 282328 111732
rect 282288 110809 282316 111726
rect 282274 110800 282330 110809
rect 282274 110735 282330 110744
rect 282828 110424 282880 110430
rect 282828 110366 282880 110372
rect 282840 109313 282868 110366
rect 282826 109304 282882 109313
rect 282826 109239 282882 109248
rect 282368 108996 282420 109002
rect 282368 108938 282420 108944
rect 282182 108488 282238 108497
rect 282182 108423 282238 108432
rect 282380 107817 282408 108938
rect 282366 107808 282422 107817
rect 282366 107743 282422 107752
rect 281630 106992 281686 107001
rect 281630 106927 281686 106936
rect 281644 91089 281672 106927
rect 281814 106176 281870 106185
rect 281814 106111 281870 106120
rect 281724 103216 281776 103222
rect 281722 103184 281724 103193
rect 281776 103184 281778 103193
rect 281722 103119 281778 103128
rect 281722 100872 281778 100881
rect 281722 100807 281778 100816
rect 281736 95198 281764 100807
rect 281724 95192 281776 95198
rect 281724 95134 281776 95140
rect 281828 92478 281856 106111
rect 281908 104848 281960 104854
rect 281908 104790 281960 104796
rect 281920 104009 281948 104790
rect 281906 104000 281962 104009
rect 281906 103935 281962 103944
rect 282828 103488 282880 103494
rect 282828 103430 282880 103436
rect 282840 102377 282868 103430
rect 283576 103222 283604 156674
rect 284404 104854 284432 204886
rect 284496 164150 284524 224946
rect 284956 178022 284984 299474
rect 285600 207641 285628 367095
rect 285692 225010 285720 377590
rect 287072 367577 287100 377590
rect 287058 367568 287114 367577
rect 287058 367503 287114 367512
rect 287058 327176 287114 327185
rect 287058 327111 287114 327120
rect 285772 320884 285824 320890
rect 285772 320826 285824 320832
rect 286968 320884 287020 320890
rect 286968 320826 287020 320832
rect 285784 320210 285812 320826
rect 285772 320204 285824 320210
rect 285772 320146 285824 320152
rect 285680 225004 285732 225010
rect 285680 224946 285732 224952
rect 285680 224256 285732 224262
rect 285680 224198 285732 224204
rect 285586 207632 285642 207641
rect 285586 207567 285642 207576
rect 285034 192672 285090 192681
rect 285034 192607 285090 192616
rect 285048 178702 285076 192607
rect 285036 178696 285088 178702
rect 285036 178638 285088 178644
rect 284944 178016 284996 178022
rect 284944 177958 284996 177964
rect 284574 176488 284630 176497
rect 284574 176423 284630 176432
rect 284484 164144 284536 164150
rect 284484 164086 284536 164092
rect 284588 138990 284616 176423
rect 284576 138984 284628 138990
rect 284576 138926 284628 138932
rect 285692 114170 285720 224198
rect 285864 196716 285916 196722
rect 285864 196658 285916 196664
rect 285772 188352 285824 188358
rect 285772 188294 285824 188300
rect 285784 116754 285812 188294
rect 285876 134978 285904 196658
rect 286980 193866 287008 320826
rect 286968 193860 287020 193866
rect 286968 193802 287020 193808
rect 285956 179784 286008 179790
rect 285956 179726 286008 179732
rect 285968 155718 285996 179726
rect 287072 165238 287100 327111
rect 287704 287700 287756 287706
rect 287704 287642 287756 287648
rect 287152 259480 287204 259486
rect 287152 259422 287204 259428
rect 287060 165232 287112 165238
rect 287060 165174 287112 165180
rect 285956 155712 286008 155718
rect 285956 155654 286008 155660
rect 285864 134972 285916 134978
rect 285864 134914 285916 134920
rect 285772 116748 285824 116754
rect 285772 116690 285824 116696
rect 285680 114164 285732 114170
rect 285680 114106 285732 114112
rect 287164 112674 287192 259422
rect 287716 237386 287744 287642
rect 288348 260160 288400 260166
rect 288348 260102 288400 260108
rect 288360 259486 288388 260102
rect 288348 259480 288400 259486
rect 288348 259422 288400 259428
rect 287704 237380 287756 237386
rect 287704 237322 287756 237328
rect 287244 214600 287296 214606
rect 287244 214542 287296 214548
rect 287256 118114 287284 214542
rect 288452 194449 288480 377590
rect 289728 342916 289780 342922
rect 289728 342858 289780 342864
rect 289740 322833 289768 342858
rect 289726 322824 289782 322833
rect 289726 322759 289782 322768
rect 289740 322250 289768 322759
rect 289728 322244 289780 322250
rect 289728 322186 289780 322192
rect 289820 306400 289872 306406
rect 289820 306342 289872 306348
rect 288530 289912 288586 289921
rect 288530 289847 288586 289856
rect 288438 194440 288494 194449
rect 288438 194375 288494 194384
rect 287336 181484 287388 181490
rect 287336 181426 287388 181432
rect 287348 142458 287376 181426
rect 288440 178016 288492 178022
rect 288440 177958 288492 177964
rect 288452 168026 288480 177958
rect 288440 168020 288492 168026
rect 288440 167962 288492 167968
rect 287336 142452 287388 142458
rect 287336 142394 287388 142400
rect 288544 120086 288572 289847
rect 288624 258732 288676 258738
rect 288624 258674 288676 258680
rect 288636 258126 288664 258674
rect 288624 258120 288676 258126
rect 288624 258062 288676 258068
rect 288636 158710 288664 258062
rect 288714 202192 288770 202201
rect 288714 202127 288770 202136
rect 288728 201550 288756 202127
rect 288716 201544 288768 201550
rect 288714 201512 288716 201521
rect 288768 201512 288770 201521
rect 288714 201447 288770 201456
rect 288714 178800 288770 178809
rect 288714 178735 288770 178744
rect 288624 158704 288676 158710
rect 288624 158646 288676 158652
rect 288728 121650 288756 178735
rect 289832 140758 289860 306342
rect 291212 298761 291240 377590
rect 291842 341592 291898 341601
rect 291842 341527 291898 341536
rect 291198 298752 291254 298761
rect 291198 298687 291254 298696
rect 291292 289128 291344 289134
rect 291292 289070 291344 289076
rect 291304 288561 291332 289070
rect 291290 288552 291346 288561
rect 291290 288487 291346 288496
rect 291200 269816 291252 269822
rect 291200 269758 291252 269764
rect 289912 240236 289964 240242
rect 289912 240178 289964 240184
rect 289924 153882 289952 240178
rect 290096 191140 290148 191146
rect 290096 191082 290148 191088
rect 290002 177440 290058 177449
rect 290002 177375 290058 177384
rect 289912 153876 289964 153882
rect 289912 153818 289964 153824
rect 289820 140752 289872 140758
rect 289820 140694 289872 140700
rect 288716 121644 288768 121650
rect 288716 121586 288768 121592
rect 288532 120080 288584 120086
rect 288532 120022 288584 120028
rect 287244 118108 287296 118114
rect 287244 118050 287296 118056
rect 290016 117298 290044 177375
rect 290108 168366 290136 191082
rect 290096 168360 290148 168366
rect 290096 168302 290148 168308
rect 291212 126954 291240 269758
rect 291304 153785 291332 288487
rect 291382 178664 291438 178673
rect 291382 178599 291438 178608
rect 291290 153776 291346 153785
rect 291290 153711 291346 153720
rect 291200 126948 291252 126954
rect 291200 126890 291252 126896
rect 290004 117292 290056 117298
rect 290004 117234 290056 117240
rect 291108 117292 291160 117298
rect 291108 117234 291160 117240
rect 291120 117201 291148 117234
rect 291106 117192 291162 117201
rect 291106 117127 291162 117136
rect 287152 112668 287204 112674
rect 287152 112610 287204 112616
rect 284392 104848 284444 104854
rect 284392 104790 284444 104796
rect 283564 103216 283616 103222
rect 283564 103158 283616 103164
rect 282826 102368 282882 102377
rect 282826 102303 282882 102312
rect 282826 99376 282882 99385
rect 282000 99340 282052 99346
rect 282826 99311 282882 99320
rect 282000 99282 282052 99288
rect 282012 98569 282040 99282
rect 282840 99278 282868 99311
rect 282828 99272 282880 99278
rect 282828 99214 282880 99220
rect 281998 98560 282054 98569
rect 281998 98495 282054 98504
rect 282828 97980 282880 97986
rect 282828 97922 282880 97928
rect 282736 97912 282788 97918
rect 282840 97889 282868 97922
rect 291396 97918 291424 178599
rect 291384 97912 291436 97918
rect 282736 97854 282788 97860
rect 282826 97880 282882 97889
rect 282748 97073 282776 97854
rect 291384 97854 291436 97860
rect 282826 97815 282882 97824
rect 282734 97064 282790 97073
rect 282734 96999 282790 97008
rect 282828 96620 282880 96626
rect 282828 96562 282880 96568
rect 282840 96393 282868 96562
rect 282826 96384 282882 96393
rect 282826 96319 282882 96328
rect 281816 92472 281868 92478
rect 281816 92414 281868 92420
rect 281630 91080 281686 91089
rect 281630 91015 281686 91024
rect 281630 90400 281686 90409
rect 281630 90335 281686 90344
rect 281540 81388 281592 81394
rect 281540 81330 281592 81336
rect 278688 75200 278740 75206
rect 278688 75142 278740 75148
rect 278044 31068 278096 31074
rect 278044 31010 278096 31016
rect 277400 29640 277452 29646
rect 277400 29582 277452 29588
rect 276112 12436 276164 12442
rect 276112 12378 276164 12384
rect 276020 3596 276072 3602
rect 276020 3538 276072 3544
rect 274824 3528 274876 3534
rect 274824 3470 274876 3476
rect 275284 3528 275336 3534
rect 276124 3482 276152 12378
rect 277412 6914 277440 29582
rect 277490 22672 277546 22681
rect 277490 22607 277546 22616
rect 277504 12442 277532 22607
rect 277492 12436 277544 12442
rect 277492 12378 277544 12384
rect 277412 6886 278360 6914
rect 277124 3596 277176 3602
rect 277124 3538 277176 3544
rect 275284 3470 275336 3476
rect 273996 2984 274048 2990
rect 273996 2926 274048 2932
rect 273456 598 273668 626
rect 273456 490 273484 598
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273272 462 273484 490
rect 273640 480 273668 598
rect 274836 480 274864 3470
rect 276032 3454 276152 3482
rect 276032 480 276060 3454
rect 277136 480 277164 3538
rect 278332 480 278360 6886
rect 278700 4214 278728 75142
rect 280804 47592 280856 47598
rect 280804 47534 280856 47540
rect 279424 43444 279476 43450
rect 279424 43386 279476 43392
rect 279436 31754 279464 43386
rect 278780 31748 278832 31754
rect 278780 31690 278832 31696
rect 279424 31748 279476 31754
rect 279424 31690 279476 31696
rect 278792 16574 278820 31690
rect 280816 19310 280844 47534
rect 280896 33856 280948 33862
rect 280896 33798 280948 33804
rect 280804 19304 280856 19310
rect 280804 19246 280856 19252
rect 280908 17950 280936 33798
rect 281540 31068 281592 31074
rect 281540 31010 281592 31016
rect 280896 17944 280948 17950
rect 280896 17886 280948 17892
rect 280908 17338 280936 17886
rect 280160 17332 280212 17338
rect 280160 17274 280212 17280
rect 280896 17332 280948 17338
rect 280896 17274 280948 17280
rect 280172 16574 280200 17274
rect 278792 16546 279096 16574
rect 280172 16546 280752 16574
rect 278688 4208 278740 4214
rect 278688 4150 278740 4156
rect 278700 2689 278728 4150
rect 278686 2680 278742 2689
rect 278686 2615 278742 2624
rect 279068 490 279096 16546
rect 279344 598 279556 626
rect 279344 490 279372 598
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279068 462 279372 490
rect 279528 480 279556 598
rect 280724 480 280752 16546
rect 281552 490 281580 31010
rect 281644 3330 281672 90335
rect 289084 69692 289136 69698
rect 289084 69634 289136 69640
rect 288348 61396 288400 61402
rect 288348 61338 288400 61344
rect 288360 60489 288388 61338
rect 288346 60480 288402 60489
rect 288346 60415 288402 60424
rect 285680 47592 285732 47598
rect 285680 47534 285732 47540
rect 284944 21412 284996 21418
rect 284944 21354 284996 21360
rect 284956 20641 284984 21354
rect 284390 20632 284446 20641
rect 284390 20567 284446 20576
rect 284942 20632 284998 20641
rect 284942 20567 284998 20576
rect 284404 6914 284432 20567
rect 284944 19304 284996 19310
rect 284944 19246 284996 19252
rect 284956 18698 284984 19246
rect 284944 18692 284996 18698
rect 284944 18634 284996 18640
rect 284956 16574 284984 18634
rect 285692 16574 285720 47534
rect 284956 16546 285076 16574
rect 285692 16546 286640 16574
rect 284404 6886 284984 6914
rect 283104 4208 283156 4214
rect 283104 4150 283156 4156
rect 281632 3324 281684 3330
rect 281632 3266 281684 3272
rect 281736 598 281948 626
rect 281736 490 281764 598
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281552 462 281764 490
rect 281920 480 281948 598
rect 283116 480 283144 4150
rect 284300 3528 284352 3534
rect 284300 3470 284352 3476
rect 284312 480 284340 3470
rect 284956 490 284984 6886
rect 285048 3534 285076 16546
rect 285036 3528 285088 3534
rect 285036 3470 285088 3476
rect 285232 598 285444 626
rect 285232 490 285260 598
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 284956 462 285260 490
rect 285416 480 285444 598
rect 286612 480 286640 16546
rect 288360 5681 288388 60415
rect 288440 18624 288492 18630
rect 288440 18566 288492 18572
rect 288452 11014 288480 18566
rect 288440 11008 288492 11014
rect 288440 10950 288492 10956
rect 288992 11008 289044 11014
rect 288992 10950 289044 10956
rect 287794 5672 287850 5681
rect 287794 5607 287850 5616
rect 288346 5672 288402 5681
rect 288346 5607 288402 5616
rect 287808 480 287836 5607
rect 289004 480 289032 10950
rect 289096 6769 289124 69634
rect 289082 6760 289138 6769
rect 289082 6695 289138 6704
rect 289096 4078 289124 6695
rect 291856 4146 291884 341527
rect 292592 310282 292620 377590
rect 294616 374678 294644 377604
rect 296272 374746 296300 377604
rect 295248 374740 295300 374746
rect 295248 374682 295300 374688
rect 296260 374740 296312 374746
rect 296260 374682 296312 374688
rect 294604 374672 294656 374678
rect 294604 374614 294656 374620
rect 292580 310276 292632 310282
rect 292580 310218 292632 310224
rect 293224 310276 293276 310282
rect 293224 310218 293276 310224
rect 292592 309806 292620 310218
rect 292580 309800 292632 309806
rect 292580 309742 292632 309748
rect 293236 280838 293264 310218
rect 293224 280832 293276 280838
rect 293224 280774 293276 280780
rect 293960 271176 294012 271182
rect 293960 271118 294012 271124
rect 292580 258800 292632 258806
rect 292580 258742 292632 258748
rect 292488 225616 292540 225622
rect 292488 225558 292540 225564
rect 292500 213897 292528 225558
rect 292486 213888 292542 213897
rect 292486 213823 292542 213832
rect 292592 149054 292620 258742
rect 293222 213888 293278 213897
rect 293222 213823 293278 213832
rect 292672 195288 292724 195294
rect 292672 195230 292724 195236
rect 292580 149048 292632 149054
rect 292580 148990 292632 148996
rect 292684 136610 292712 195230
rect 292764 180124 292816 180130
rect 292764 180066 292816 180072
rect 292776 147558 292804 180066
rect 292764 147552 292816 147558
rect 292764 147494 292816 147500
rect 292672 136604 292724 136610
rect 292672 136546 292724 136552
rect 293236 99385 293264 213823
rect 293972 111790 294000 271118
rect 295260 238377 295288 374682
rect 297928 374066 297956 377604
rect 299492 377590 299598 377618
rect 298836 375352 298888 375358
rect 298836 375294 298888 375300
rect 295984 374060 296036 374066
rect 295984 374002 296036 374008
rect 297916 374060 297968 374066
rect 297916 374002 297968 374008
rect 295996 354074 296024 374002
rect 295984 354068 296036 354074
rect 295984 354010 296036 354016
rect 297362 331256 297418 331265
rect 297362 331191 297418 331200
rect 298006 331256 298062 331265
rect 298006 331191 298008 331200
rect 295340 294636 295392 294642
rect 295340 294578 295392 294584
rect 295352 294545 295380 294578
rect 295338 294536 295394 294545
rect 295338 294471 295394 294480
rect 295246 238368 295302 238377
rect 295246 238303 295302 238312
rect 295260 238066 295288 238303
rect 295248 238060 295300 238066
rect 295248 238002 295300 238008
rect 294052 220108 294104 220114
rect 294052 220050 294104 220056
rect 293960 111784 294012 111790
rect 293960 111726 294012 111732
rect 292670 99376 292726 99385
rect 292670 99311 292726 99320
rect 293222 99376 293278 99385
rect 293222 99311 293278 99320
rect 292684 16574 292712 99311
rect 294064 99278 294092 220050
rect 294144 193860 294196 193866
rect 294144 193802 294196 193808
rect 294156 146198 294184 193802
rect 294234 180024 294290 180033
rect 294234 179959 294290 179968
rect 294248 156738 294276 179959
rect 294236 156732 294288 156738
rect 294236 156674 294288 156680
rect 294144 146192 294196 146198
rect 294144 146134 294196 146140
rect 295352 115870 295380 294471
rect 297376 281518 297404 331191
rect 298060 331191 298062 331200
rect 298008 331162 298060 331168
rect 298744 307080 298796 307086
rect 298744 307022 298796 307028
rect 298756 282878 298784 307022
rect 298100 282872 298152 282878
rect 298100 282814 298152 282820
rect 298744 282872 298796 282878
rect 298744 282814 298796 282820
rect 297364 281512 297416 281518
rect 297364 281454 297416 281460
rect 296720 276684 296772 276690
rect 296720 276626 296772 276632
rect 295432 257372 295484 257378
rect 295432 257314 295484 257320
rect 295444 142050 295472 257314
rect 295524 198008 295576 198014
rect 295524 197950 295576 197956
rect 295536 169726 295564 197950
rect 295982 184376 296038 184385
rect 295982 184311 296038 184320
rect 295524 169720 295576 169726
rect 295524 169662 295576 169668
rect 295432 142044 295484 142050
rect 295432 141986 295484 141992
rect 295340 115864 295392 115870
rect 295340 115806 295392 115812
rect 294052 99272 294104 99278
rect 294052 99214 294104 99220
rect 295338 33144 295394 33153
rect 295338 33079 295394 33088
rect 295352 16574 295380 33079
rect 292684 16546 293264 16574
rect 295352 16546 295656 16574
rect 291844 4140 291896 4146
rect 291844 4082 291896 4088
rect 289084 4072 289136 4078
rect 289084 4014 289136 4020
rect 291856 3738 291884 4082
rect 292580 4072 292632 4078
rect 292580 4014 292632 4020
rect 291384 3732 291436 3738
rect 291384 3674 291436 3680
rect 291844 3732 291896 3738
rect 291844 3674 291896 3680
rect 290186 3496 290242 3505
rect 290186 3431 290242 3440
rect 290200 480 290228 3431
rect 291396 480 291424 3674
rect 292592 480 292620 4014
rect 293236 490 293264 16546
rect 295340 13796 295392 13802
rect 295340 13738 295392 13744
rect 295352 12510 295380 13738
rect 295340 12504 295392 12510
rect 295340 12446 295392 12452
rect 294878 3496 294934 3505
rect 294878 3431 294934 3440
rect 293512 598 293724 626
rect 293512 490 293540 598
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293236 462 293540 490
rect 293696 480 293724 598
rect 294892 480 294920 3431
rect 295628 490 295656 16546
rect 295892 13796 295944 13802
rect 295892 13738 295944 13744
rect 295904 13705 295932 13738
rect 295890 13696 295946 13705
rect 295890 13631 295946 13640
rect 295996 3913 296024 184311
rect 296074 44840 296130 44849
rect 296074 44775 296130 44784
rect 296088 33153 296116 44775
rect 296074 33144 296130 33153
rect 296074 33079 296130 33088
rect 296732 27606 296760 276626
rect 297362 231976 297418 231985
rect 297362 231911 297418 231920
rect 296902 196752 296958 196761
rect 296902 196687 296958 196696
rect 296812 186992 296864 186998
rect 296812 186934 296864 186940
rect 296824 99346 296852 186934
rect 296916 160002 296944 196687
rect 296904 159996 296956 160002
rect 296904 159938 296956 159944
rect 297376 152522 297404 231911
rect 297364 152516 297416 152522
rect 297364 152458 297416 152464
rect 298112 110430 298140 282814
rect 298744 264240 298796 264246
rect 298744 264182 298796 264188
rect 298284 227044 298336 227050
rect 298284 226986 298336 226992
rect 298192 192568 298244 192574
rect 298192 192510 298244 192516
rect 298204 118658 298232 192510
rect 298296 153202 298324 226986
rect 298284 153196 298336 153202
rect 298284 153138 298336 153144
rect 298192 118652 298244 118658
rect 298192 118594 298244 118600
rect 298100 110424 298152 110430
rect 298100 110366 298152 110372
rect 298756 101425 298784 264182
rect 298848 240242 298876 375294
rect 299388 249076 299440 249082
rect 299388 249018 299440 249024
rect 299400 248402 299428 249018
rect 299388 248396 299440 248402
rect 299388 248338 299440 248344
rect 298836 240236 298888 240242
rect 298836 240178 298888 240184
rect 299492 208185 299520 377590
rect 301240 375358 301268 377604
rect 302252 377590 302910 377618
rect 303632 377590 304566 377618
rect 305012 377590 306222 377618
rect 307772 377590 307878 377618
rect 309152 377590 309534 377618
rect 310532 377590 311190 377618
rect 301228 375352 301280 375358
rect 301228 375294 301280 375300
rect 300216 374128 300268 374134
rect 300216 374070 300268 374076
rect 300124 356788 300176 356794
rect 300124 356730 300176 356736
rect 299572 261520 299624 261526
rect 299572 261462 299624 261468
rect 299584 261361 299612 261462
rect 299570 261352 299626 261361
rect 299570 261287 299626 261296
rect 299478 208176 299534 208185
rect 299478 208111 299534 208120
rect 299492 207641 299520 208111
rect 299478 207632 299534 207641
rect 299478 207567 299534 207576
rect 299386 147792 299442 147801
rect 299386 147727 299442 147736
rect 299400 147694 299428 147727
rect 299388 147688 299440 147694
rect 299388 147630 299440 147636
rect 298742 101416 298798 101425
rect 298742 101351 298798 101360
rect 296812 99340 296864 99346
rect 296812 99282 296864 99288
rect 298100 91792 298152 91798
rect 298100 91734 298152 91740
rect 298112 87009 298140 91734
rect 298098 87000 298154 87009
rect 298098 86935 298154 86944
rect 297362 72448 297418 72457
rect 297362 72383 297418 72392
rect 296720 27600 296772 27606
rect 296720 27542 296772 27548
rect 296732 26926 296760 27542
rect 296720 26920 296772 26926
rect 296720 26862 296772 26868
rect 297376 8265 297404 72383
rect 297362 8256 297418 8265
rect 297362 8191 297418 8200
rect 297376 6914 297404 8191
rect 297284 6886 297404 6914
rect 295982 3904 296038 3913
rect 295982 3839 296038 3848
rect 295904 598 296116 626
rect 295904 490 295932 598
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 295628 462 295932 490
rect 296088 480 296116 598
rect 297284 480 297312 6886
rect 298468 6180 298520 6186
rect 298468 6122 298520 6128
rect 298480 480 298508 6122
rect 299400 3194 299428 147630
rect 299584 119406 299612 261287
rect 300136 240854 300164 356730
rect 300228 355366 300256 374070
rect 300216 355360 300268 355366
rect 300216 355302 300268 355308
rect 301320 344344 301372 344350
rect 301320 344286 301372 344292
rect 301332 343670 301360 344286
rect 300952 343664 301004 343670
rect 300952 343606 301004 343612
rect 301320 343664 301372 343670
rect 301320 343606 301372 343612
rect 300860 336048 300912 336054
rect 300860 335990 300912 335996
rect 300216 248396 300268 248402
rect 300216 248338 300268 248344
rect 300228 247722 300256 248338
rect 300216 247716 300268 247722
rect 300216 247658 300268 247664
rect 300124 240848 300176 240854
rect 300124 240790 300176 240796
rect 299754 207768 299810 207777
rect 299754 207703 299810 207712
rect 299664 178696 299716 178702
rect 299664 178638 299716 178644
rect 299676 146266 299704 178638
rect 299768 150346 299796 207703
rect 300122 203688 300178 203697
rect 300122 203623 300178 203632
rect 299756 150340 299808 150346
rect 299756 150282 299808 150288
rect 299664 146260 299716 146266
rect 299664 146202 299716 146208
rect 299572 119400 299624 119406
rect 299572 119342 299624 119348
rect 300136 97306 300164 203623
rect 300228 178702 300256 247658
rect 300216 178696 300268 178702
rect 300216 178638 300268 178644
rect 300124 97300 300176 97306
rect 300124 97242 300176 97248
rect 300122 33824 300178 33833
rect 300122 33759 300178 33768
rect 299662 13152 299718 13161
rect 299662 13087 299664 13096
rect 299716 13087 299718 13096
rect 299664 13058 299716 13064
rect 300136 3913 300164 33759
rect 300872 30326 300900 335990
rect 300964 175166 300992 343606
rect 302252 261594 302280 377590
rect 302882 299568 302938 299577
rect 302882 299503 302938 299512
rect 302896 282198 302924 299503
rect 303632 291145 303660 377590
rect 305012 342281 305040 377590
rect 307772 374066 307800 377590
rect 307760 374060 307812 374066
rect 307760 374002 307812 374008
rect 307772 369073 307800 374002
rect 307758 369064 307814 369073
rect 307758 368999 307814 369008
rect 309152 363662 309180 377590
rect 309140 363656 309192 363662
rect 309140 363598 309192 363604
rect 307024 358080 307076 358086
rect 307024 358022 307076 358028
rect 304998 342272 305054 342281
rect 304998 342207 305054 342216
rect 305642 342272 305698 342281
rect 305642 342207 305698 342216
rect 304998 306504 305054 306513
rect 304998 306439 305054 306448
rect 304264 295996 304316 296002
rect 304264 295938 304316 295944
rect 304276 295458 304304 295938
rect 303712 295452 303764 295458
rect 303712 295394 303764 295400
rect 304264 295452 304316 295458
rect 304264 295394 304316 295400
rect 303618 291136 303674 291145
rect 303618 291071 303674 291080
rect 302884 282192 302936 282198
rect 302884 282134 302936 282140
rect 302884 267028 302936 267034
rect 302884 266970 302936 266976
rect 302240 261588 302292 261594
rect 302240 261530 302292 261536
rect 302240 256012 302292 256018
rect 302240 255954 302292 255960
rect 301044 250572 301096 250578
rect 301044 250514 301096 250520
rect 300952 175160 301004 175166
rect 300952 175102 301004 175108
rect 301056 96626 301084 250514
rect 301136 184204 301188 184210
rect 301136 184146 301188 184152
rect 301148 139398 301176 184146
rect 301136 139392 301188 139398
rect 301136 139334 301188 139340
rect 302252 97986 302280 255954
rect 302332 222896 302384 222902
rect 302332 222838 302384 222844
rect 302344 115938 302372 222838
rect 302332 115932 302384 115938
rect 302332 115874 302384 115880
rect 302896 108322 302924 266970
rect 303618 266384 303674 266393
rect 303618 266319 303674 266328
rect 302976 242956 303028 242962
rect 302976 242898 303028 242904
rect 302988 144294 303016 242898
rect 303632 144906 303660 266319
rect 303620 144900 303672 144906
rect 303620 144842 303672 144848
rect 302976 144288 303028 144294
rect 302976 144230 303028 144236
rect 303618 140856 303674 140865
rect 303618 140791 303620 140800
rect 303672 140791 303674 140800
rect 303620 140762 303672 140768
rect 302884 108316 302936 108322
rect 302884 108258 302936 108264
rect 302240 97980 302292 97986
rect 302240 97922 302292 97928
rect 301044 96620 301096 96626
rect 301044 96562 301096 96568
rect 301504 72480 301556 72486
rect 301504 72422 301556 72428
rect 300860 30320 300912 30326
rect 300860 30262 300912 30268
rect 301320 30320 301372 30326
rect 301320 30262 301372 30268
rect 301332 29646 301360 30262
rect 301320 29640 301372 29646
rect 301320 29582 301372 29588
rect 301516 4146 301544 72422
rect 302882 64152 302938 64161
rect 302882 64087 302938 64096
rect 302896 23361 302924 64087
rect 302974 35184 303030 35193
rect 302974 35119 303030 35128
rect 302988 34649 303016 35119
rect 302974 34640 303030 34649
rect 302974 34575 303030 34584
rect 302882 23352 302938 23361
rect 302882 23287 302938 23296
rect 302988 16574 303016 34575
rect 303526 23352 303582 23361
rect 303526 23287 303582 23296
rect 302988 16546 303200 16574
rect 301504 4140 301556 4146
rect 301504 4082 301556 4088
rect 300122 3904 300178 3913
rect 300122 3839 300178 3848
rect 299388 3188 299440 3194
rect 299388 3130 299440 3136
rect 299676 598 299888 626
rect 299676 480 299704 598
rect 299860 490 299888 598
rect 300136 490 300164 3839
rect 300766 3496 300822 3505
rect 300766 3431 300822 3440
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 299860 462 300164 490
rect 300780 480 300808 3431
rect 301964 3188 302016 3194
rect 301964 3130 302016 3136
rect 301976 480 302004 3130
rect 303172 480 303200 16546
rect 303540 3534 303568 23287
rect 303632 16574 303660 140762
rect 303724 125594 303752 295394
rect 304262 291136 304318 291145
rect 304262 291071 304318 291080
rect 304276 290465 304304 291071
rect 304262 290456 304318 290465
rect 304262 290391 304318 290400
rect 304276 264246 304304 290391
rect 304448 267028 304500 267034
rect 304448 266970 304500 266976
rect 304460 266393 304488 266970
rect 304446 266384 304502 266393
rect 304446 266319 304502 266328
rect 304264 264240 304316 264246
rect 304264 264182 304316 264188
rect 304264 218816 304316 218822
rect 304264 218758 304316 218764
rect 303804 180872 303856 180878
rect 303804 180814 303856 180820
rect 303816 156670 303844 180814
rect 303804 156664 303856 156670
rect 303804 156606 303856 156612
rect 303712 125588 303764 125594
rect 303712 125530 303764 125536
rect 304276 107642 304304 218758
rect 305012 156097 305040 306439
rect 305092 239488 305144 239494
rect 305092 239430 305144 239436
rect 305104 238785 305132 239430
rect 305090 238776 305146 238785
rect 305090 238711 305146 238720
rect 304998 156088 305054 156097
rect 304998 156023 305054 156032
rect 305104 109002 305132 238711
rect 305092 108996 305144 109002
rect 305092 108938 305144 108944
rect 304264 107636 304316 107642
rect 304264 107578 304316 107584
rect 304264 87644 304316 87650
rect 304264 87586 304316 87592
rect 304276 34649 304304 87586
rect 304262 34640 304318 34649
rect 304262 34575 304318 34584
rect 305656 20602 305684 342207
rect 305736 330608 305788 330614
rect 305736 330550 305788 330556
rect 305748 131782 305776 330550
rect 306380 253224 306432 253230
rect 306380 253166 306432 253172
rect 306392 137970 306420 253166
rect 306470 214568 306526 214577
rect 306470 214503 306526 214512
rect 306484 158030 306512 214503
rect 306472 158024 306524 158030
rect 306472 157966 306524 157972
rect 306380 137964 306432 137970
rect 306380 137906 306432 137912
rect 305736 131776 305788 131782
rect 305736 131718 305788 131724
rect 305644 20596 305696 20602
rect 305644 20538 305696 20544
rect 303632 16546 303936 16574
rect 303528 3528 303580 3534
rect 303528 3470 303580 3476
rect 303908 490 303936 16546
rect 307036 6914 307064 358022
rect 309876 355360 309928 355366
rect 309876 355302 309928 355308
rect 307116 337408 307168 337414
rect 307116 337350 307168 337356
rect 307128 225622 307156 337350
rect 309140 297492 309192 297498
rect 309140 297434 309192 297440
rect 308404 295384 308456 295390
rect 308404 295326 308456 295332
rect 308416 276690 308444 295326
rect 308404 276684 308456 276690
rect 308404 276626 308456 276632
rect 308404 262948 308456 262954
rect 308404 262890 308456 262896
rect 308416 257378 308444 262890
rect 309046 260128 309102 260137
rect 309046 260063 309102 260072
rect 309060 259457 309088 260063
rect 309046 259448 309102 259457
rect 309046 259383 309102 259392
rect 308404 257372 308456 257378
rect 308404 257314 308456 257320
rect 307760 253292 307812 253298
rect 307760 253234 307812 253240
rect 307116 225616 307168 225622
rect 307116 225558 307168 225564
rect 307114 223680 307170 223689
rect 307114 223615 307170 223624
rect 306760 6886 307064 6914
rect 306760 4078 306788 6886
rect 307128 4146 307156 223615
rect 307772 124166 307800 253234
rect 307852 199436 307904 199442
rect 307852 199378 307904 199384
rect 307864 131034 307892 199378
rect 309060 159390 309088 259383
rect 309152 164218 309180 297434
rect 309784 278792 309836 278798
rect 309784 278734 309836 278740
rect 309140 164212 309192 164218
rect 309140 164154 309192 164160
rect 309048 159384 309100 159390
rect 309048 159326 309100 159332
rect 309796 149734 309824 278734
rect 309888 259457 309916 355302
rect 309874 259448 309930 259457
rect 309874 259383 309930 259392
rect 309876 240848 309928 240854
rect 309876 240790 309928 240796
rect 309784 149728 309836 149734
rect 309784 149670 309836 149676
rect 307852 131028 307904 131034
rect 307852 130970 307904 130976
rect 307760 124160 307812 124166
rect 307760 124102 307812 124108
rect 309888 122806 309916 240790
rect 309968 209840 310020 209846
rect 309968 209782 310020 209788
rect 309980 124166 310008 209782
rect 309968 124160 310020 124166
rect 309968 124102 310020 124108
rect 309876 122800 309928 122806
rect 309876 122742 309928 122748
rect 309888 121514 309916 122742
rect 309140 121508 309192 121514
rect 309140 121450 309192 121456
rect 309876 121508 309928 121514
rect 309876 121450 309928 121456
rect 308404 62824 308456 62830
rect 308404 62766 308456 62772
rect 308416 24818 308444 62766
rect 307760 24812 307812 24818
rect 307760 24754 307812 24760
rect 308404 24812 308456 24818
rect 308404 24754 308456 24760
rect 307116 4140 307168 4146
rect 307116 4082 307168 4088
rect 306748 4072 306800 4078
rect 306748 4014 306800 4020
rect 305552 3528 305604 3534
rect 305552 3470 305604 3476
rect 304184 598 304396 626
rect 304184 490 304212 598
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 303908 462 304212 490
rect 304368 480 304396 598
rect 305564 480 305592 3470
rect 306760 480 306788 4014
rect 307772 610 307800 24754
rect 309152 6914 309180 121450
rect 309784 84856 309836 84862
rect 309784 84798 309836 84804
rect 309796 16574 309824 84798
rect 310532 17921 310560 377590
rect 312832 375222 312860 377604
rect 313292 377590 314502 377618
rect 316052 377590 316158 377618
rect 317616 377590 317998 377618
rect 311900 375216 311952 375222
rect 311900 375158 311952 375164
rect 312820 375216 312872 375222
rect 312820 375158 312872 375164
rect 311912 374134 311940 375158
rect 311900 374128 311952 374134
rect 311900 374070 311952 374076
rect 310612 250504 310664 250510
rect 310612 250446 310664 250452
rect 310624 131102 310652 250446
rect 310612 131096 310664 131102
rect 310612 131038 310664 131044
rect 311912 55214 311940 374070
rect 313292 337385 313320 377590
rect 313924 374060 313976 374066
rect 313924 374002 313976 374008
rect 313278 337376 313334 337385
rect 313278 337311 313334 337320
rect 313280 322244 313332 322250
rect 313280 322186 313332 322192
rect 311992 242208 312044 242214
rect 311992 242150 312044 242156
rect 312004 241602 312032 242150
rect 311992 241596 312044 241602
rect 311992 241538 312044 241544
rect 312004 151094 312032 241538
rect 311992 151088 312044 151094
rect 311992 151030 312044 151036
rect 313292 142118 313320 322186
rect 313372 272536 313424 272542
rect 313372 272478 313424 272484
rect 313280 142112 313332 142118
rect 313280 142054 313332 142060
rect 313384 126274 313412 272478
rect 313936 239426 313964 374002
rect 315120 293276 315172 293282
rect 315120 293218 315172 293224
rect 315132 292641 315160 293218
rect 314658 292632 314714 292641
rect 314658 292567 314714 292576
rect 315118 292632 315174 292641
rect 315118 292567 315174 292576
rect 313924 239420 313976 239426
rect 313924 239362 313976 239368
rect 313462 231160 313518 231169
rect 313462 231095 313518 231104
rect 313476 154562 313504 231095
rect 314016 175976 314068 175982
rect 314016 175918 314068 175924
rect 314028 175302 314056 175918
rect 314016 175296 314068 175302
rect 314016 175238 314068 175244
rect 314028 161474 314056 175238
rect 313936 161446 314056 161474
rect 313464 154556 313516 154562
rect 313464 154498 313516 154504
rect 313372 126268 313424 126274
rect 313372 126210 313424 126216
rect 313936 82822 313964 161446
rect 314672 103494 314700 292567
rect 316052 264314 316080 377590
rect 317616 373994 317644 377590
rect 319640 376689 319668 377604
rect 320192 377590 321310 377618
rect 319626 376680 319682 376689
rect 319626 376615 319682 376624
rect 319640 373994 319668 376615
rect 317340 373966 317644 373994
rect 319456 373966 319668 373994
rect 316040 264308 316092 264314
rect 316040 264250 316092 264256
rect 317236 246356 317288 246362
rect 317236 246298 317288 246304
rect 317248 245682 317276 246298
rect 316040 245676 316092 245682
rect 316040 245618 316092 245624
rect 317236 245676 317288 245682
rect 317236 245618 317288 245624
rect 315302 213208 315358 213217
rect 315302 213143 315358 213152
rect 315316 125594 315344 213143
rect 316052 128246 316080 245618
rect 316682 228304 316738 228313
rect 316682 228239 316738 228248
rect 316040 128240 316092 128246
rect 316040 128182 316092 128188
rect 315304 125588 315356 125594
rect 315304 125530 315356 125536
rect 314660 103488 314712 103494
rect 314660 103430 314712 103436
rect 314014 84824 314070 84833
rect 314014 84759 314070 84768
rect 313924 82816 313976 82822
rect 313922 82784 313924 82793
rect 313976 82784 313978 82793
rect 313922 82719 313978 82728
rect 313936 82693 313964 82719
rect 311900 55208 311952 55214
rect 311900 55150 311952 55156
rect 311912 54602 311940 55150
rect 311900 54596 311952 54602
rect 311900 54538 311952 54544
rect 310518 17912 310574 17921
rect 310518 17847 310574 17856
rect 309796 16546 309916 16574
rect 309152 6886 309824 6914
rect 307944 4140 307996 4146
rect 307944 4082 307996 4088
rect 307760 604 307812 610
rect 307760 546 307812 552
rect 307956 480 307984 4082
rect 309048 604 309100 610
rect 309048 546 309100 552
rect 309060 480 309088 546
rect 309796 490 309824 6886
rect 309888 4146 309916 16546
rect 310532 15162 310560 17847
rect 310520 15156 310572 15162
rect 310520 15098 310572 15104
rect 311440 14544 311492 14550
rect 311440 14486 311492 14492
rect 309876 4140 309928 4146
rect 309876 4082 309928 4088
rect 310072 598 310284 626
rect 310072 490 310100 598
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 309796 462 310100 490
rect 310256 480 310284 598
rect 311452 480 311480 14486
rect 314028 9625 314056 84759
rect 314660 44872 314712 44878
rect 314660 44814 314712 44820
rect 314014 9616 314070 9625
rect 314014 9551 314070 9560
rect 314028 6914 314056 9551
rect 313844 6886 314056 6914
rect 312636 4004 312688 4010
rect 312636 3946 312688 3952
rect 312648 480 312676 3946
rect 313844 480 313872 6886
rect 314672 490 314700 44814
rect 316040 20664 316092 20670
rect 316040 20606 316092 20612
rect 316052 16574 316080 20606
rect 316052 16546 316264 16574
rect 314856 598 315068 626
rect 314856 490 314884 598
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314672 462 314884 490
rect 315040 480 315068 598
rect 316236 480 316264 16546
rect 316696 5506 316724 228239
rect 317340 215121 317368 373966
rect 319456 351257 319484 373966
rect 320192 361729 320220 377590
rect 322204 374672 322256 374678
rect 322204 374614 322256 374620
rect 320178 361720 320234 361729
rect 320178 361655 320234 361664
rect 320822 361720 320878 361729
rect 320822 361655 320878 361664
rect 319442 351248 319498 351257
rect 319442 351183 319498 351192
rect 320180 316736 320232 316742
rect 320180 316678 320232 316684
rect 320192 316130 320220 316678
rect 320180 316124 320232 316130
rect 320180 316066 320232 316072
rect 317418 313304 317474 313313
rect 317418 313239 317474 313248
rect 317326 215112 317382 215121
rect 317326 215047 317382 215056
rect 317340 214606 317368 215047
rect 317328 214600 317380 214606
rect 317328 214542 317380 214548
rect 316774 195392 316830 195401
rect 316774 195327 316830 195336
rect 316788 20670 316816 195327
rect 317432 150414 317460 313239
rect 318798 307864 318854 307873
rect 318798 307799 318854 307808
rect 318154 302288 318210 302297
rect 318154 302223 318210 302232
rect 318168 195362 318196 302223
rect 318246 211168 318302 211177
rect 318246 211103 318302 211112
rect 318156 195356 318208 195362
rect 318156 195298 318208 195304
rect 318062 195256 318118 195265
rect 318062 195191 318118 195200
rect 317420 150408 317472 150414
rect 317420 150350 317472 150356
rect 316776 20664 316828 20670
rect 316776 20606 316828 20612
rect 318076 6798 318104 195191
rect 318260 129062 318288 211103
rect 318812 135250 318840 307799
rect 319444 282940 319496 282946
rect 319444 282882 319496 282888
rect 319456 163538 319484 282882
rect 319444 163532 319496 163538
rect 319444 163474 319496 163480
rect 320192 160070 320220 316066
rect 320180 160064 320232 160070
rect 320180 160006 320232 160012
rect 318800 135244 318852 135250
rect 318800 135186 318852 135192
rect 318248 129056 318300 129062
rect 318248 128998 318300 129004
rect 319442 73808 319498 73817
rect 319442 73743 319498 73752
rect 318156 64184 318208 64190
rect 318156 64126 318208 64132
rect 318064 6792 318116 6798
rect 318064 6734 318116 6740
rect 316684 5500 316736 5506
rect 316684 5442 316736 5448
rect 317328 5500 317380 5506
rect 317328 5442 317380 5448
rect 317340 480 317368 5442
rect 318168 4010 318196 64126
rect 319456 6798 319484 73743
rect 320836 35902 320864 361655
rect 322216 291854 322244 374614
rect 322294 358048 322350 358057
rect 322294 357983 322350 357992
rect 322204 291848 322256 291854
rect 322204 291790 322256 291796
rect 322308 276758 322336 357983
rect 322296 276752 322348 276758
rect 322296 276694 322348 276700
rect 322204 251864 322256 251870
rect 322204 251806 322256 251812
rect 321560 215960 321612 215966
rect 321560 215902 321612 215908
rect 320914 185736 320970 185745
rect 320914 185671 320970 185680
rect 320928 106282 320956 185671
rect 321572 113150 321600 215902
rect 322216 145586 322244 251806
rect 322952 239494 322980 377604
rect 324332 377590 324622 377618
rect 326278 377590 326384 377618
rect 324332 345681 324360 377590
rect 326356 374066 326384 377590
rect 327092 377590 327934 377618
rect 328472 377590 329590 377618
rect 326344 374060 326396 374066
rect 326344 374002 326396 374008
rect 324686 358184 324742 358193
rect 324686 358119 324742 358128
rect 325606 358184 325662 358193
rect 325606 358119 325662 358128
rect 324700 357513 324728 358119
rect 324686 357504 324742 357513
rect 324686 357439 324742 357448
rect 324318 345672 324374 345681
rect 324318 345607 324374 345616
rect 323030 321600 323086 321609
rect 323030 321535 323086 321544
rect 322940 239488 322992 239494
rect 322940 239430 322992 239436
rect 322296 233912 322348 233918
rect 322296 233854 322348 233860
rect 322204 145580 322256 145586
rect 322204 145522 322256 145528
rect 322202 139496 322258 139505
rect 322202 139431 322258 139440
rect 321560 113144 321612 113150
rect 321560 113086 321612 113092
rect 320916 106276 320968 106282
rect 320916 106218 320968 106224
rect 321560 46232 321612 46238
rect 321560 46174 321612 46180
rect 320824 35896 320876 35902
rect 320824 35838 320876 35844
rect 320836 34542 320864 35838
rect 320180 34536 320232 34542
rect 320180 34478 320232 34484
rect 320824 34536 320876 34542
rect 320824 34478 320876 34484
rect 320192 16574 320220 34478
rect 321572 16574 321600 46174
rect 320192 16546 320496 16574
rect 321572 16546 322152 16574
rect 319444 6792 319496 6798
rect 319444 6734 319496 6740
rect 319456 4570 319484 6734
rect 319456 4542 319760 4570
rect 318156 4004 318208 4010
rect 318156 3946 318208 3952
rect 318522 3360 318578 3369
rect 318522 3295 318578 3304
rect 318536 480 318564 3295
rect 319732 480 319760 4542
rect 320468 490 320496 16546
rect 320744 598 320956 626
rect 320744 490 320772 598
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320468 462 320772 490
rect 320928 480 320956 598
rect 322124 480 322152 16546
rect 322216 3777 322244 139431
rect 322308 103494 322336 233854
rect 323044 147626 323072 321535
rect 324320 298784 324372 298790
rect 324320 298726 324372 298732
rect 324332 298178 324360 298726
rect 324320 298172 324372 298178
rect 324320 298114 324372 298120
rect 323584 268388 323636 268394
rect 323584 268330 323636 268336
rect 323032 147620 323084 147626
rect 323032 147562 323084 147568
rect 323596 114510 323624 268330
rect 323674 221504 323730 221513
rect 323674 221439 323730 221448
rect 323584 114504 323636 114510
rect 323584 114446 323636 114452
rect 322296 103488 322348 103494
rect 322296 103430 322348 103436
rect 323688 69018 323716 221439
rect 324332 132462 324360 298114
rect 325620 195294 325648 358119
rect 326356 352617 326384 374002
rect 326342 352608 326398 352617
rect 326342 352543 326398 352552
rect 326988 326392 327040 326398
rect 326988 326334 327040 326340
rect 327000 325718 327028 326334
rect 325700 325712 325752 325718
rect 325700 325654 325752 325660
rect 326988 325712 327040 325718
rect 326988 325654 327040 325660
rect 325608 195288 325660 195294
rect 325608 195230 325660 195236
rect 324962 191176 325018 191185
rect 324962 191111 325018 191120
rect 324320 132456 324372 132462
rect 324320 132398 324372 132404
rect 324976 83502 325004 191111
rect 325712 161430 325740 325654
rect 327092 228993 327120 377590
rect 328472 358193 328500 377590
rect 329104 374060 329156 374066
rect 329104 374002 329156 374008
rect 328458 358184 328514 358193
rect 328458 358119 328514 358128
rect 327724 311908 327776 311914
rect 327724 311850 327776 311856
rect 327172 244316 327224 244322
rect 327172 244258 327224 244264
rect 327078 228984 327134 228993
rect 327078 228919 327134 228928
rect 327092 228410 327120 228919
rect 327080 228404 327132 228410
rect 327080 228346 327132 228352
rect 326344 195356 326396 195362
rect 326344 195298 326396 195304
rect 325700 161424 325752 161430
rect 325700 161366 325752 161372
rect 324964 83496 325016 83502
rect 324964 83438 325016 83444
rect 322940 69012 322992 69018
rect 322940 68954 322992 68960
rect 323676 69012 323728 69018
rect 323676 68954 323728 68960
rect 322202 3768 322258 3777
rect 322202 3703 322258 3712
rect 322952 490 322980 68954
rect 324412 5568 324464 5574
rect 324412 5510 324464 5516
rect 323136 598 323348 626
rect 323136 490 323164 598
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 322952 462 323164 490
rect 323320 480 323348 598
rect 324424 480 324452 5510
rect 324976 3262 325004 83438
rect 325054 37904 325110 37913
rect 325054 37839 325110 37848
rect 325068 6866 325096 37839
rect 325056 6860 325108 6866
rect 325056 6802 325108 6808
rect 325068 5574 325096 6802
rect 325056 5568 325108 5574
rect 325056 5510 325108 5516
rect 326356 4049 326384 195298
rect 327184 135930 327212 244258
rect 327172 135924 327224 135930
rect 327172 135866 327224 135872
rect 327080 131776 327132 131782
rect 327080 131718 327132 131724
rect 327092 16574 327120 131718
rect 327736 104854 327764 311850
rect 328368 244996 328420 245002
rect 328368 244938 328420 244944
rect 328380 244322 328408 244938
rect 328368 244316 328420 244322
rect 328368 244258 328420 244264
rect 329116 143546 329144 374002
rect 330300 323604 330352 323610
rect 330300 323546 330352 323552
rect 330312 322998 330340 323546
rect 329840 322992 329892 322998
rect 329840 322934 329892 322940
rect 330300 322992 330352 322998
rect 330300 322934 330352 322940
rect 329852 162790 329880 322934
rect 331232 246362 331260 377604
rect 332612 377590 332902 377618
rect 331862 371920 331918 371929
rect 331862 371855 331918 371864
rect 331220 246356 331272 246362
rect 331220 246298 331272 246304
rect 329840 162784 329892 162790
rect 329840 162726 329892 162732
rect 329104 143540 329156 143546
rect 329104 143482 329156 143488
rect 330484 143540 330536 143546
rect 330484 143482 330536 143488
rect 329102 140856 329158 140865
rect 329102 140791 329158 140800
rect 327724 104848 327776 104854
rect 327724 104790 327776 104796
rect 327092 16546 328040 16574
rect 326342 4040 326398 4049
rect 326342 3975 326398 3984
rect 324964 3256 325016 3262
rect 324964 3198 325016 3204
rect 325608 3256 325660 3262
rect 325608 3198 325660 3204
rect 325620 480 325648 3198
rect 326356 490 326384 3975
rect 326632 598 326844 626
rect 326632 490 326660 598
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326356 462 326660 490
rect 326816 480 326844 598
rect 328012 480 328040 16546
rect 328736 14476 328788 14482
rect 328736 14418 328788 14424
rect 328748 490 328776 14418
rect 329116 3369 329144 140791
rect 330496 66910 330524 143482
rect 331220 80708 331272 80714
rect 331220 80650 331272 80656
rect 330484 66904 330536 66910
rect 330484 66846 330536 66852
rect 330496 6914 330524 66846
rect 330404 6886 330524 6914
rect 329102 3360 329158 3369
rect 329102 3295 329158 3304
rect 329024 598 329236 626
rect 329024 490 329052 598
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 328748 462 329052 490
rect 329208 480 329236 598
rect 330404 480 330432 6886
rect 331232 490 331260 80650
rect 331876 64870 331904 371855
rect 332612 345030 332640 377590
rect 334544 374678 334572 377604
rect 335372 377590 336214 377618
rect 334532 374672 334584 374678
rect 334532 374614 334584 374620
rect 334716 374672 334768 374678
rect 334716 374614 334768 374620
rect 332600 345024 332652 345030
rect 332600 344966 332652 344972
rect 334624 254652 334676 254658
rect 334624 254594 334676 254600
rect 331956 251184 332008 251190
rect 331956 251126 332008 251132
rect 331968 235385 331996 251126
rect 331954 235376 332010 235385
rect 331954 235311 332010 235320
rect 331968 153882 331996 235311
rect 331956 153876 332008 153882
rect 331956 153818 332008 153824
rect 331956 135924 332008 135930
rect 331956 135866 332008 135872
rect 331968 94518 331996 135866
rect 334636 96626 334664 254594
rect 334728 251190 334756 374614
rect 335372 349858 335400 377590
rect 337856 375358 337884 377604
rect 339512 375358 339540 377604
rect 336004 375352 336056 375358
rect 336004 375294 336056 375300
rect 337844 375352 337896 375358
rect 337844 375294 337896 375300
rect 339500 375352 339552 375358
rect 339500 375294 339552 375300
rect 335360 349852 335412 349858
rect 335360 349794 335412 349800
rect 334716 251184 334768 251190
rect 334716 251126 334768 251132
rect 336016 175982 336044 375294
rect 339512 374678 339540 375294
rect 339500 374672 339552 374678
rect 341168 374649 341196 377604
rect 342272 377590 342838 377618
rect 343652 377590 344494 377618
rect 345032 377590 346150 377618
rect 339500 374614 339552 374620
rect 341154 374640 341210 374649
rect 341154 374575 341210 374584
rect 340144 366444 340196 366450
rect 340144 366386 340196 366392
rect 340156 365770 340184 366386
rect 341616 366376 341668 366382
rect 341616 366318 341668 366324
rect 340144 365764 340196 365770
rect 340144 365706 340196 365712
rect 338764 362228 338816 362234
rect 338764 362170 338816 362176
rect 338026 361040 338082 361049
rect 338026 360975 338082 360984
rect 338040 360233 338068 360975
rect 337382 360224 337438 360233
rect 337382 360159 337438 360168
rect 338026 360224 338082 360233
rect 338026 360159 338082 360168
rect 336094 236056 336150 236065
rect 336094 235991 336150 236000
rect 336004 175976 336056 175982
rect 336004 175918 336056 175924
rect 334716 150476 334768 150482
rect 334716 150418 334768 150424
rect 334624 96620 334676 96626
rect 334624 96562 334676 96568
rect 331956 94512 332008 94518
rect 331956 94454 332008 94460
rect 332600 65544 332652 65550
rect 332600 65486 332652 65492
rect 331864 64864 331916 64870
rect 331864 64806 331916 64812
rect 331876 64190 331904 64806
rect 331864 64184 331916 64190
rect 331864 64126 331916 64132
rect 332612 3534 332640 65486
rect 334728 47598 334756 150418
rect 335358 137728 335414 137737
rect 335358 137663 335414 137672
rect 334716 47592 334768 47598
rect 334716 47534 334768 47540
rect 333980 37936 334032 37942
rect 333980 37878 334032 37884
rect 333992 16574 334020 37878
rect 335372 16574 335400 137663
rect 336108 111790 336136 235991
rect 336096 111784 336148 111790
rect 336096 111726 336148 111732
rect 337396 48278 337424 360159
rect 338118 335472 338174 335481
rect 338118 335407 338174 335416
rect 337476 79348 337528 79354
rect 337476 79290 337528 79296
rect 337384 48272 337436 48278
rect 337384 48214 337436 48220
rect 337396 48074 337424 48214
rect 336004 48068 336056 48074
rect 336004 48010 336056 48016
rect 337384 48068 337436 48074
rect 337384 48010 337436 48016
rect 333992 16546 334664 16574
rect 335372 16546 335952 16574
rect 332692 4072 332744 4078
rect 332692 4014 332744 4020
rect 332600 3528 332652 3534
rect 332600 3470 332652 3476
rect 331416 598 331628 626
rect 331416 490 331444 598
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331232 462 331444 490
rect 331600 480 331628 598
rect 332704 480 332732 4014
rect 333888 3528 333940 3534
rect 333888 3470 333940 3476
rect 333900 480 333928 3470
rect 334636 490 334664 16546
rect 335924 3482 335952 16546
rect 336016 4078 336044 48010
rect 337488 20602 337516 79290
rect 338132 37942 338160 335407
rect 338776 222902 338804 362170
rect 338764 222896 338816 222902
rect 338764 222838 338816 222844
rect 338212 119400 338264 119406
rect 338212 119342 338264 119348
rect 338120 37936 338172 37942
rect 338120 37878 338172 37884
rect 336740 20596 336792 20602
rect 336740 20538 336792 20544
rect 337476 20596 337528 20602
rect 337476 20538 337528 20544
rect 336752 16574 336780 20538
rect 338224 16574 338252 119342
rect 340156 80714 340184 365706
rect 341524 324964 341576 324970
rect 341524 324906 341576 324912
rect 340236 244928 340288 244934
rect 340236 244870 340288 244876
rect 340248 128314 340276 244870
rect 340236 128308 340288 128314
rect 340236 128250 340288 128256
rect 340144 80708 340196 80714
rect 340144 80650 340196 80656
rect 339500 51740 339552 51746
rect 339500 51682 339552 51688
rect 339408 38616 339460 38622
rect 339408 38558 339460 38564
rect 339420 37942 339448 38558
rect 339408 37936 339460 37942
rect 339408 37878 339460 37884
rect 336752 16546 337056 16574
rect 338224 16546 338712 16574
rect 336004 4072 336056 4078
rect 336004 4014 336056 4020
rect 335924 3454 336320 3482
rect 334912 598 335124 626
rect 334912 490 334940 598
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 334636 462 334940 490
rect 335096 480 335124 598
rect 336292 480 336320 3454
rect 337028 490 337056 16546
rect 337304 598 337516 626
rect 337304 490 337332 598
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337028 462 337332 490
rect 337488 480 337516 598
rect 338684 480 338712 16546
rect 339512 490 339540 51682
rect 341536 19378 341564 324906
rect 341628 298790 341656 366318
rect 342272 318102 342300 377590
rect 342904 376100 342956 376106
rect 342904 376042 342956 376048
rect 342260 318096 342312 318102
rect 342260 318038 342312 318044
rect 341616 298784 341668 298790
rect 341616 298726 341668 298732
rect 342916 243574 342944 376042
rect 343652 369850 343680 377590
rect 345032 370530 345060 377590
rect 345664 377460 345716 377466
rect 345664 377402 345716 377408
rect 345020 370524 345072 370530
rect 345020 370466 345072 370472
rect 343640 369844 343692 369850
rect 343640 369786 343692 369792
rect 344284 369844 344336 369850
rect 344284 369786 344336 369792
rect 344296 332586 344324 369786
rect 344284 332580 344336 332586
rect 344284 332522 344336 332528
rect 344282 319424 344338 319433
rect 344282 319359 344338 319368
rect 342904 243568 342956 243574
rect 342904 243510 342956 243516
rect 342994 235240 343050 235249
rect 342994 235175 343050 235184
rect 342904 139528 342956 139534
rect 342904 139470 342956 139476
rect 341524 19372 341576 19378
rect 341524 19314 341576 19320
rect 340970 3496 341026 3505
rect 340970 3431 341026 3440
rect 339696 598 339908 626
rect 339696 490 339724 598
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339512 462 339724 490
rect 339880 480 339908 598
rect 340984 480 341012 3431
rect 341536 3262 341564 19314
rect 342168 7608 342220 7614
rect 342168 7550 342220 7556
rect 341524 3256 341576 3262
rect 341524 3198 341576 3204
rect 342180 480 342208 7550
rect 342916 4146 342944 139470
rect 343008 121446 343036 235175
rect 342996 121440 343048 121446
rect 342996 121382 343048 121388
rect 344296 27538 344324 319359
rect 345676 242214 345704 377402
rect 345756 367804 345808 367810
rect 345756 367746 345808 367752
rect 345768 307086 345796 367746
rect 347042 340096 347098 340105
rect 347042 340031 347098 340040
rect 345756 307080 345808 307086
rect 345756 307022 345808 307028
rect 345664 242208 345716 242214
rect 345664 242150 345716 242156
rect 345664 239420 345716 239426
rect 345664 239362 345716 239368
rect 344284 27532 344336 27538
rect 344284 27474 344336 27480
rect 343364 15904 343416 15910
rect 343364 15846 343416 15852
rect 342904 4140 342956 4146
rect 342904 4082 342956 4088
rect 343376 480 343404 15846
rect 344296 3505 344324 27474
rect 345676 8294 345704 239362
rect 347056 81394 347084 340031
rect 347792 287706 347820 377604
rect 349172 377590 349462 377618
rect 350552 377590 351118 377618
rect 351932 377590 352774 377618
rect 353312 377590 354430 377618
rect 348424 367872 348476 367878
rect 348424 367814 348476 367820
rect 348436 326398 348464 367814
rect 349172 328438 349200 377590
rect 350552 373318 350580 377590
rect 351182 377360 351238 377369
rect 351182 377295 351238 377304
rect 350540 373312 350592 373318
rect 350540 373254 350592 373260
rect 349160 328432 349212 328438
rect 349160 328374 349212 328380
rect 348424 326392 348476 326398
rect 348424 326334 348476 326340
rect 351196 323610 351224 377295
rect 351184 323604 351236 323610
rect 351184 323546 351236 323552
rect 351932 316810 351960 377590
rect 353312 360097 353340 377590
rect 355322 377567 355378 377576
rect 354036 374060 354088 374066
rect 354036 374002 354088 374008
rect 353942 366344 353998 366353
rect 353942 366279 353998 366288
rect 353298 360088 353354 360097
rect 353298 360023 353354 360032
rect 353956 338774 353984 366279
rect 353944 338768 353996 338774
rect 353944 338710 353996 338716
rect 351920 316804 351972 316810
rect 351920 316746 351972 316752
rect 352564 316804 352616 316810
rect 352564 316746 352616 316752
rect 352576 316062 352604 316746
rect 352564 316056 352616 316062
rect 352564 315998 352616 316004
rect 349802 315344 349858 315353
rect 349802 315279 349858 315288
rect 347780 287700 347832 287706
rect 347780 287642 347832 287648
rect 348424 249144 348476 249150
rect 348424 249086 348476 249092
rect 347044 81388 347096 81394
rect 347044 81330 347096 81336
rect 346400 21480 346452 21486
rect 346400 21422 346452 21428
rect 346412 19378 346440 21422
rect 346400 19372 346452 19378
rect 346400 19314 346452 19320
rect 345664 8288 345716 8294
rect 345664 8230 345716 8236
rect 345676 6914 345704 8230
rect 345676 6886 345796 6914
rect 344282 3496 344338 3505
rect 344282 3431 344338 3440
rect 344560 3256 344612 3262
rect 344560 3198 344612 3204
rect 344572 480 344600 3198
rect 345768 480 345796 6886
rect 348436 4146 348464 249086
rect 349816 94489 349844 315279
rect 352576 285025 352604 315998
rect 352562 285016 352618 285025
rect 352562 284951 352618 284960
rect 352564 283620 352616 283626
rect 352564 283562 352616 283568
rect 351182 196616 351238 196625
rect 351182 196551 351238 196560
rect 349896 195288 349948 195294
rect 349896 195230 349948 195236
rect 349802 94480 349858 94489
rect 349802 94415 349858 94424
rect 349908 89010 349936 195230
rect 349896 89004 349948 89010
rect 349896 88946 349948 88952
rect 348424 4140 348476 4146
rect 348424 4082 348476 4088
rect 346950 3360 347006 3369
rect 346950 3295 347006 3304
rect 346964 480 346992 3295
rect 348068 598 348280 626
rect 348068 480 348096 598
rect 348252 490 348280 598
rect 348436 490 348464 4082
rect 351196 3670 351224 196551
rect 352576 118658 352604 283562
rect 353944 275392 353996 275398
rect 353944 275334 353996 275340
rect 353956 158030 353984 275334
rect 354048 261526 354076 374002
rect 354588 362296 354640 362302
rect 354588 362238 354640 362244
rect 354036 261520 354088 261526
rect 354036 261462 354088 261468
rect 353944 158024 353996 158030
rect 353944 157966 353996 157972
rect 352654 138680 352710 138689
rect 352654 138615 352710 138624
rect 352564 118652 352616 118658
rect 352564 118594 352616 118600
rect 352668 65550 352696 138615
rect 354600 126274 354628 362238
rect 355336 344350 355364 377567
rect 356072 374066 356100 377604
rect 356060 374060 356112 374066
rect 356060 374002 356112 374008
rect 355324 344344 355376 344350
rect 355324 344286 355376 344292
rect 356164 311137 356192 489886
rect 356242 423736 356298 423745
rect 356242 423671 356298 423680
rect 356256 366450 356284 423671
rect 356334 382392 356390 382401
rect 356334 382327 356390 382336
rect 356348 377641 356376 382327
rect 356334 377632 356390 377641
rect 356334 377567 356390 377576
rect 356244 366444 356296 366450
rect 356244 366386 356296 366392
rect 356716 349178 356744 507583
rect 357164 496800 357216 496806
rect 357164 496742 357216 496748
rect 357176 495553 357204 496742
rect 357162 495544 357218 495553
rect 357162 495479 357218 495488
rect 358096 487257 358124 514927
rect 358726 510096 358782 510105
rect 358726 510031 358782 510040
rect 358740 509726 358768 510031
rect 358728 509720 358780 509726
rect 358728 509662 358780 509668
rect 358726 505200 358782 505209
rect 358726 505135 358728 505144
rect 358780 505135 358782 505144
rect 358728 505106 358780 505112
rect 358726 502752 358782 502761
rect 358726 502687 358782 502696
rect 358740 502382 358768 502687
rect 358728 502376 358780 502382
rect 358728 502318 358780 502324
rect 358636 494012 358688 494018
rect 358636 493954 358688 493960
rect 358648 493105 358676 493954
rect 358634 493096 358690 493105
rect 358634 493031 358690 493040
rect 358726 487792 358782 487801
rect 358726 487727 358782 487736
rect 358082 487248 358138 487257
rect 358082 487183 358138 487192
rect 358740 486470 358768 487727
rect 358728 486464 358780 486470
rect 358728 486406 358780 486412
rect 358082 485344 358138 485353
rect 358082 485279 358138 485288
rect 357898 470656 357954 470665
rect 357898 470591 357900 470600
rect 357952 470591 357954 470600
rect 357900 470562 357952 470568
rect 357438 458416 357494 458425
rect 357438 458351 357494 458360
rect 357452 373289 357480 458351
rect 357530 438968 357586 438977
rect 357530 438903 357586 438912
rect 357438 373280 357494 373289
rect 357438 373215 357494 373224
rect 357544 362273 357572 438903
rect 357898 436384 357954 436393
rect 357898 436319 357954 436328
rect 357912 436150 357940 436319
rect 357900 436144 357952 436150
rect 357900 436086 357952 436092
rect 358096 420238 358124 485279
rect 358726 482896 358782 482905
rect 358726 482831 358782 482840
rect 358740 481710 358768 482831
rect 358728 481704 358780 481710
rect 358728 481646 358780 481652
rect 358726 480448 358782 480457
rect 358726 480383 358782 480392
rect 358740 480282 358768 480383
rect 358728 480276 358780 480282
rect 358728 480218 358780 480224
rect 358726 478000 358782 478009
rect 358726 477935 358782 477944
rect 358740 477562 358768 477935
rect 358728 477556 358780 477562
rect 358728 477498 358780 477504
rect 358542 473104 358598 473113
rect 358542 473039 358598 473048
rect 358556 472054 358584 473039
rect 358544 472048 358596 472054
rect 358544 471990 358596 471996
rect 358726 465760 358782 465769
rect 358726 465695 358782 465704
rect 358740 465118 358768 465695
rect 358728 465112 358780 465118
rect 358728 465054 358780 465060
rect 358450 460864 358506 460873
rect 358450 460799 358506 460808
rect 358464 459610 358492 460799
rect 358452 459604 358504 459610
rect 358452 459546 358504 459552
rect 358726 455968 358782 455977
rect 358726 455903 358782 455912
rect 358740 455462 358768 455903
rect 358728 455456 358780 455462
rect 358728 455398 358780 455404
rect 358726 453520 358782 453529
rect 358726 453455 358782 453464
rect 358740 452674 358768 453455
rect 358728 452668 358780 452674
rect 358728 452610 358780 452616
rect 358726 451072 358782 451081
rect 358726 451007 358782 451016
rect 358740 449954 358768 451007
rect 358728 449948 358780 449954
rect 358728 449890 358780 449896
rect 358728 449200 358780 449206
rect 358728 449142 358780 449148
rect 358740 448769 358768 449142
rect 358726 448760 358782 448769
rect 358726 448695 358782 448704
rect 358726 446176 358782 446185
rect 358726 446111 358782 446120
rect 358740 445806 358768 446111
rect 358728 445800 358780 445806
rect 358728 445742 358780 445748
rect 358726 443728 358782 443737
rect 358726 443663 358782 443672
rect 358740 443018 358768 443663
rect 358728 443012 358780 443018
rect 358728 442954 358780 442960
rect 358726 441280 358782 441289
rect 358726 441215 358782 441224
rect 358740 440298 358768 441215
rect 358728 440292 358780 440298
rect 358728 440234 358780 440240
rect 358726 438968 358782 438977
rect 358726 438903 358728 438912
rect 358780 438903 358782 438912
rect 358728 438874 358780 438880
rect 358726 433936 358782 433945
rect 358726 433871 358782 433880
rect 358740 433362 358768 433871
rect 358728 433356 358780 433362
rect 358728 433298 358780 433304
rect 358726 431488 358782 431497
rect 358726 431423 358782 431432
rect 358740 430642 358768 431423
rect 358728 430636 358780 430642
rect 358728 430578 358780 430584
rect 358726 429040 358782 429049
rect 358726 428975 358782 428984
rect 358740 427854 358768 428975
rect 358728 427848 358780 427854
rect 358728 427790 358780 427796
rect 358726 426592 358782 426601
rect 358726 426527 358782 426536
rect 358740 426494 358768 426527
rect 358728 426488 358780 426494
rect 358728 426430 358780 426436
rect 358726 421696 358782 421705
rect 358726 421631 358782 421640
rect 358740 420986 358768 421631
rect 358728 420980 358780 420986
rect 358728 420922 358780 420928
rect 358084 420232 358136 420238
rect 358084 420174 358136 420180
rect 358726 419248 358782 419257
rect 358726 419183 358782 419192
rect 358740 418198 358768 419183
rect 358728 418192 358780 418198
rect 358728 418134 358780 418140
rect 358728 416832 358780 416838
rect 358726 416800 358728 416809
rect 358780 416800 358782 416809
rect 358726 416735 358782 416744
rect 358726 414352 358782 414361
rect 358726 414287 358782 414296
rect 358740 414050 358768 414287
rect 358728 414044 358780 414050
rect 358728 413986 358780 413992
rect 358726 411904 358782 411913
rect 358726 411839 358782 411848
rect 358740 411330 358768 411839
rect 358728 411324 358780 411330
rect 358728 411266 358780 411272
rect 358726 409456 358782 409465
rect 358726 409391 358782 409400
rect 358740 408542 358768 409391
rect 358728 408536 358780 408542
rect 358728 408478 358780 408484
rect 358726 407008 358782 407017
rect 358726 406943 358782 406952
rect 358740 405754 358768 406943
rect 358728 405748 358780 405754
rect 358728 405690 358780 405696
rect 358726 404288 358782 404297
rect 358726 404223 358782 404232
rect 358740 403510 358768 404223
rect 358728 403504 358780 403510
rect 358728 403446 358780 403452
rect 358726 401840 358782 401849
rect 358726 401775 358782 401784
rect 358740 401674 358768 401775
rect 358728 401668 358780 401674
rect 358728 401610 358780 401616
rect 358634 399392 358690 399401
rect 358634 399327 358690 399336
rect 358648 398886 358676 399327
rect 358636 398880 358688 398886
rect 358636 398822 358688 398828
rect 358726 394496 358782 394505
rect 358726 394431 358782 394440
rect 358740 393378 358768 394431
rect 358728 393372 358780 393378
rect 358728 393314 358780 393320
rect 357622 392048 357678 392057
rect 357622 391983 357678 391992
rect 357636 376106 357664 391983
rect 357714 389600 357770 389609
rect 357714 389535 357770 389544
rect 357728 377466 357756 389535
rect 358726 387152 358782 387161
rect 358726 387087 358782 387096
rect 358740 386442 358768 387087
rect 358728 386436 358780 386442
rect 358728 386378 358780 386384
rect 358726 384704 358782 384713
rect 358726 384639 358782 384648
rect 358740 383722 358768 384639
rect 358728 383716 358780 383722
rect 358728 383658 358780 383664
rect 358634 379808 358690 379817
rect 358634 379743 358690 379752
rect 358648 379574 358676 379743
rect 358636 379568 358688 379574
rect 358636 379510 358688 379516
rect 357716 377460 357768 377466
rect 357716 377402 357768 377408
rect 357624 376100 357676 376106
rect 357624 376042 357676 376048
rect 358082 375184 358138 375193
rect 358082 375119 358138 375128
rect 357530 362264 357586 362273
rect 357530 362199 357586 362208
rect 356704 349172 356756 349178
rect 356704 349114 356756 349120
rect 357348 349172 357400 349178
rect 357348 349114 357400 349120
rect 357360 348498 357388 349114
rect 357348 348492 357400 348498
rect 357348 348434 357400 348440
rect 358096 327078 358124 375119
rect 358176 371272 358228 371278
rect 358176 371214 358228 371220
rect 358188 337414 358216 371214
rect 358728 365016 358780 365022
rect 358728 364958 358780 364964
rect 358176 337408 358228 337414
rect 358176 337350 358228 337356
rect 358084 327072 358136 327078
rect 358084 327014 358136 327020
rect 356150 311128 356206 311137
rect 356150 311063 356206 311072
rect 356794 311128 356850 311137
rect 356794 311063 356850 311072
rect 355324 268388 355376 268394
rect 355324 268330 355376 268336
rect 355336 233209 355364 268330
rect 356704 251252 356756 251258
rect 356704 251194 356756 251200
rect 355322 233200 355378 233209
rect 355322 233135 355378 233144
rect 356716 148374 356744 251194
rect 356808 244934 356836 311063
rect 358084 309188 358136 309194
rect 358084 309130 358136 309136
rect 356796 244928 356848 244934
rect 356796 244870 356848 244876
rect 356794 204912 356850 204921
rect 356794 204847 356850 204856
rect 356704 148368 356756 148374
rect 356704 148310 356756 148316
rect 356702 142488 356758 142497
rect 356702 142423 356758 142432
rect 353944 126268 353996 126274
rect 353944 126210 353996 126216
rect 354588 126268 354640 126274
rect 354588 126210 354640 126216
rect 352656 65544 352708 65550
rect 352562 65512 352618 65521
rect 352656 65486 352708 65492
rect 352562 65447 352618 65456
rect 352576 4049 352604 65447
rect 353956 62830 353984 126210
rect 355324 80708 355376 80714
rect 355324 80650 355376 80656
rect 355336 63510 355364 80650
rect 355324 63504 355376 63510
rect 355324 63446 355376 63452
rect 353944 62824 353996 62830
rect 353944 62766 353996 62772
rect 356716 7614 356744 142423
rect 356808 115938 356836 204847
rect 356796 115932 356848 115938
rect 356796 115874 356848 115880
rect 358096 98666 358124 309130
rect 358740 274650 358768 364958
rect 358832 296002 358860 538319
rect 359476 536110 359504 702578
rect 372620 547936 372672 547942
rect 372620 547878 372672 547884
rect 361856 546508 361908 546514
rect 361856 546450 361908 546456
rect 360476 539708 360528 539714
rect 360476 539650 360528 539656
rect 360200 538348 360252 538354
rect 360200 538290 360252 538296
rect 359464 536104 359516 536110
rect 359464 536046 359516 536052
rect 358910 497856 358966 497865
rect 358910 497791 358966 497800
rect 358820 295996 358872 296002
rect 358820 295938 358872 295944
rect 358728 274644 358780 274650
rect 358728 274586 358780 274592
rect 358740 273290 358768 274586
rect 358728 273284 358780 273290
rect 358728 273226 358780 273232
rect 358924 272542 358952 497791
rect 359002 463312 359058 463321
rect 359002 463247 359058 463256
rect 359016 355366 359044 463247
rect 359094 396944 359150 396953
rect 359094 396879 359150 396888
rect 359108 365702 359136 396879
rect 359096 365696 359148 365702
rect 359096 365638 359148 365644
rect 359004 355360 359056 355366
rect 359004 355302 359056 355308
rect 360212 320890 360240 538290
rect 360292 509720 360344 509726
rect 360292 509662 360344 509668
rect 360200 320884 360252 320890
rect 360200 320826 360252 320832
rect 360304 316742 360332 509662
rect 360384 436144 360436 436150
rect 360384 436086 360436 436092
rect 360292 316736 360344 316742
rect 360292 316678 360344 316684
rect 359462 308408 359518 308417
rect 359462 308343 359518 308352
rect 358912 272536 358964 272542
rect 358912 272478 358964 272484
rect 358176 254584 358228 254590
rect 358176 254526 358228 254532
rect 358188 133210 358216 254526
rect 358176 133204 358228 133210
rect 358176 133146 358228 133152
rect 359476 111110 359504 308343
rect 360396 256018 360424 436086
rect 360488 371278 360516 539650
rect 361672 418192 361724 418198
rect 361672 418134 361724 418140
rect 361580 379568 361632 379574
rect 361580 379510 361632 379516
rect 360476 371272 360528 371278
rect 360476 371214 360528 371220
rect 361592 362234 361620 379510
rect 361684 369170 361712 418134
rect 361764 398880 361816 398886
rect 361764 398822 361816 398828
rect 361672 369164 361724 369170
rect 361672 369106 361724 369112
rect 361776 364993 361804 398822
rect 361868 377369 361896 546450
rect 363052 545216 363104 545222
rect 363052 545158 363104 545164
rect 362958 538248 363014 538257
rect 362958 538183 363014 538192
rect 361854 377360 361910 377369
rect 361854 377295 361910 377304
rect 361762 364984 361818 364993
rect 361762 364919 361818 364928
rect 361580 362228 361632 362234
rect 361580 362170 361632 362176
rect 360844 305108 360896 305114
rect 360844 305050 360896 305056
rect 360384 256012 360436 256018
rect 360384 255954 360436 255960
rect 360856 118590 360884 305050
rect 362972 293282 363000 538183
rect 363064 362302 363092 545158
rect 364432 545148 364484 545154
rect 364432 545090 364484 545096
rect 364340 481704 364392 481710
rect 364340 481646 364392 481652
rect 363236 455456 363288 455462
rect 363236 455398 363288 455404
rect 363144 403504 363196 403510
rect 363144 403446 363196 403452
rect 363052 362296 363104 362302
rect 363052 362238 363104 362244
rect 362960 293276 363012 293282
rect 362960 293218 363012 293224
rect 361486 245712 361542 245721
rect 361486 245647 361542 245656
rect 360844 118584 360896 118590
rect 360844 118526 360896 118532
rect 359556 111852 359608 111858
rect 359556 111794 359608 111800
rect 359464 111104 359516 111110
rect 359464 111046 359516 111052
rect 358084 98660 358136 98666
rect 358084 98602 358136 98608
rect 357440 89004 357492 89010
rect 357440 88946 357492 88952
rect 356704 7608 356756 7614
rect 356704 7550 356756 7556
rect 352562 4040 352618 4049
rect 352562 3975 352618 3984
rect 351642 3904 351698 3913
rect 351642 3839 351698 3848
rect 351656 3670 351684 3839
rect 351184 3664 351236 3670
rect 351184 3606 351236 3612
rect 351644 3664 351696 3670
rect 351644 3606 351696 3612
rect 349252 3460 349304 3466
rect 349252 3402 349304 3408
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 348252 462 348464 490
rect 349264 480 349292 3402
rect 350448 2100 350500 2106
rect 350448 2042 350500 2048
rect 350460 480 350488 2042
rect 351656 480 351684 3606
rect 357452 3466 357480 88946
rect 359464 82136 359516 82142
rect 359464 82078 359516 82084
rect 357440 3460 357492 3466
rect 357440 3402 357492 3408
rect 359476 3369 359504 82078
rect 359568 60722 359596 111794
rect 360844 109744 360896 109750
rect 360844 109686 360896 109692
rect 359556 60716 359608 60722
rect 359556 60658 359608 60664
rect 360856 14550 360884 109686
rect 361500 96529 361528 245647
rect 363156 245002 363184 403446
rect 363248 370705 363276 455398
rect 363234 370696 363290 370705
rect 363234 370631 363290 370640
rect 363604 273284 363656 273290
rect 363604 273226 363656 273232
rect 363144 244996 363196 245002
rect 363144 244938 363196 244944
rect 363616 134570 363644 273226
rect 364352 269793 364380 481646
rect 364444 367878 364472 545090
rect 365720 543856 365772 543862
rect 365720 543798 365772 543804
rect 364524 405748 364576 405754
rect 364524 405690 364576 405696
rect 364432 367872 364484 367878
rect 364432 367814 364484 367820
rect 364536 354006 364564 405690
rect 365732 367810 365760 543798
rect 367284 542496 367336 542502
rect 367284 542438 367336 542444
rect 367192 477556 367244 477562
rect 367192 477498 367244 477504
rect 365904 449200 365956 449206
rect 365904 449142 365956 449148
rect 365812 416832 365864 416838
rect 365812 416774 365864 416780
rect 365720 367804 365772 367810
rect 365720 367746 365772 367752
rect 364524 354000 364576 354006
rect 364524 353942 364576 353948
rect 364338 269784 364394 269793
rect 364338 269719 364394 269728
rect 365824 250510 365852 416774
rect 365916 372609 365944 449142
rect 367100 440292 367152 440298
rect 367100 440234 367152 440240
rect 365996 414044 366048 414050
rect 365996 413986 366048 413992
rect 366008 376009 366036 413986
rect 365994 376000 366050 376009
rect 365994 375935 366050 375944
rect 365902 372600 365958 372609
rect 365902 372535 365958 372544
rect 365812 250504 365864 250510
rect 365812 250446 365864 250452
rect 363694 226944 363750 226953
rect 363694 226879 363750 226888
rect 363604 134564 363656 134570
rect 363604 134506 363656 134512
rect 363604 127016 363656 127022
rect 363604 126958 363656 126964
rect 361486 96520 361542 96529
rect 361486 96455 361542 96464
rect 363616 17950 363644 126958
rect 363708 115258 363736 226879
rect 363696 115252 363748 115258
rect 363696 115194 363748 115200
rect 367112 113150 367140 440234
rect 367204 267034 367232 477498
rect 367296 366382 367324 542438
rect 371240 528624 371292 528630
rect 371240 528566 371292 528572
rect 369860 502376 369912 502382
rect 369860 502318 369912 502324
rect 368572 470620 368624 470626
rect 368572 470562 368624 470568
rect 368480 445800 368532 445806
rect 368480 445742 368532 445748
rect 367376 408536 367428 408542
rect 367376 408478 367428 408484
rect 367284 366376 367336 366382
rect 367284 366318 367336 366324
rect 367388 341465 367416 408478
rect 367374 341456 367430 341465
rect 367374 341391 367430 341400
rect 367742 284880 367798 284889
rect 367742 284815 367798 284824
rect 367192 267028 367244 267034
rect 367192 266970 367244 266976
rect 367100 113144 367152 113150
rect 367100 113086 367152 113092
rect 367756 101289 367784 284815
rect 368492 258806 368520 445742
rect 368584 366353 368612 470562
rect 368676 393417 368704 393443
rect 368662 393408 368718 393417
rect 368662 393343 368664 393352
rect 368716 393343 368718 393352
rect 368664 393314 368716 393320
rect 368676 370569 368704 393314
rect 368662 370560 368718 370569
rect 368662 370495 368718 370504
rect 368570 366344 368626 366353
rect 368570 366279 368626 366288
rect 369872 289134 369900 502318
rect 370044 433356 370096 433362
rect 370044 433298 370096 433304
rect 369952 426488 370004 426494
rect 369952 426430 370004 426436
rect 369860 289128 369912 289134
rect 369860 289070 369912 289076
rect 368480 258800 368532 258806
rect 368480 258742 368532 258748
rect 369964 253230 369992 426430
rect 370056 365022 370084 433298
rect 370044 365016 370096 365022
rect 370044 364958 370096 364964
rect 371252 331226 371280 528566
rect 371332 430636 371384 430642
rect 371332 430578 371384 430584
rect 371240 331220 371292 331226
rect 371240 331162 371292 331168
rect 370504 273964 370556 273970
rect 370504 273906 370556 273912
rect 369952 253224 370004 253230
rect 369952 253166 370004 253172
rect 370516 166326 370544 273906
rect 371344 253298 371372 430578
rect 371424 420980 371476 420986
rect 371424 420922 371476 420928
rect 371436 371929 371464 420922
rect 371422 371920 371478 371929
rect 371422 371855 371478 371864
rect 371884 265668 371936 265674
rect 371884 265610 371936 265616
rect 371332 253292 371384 253298
rect 371332 253234 371384 253240
rect 370596 202156 370648 202162
rect 370596 202098 370648 202104
rect 370504 166320 370556 166326
rect 370504 166262 370556 166268
rect 370504 129736 370556 129742
rect 370504 129678 370556 129684
rect 367836 107704 367888 107710
rect 367836 107646 367888 107652
rect 367742 101280 367798 101289
rect 367742 101215 367798 101224
rect 363604 17944 363656 17950
rect 363604 17886 363656 17892
rect 367848 16590 367876 107646
rect 370516 18698 370544 129678
rect 370608 95198 370636 202098
rect 371896 132462 371924 265610
rect 371974 229120 372030 229129
rect 371974 229055 372030 229064
rect 371988 170406 372016 229055
rect 371976 170400 372028 170406
rect 371976 170342 372028 170348
rect 371976 163532 372028 163538
rect 371976 163474 372028 163480
rect 371884 132456 371936 132462
rect 371884 132398 371936 132404
rect 371988 105602 372016 163474
rect 372632 129742 372660 547878
rect 376852 543788 376904 543794
rect 376852 543730 376904 543736
rect 376760 527196 376812 527202
rect 376760 527138 376812 527144
rect 375472 524476 375524 524482
rect 375472 524418 375524 524424
rect 374736 516180 374788 516186
rect 374736 516122 374788 516128
rect 374092 459604 374144 459610
rect 374092 459546 374144 459552
rect 372712 443012 372764 443018
rect 372712 442954 372764 442960
rect 372724 258738 372752 442954
rect 374000 411324 374052 411330
rect 374000 411266 374052 411272
rect 374012 278050 374040 411266
rect 374104 329798 374132 459546
rect 374092 329792 374144 329798
rect 374092 329734 374144 329740
rect 374748 329118 374776 516122
rect 375288 460216 375340 460222
rect 375288 460158 375340 460164
rect 375300 459610 375328 460158
rect 375288 459604 375340 459610
rect 375288 459546 375340 459552
rect 375380 449948 375432 449954
rect 375380 449890 375432 449896
rect 374736 329112 374788 329118
rect 374736 329054 374788 329060
rect 374642 328808 374698 328817
rect 374642 328743 374698 328752
rect 374000 278044 374052 278050
rect 374000 277986 374052 277992
rect 372712 258732 372764 258738
rect 372712 258674 372764 258680
rect 374656 142118 374684 328743
rect 375392 260166 375420 449890
rect 375484 342922 375512 524418
rect 375472 342916 375524 342922
rect 375472 342858 375524 342864
rect 376024 278044 376076 278050
rect 376024 277986 376076 277992
rect 375380 260160 375432 260166
rect 375380 260102 375432 260108
rect 374734 208992 374790 209001
rect 374734 208927 374790 208936
rect 374748 151094 374776 208927
rect 374736 151088 374788 151094
rect 374736 151030 374788 151036
rect 374644 142112 374696 142118
rect 374644 142054 374696 142060
rect 374736 135312 374788 135318
rect 374736 135254 374788 135260
rect 372620 129736 372672 129742
rect 372620 129678 372672 129684
rect 374748 122806 374776 135254
rect 374736 122800 374788 122806
rect 374736 122742 374788 122748
rect 374644 121508 374696 121514
rect 374644 121450 374696 121456
rect 371976 105596 372028 105602
rect 371976 105538 372028 105544
rect 370596 95192 370648 95198
rect 370596 95134 370648 95140
rect 374656 27606 374684 121450
rect 376036 99346 376064 277986
rect 376772 142118 376800 527138
rect 376864 273222 376892 543730
rect 378140 480276 378192 480282
rect 378140 480218 378192 480224
rect 376944 465112 376996 465118
rect 376944 465054 376996 465060
rect 376956 356726 376984 465054
rect 376944 356720 376996 356726
rect 376944 356662 376996 356668
rect 378152 351121 378180 480218
rect 378796 375358 378824 702646
rect 382924 700324 382976 700330
rect 382924 700266 382976 700272
rect 380990 541240 381046 541249
rect 380990 541175 381046 541184
rect 380898 535664 380954 535673
rect 380898 535599 380954 535608
rect 379520 420232 379572 420238
rect 379520 420174 379572 420180
rect 378784 375352 378836 375358
rect 378784 375294 378836 375300
rect 378874 374640 378930 374649
rect 378874 374575 378930 374584
rect 378138 351112 378194 351121
rect 378138 351047 378194 351056
rect 376852 273216 376904 273222
rect 376852 273158 376904 273164
rect 378782 266248 378838 266257
rect 378782 266183 378838 266192
rect 378796 262886 378824 266183
rect 378784 262880 378836 262886
rect 378784 262822 378836 262828
rect 377404 247104 377456 247110
rect 377404 247046 377456 247052
rect 376760 142112 376812 142118
rect 376760 142054 376812 142060
rect 376772 134473 376800 142054
rect 376758 134464 376814 134473
rect 376758 134399 376814 134408
rect 377416 102785 377444 247046
rect 378796 120086 378824 262822
rect 378888 162178 378916 374575
rect 378876 162172 378928 162178
rect 378876 162114 378928 162120
rect 378876 133952 378928 133958
rect 378876 133894 378928 133900
rect 378784 120080 378836 120086
rect 378784 120022 378836 120028
rect 377496 111920 377548 111926
rect 377496 111862 377548 111868
rect 377402 102776 377458 102785
rect 377402 102711 377458 102720
rect 376024 99340 376076 99346
rect 376024 99282 376076 99288
rect 376024 93220 376076 93226
rect 376024 93162 376076 93168
rect 374644 27600 374696 27606
rect 374644 27542 374696 27548
rect 370504 18692 370556 18698
rect 370504 18634 370556 18640
rect 367836 16584 367888 16590
rect 367836 16526 367888 16532
rect 360844 14544 360896 14550
rect 360844 14486 360896 14492
rect 376036 3913 376064 93162
rect 377508 11014 377536 111862
rect 377496 11008 377548 11014
rect 377496 10950 377548 10956
rect 378888 6186 378916 133894
rect 379532 88262 379560 420174
rect 380164 211812 380216 211818
rect 380164 211754 380216 211760
rect 380176 163538 380204 211754
rect 380912 194585 380940 535599
rect 381004 246265 381032 541175
rect 382280 427848 382332 427854
rect 382280 427790 382332 427796
rect 382292 294642 382320 427790
rect 382936 376038 382964 700266
rect 393964 539640 394016 539646
rect 393964 539582 394016 539588
rect 388444 519580 388496 519586
rect 388444 519522 388496 519528
rect 385040 486464 385092 486470
rect 385040 486406 385092 486412
rect 382924 376032 382976 376038
rect 382924 375974 382976 375980
rect 382280 294636 382332 294642
rect 382280 294578 382332 294584
rect 380990 246256 381046 246265
rect 380990 246191 381046 246200
rect 380898 194576 380954 194585
rect 380898 194511 380954 194520
rect 380164 163532 380216 163538
rect 380164 163474 380216 163480
rect 380912 139369 380940 194511
rect 382936 145654 382964 375974
rect 385052 271862 385080 486406
rect 385132 386436 385184 386442
rect 385132 386378 385184 386384
rect 385144 372745 385172 386378
rect 385130 372736 385186 372745
rect 385130 372671 385186 372680
rect 385682 372736 385738 372745
rect 385682 372671 385738 372680
rect 385040 271856 385092 271862
rect 385040 271798 385092 271804
rect 383016 257372 383068 257378
rect 383016 257314 383068 257320
rect 382924 145648 382976 145654
rect 382924 145590 382976 145596
rect 381544 142180 381596 142186
rect 381544 142122 381596 142128
rect 380898 139360 380954 139369
rect 380898 139295 380954 139304
rect 380912 138689 380940 139295
rect 380898 138680 380954 138689
rect 380898 138615 380954 138624
rect 379520 88256 379572 88262
rect 379520 88198 379572 88204
rect 379532 87650 379560 88198
rect 379520 87644 379572 87650
rect 379520 87586 379572 87592
rect 381556 55894 381584 142122
rect 381636 134564 381688 134570
rect 381636 134506 381688 134512
rect 381648 107574 381676 134506
rect 381636 107568 381688 107574
rect 381636 107510 381688 107516
rect 383028 104174 383056 257314
rect 384304 238060 384356 238066
rect 384304 238002 384356 238008
rect 383108 140888 383160 140894
rect 383108 140830 383160 140836
rect 383016 104168 383068 104174
rect 382922 104136 382978 104145
rect 383016 104110 383068 104116
rect 382922 104071 382978 104080
rect 381636 98660 381688 98666
rect 381636 98602 381688 98608
rect 381648 91050 381676 98602
rect 381636 91044 381688 91050
rect 381636 90986 381688 90992
rect 381544 55888 381596 55894
rect 381544 55830 381596 55836
rect 381636 55888 381688 55894
rect 381636 55830 381688 55836
rect 378876 6180 378928 6186
rect 378876 6122 378928 6128
rect 376022 3904 376078 3913
rect 376022 3839 376078 3848
rect 359462 3360 359518 3369
rect 359462 3295 359518 3304
rect 381648 2106 381676 55830
rect 382936 14482 382964 104071
rect 383120 69698 383148 140830
rect 384316 99278 384344 238002
rect 385696 99657 385724 372671
rect 387064 221468 387116 221474
rect 387064 221410 387116 221416
rect 385776 153876 385828 153882
rect 385776 153818 385828 153824
rect 385788 113830 385816 153818
rect 385776 113824 385828 113830
rect 385776 113766 385828 113772
rect 385776 109064 385828 109070
rect 385776 109006 385828 109012
rect 385682 99648 385738 99657
rect 385682 99583 385738 99592
rect 384304 99272 384356 99278
rect 384304 99214 384356 99220
rect 383108 69692 383160 69698
rect 383108 69634 383160 69640
rect 382924 14476 382976 14482
rect 382924 14418 382976 14424
rect 385788 12374 385816 109006
rect 387076 99521 387104 221410
rect 387156 146328 387208 146334
rect 387156 146270 387208 146276
rect 387168 135930 387196 146270
rect 387156 135924 387208 135930
rect 387156 135866 387208 135872
rect 387062 99512 387118 99521
rect 387062 99447 387118 99456
rect 388456 99249 388484 519522
rect 389180 472048 389232 472054
rect 389180 471990 389232 471996
rect 389192 294001 389220 471990
rect 392584 438932 392636 438938
rect 392584 438874 392636 438880
rect 389822 317520 389878 317529
rect 389822 317455 389878 317464
rect 389178 293992 389234 294001
rect 389178 293927 389234 293936
rect 389192 291854 389220 293927
rect 389180 291848 389232 291854
rect 389180 291790 389232 291796
rect 388536 135380 388588 135386
rect 388536 135322 388588 135328
rect 388442 99240 388498 99249
rect 388442 99175 388498 99184
rect 388548 31074 388576 135322
rect 389836 96558 389864 317455
rect 389916 297424 389968 297430
rect 389916 297366 389968 297372
rect 389928 153882 389956 297366
rect 391202 198112 391258 198121
rect 391202 198047 391258 198056
rect 391216 167686 391244 198047
rect 391204 167680 391256 167686
rect 391204 167622 391256 167628
rect 389916 153876 389968 153882
rect 389916 153818 389968 153824
rect 391204 133204 391256 133210
rect 391204 133146 391256 133152
rect 389916 129804 389968 129810
rect 389916 129746 389968 129752
rect 389824 96552 389876 96558
rect 389824 96494 389876 96500
rect 388536 31068 388588 31074
rect 388536 31010 388588 31016
rect 389928 22778 389956 129746
rect 391216 117298 391244 133146
rect 391204 117292 391256 117298
rect 391204 117234 391256 117240
rect 392596 99793 392624 438874
rect 392674 310584 392730 310593
rect 392674 310519 392730 310528
rect 392688 125526 392716 310519
rect 392768 132524 392820 132530
rect 392768 132466 392820 132472
rect 392676 125520 392728 125526
rect 392676 125462 392728 125468
rect 392582 99784 392638 99793
rect 392582 99719 392638 99728
rect 391940 97300 391992 97306
rect 391940 97242 391992 97248
rect 391952 95130 391980 97242
rect 391940 95124 391992 95130
rect 391940 95066 391992 95072
rect 392780 28286 392808 132466
rect 393976 95169 394004 539582
rect 395988 520940 396040 520946
rect 395988 520882 396040 520888
rect 396000 520334 396028 520882
rect 395988 520328 396040 520334
rect 395988 520270 396040 520276
rect 395344 276684 395396 276690
rect 395344 276626 395396 276632
rect 394056 216708 394108 216714
rect 394056 216650 394108 216656
rect 394068 97753 394096 216650
rect 395356 99414 395384 276626
rect 395436 151088 395488 151094
rect 395436 151030 395488 151036
rect 395448 139398 395476 151030
rect 396000 145625 396028 520270
rect 412652 494018 412680 703582
rect 413480 703474 413508 703582
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 413664 703474 413692 703520
rect 413480 703446 413692 703474
rect 429856 700330 429884 703520
rect 462332 702710 462360 703520
rect 478524 702914 478552 703520
rect 478512 702908 478564 702914
rect 478512 702850 478564 702856
rect 494808 702846 494836 703520
rect 494796 702840 494848 702846
rect 494796 702782 494848 702788
rect 462320 702704 462372 702710
rect 462320 702646 462372 702652
rect 527192 702506 527220 703520
rect 543476 702642 543504 703520
rect 543464 702636 543516 702642
rect 543464 702578 543516 702584
rect 559668 702574 559696 703520
rect 559656 702568 559708 702574
rect 559656 702510 559708 702516
rect 527180 702500 527232 702506
rect 527180 702442 527232 702448
rect 429844 700324 429896 700330
rect 429844 700266 429896 700272
rect 582654 697232 582710 697241
rect 582654 697167 582710 697176
rect 582562 683904 582618 683913
rect 582562 683839 582618 683848
rect 582378 670712 582434 670721
rect 582378 670647 582434 670656
rect 580354 554840 580410 554849
rect 580354 554775 580410 554784
rect 579896 538212 579948 538218
rect 579896 538154 579948 538160
rect 579908 537849 579936 538154
rect 579894 537840 579950 537849
rect 579894 537775 579950 537784
rect 580264 535492 580316 535498
rect 580264 535434 580316 535440
rect 427820 534812 427872 534818
rect 427820 534754 427872 534760
rect 414664 505164 414716 505170
rect 414664 505106 414716 505112
rect 412640 494012 412692 494018
rect 412640 493954 412692 493960
rect 398840 452668 398892 452674
rect 398840 452610 398892 452616
rect 397458 188320 397514 188329
rect 397458 188255 397514 188264
rect 395986 145616 396042 145625
rect 395986 145551 396042 145560
rect 396722 142352 396778 142361
rect 396722 142287 396778 142296
rect 395526 142216 395582 142225
rect 395526 142151 395582 142160
rect 395436 139392 395488 139398
rect 395436 139334 395488 139340
rect 395434 134464 395490 134473
rect 395434 134399 395490 134408
rect 395448 132705 395476 134399
rect 395434 132696 395490 132705
rect 395434 132631 395490 132640
rect 395448 119406 395476 132631
rect 395436 119400 395488 119406
rect 395436 119342 395488 119348
rect 395436 100768 395488 100774
rect 395436 100710 395488 100716
rect 395344 99408 395396 99414
rect 395344 99350 395396 99356
rect 394054 97744 394110 97753
rect 394054 97679 394110 97688
rect 394148 96960 394200 96966
rect 394148 96902 394200 96908
rect 393962 95160 394018 95169
rect 393962 95095 394018 95104
rect 393318 94480 393374 94489
rect 393318 94415 393374 94424
rect 393332 88233 393360 94415
rect 393318 88224 393374 88233
rect 393318 88159 393374 88168
rect 392768 28280 392820 28286
rect 392768 28222 392820 28228
rect 389916 22772 389968 22778
rect 389916 22714 389968 22720
rect 385776 12368 385828 12374
rect 385776 12310 385828 12316
rect 394160 8294 394188 96902
rect 395448 35902 395476 100710
rect 395540 93158 395568 142151
rect 395620 136672 395672 136678
rect 395620 136614 395672 136620
rect 395632 131782 395660 136614
rect 395620 131776 395672 131782
rect 395620 131718 395672 131724
rect 395528 93152 395580 93158
rect 395528 93094 395580 93100
rect 395436 35896 395488 35902
rect 395436 35838 395488 35844
rect 396736 20670 396764 142287
rect 397366 115832 397422 115841
rect 397366 115767 397422 115776
rect 397380 115258 397408 115767
rect 397368 115252 397420 115258
rect 397368 115194 397420 115200
rect 397380 86290 397408 115194
rect 397472 111874 397500 188255
rect 398748 156664 398800 156670
rect 398748 156606 398800 156612
rect 398656 155236 398708 155242
rect 398656 155178 398708 155184
rect 398472 146940 398524 146946
rect 398472 146882 398524 146888
rect 397552 139392 397604 139398
rect 397550 139360 397552 139369
rect 397604 139360 397606 139369
rect 397550 139295 397606 139304
rect 397918 137320 397974 137329
rect 397918 137255 397974 137264
rect 397932 136678 397960 137255
rect 397920 136672 397972 136678
rect 397920 136614 397972 136620
rect 397642 136232 397698 136241
rect 397642 136167 397698 136176
rect 397550 135416 397606 135425
rect 397656 135386 397684 136167
rect 397550 135351 397606 135360
rect 397644 135380 397696 135386
rect 397564 135318 397592 135351
rect 397644 135322 397696 135328
rect 397552 135312 397604 135318
rect 397552 135254 397604 135260
rect 397642 134736 397698 134745
rect 397642 134671 397698 134680
rect 397656 133958 397684 134671
rect 397644 133952 397696 133958
rect 397644 133894 397696 133900
rect 397550 133512 397606 133521
rect 397550 133447 397606 133456
rect 397564 132530 397592 133447
rect 397552 132524 397604 132530
rect 397552 132466 397604 132472
rect 398484 132462 398512 146882
rect 398472 132456 398524 132462
rect 398472 132398 398524 132404
rect 398484 131753 398512 132398
rect 398470 131744 398526 131753
rect 398470 131679 398526 131688
rect 397552 129736 397604 129742
rect 398668 129713 398696 155178
rect 397552 129678 397604 129684
rect 398654 129704 398710 129713
rect 397564 129033 397592 129678
rect 398654 129639 398710 129648
rect 398196 129056 398248 129062
rect 397550 129024 397606 129033
rect 398196 128998 398248 129004
rect 397550 128959 397606 128968
rect 397552 128308 397604 128314
rect 397552 128250 397604 128256
rect 397564 128217 397592 128250
rect 397550 128208 397606 128217
rect 397550 128143 397606 128152
rect 397550 127120 397606 127129
rect 397550 127055 397606 127064
rect 397564 127022 397592 127055
rect 397552 127016 397604 127022
rect 397552 126958 397604 126964
rect 397550 126304 397606 126313
rect 397550 126239 397552 126248
rect 397604 126239 397606 126248
rect 397552 126210 397604 126216
rect 397644 125588 397696 125594
rect 397644 125530 397696 125536
rect 397552 125520 397604 125526
rect 397552 125462 397604 125468
rect 397564 125225 397592 125462
rect 397550 125216 397606 125225
rect 397550 125151 397606 125160
rect 397656 124409 397684 125530
rect 397642 124400 397698 124409
rect 397642 124335 397698 124344
rect 397552 124160 397604 124166
rect 397552 124102 397604 124108
rect 397564 123321 397592 124102
rect 397550 123312 397606 123321
rect 397550 123247 397606 123256
rect 397550 122360 397606 122369
rect 397550 122295 397606 122304
rect 397564 121514 397592 122295
rect 397552 121508 397604 121514
rect 397552 121450 397604 121456
rect 398208 121417 398236 128998
rect 398760 121446 398788 156606
rect 398852 130937 398880 452610
rect 406384 401668 406436 401674
rect 406384 401610 406436 401616
rect 403624 383716 403676 383722
rect 403624 383658 403676 383664
rect 400220 349172 400272 349178
rect 400220 349114 400272 349120
rect 398932 231124 398984 231130
rect 398932 231066 398984 231072
rect 398944 151814 398972 231066
rect 398944 151786 399616 151814
rect 399588 139890 399616 151786
rect 400232 140350 400260 349114
rect 401600 291236 401652 291242
rect 401600 291178 401652 291184
rect 400770 142216 400826 142225
rect 400770 142151 400826 142160
rect 400220 140344 400272 140350
rect 400220 140286 400272 140292
rect 399588 139862 400062 139890
rect 400784 139876 400812 142151
rect 401324 140344 401376 140350
rect 401324 140286 401376 140292
rect 401336 139890 401364 140286
rect 401612 139890 401640 291178
rect 403072 228404 403124 228410
rect 403072 228346 403124 228352
rect 401690 180840 401746 180849
rect 401690 180775 401746 180784
rect 401704 151814 401732 180775
rect 403084 151814 403112 228346
rect 401704 151786 402192 151814
rect 403084 151786 403480 151814
rect 402164 139890 402192 151786
rect 403452 139890 403480 151786
rect 403636 144226 403664 383658
rect 405738 206408 405794 206417
rect 405738 206343 405794 206352
rect 404358 184240 404414 184249
rect 404358 184175 404414 184184
rect 404372 151814 404400 184175
rect 404372 151786 404492 151814
rect 403624 144220 403676 144226
rect 403624 144162 403676 144168
rect 401336 139876 401548 139890
rect 401350 139862 401548 139876
rect 401612 139862 401902 139890
rect 402164 139862 402638 139890
rect 403452 139862 403926 139890
rect 401520 139602 401548 139862
rect 401508 139596 401560 139602
rect 401508 139538 401560 139544
rect 402992 139466 403190 139482
rect 399484 139460 399536 139466
rect 399484 139402 399536 139408
rect 402980 139460 403190 139466
rect 403032 139454 403190 139460
rect 402980 139402 403032 139408
rect 398838 130928 398894 130937
rect 398838 130863 398894 130872
rect 398852 129810 398880 130863
rect 398840 129804 398892 129810
rect 398840 129746 398892 129752
rect 398748 121440 398800 121446
rect 398194 121408 398250 121417
rect 398748 121382 398800 121388
rect 398194 121343 398250 121352
rect 398760 120601 398788 121382
rect 398746 120592 398802 120601
rect 398746 120527 398802 120536
rect 397552 120080 397604 120086
rect 397552 120022 397604 120028
rect 397564 119785 397592 120022
rect 397550 119776 397606 119785
rect 397550 119711 397606 119720
rect 397644 118652 397696 118658
rect 397644 118594 397696 118600
rect 397552 118584 397604 118590
rect 397550 118552 397552 118561
rect 397604 118552 397606 118561
rect 397550 118487 397606 118496
rect 397656 117881 397684 118594
rect 397642 117872 397698 117881
rect 397642 117807 397698 117816
rect 397552 117292 397604 117298
rect 397552 117234 397604 117240
rect 397564 116793 397592 117234
rect 397550 116784 397606 116793
rect 397550 116719 397606 116728
rect 397552 115932 397604 115938
rect 397552 115874 397604 115880
rect 397564 114889 397592 115874
rect 397550 114880 397606 114889
rect 397550 114815 397606 114824
rect 397552 114504 397604 114510
rect 397552 114446 397604 114452
rect 397564 114073 397592 114446
rect 397550 114064 397606 114073
rect 397550 113999 397606 114008
rect 397920 113824 397972 113830
rect 397920 113766 397972 113772
rect 397932 113174 397960 113766
rect 397932 113146 398144 113174
rect 397642 113112 397698 113121
rect 397642 113047 397698 113056
rect 397656 111926 397684 113047
rect 397734 112024 397790 112033
rect 397734 111959 397790 111968
rect 397644 111920 397696 111926
rect 397472 111846 397592 111874
rect 397644 111862 397696 111868
rect 397748 111858 397776 111959
rect 397460 111784 397512 111790
rect 397460 111726 397512 111732
rect 397472 111353 397500 111726
rect 397458 111344 397514 111353
rect 397458 111279 397514 111288
rect 397564 110265 397592 111846
rect 397736 111852 397788 111858
rect 397736 111794 397788 111800
rect 397644 111104 397696 111110
rect 397644 111046 397696 111052
rect 397550 110256 397606 110265
rect 397550 110191 397606 110200
rect 397564 109750 397592 110191
rect 397552 109744 397604 109750
rect 397552 109686 397604 109692
rect 397458 109304 397514 109313
rect 397458 109239 397514 109248
rect 397472 109070 397500 109239
rect 397460 109064 397512 109070
rect 397460 109006 397512 109012
rect 397458 108216 397514 108225
rect 397458 108151 397514 108160
rect 397472 107710 397500 108151
rect 397460 107704 397512 107710
rect 397460 107646 397512 107652
rect 397552 107636 397604 107642
rect 397552 107578 397604 107584
rect 397460 107568 397512 107574
rect 397564 107545 397592 107578
rect 397460 107510 397512 107516
rect 397550 107536 397606 107545
rect 397472 106729 397500 107510
rect 397550 107471 397606 107480
rect 397458 106720 397514 106729
rect 397458 106655 397514 106664
rect 397460 106276 397512 106282
rect 397460 106218 397512 106224
rect 397472 105641 397500 106218
rect 397458 105632 397514 105641
rect 397458 105567 397514 105576
rect 397460 104848 397512 104854
rect 397458 104816 397460 104825
rect 397512 104816 397514 104825
rect 397458 104751 397514 104760
rect 397656 104145 397684 111046
rect 397642 104136 397698 104145
rect 397642 104071 397698 104080
rect 397460 103488 397512 103494
rect 397460 103430 397512 103436
rect 397472 102921 397500 103430
rect 397458 102912 397514 102921
rect 397458 102847 397514 102856
rect 397458 101688 397514 101697
rect 397458 101623 397514 101632
rect 397472 99385 397500 101623
rect 397550 100872 397606 100881
rect 397550 100807 397606 100816
rect 397564 100774 397592 100807
rect 397552 100768 397604 100774
rect 397552 100710 397604 100716
rect 397458 99376 397514 99385
rect 397458 99311 397514 99320
rect 398116 93838 398144 113146
rect 398196 108316 398248 108322
rect 398196 108258 398248 108264
rect 398208 100774 398236 108258
rect 398196 100768 398248 100774
rect 398196 100710 398248 100716
rect 398840 94172 398892 94178
rect 398840 94114 398892 94120
rect 398104 93832 398156 93838
rect 398104 93774 398156 93780
rect 397368 86284 397420 86290
rect 397368 86226 397420 86232
rect 398852 72486 398880 94114
rect 398840 72480 398892 72486
rect 398840 72422 398892 72428
rect 399496 39273 399524 139402
rect 399852 139392 399904 139398
rect 399852 139334 399904 139340
rect 404084 139392 404136 139398
rect 404464 139346 404492 151786
rect 405188 142180 405240 142186
rect 405188 142122 405240 142128
rect 405200 139876 405228 142122
rect 405752 140758 405780 206343
rect 405830 185600 405886 185609
rect 405830 185535 405886 185544
rect 405844 151814 405872 185535
rect 406396 164898 406424 401610
rect 413284 363724 413336 363730
rect 413284 363666 413336 363672
rect 409880 329112 409932 329118
rect 409880 329054 409932 329060
rect 407120 291848 407172 291854
rect 407120 291790 407172 291796
rect 406384 164892 406436 164898
rect 406384 164834 406436 164840
rect 405844 151786 406332 151814
rect 405922 145616 405978 145625
rect 405922 145551 405978 145560
rect 405740 140752 405792 140758
rect 405740 140694 405792 140700
rect 405936 139890 405964 145551
rect 406304 142497 406332 151786
rect 406290 142488 406346 142497
rect 406290 142423 406346 142432
rect 405766 139862 405964 139890
rect 406304 139876 406332 142423
rect 406660 140752 406712 140758
rect 406660 140694 406712 140700
rect 406672 139890 406700 140694
rect 407132 139890 407160 291790
rect 407210 224224 407266 224233
rect 407210 224159 407266 224168
rect 407224 150482 407252 224159
rect 407212 150476 407264 150482
rect 407212 150418 407264 150424
rect 407224 143546 407252 150418
rect 407672 147688 407724 147694
rect 407672 147630 407724 147636
rect 407212 143540 407264 143546
rect 407212 143482 407264 143488
rect 407684 139890 407712 147630
rect 408868 143540 408920 143546
rect 408868 143482 408920 143488
rect 406672 139862 407054 139890
rect 407132 139862 407606 139890
rect 407684 139862 408342 139890
rect 408880 139876 408908 143482
rect 409892 143449 409920 329054
rect 411904 300892 411956 300898
rect 411904 300834 411956 300840
rect 410524 236700 410576 236706
rect 410524 236642 410576 236648
rect 409972 145580 410024 145586
rect 409972 145522 410024 145528
rect 409878 143440 409934 143449
rect 409878 143375 409934 143384
rect 409604 140820 409656 140826
rect 409604 140762 409656 140768
rect 409616 139876 409644 140762
rect 409984 139890 410012 145522
rect 410536 143546 410564 236642
rect 411916 148442 411944 300834
rect 412638 220144 412694 220153
rect 412638 220079 412694 220088
rect 411994 199336 412050 199345
rect 411994 199271 412050 199280
rect 411904 148436 411956 148442
rect 411904 148378 411956 148384
rect 411442 145616 411498 145625
rect 412008 145586 412036 199271
rect 411442 145551 411498 145560
rect 411996 145580 412048 145586
rect 410524 143540 410576 143546
rect 410524 143482 410576 143488
rect 410890 143440 410946 143449
rect 410890 143375 410946 143384
rect 409984 139862 410182 139890
rect 410904 139876 410932 143375
rect 411456 139876 411484 145551
rect 411996 145522 412048 145528
rect 411996 143540 412048 143546
rect 411996 143482 412048 143488
rect 412008 139876 412036 143482
rect 412652 140758 412680 220079
rect 412732 145648 412784 145654
rect 412732 145590 412784 145596
rect 412640 140752 412692 140758
rect 412640 140694 412692 140700
rect 412744 139876 412772 145590
rect 413296 143478 413324 363666
rect 414676 282266 414704 505106
rect 420920 370524 420972 370530
rect 420920 370466 420972 370472
rect 418802 367160 418858 367169
rect 418802 367095 418858 367104
rect 414664 282260 414716 282266
rect 414664 282202 414716 282208
rect 414756 282192 414808 282198
rect 414756 282134 414808 282140
rect 414020 218748 414072 218754
rect 414020 218690 414072 218696
rect 413284 143472 413336 143478
rect 413284 143414 413336 143420
rect 412916 140752 412968 140758
rect 412916 140694 412968 140700
rect 412928 139890 412956 140694
rect 412928 139862 413310 139890
rect 414032 139876 414060 218690
rect 414112 178696 414164 178702
rect 414112 178638 414164 178644
rect 414124 139890 414152 178638
rect 414204 158024 414256 158030
rect 414204 157966 414256 157972
rect 414216 142154 414244 157966
rect 414768 143546 414796 282134
rect 417424 275324 417476 275330
rect 417424 275266 417476 275272
rect 416778 233336 416834 233345
rect 416778 233271 416834 233280
rect 414756 143540 414808 143546
rect 414756 143482 414808 143488
rect 416412 143540 416464 143546
rect 416412 143482 416464 143488
rect 415860 142860 415912 142866
rect 415860 142802 415912 142808
rect 414216 142126 414888 142154
rect 414860 139890 414888 142126
rect 414124 139862 414598 139890
rect 414860 139862 415334 139890
rect 415872 139876 415900 142802
rect 416424 139876 416452 143482
rect 416792 142866 416820 233271
rect 416780 142860 416832 142866
rect 416780 142802 416832 142808
rect 417148 140888 417200 140894
rect 417148 140830 417200 140836
rect 417160 139876 417188 140830
rect 417436 140078 417464 275266
rect 418252 162172 418304 162178
rect 418252 162114 418304 162120
rect 418264 151814 418292 162114
rect 418264 151786 418568 151814
rect 418436 143472 418488 143478
rect 418436 143414 418488 143420
rect 417424 140072 417476 140078
rect 417424 140014 417476 140020
rect 418448 139876 418476 143414
rect 417332 139664 417384 139670
rect 417384 139612 417726 139618
rect 417332 139606 417726 139612
rect 417344 139590 417726 139606
rect 418540 139482 418568 151786
rect 418816 142186 418844 367095
rect 420184 240780 420236 240786
rect 420184 240722 420236 240728
rect 420196 146266 420224 240722
rect 420276 164892 420328 164898
rect 420276 164834 420328 164840
rect 420184 146260 420236 146266
rect 420184 146202 420236 146208
rect 419724 144220 419776 144226
rect 419724 144162 419776 144168
rect 418804 142180 418856 142186
rect 418804 142122 418856 142128
rect 419736 139618 419764 144162
rect 419906 139632 419962 139641
rect 419736 139604 419906 139618
rect 419750 139590 419906 139604
rect 419906 139567 419962 139576
rect 418710 139496 418766 139505
rect 418540 139454 418710 139482
rect 420288 139482 420316 164834
rect 420932 143449 420960 370466
rect 421564 280832 421616 280838
rect 421564 280774 421616 280780
rect 421576 150414 421604 280774
rect 425702 200832 425758 200841
rect 425702 200767 425758 200776
rect 425060 159384 425112 159390
rect 425060 159326 425112 159332
rect 425072 151814 425100 159326
rect 425072 151786 425560 151814
rect 421104 150408 421156 150414
rect 421104 150350 421156 150356
rect 421564 150408 421616 150414
rect 421564 150350 421616 150356
rect 420918 143440 420974 143449
rect 420918 143375 420974 143384
rect 421116 139890 421144 150350
rect 422944 146260 422996 146266
rect 422944 146202 422996 146208
rect 422392 145580 422444 145586
rect 422392 145522 422444 145528
rect 422114 143440 422170 143449
rect 422114 143375 422170 143384
rect 421116 139862 421590 139890
rect 422128 139876 422156 143375
rect 422404 139890 422432 145522
rect 422956 139890 422984 146202
rect 424692 144220 424744 144226
rect 424692 144162 424744 144168
rect 424140 142180 424192 142186
rect 424140 142122 424192 142128
rect 422404 139862 422878 139890
rect 422956 139862 423430 139890
rect 424152 139876 424180 142122
rect 424704 139876 424732 144162
rect 425428 140888 425480 140894
rect 425428 140830 425480 140836
rect 425440 139876 425468 140830
rect 425532 139890 425560 151786
rect 425716 142186 425744 200767
rect 426438 197976 426494 197985
rect 426438 197911 426494 197920
rect 426452 151814 426480 197911
rect 426452 151786 426572 151814
rect 425796 149728 425848 149734
rect 425796 149670 425848 149676
rect 425704 142180 425756 142186
rect 425704 142122 425756 142128
rect 425808 140894 425836 149670
rect 425796 140888 425848 140894
rect 426544 140865 426572 151786
rect 427832 142361 427860 534754
rect 580276 484673 580304 535434
rect 580368 524521 580396 554775
rect 580354 524512 580410 524521
rect 580354 524447 580410 524456
rect 580262 484664 580318 484673
rect 580262 484599 580318 484608
rect 580262 471472 580318 471481
rect 580262 471407 580318 471416
rect 580276 378049 580304 471407
rect 580354 378448 580410 378457
rect 580354 378383 580410 378392
rect 580262 378040 580318 378049
rect 580262 377975 580318 377984
rect 452660 373312 452712 373318
rect 452660 373254 452712 373260
rect 447140 305040 447192 305046
rect 447140 304982 447192 304988
rect 435364 303680 435416 303686
rect 435364 303622 435416 303628
rect 431960 282260 432012 282266
rect 431960 282202 432012 282208
rect 429198 222864 429254 222873
rect 429198 222799 429254 222808
rect 428462 206272 428518 206281
rect 428462 206207 428518 206216
rect 428476 151814 428504 206207
rect 429212 151814 429240 222799
rect 430578 181384 430634 181393
rect 430578 181319 430634 181328
rect 428476 151786 428596 151814
rect 429212 151786 429976 151814
rect 427818 142352 427874 142361
rect 427818 142287 427874 142296
rect 425796 140830 425848 140836
rect 426530 140856 426586 140865
rect 426530 140791 426586 140800
rect 425532 139862 426006 139890
rect 426544 139876 426572 140791
rect 427832 139876 427860 142287
rect 428568 140826 428596 151786
rect 428556 140820 428608 140826
rect 428556 140762 428608 140768
rect 428568 139876 428596 140762
rect 429948 139890 429976 151786
rect 430592 143546 430620 181319
rect 430672 167680 430724 167686
rect 430672 167622 430724 167628
rect 430580 143540 430632 143546
rect 430580 143482 430632 143488
rect 430684 139890 430712 167622
rect 431316 143540 431368 143546
rect 431316 143482 431368 143488
rect 431328 139890 431356 143482
rect 431972 142225 432000 282202
rect 434718 225040 434774 225049
rect 434718 224975 434774 224984
rect 432052 182844 432104 182850
rect 432052 182786 432104 182792
rect 431958 142216 432014 142225
rect 431958 142151 432014 142160
rect 432064 139890 432092 182786
rect 433984 170400 434036 170406
rect 433984 170342 434036 170348
rect 432970 142216 433026 142225
rect 432970 142151 433026 142160
rect 433524 142180 433576 142186
rect 429948 139862 430422 139890
rect 430684 139862 430974 139890
rect 431328 139862 431710 139890
rect 432064 139862 432262 139890
rect 432984 139876 433012 142151
rect 433524 142122 433576 142128
rect 433536 139876 433564 142122
rect 433996 140049 434024 170342
rect 434732 151814 434760 224975
rect 434732 151786 434944 151814
rect 434076 148436 434128 148442
rect 434076 148378 434128 148384
rect 434088 142186 434116 148378
rect 434076 142180 434128 142186
rect 434076 142122 434128 142128
rect 433982 140040 434038 140049
rect 433982 139975 434038 139984
rect 434088 139890 434116 142122
rect 434916 139890 434944 151786
rect 435376 140865 435404 303622
rect 445760 290012 445812 290018
rect 445760 289954 445812 289960
rect 442998 287192 443054 287201
rect 442998 287127 443054 287136
rect 436284 244928 436336 244934
rect 436284 244870 436336 244876
rect 436190 204368 436246 204377
rect 436190 204303 436246 204312
rect 435362 140856 435418 140865
rect 435362 140791 435418 140800
rect 436204 139890 436232 204303
rect 436296 151814 436324 244870
rect 437480 201544 437532 201550
rect 437480 201486 437532 201492
rect 436296 151786 436968 151814
rect 436652 146328 436704 146334
rect 436652 146270 436704 146276
rect 434088 139862 434286 139890
rect 434916 139862 435390 139890
rect 436126 139862 436232 139890
rect 436664 139876 436692 146270
rect 436940 139890 436968 151786
rect 437492 139890 437520 201486
rect 440238 200696 440294 200705
rect 440238 200631 440294 200640
rect 439872 166320 439924 166326
rect 439872 166262 439924 166268
rect 438952 153876 439004 153882
rect 438952 153818 439004 153824
rect 438964 151814 438992 153818
rect 439884 151814 439912 166262
rect 438964 151786 439360 151814
rect 439884 151786 440004 151814
rect 438676 142860 438728 142866
rect 438676 142802 438728 142808
rect 436940 139862 437414 139890
rect 437492 139862 437966 139890
rect 438688 139876 438716 142802
rect 439332 139890 439360 151786
rect 439332 139862 439806 139890
rect 420550 139768 420606 139777
rect 420606 139726 420854 139754
rect 420550 139703 420606 139712
rect 420550 139496 420606 139505
rect 418766 139454 419014 139482
rect 420288 139468 420550 139482
rect 420302 139454 420550 139468
rect 418710 139431 418766 139440
rect 420550 139431 420606 139440
rect 426898 139496 426954 139505
rect 428738 139496 428794 139505
rect 426954 139454 427294 139482
rect 426898 139431 426954 139440
rect 429474 139496 429530 139505
rect 428794 139454 429134 139482
rect 428738 139431 428794 139440
rect 434994 139496 435050 139505
rect 429530 139454 429870 139482
rect 434838 139454 434994 139482
rect 429474 139431 429530 139440
rect 434994 139431 435050 139440
rect 439042 139496 439098 139505
rect 439098 139454 439254 139482
rect 439042 139431 439098 139440
rect 404136 139340 404492 139346
rect 404084 139334 404492 139340
rect 399864 137737 399892 139334
rect 404096 139332 404492 139334
rect 404096 139318 404478 139332
rect 399850 137728 399906 137737
rect 399850 137663 399906 137672
rect 439976 132025 440004 151786
rect 439962 132016 440018 132025
rect 439962 131951 440018 131960
rect 440252 106457 440280 200631
rect 441710 179752 441766 179761
rect 441710 179687 441766 179696
rect 440330 177304 440386 177313
rect 440330 177239 440386 177248
rect 440344 109177 440372 177239
rect 441618 160712 441674 160721
rect 441618 160647 441674 160656
rect 440514 140856 440570 140865
rect 440514 140791 440570 140800
rect 440422 140040 440478 140049
rect 440422 139975 440478 139984
rect 440436 128761 440464 139975
rect 440422 128752 440478 128761
rect 440422 128687 440478 128696
rect 440422 125896 440478 125905
rect 440422 125831 440478 125840
rect 440330 109168 440386 109177
rect 440330 109103 440386 109112
rect 440238 106448 440294 106457
rect 440238 106383 440294 106392
rect 399760 105596 399812 105602
rect 399760 105538 399812 105544
rect 399772 100638 399800 105538
rect 399852 104168 399904 104174
rect 399852 104110 399904 104116
rect 399864 100706 399892 104110
rect 439964 101448 440016 101454
rect 439964 101390 440016 101396
rect 439976 100774 440004 101390
rect 439964 100768 440016 100774
rect 401414 100736 401470 100745
rect 399852 100700 399904 100706
rect 421654 100736 421710 100745
rect 403360 100706 403742 100722
rect 401414 100671 401470 100680
rect 403348 100700 403742 100706
rect 399852 100642 399904 100648
rect 399760 100632 399812 100638
rect 399760 100574 399812 100580
rect 399680 100014 400062 100042
rect 400324 100014 400614 100042
rect 399680 94178 399708 100014
rect 399668 94172 399720 94178
rect 399668 94114 399720 94120
rect 399482 39264 399538 39273
rect 399482 39199 399538 39208
rect 396724 20664 396776 20670
rect 396724 20606 396776 20612
rect 400324 13802 400352 100014
rect 401152 96966 401180 100028
rect 401428 97918 401456 100671
rect 403400 100694 403742 100700
rect 404636 100700 404688 100706
rect 403348 100642 403400 100648
rect 421406 100694 421654 100722
rect 421654 100671 421710 100680
rect 425058 100736 425114 100745
rect 428646 100736 428702 100745
rect 425114 100694 425270 100722
rect 425058 100671 425114 100680
rect 428702 100694 428950 100722
rect 439070 100706 439360 100722
rect 439964 100710 440016 100716
rect 439070 100700 439372 100706
rect 439070 100694 439320 100700
rect 428646 100671 428702 100680
rect 404636 100642 404688 100648
rect 439320 100642 439372 100648
rect 402980 100632 403032 100638
rect 403032 100580 403190 100586
rect 402980 100574 403190 100580
rect 402992 100558 403190 100574
rect 404648 100042 404676 100642
rect 401612 100014 401902 100042
rect 402072 100014 402454 100042
rect 401416 97912 401468 97918
rect 401416 97854 401468 97860
rect 401140 96960 401192 96966
rect 401140 96902 401192 96908
rect 401612 64870 401640 100014
rect 402072 86970 402100 100014
rect 404464 99793 404492 100028
rect 404648 100026 405320 100042
rect 404648 100020 405332 100026
rect 404648 100014 405280 100020
rect 405280 99962 405332 99968
rect 404450 99784 404506 99793
rect 404450 99719 404506 99728
rect 404464 97850 404492 99719
rect 405568 99657 405596 100028
rect 405844 100014 406318 100042
rect 406488 100014 406870 100042
rect 404542 99648 404598 99657
rect 404542 99583 404598 99592
rect 405554 99648 405610 99657
rect 405554 99583 405610 99592
rect 403624 97844 403676 97850
rect 403624 97786 403676 97792
rect 404452 97844 404504 97850
rect 404452 97786 404504 97792
rect 402060 86964 402112 86970
rect 402060 86906 402112 86912
rect 401600 64864 401652 64870
rect 401600 64806 401652 64812
rect 403636 15910 403664 97786
rect 404556 84194 404584 99583
rect 405740 93968 405792 93974
rect 405740 93910 405792 93916
rect 404464 84166 404584 84194
rect 404464 76566 404492 84166
rect 404452 76560 404504 76566
rect 404452 76502 404504 76508
rect 405752 27538 405780 93910
rect 405844 55214 405872 100014
rect 406488 93974 406516 100014
rect 407592 99385 407620 100028
rect 407684 100014 408158 100042
rect 408512 100014 408894 100042
rect 408972 100014 409446 100042
rect 407578 99376 407634 99385
rect 407578 99311 407634 99320
rect 406476 93968 406528 93974
rect 406476 93910 406528 93916
rect 407684 84194 407712 100014
rect 407132 84166 407712 84194
rect 405832 55208 405884 55214
rect 405832 55150 405884 55156
rect 405740 27532 405792 27538
rect 405740 27474 405792 27480
rect 403624 15904 403676 15910
rect 403624 15846 403676 15852
rect 400312 13796 400364 13802
rect 400312 13738 400364 13744
rect 394148 8288 394200 8294
rect 394148 8230 394200 8236
rect 407132 4826 407160 84166
rect 408512 81394 408540 100014
rect 408972 96914 409000 100014
rect 408604 96886 409000 96914
rect 408604 93809 408632 96886
rect 408590 93800 408646 93809
rect 408590 93735 408646 93744
rect 409984 84194 410012 100028
rect 410076 100014 410734 100042
rect 411286 100014 411392 100042
rect 410076 95305 410104 100014
rect 410062 95296 410118 95305
rect 410062 95231 410118 95240
rect 410076 88330 410104 95231
rect 411364 91118 411392 100014
rect 412008 99278 412036 100028
rect 412100 100014 412574 100042
rect 411996 99272 412048 99278
rect 411996 99214 412048 99220
rect 412100 93854 412128 100014
rect 413296 95198 413324 100028
rect 413388 100014 413862 100042
rect 414124 100014 414414 100042
rect 414768 100014 415150 100042
rect 415412 100014 415702 100042
rect 413284 95192 413336 95198
rect 413284 95134 413336 95140
rect 411456 93826 412128 93854
rect 411352 91112 411404 91118
rect 411352 91054 411404 91060
rect 410064 88324 410116 88330
rect 410064 88266 410116 88272
rect 409892 84166 410012 84194
rect 408500 81388 408552 81394
rect 408500 81330 408552 81336
rect 408512 46238 408540 81330
rect 408500 46232 408552 46238
rect 408500 46174 408552 46180
rect 409892 6866 409920 84166
rect 411456 21486 411484 93826
rect 411904 91112 411956 91118
rect 411904 91054 411956 91060
rect 411916 80034 411944 91054
rect 413388 84194 413416 100014
rect 414020 96960 414072 96966
rect 414020 96902 414072 96908
rect 412652 84166 413416 84194
rect 411904 80028 411956 80034
rect 411904 79970 411956 79976
rect 411444 21480 411496 21486
rect 411444 21422 411496 21428
rect 409880 6860 409932 6866
rect 409880 6802 409932 6808
rect 407120 4820 407172 4826
rect 407120 4762 407172 4768
rect 412652 2786 412680 84166
rect 414032 36582 414060 96902
rect 414124 49026 414152 100014
rect 414768 96966 414796 100014
rect 414756 96960 414808 96966
rect 414756 96902 414808 96908
rect 414112 49020 414164 49026
rect 414112 48962 414164 48968
rect 415412 43450 415440 100014
rect 416424 96529 416452 100028
rect 416410 96520 416466 96529
rect 416410 96455 416466 96464
rect 416976 84194 417004 100028
rect 417712 99346 417740 100028
rect 417700 99340 417752 99346
rect 417700 99282 417752 99288
rect 418264 95130 418292 100028
rect 418804 96756 418856 96762
rect 418804 96698 418856 96704
rect 418252 95124 418304 95130
rect 418252 95066 418304 95072
rect 418264 94518 418292 95066
rect 418252 94512 418304 94518
rect 418252 94454 418304 94460
rect 416884 84166 417004 84194
rect 416884 69018 416912 84166
rect 416872 69012 416924 69018
rect 416872 68954 416924 68960
rect 415400 43444 415452 43450
rect 415400 43386 415452 43392
rect 418816 38622 418844 96698
rect 419000 96558 419028 100028
rect 419566 100014 419672 100042
rect 418988 96552 419040 96558
rect 418988 96494 419040 96500
rect 419644 93226 419672 100014
rect 420104 96762 420132 100028
rect 420472 100014 420854 100042
rect 420092 96756 420144 96762
rect 420092 96698 420144 96704
rect 419632 93220 419684 93226
rect 419632 93162 419684 93168
rect 420472 84194 420500 100014
rect 422128 99521 422156 100028
rect 422114 99512 422170 99521
rect 422114 99447 422170 99456
rect 421564 96892 421616 96898
rect 421564 96834 421616 96840
rect 419736 84166 420500 84194
rect 419736 61402 419764 84166
rect 419724 61396 419776 61402
rect 419724 61338 419776 61344
rect 418804 38616 418856 38622
rect 418804 38558 418856 38564
rect 414020 36576 414072 36582
rect 414020 36518 414072 36524
rect 421576 21418 421604 96834
rect 422680 96626 422708 100028
rect 423416 96898 423444 100028
rect 423692 100014 423982 100042
rect 424152 100014 424534 100042
rect 425440 100014 425822 100042
rect 423404 96892 423456 96898
rect 423404 96834 423456 96840
rect 422668 96620 422720 96626
rect 422668 96562 422720 96568
rect 423692 58682 423720 100014
rect 424152 91798 424180 100014
rect 425440 92449 425468 100014
rect 425886 99512 425942 99521
rect 425886 99447 425942 99456
rect 425426 92440 425482 92449
rect 425426 92375 425482 92384
rect 424140 91792 424192 91798
rect 424140 91734 424192 91740
rect 423680 58676 423732 58682
rect 423680 58618 423732 58624
rect 421564 21412 421616 21418
rect 421564 21354 421616 21360
rect 425900 5506 425928 99447
rect 426544 89010 426572 100028
rect 426636 100014 427110 100042
rect 426636 92546 426664 100014
rect 427832 97753 427860 100028
rect 428016 100014 428398 100042
rect 427818 97744 427874 97753
rect 427818 97679 427874 97688
rect 426624 92540 426676 92546
rect 426624 92482 426676 92488
rect 426636 91050 426664 92482
rect 426624 91044 426676 91050
rect 426624 90986 426676 90992
rect 426532 89004 426584 89010
rect 426532 88946 426584 88952
rect 428016 84182 428044 100014
rect 429672 99249 429700 100028
rect 429764 100014 430238 100042
rect 430684 100014 430974 100042
rect 431144 100014 431526 100042
rect 429658 99240 429714 99249
rect 429658 99175 429714 99184
rect 429764 88262 429792 100014
rect 430580 96960 430632 96966
rect 430580 96902 430632 96908
rect 429842 95840 429898 95849
rect 429842 95775 429898 95784
rect 429752 88256 429804 88262
rect 429752 88198 429804 88204
rect 428004 84176 428056 84182
rect 428004 84118 428056 84124
rect 425888 5500 425940 5506
rect 425888 5442 425940 5448
rect 429856 4146 429884 95775
rect 430592 40798 430620 96902
rect 430684 88233 430712 100014
rect 431144 96966 431172 100014
rect 432248 97918 432276 100028
rect 432800 99414 432828 100028
rect 432788 99408 432840 99414
rect 432788 99350 432840 99356
rect 433536 99278 433564 100028
rect 433720 100014 434102 100042
rect 433524 99272 433576 99278
rect 433524 99214 433576 99220
rect 432236 97912 432288 97918
rect 432236 97854 432288 97860
rect 431132 96960 431184 96966
rect 431132 96902 431184 96908
rect 432602 96928 432658 96937
rect 432602 96863 432658 96872
rect 430670 88224 430726 88233
rect 430670 88159 430726 88168
rect 430684 51746 430712 88159
rect 430672 51740 430724 51746
rect 430672 51682 430724 51688
rect 430580 40792 430632 40798
rect 430580 40734 430632 40740
rect 432616 30326 432644 96863
rect 433720 84194 433748 100014
rect 434640 97986 434668 100028
rect 434628 97980 434680 97986
rect 434628 97922 434680 97928
rect 435376 97918 435404 100028
rect 435468 100014 435942 100042
rect 436112 100014 436678 100042
rect 435364 97912 435416 97918
rect 435364 97854 435416 97860
rect 435468 96914 435496 100014
rect 435548 99408 435600 99414
rect 435548 99350 435600 99356
rect 434732 96886 435496 96914
rect 434732 93838 434760 96886
rect 434720 93832 434772 93838
rect 434720 93774 434772 93780
rect 435560 84194 435588 99350
rect 433352 84166 433748 84194
rect 435468 84166 435588 84194
rect 433352 51066 433380 84166
rect 435468 82822 435496 84166
rect 435456 82816 435508 82822
rect 435456 82758 435508 82764
rect 436112 63510 436140 100014
rect 437216 95169 437244 100028
rect 437492 100014 437966 100042
rect 437202 95160 437258 95169
rect 437202 95095 437258 95104
rect 436100 63504 436152 63510
rect 436100 63446 436152 63452
rect 433340 51060 433392 51066
rect 433340 51002 433392 51008
rect 437492 48278 437520 100014
rect 438504 96937 438532 100028
rect 439332 100014 439806 100042
rect 438490 96928 438546 96937
rect 438490 96863 438546 96872
rect 439332 84194 439360 100014
rect 438872 84166 439360 84194
rect 438872 78674 438900 84166
rect 440436 79354 440464 125831
rect 440528 117609 440556 140791
rect 441632 121446 441660 160647
rect 441724 140865 441752 179687
rect 442264 148368 442316 148374
rect 442264 148310 442316 148316
rect 441988 144288 442040 144294
rect 441988 144230 442040 144236
rect 441710 140856 441766 140865
rect 441710 140791 441766 140800
rect 441712 140072 441764 140078
rect 441712 140014 441764 140020
rect 441620 121440 441672 121446
rect 441620 121382 441672 121388
rect 441724 118697 441752 140014
rect 442000 130665 442028 144230
rect 442172 139392 442224 139398
rect 442172 139334 442224 139340
rect 442184 138281 442212 139334
rect 442170 138272 442226 138281
rect 442170 138207 442226 138216
rect 441986 130656 442042 130665
rect 441986 130591 442042 130600
rect 442276 122806 442304 148310
rect 442908 137284 442960 137290
rect 442908 137226 442960 137232
rect 442920 137193 442948 137226
rect 442906 137184 442962 137193
rect 442906 137119 442962 137128
rect 442906 136232 442962 136241
rect 442906 136167 442962 136176
rect 442920 135522 442948 136167
rect 442908 135516 442960 135522
rect 442908 135458 442960 135464
rect 442906 135144 442962 135153
rect 443012 135130 443040 287127
rect 443092 192500 443144 192506
rect 443092 192442 443144 192448
rect 442962 135102 443040 135130
rect 442906 135079 442962 135088
rect 442908 133272 442960 133278
rect 442906 133240 442908 133249
rect 442960 133240 442962 133249
rect 442906 133175 442962 133184
rect 443104 132494 443132 192442
rect 444470 189816 444526 189825
rect 444470 189751 444526 189760
rect 443184 152516 443236 152522
rect 443184 152458 443236 152464
rect 443196 134473 443224 152458
rect 443182 134464 443238 134473
rect 443182 134399 443238 134408
rect 444380 133884 444432 133890
rect 444380 133826 444432 133832
rect 444392 133278 444420 133826
rect 444380 133272 444432 133278
rect 444380 133214 444432 133220
rect 443012 132466 443132 132494
rect 442908 132456 442960 132462
rect 442906 132424 442908 132433
rect 442960 132424 442962 132433
rect 442906 132359 442962 132368
rect 442906 129704 442962 129713
rect 443012 129690 443040 132466
rect 442962 129662 443040 129690
rect 442906 129639 442962 129648
rect 442906 127800 442962 127809
rect 442906 127735 442962 127744
rect 442920 127634 442948 127735
rect 442908 127628 442960 127634
rect 442908 127570 442960 127576
rect 442906 126712 442962 126721
rect 442906 126647 442962 126656
rect 442920 125662 442948 126647
rect 442908 125656 442960 125662
rect 442908 125598 442960 125604
rect 442908 124160 442960 124166
rect 442906 124128 442908 124137
rect 442960 124128 442962 124137
rect 442816 124092 442868 124098
rect 442906 124063 442962 124072
rect 442816 124034 442868 124040
rect 442828 123321 442856 124034
rect 442814 123312 442870 123321
rect 442814 123247 442870 123256
rect 442264 122800 442316 122806
rect 442264 122742 442316 122748
rect 442908 122800 442960 122806
rect 442908 122742 442960 122748
rect 442632 121440 442684 121446
rect 442920 121417 442948 122742
rect 442998 122088 443054 122097
rect 442998 122023 443054 122032
rect 442632 121382 442684 121388
rect 442906 121408 442962 121417
rect 442644 120329 442672 121382
rect 442906 121343 442962 121352
rect 442630 120320 442686 120329
rect 442630 120255 442686 120264
rect 442908 119740 442960 119746
rect 442908 119682 442960 119688
rect 442920 119513 442948 119682
rect 442906 119504 442962 119513
rect 442906 119439 442962 119448
rect 441710 118688 441766 118697
rect 441710 118623 441766 118632
rect 440514 117600 440570 117609
rect 440514 117535 440570 117544
rect 441710 116648 441766 116657
rect 441710 116583 441766 116592
rect 440514 114744 440570 114753
rect 440514 114679 440570 114688
rect 440528 99414 440556 114679
rect 441618 101688 441674 101697
rect 441618 101623 441674 101632
rect 440516 99408 440568 99414
rect 440516 99350 440568 99356
rect 440424 79348 440476 79354
rect 440424 79290 440476 79296
rect 438860 78668 438912 78674
rect 438860 78610 438912 78616
rect 441632 66910 441660 101623
rect 441724 84862 441752 116583
rect 442906 115560 442962 115569
rect 442906 115495 442962 115504
rect 442920 114578 442948 115495
rect 442908 114572 442960 114578
rect 442908 114514 442960 114520
rect 442356 113960 442408 113966
rect 442356 113902 442408 113908
rect 442368 113801 442396 113902
rect 442354 113792 442410 113801
rect 442354 113727 442410 113736
rect 443012 113174 443040 122023
rect 443012 113146 443132 113174
rect 442170 111752 442226 111761
rect 442170 111687 442226 111696
rect 442184 111110 442212 111687
rect 442356 111580 442408 111586
rect 442356 111522 442408 111528
rect 442172 111104 442224 111110
rect 442368 111081 442396 111522
rect 442172 111046 442224 111052
rect 442354 111072 442410 111081
rect 442354 111007 442410 111016
rect 441802 110120 441858 110129
rect 441802 110055 441858 110064
rect 441712 84856 441764 84862
rect 441712 84798 441764 84804
rect 441816 83502 441844 110055
rect 442906 108216 442962 108225
rect 442906 108151 442962 108160
rect 442920 107710 442948 108151
rect 442908 107704 442960 107710
rect 442908 107646 442960 107652
rect 442540 107636 442592 107642
rect 442540 107578 442592 107584
rect 442552 107273 442580 107578
rect 442538 107264 442594 107273
rect 442538 107199 442594 107208
rect 441986 104408 442042 104417
rect 441986 104343 442042 104352
rect 442000 104174 442028 104343
rect 441988 104168 442040 104174
rect 441988 104110 442040 104116
rect 442000 84194 442028 104110
rect 442906 103592 442962 103601
rect 442962 103550 443040 103578
rect 442906 103527 442962 103536
rect 442724 102808 442776 102814
rect 442724 102750 442776 102756
rect 442736 102649 442764 102750
rect 442722 102640 442778 102649
rect 442722 102575 442778 102584
rect 441908 84166 442028 84194
rect 441804 83496 441856 83502
rect 441804 83438 441856 83444
rect 441908 82142 441936 84166
rect 441896 82136 441948 82142
rect 441896 82078 441948 82084
rect 441620 66904 441672 66910
rect 441620 66846 441672 66852
rect 437480 48272 437532 48278
rect 437480 48214 437532 48220
rect 432604 30320 432656 30326
rect 432604 30262 432656 30268
rect 443012 12442 443040 103550
rect 443104 71777 443132 113146
rect 443090 71768 443146 71777
rect 443090 71703 443146 71712
rect 444392 44878 444420 133214
rect 444484 102814 444512 189751
rect 444472 102808 444524 102814
rect 444472 102750 444524 102756
rect 445772 99278 445800 289954
rect 445852 209092 445904 209098
rect 445852 209034 445904 209040
rect 445864 111586 445892 209034
rect 447152 137290 447180 304982
rect 450544 264240 450596 264246
rect 450544 264182 450596 264188
rect 448518 229800 448574 229809
rect 448518 229735 448574 229744
rect 447232 214600 447284 214606
rect 447232 214542 447284 214548
rect 447140 137284 447192 137290
rect 447140 137226 447192 137232
rect 447244 124098 447272 214542
rect 447416 163532 447468 163538
rect 447416 163474 447468 163480
rect 447322 138680 447378 138689
rect 447322 138615 447378 138624
rect 447232 124092 447284 124098
rect 447232 124034 447284 124040
rect 445944 114572 445996 114578
rect 445944 114514 445996 114520
rect 445852 111580 445904 111586
rect 445852 111522 445904 111528
rect 445760 99272 445812 99278
rect 445760 99214 445812 99220
rect 444380 44872 444432 44878
rect 444380 44814 444432 44820
rect 445956 25566 445984 114514
rect 447140 111104 447192 111110
rect 447140 111046 447192 111052
rect 445944 25560 445996 25566
rect 445944 25502 445996 25508
rect 443000 12436 443052 12442
rect 443000 12378 443052 12384
rect 447152 9654 447180 111046
rect 447336 55894 447364 138615
rect 447428 119746 447456 163474
rect 447416 119740 447468 119746
rect 447416 119682 447468 119688
rect 448532 97918 448560 229735
rect 449898 203552 449954 203561
rect 449898 203487 449954 203496
rect 448610 189680 448666 189689
rect 448610 189615 448666 189624
rect 448624 133890 448652 189615
rect 448704 135516 448756 135522
rect 448704 135458 448756 135464
rect 448612 133884 448664 133890
rect 448612 133826 448664 133832
rect 448520 97912 448572 97918
rect 448520 97854 448572 97860
rect 448716 75206 448744 135458
rect 449912 113966 449940 203487
rect 450556 149054 450584 264182
rect 451278 191040 451334 191049
rect 451278 190975 451334 190984
rect 449992 149048 450044 149054
rect 449992 148990 450044 148996
rect 450544 149048 450596 149054
rect 450544 148990 450596 148996
rect 450004 142866 450032 148990
rect 449992 142860 450044 142866
rect 449992 142802 450044 142808
rect 449992 127628 450044 127634
rect 449992 127570 450044 127576
rect 449900 113960 449952 113966
rect 449900 113902 449952 113908
rect 448704 75200 448756 75206
rect 448704 75142 448756 75148
rect 447324 55888 447376 55894
rect 447324 55830 447376 55836
rect 450004 42090 450032 127570
rect 451292 104174 451320 190975
rect 452672 114578 452700 373254
rect 580368 369850 580396 378383
rect 582392 375329 582420 670647
rect 582470 644056 582526 644065
rect 582470 643991 582526 644000
rect 582484 551313 582512 643991
rect 582470 551304 582526 551313
rect 582470 551239 582526 551248
rect 582472 520328 582524 520334
rect 582472 520270 582524 520276
rect 582484 511329 582512 520270
rect 582470 511320 582526 511329
rect 582470 511255 582526 511264
rect 582576 460222 582604 683839
rect 582564 460216 582616 460222
rect 582564 460158 582616 460164
rect 582562 458144 582618 458153
rect 582562 458079 582618 458088
rect 582472 455456 582524 455462
rect 582472 455398 582524 455404
rect 582484 431633 582512 455398
rect 582470 431624 582526 431633
rect 582470 431559 582526 431568
rect 582378 375320 582434 375329
rect 582378 375255 582434 375264
rect 580356 369844 580408 369850
rect 580356 369786 580408 369792
rect 582378 365120 582434 365129
rect 582378 365055 582434 365064
rect 582392 333266 582420 365055
rect 582380 333260 582432 333266
rect 582380 333202 582432 333208
rect 460940 312588 460992 312594
rect 460940 312530 460992 312536
rect 456800 212560 456852 212566
rect 456800 212502 456852 212508
rect 454040 125656 454092 125662
rect 454040 125598 454092 125604
rect 452660 114572 452712 114578
rect 452660 114514 452712 114520
rect 452660 107704 452712 107710
rect 452660 107646 452712 107652
rect 451280 104168 451332 104174
rect 451280 104110 451332 104116
rect 449992 42084 450044 42090
rect 449992 42026 450044 42032
rect 447140 9648 447192 9654
rect 447140 9590 447192 9596
rect 452672 8265 452700 107646
rect 454052 13122 454080 125598
rect 456812 107642 456840 212502
rect 460952 139398 460980 312530
rect 580170 272232 580226 272241
rect 580170 272167 580226 272176
rect 580184 268394 580212 272167
rect 580172 268388 580224 268394
rect 580172 268330 580224 268336
rect 463700 241528 463752 241534
rect 463700 241470 463752 241476
rect 460940 139392 460992 139398
rect 460940 139334 460992 139340
rect 456800 107636 456852 107642
rect 456800 107578 456852 107584
rect 463712 101454 463740 241470
rect 465080 232552 465132 232558
rect 465080 232494 465132 232500
rect 464344 140888 464396 140894
rect 464344 140830 464396 140836
rect 464356 126954 464384 140830
rect 464344 126948 464396 126954
rect 464344 126890 464396 126896
rect 463700 101448 463752 101454
rect 463700 101390 463752 101396
rect 465092 97986 465120 232494
rect 580906 179208 580962 179217
rect 580906 179143 580962 179152
rect 580920 147694 580948 179143
rect 582470 165880 582526 165889
rect 582470 165815 582526 165824
rect 580908 147688 580960 147694
rect 580908 147630 580960 147636
rect 582380 147688 582432 147694
rect 582380 147630 582432 147636
rect 580172 139460 580224 139466
rect 580172 139402 580224 139408
rect 580184 139369 580212 139402
rect 580170 139360 580226 139369
rect 580170 139295 580226 139304
rect 580172 126948 580224 126954
rect 580172 126890 580224 126896
rect 580184 126041 580212 126890
rect 580170 126032 580226 126041
rect 580170 125967 580226 125976
rect 582392 121446 582420 147630
rect 582484 122806 582512 165815
rect 582576 144226 582604 458079
rect 582668 449206 582696 697167
rect 582930 630864 582986 630873
rect 582930 630799 582986 630808
rect 582746 617536 582802 617545
rect 582746 617471 582802 617480
rect 582760 541657 582788 617471
rect 582838 577688 582894 577697
rect 582838 577623 582894 577632
rect 582746 541648 582802 541657
rect 582746 541583 582802 541592
rect 582746 535528 582802 535537
rect 582746 535463 582802 535472
rect 582656 449200 582708 449206
rect 582656 449142 582708 449148
rect 582654 404968 582710 404977
rect 582654 404903 582710 404912
rect 582668 145625 582696 404903
rect 582760 298761 582788 535463
rect 582852 376689 582880 577623
rect 582944 558210 582972 630799
rect 583022 591016 583078 591025
rect 583022 590951 583078 590960
rect 582932 558204 582984 558210
rect 582932 558146 582984 558152
rect 582932 532024 582984 532030
rect 582932 531966 582984 531972
rect 582944 404977 582972 531966
rect 583036 496806 583064 590951
rect 583114 564360 583170 564369
rect 583114 564295 583170 564304
rect 583128 556209 583156 564295
rect 583114 556200 583170 556209
rect 583114 556135 583170 556144
rect 583758 556200 583814 556209
rect 583758 556135 583814 556144
rect 583114 536888 583170 536897
rect 583114 536823 583170 536832
rect 583024 496800 583076 496806
rect 583024 496742 583076 496748
rect 583024 465112 583076 465118
rect 583024 465054 583076 465060
rect 583036 418305 583064 465054
rect 583128 458153 583156 536823
rect 583114 458144 583170 458153
rect 583114 458079 583170 458088
rect 583022 418296 583078 418305
rect 583022 418231 583078 418240
rect 582930 404968 582986 404977
rect 582930 404903 582986 404912
rect 582838 376680 582894 376689
rect 582838 376615 582894 376624
rect 582930 351928 582986 351937
rect 582930 351863 582986 351872
rect 582944 347070 582972 351863
rect 582932 347064 582984 347070
rect 582932 347006 582984 347012
rect 582838 325272 582894 325281
rect 582838 325207 582894 325216
rect 582746 298752 582802 298761
rect 582746 298687 582802 298696
rect 582760 156670 582788 298687
rect 582852 249082 582880 325207
rect 582840 249076 582892 249082
rect 582840 249018 582892 249024
rect 582838 234696 582894 234705
rect 582838 234631 582894 234640
rect 582748 156664 582800 156670
rect 582748 156606 582800 156612
rect 582746 152688 582802 152697
rect 582746 152623 582802 152632
rect 582654 145616 582710 145625
rect 582654 145551 582710 145560
rect 582564 144220 582616 144226
rect 582564 144162 582616 144168
rect 582656 140820 582708 140826
rect 582656 140762 582708 140768
rect 582564 137284 582616 137290
rect 582564 137226 582616 137232
rect 582472 122800 582524 122806
rect 582472 122742 582524 122748
rect 582380 121440 582432 121446
rect 582380 121382 582432 121388
rect 580172 100020 580224 100026
rect 580172 99962 580224 99968
rect 580184 99521 580212 99962
rect 580170 99512 580226 99521
rect 580170 99447 580226 99456
rect 465080 97980 465132 97986
rect 465080 97922 465132 97928
rect 582470 95296 582526 95305
rect 582470 95231 582526 95240
rect 582380 91112 582432 91118
rect 582380 91054 582432 91060
rect 582392 86193 582420 91054
rect 582378 86184 582434 86193
rect 582378 86119 582434 86128
rect 582380 86080 582432 86086
rect 582380 86022 582432 86028
rect 582392 73001 582420 86022
rect 582378 72992 582434 73001
rect 582378 72927 582434 72936
rect 454040 13116 454092 13122
rect 454040 13058 454092 13064
rect 452658 8256 452714 8265
rect 452658 8191 452714 8200
rect 582484 6633 582512 95231
rect 582576 19825 582604 137226
rect 582668 59673 582696 140762
rect 582760 99346 582788 152623
rect 582748 99340 582800 99346
rect 582748 99282 582800 99288
rect 582748 94512 582800 94518
rect 582748 94454 582800 94460
rect 582654 59664 582710 59673
rect 582654 59599 582710 59608
rect 582760 33153 582788 94454
rect 582746 33144 582802 33153
rect 582746 33079 582802 33088
rect 582562 19816 582618 19825
rect 582562 19751 582618 19760
rect 582470 6624 582526 6633
rect 582470 6559 582526 6568
rect 429844 4140 429896 4146
rect 429844 4082 429896 4088
rect 582196 3528 582248 3534
rect 582196 3470 582248 3476
rect 581000 3052 581052 3058
rect 581000 2994 581052 3000
rect 412640 2780 412692 2786
rect 412640 2722 412692 2728
rect 381636 2100 381688 2106
rect 381636 2042 381688 2048
rect 581012 480 581040 2994
rect 582208 480 582236 3470
rect 582852 3058 582880 234631
rect 582944 124166 582972 347006
rect 583666 334656 583722 334665
rect 583666 334591 583722 334600
rect 583022 312080 583078 312089
rect 583022 312015 583078 312024
rect 583036 266257 583064 312015
rect 583022 266248 583078 266257
rect 583022 266183 583078 266192
rect 583022 258904 583078 258913
rect 583022 258839 583078 258848
rect 583036 149054 583064 258839
rect 583114 245576 583170 245585
rect 583114 245511 583170 245520
rect 583128 211177 583156 245511
rect 583298 232384 583354 232393
rect 583298 232319 583354 232328
rect 583114 211168 583170 211177
rect 583114 211103 583170 211112
rect 583114 192536 583170 192545
rect 583114 192471 583170 192480
rect 583024 149048 583076 149054
rect 583024 148990 583076 148996
rect 583024 142180 583076 142186
rect 583024 142122 583076 142128
rect 582932 124160 582984 124166
rect 582932 124102 582984 124108
rect 583036 112849 583064 142122
rect 583022 112840 583078 112849
rect 583022 112775 583078 112784
rect 583128 97986 583156 192471
rect 583206 186960 583262 186969
rect 583206 186895 583262 186904
rect 583116 97980 583168 97986
rect 583116 97922 583168 97928
rect 582932 92540 582984 92546
rect 582932 92482 582984 92488
rect 582944 86086 582972 92482
rect 583024 86284 583076 86290
rect 583024 86226 583076 86232
rect 582932 86080 582984 86086
rect 582932 86022 582984 86028
rect 583036 84194 583064 86226
rect 582944 84166 583064 84194
rect 582944 46345 582972 84166
rect 582930 46336 582986 46345
rect 582930 46271 582986 46280
rect 583220 3534 583248 186895
rect 583312 146946 583340 232319
rect 583390 219056 583446 219065
rect 583390 218991 583446 219000
rect 583404 150414 583432 218991
rect 583574 211168 583630 211177
rect 583574 211103 583630 211112
rect 583482 205456 583538 205465
rect 583482 205391 583538 205400
rect 583392 150408 583444 150414
rect 583392 150350 583444 150356
rect 583300 146940 583352 146946
rect 583300 146882 583352 146888
rect 583496 139398 583524 205391
rect 583588 155242 583616 211103
rect 583576 155236 583628 155242
rect 583576 155178 583628 155184
rect 583484 139392 583536 139398
rect 583484 139334 583536 139340
rect 583680 6914 583708 334591
rect 583772 132462 583800 556135
rect 583760 132456 583812 132462
rect 583760 132398 583812 132404
rect 583404 6886 583708 6914
rect 583208 3528 583260 3534
rect 583208 3470 583260 3476
rect 582840 3052 582892 3058
rect 582840 2994 582892 3000
rect 583404 480 583432 6886
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 684256 3478 684312
rect 3514 671200 3570 671256
rect 3422 658144 3478 658200
rect 3514 632068 3516 632088
rect 3516 632068 3568 632088
rect 3568 632068 3570 632088
rect 3514 632032 3570 632068
rect 3514 619112 3570 619168
rect 3514 606056 3570 606112
rect 3422 579944 3478 580000
rect 3422 566888 3478 566944
rect 3330 553832 3386 553888
rect 3422 527856 3478 527912
rect 3330 475632 3386 475688
rect 3514 514820 3570 514856
rect 3514 514800 3516 514820
rect 3516 514800 3568 514820
rect 3568 514800 3570 514820
rect 3514 501744 3570 501800
rect 14462 536016 14518 536072
rect 3514 462576 3570 462632
rect 3146 449520 3202 449576
rect 3146 423544 3202 423600
rect 3422 410488 3478 410544
rect 2778 397432 2834 397488
rect 7562 386960 7618 387016
rect 4802 385600 4858 385656
rect 3238 371356 3240 371376
rect 3240 371356 3292 371376
rect 3292 371356 3294 371376
rect 3238 371320 3294 371356
rect 3330 358944 3386 359000
rect 3422 358400 3478 358456
rect 2778 254088 2834 254144
rect 3330 214920 3386 214976
rect 3054 201864 3110 201920
rect 2778 149776 2834 149832
rect 3146 110608 3202 110664
rect 3054 58520 3110 58576
rect 2870 32408 2926 32464
rect 18 6704 74 6760
rect 3514 345344 3570 345400
rect 4066 319232 4122 319288
rect 3514 306176 3570 306232
rect 3514 293120 3570 293176
rect 3514 267144 3570 267200
rect 3514 241068 3516 241088
rect 3516 241068 3568 241088
rect 3568 241068 3570 241088
rect 3514 241032 3570 241068
rect 3514 188808 3570 188864
rect 3514 162832 3570 162888
rect 3514 136720 3570 136776
rect 3514 97552 3570 97608
rect 3514 84632 3570 84688
rect 5446 79464 5502 79520
rect 4066 21256 4122 21312
rect 3422 19352 3478 19408
rect 1674 4800 1730 4856
rect 2870 3304 2926 3360
rect 18602 372544 18658 372600
rect 18602 371320 18658 371376
rect 19246 371320 19302 371376
rect 16486 340040 16542 340096
rect 15842 193160 15898 193216
rect 16486 193160 16542 193216
rect 12346 80688 12402 80744
rect 10966 55800 11022 55856
rect 6826 37984 6882 38040
rect 17866 77832 17922 77888
rect 15106 69536 15162 69592
rect 19154 75112 19210 75168
rect 22006 72528 22062 72584
rect 20626 25472 20682 25528
rect 45466 536016 45522 536072
rect 35162 329840 35218 329896
rect 41326 240080 41382 240136
rect 50802 517520 50858 517576
rect 50802 447752 50858 447808
rect 39946 217912 40002 217968
rect 50986 518064 51042 518120
rect 50986 517520 51042 517576
rect 49606 214512 49662 214568
rect 40682 203496 40738 203552
rect 35162 178608 35218 178664
rect 36542 79328 36598 79384
rect 32402 71712 32458 71768
rect 23386 54440 23442 54496
rect 28906 50224 28962 50280
rect 27526 48864 27582 48920
rect 25318 6160 25374 6216
rect 35806 73752 35862 73808
rect 37186 42064 37242 42120
rect 52274 444624 52330 444680
rect 52182 415384 52238 415440
rect 42706 64096 42762 64152
rect 53746 533296 53802 533352
rect 53654 378664 53710 378720
rect 52182 223488 52238 223544
rect 50986 72392 51042 72448
rect 50986 71032 51042 71088
rect 48226 65456 48282 65512
rect 47582 44240 47638 44296
rect 46846 35128 46902 35184
rect 53562 216416 53618 216472
rect 56506 416608 56562 416664
rect 56506 415384 56562 415440
rect 53746 51720 53802 51776
rect 53654 46144 53710 46200
rect 54482 36488 54538 36544
rect 57702 382880 57758 382936
rect 56506 366288 56562 366344
rect 56414 340040 56470 340096
rect 56414 213832 56470 213888
rect 57794 227568 57850 227624
rect 59174 355272 59230 355328
rect 61842 453192 61898 453248
rect 60646 445712 60702 445768
rect 60554 407088 60610 407144
rect 61842 388728 61898 388784
rect 61842 388320 61898 388376
rect 60554 382336 60610 382392
rect 60462 346568 60518 346624
rect 59082 230152 59138 230208
rect 60646 331744 60702 331800
rect 60462 233144 60518 233200
rect 60554 222128 60610 222184
rect 57886 57160 57942 57216
rect 57242 17176 57298 17232
rect 58622 53080 58678 53136
rect 57150 3304 57206 3360
rect 65982 573416 66038 573472
rect 66074 559544 66130 559600
rect 65982 542272 66038 542328
rect 64602 416608 64658 416664
rect 61934 384240 61990 384296
rect 62026 374040 62082 374096
rect 61750 249872 61806 249928
rect 61842 228248 61898 228304
rect 63130 334600 63186 334656
rect 64694 391312 64750 391368
rect 64602 389136 64658 389192
rect 63406 369008 63462 369064
rect 63222 240760 63278 240816
rect 65522 380976 65578 381032
rect 64694 362208 64750 362264
rect 64602 336776 64658 336832
rect 64786 342896 64842 342952
rect 63406 284316 63408 284336
rect 63408 284316 63460 284336
rect 63460 284316 63462 284336
rect 63406 284280 63462 284316
rect 63314 231784 63370 231840
rect 64602 236544 64658 236600
rect 66810 588376 66866 588432
rect 66258 586508 66260 586528
rect 66260 586508 66312 586528
rect 66312 586508 66314 586528
rect 66258 586472 66314 586508
rect 66810 585656 66866 585712
rect 66810 582936 66866 582992
rect 66718 581712 66774 581768
rect 66810 580216 66866 580272
rect 67546 577496 67602 577552
rect 67454 576156 67510 576192
rect 67454 576136 67456 576156
rect 67456 576136 67508 576156
rect 67508 576136 67510 576156
rect 67362 574912 67418 574968
rect 66810 572056 66866 572112
rect 67362 570696 67418 570752
rect 66810 569336 66866 569392
rect 66810 567976 66866 568032
rect 66810 564984 66866 565040
rect 66810 563624 66866 563680
rect 66810 562264 66866 562320
rect 66810 560904 66866 560960
rect 66258 558320 66314 558376
rect 66810 555464 66866 555520
rect 66442 554104 66498 554160
rect 66810 550024 66866 550080
rect 66810 548664 66866 548720
rect 66902 547304 66958 547360
rect 66902 545944 66958 546000
rect 66902 544584 66958 544640
rect 66902 543224 66958 543280
rect 66994 541864 67050 541920
rect 67086 537376 67142 537432
rect 66166 536696 66222 536752
rect 66074 424224 66130 424280
rect 67086 522960 67142 523016
rect 66902 522824 66958 522880
rect 66350 439864 66406 439920
rect 66258 435396 66314 435432
rect 66258 435376 66260 435396
rect 66260 435376 66312 435396
rect 66312 435376 66314 435396
rect 66258 433236 66260 433256
rect 66260 433236 66312 433256
rect 66312 433236 66314 433256
rect 66258 433200 66314 433236
rect 66810 437688 66866 437744
rect 66074 380976 66130 381032
rect 65890 376624 65946 376680
rect 65982 357448 66038 357504
rect 65890 332696 65946 332752
rect 66534 431024 66590 431080
rect 66810 428576 66866 428632
rect 66810 426264 66866 426320
rect 66626 421912 66682 421968
rect 66810 415112 66866 415168
rect 66718 410624 66774 410680
rect 66350 406136 66406 406192
rect 66350 403688 66406 403744
rect 66350 401512 66406 401568
rect 66350 399336 66406 399392
rect 66994 396888 67050 396944
rect 67454 552744 67510 552800
rect 67362 442176 67418 442232
rect 70306 590688 70362 590744
rect 71134 590688 71190 590744
rect 70306 589872 70362 589928
rect 74906 592048 74962 592104
rect 77666 590960 77722 591016
rect 72422 588648 72478 588704
rect 82266 590824 82322 590880
rect 81346 589328 81402 589384
rect 83186 589464 83242 589520
rect 88062 588512 88118 588568
rect 67730 584296 67786 584352
rect 67638 566616 67694 566672
rect 67546 539588 67548 539608
rect 67548 539588 67600 539608
rect 67600 539588 67602 539608
rect 67546 539552 67602 539588
rect 67822 578856 67878 578912
rect 88890 560088 88946 560144
rect 88798 540096 88854 540152
rect 67730 419600 67786 419656
rect 67454 412800 67510 412856
rect 67362 396888 67418 396944
rect 67270 395936 67326 395992
rect 66810 392536 66866 392592
rect 67362 348336 67418 348392
rect 66902 326712 66958 326768
rect 66258 322360 66314 322416
rect 66810 321272 66866 321328
rect 66902 320184 66958 320240
rect 67362 341400 67418 341456
rect 66994 319096 67050 319152
rect 66810 318008 66866 318064
rect 66810 316920 66866 316976
rect 65982 305224 66038 305280
rect 65890 303048 65946 303104
rect 65982 274488 66038 274544
rect 65982 273672 66038 273728
rect 65982 255448 66038 255504
rect 65890 228928 65946 228984
rect 66534 315832 66590 315888
rect 64786 219272 64842 219328
rect 66626 314744 66682 314800
rect 66626 304136 66682 304192
rect 66718 300872 66774 300928
rect 66258 294344 66314 294400
rect 66626 288904 66682 288960
rect 66902 313928 66958 313984
rect 66902 312840 66958 312896
rect 66994 311752 67050 311808
rect 66902 309576 66958 309632
rect 66902 307400 66958 307456
rect 66902 306312 66958 306368
rect 66902 301960 66958 302016
rect 67086 310664 67142 310720
rect 66902 298696 66958 298752
rect 66902 297608 66958 297664
rect 67178 296248 67234 296304
rect 66902 295452 66958 295488
rect 66902 295432 66904 295452
rect 66904 295432 66956 295452
rect 66956 295432 66958 295452
rect 66902 293256 66958 293312
rect 66902 292168 66958 292224
rect 66902 291080 66958 291136
rect 67546 395936 67602 395992
rect 67546 394848 67602 394904
rect 69570 535472 69626 535528
rect 70490 535472 70546 535528
rect 69018 456864 69074 456920
rect 73158 536016 73214 536072
rect 72330 535472 72386 535528
rect 75182 536560 75238 536616
rect 75182 453192 75238 453248
rect 76746 536696 76802 536752
rect 72698 448568 72754 448624
rect 80058 535608 80114 535664
rect 81438 464344 81494 464400
rect 84290 535472 84346 535528
rect 82818 462848 82874 462904
rect 80886 447752 80942 447808
rect 82818 455368 82874 455424
rect 84198 447752 84254 447808
rect 86222 465704 86278 465760
rect 86866 453192 86922 453248
rect 85578 445712 85634 445768
rect 88338 457408 88394 457464
rect 87142 456048 87198 456104
rect 89718 586200 89774 586256
rect 89626 560088 89682 560144
rect 90362 589872 90418 589928
rect 89810 567296 89866 567352
rect 87050 444488 87106 444544
rect 93766 589328 93822 589384
rect 93122 588648 93178 588704
rect 91742 587560 91798 587616
rect 91374 584840 91430 584896
rect 91190 583652 91192 583672
rect 91192 583652 91244 583672
rect 91244 583652 91246 583672
rect 91190 583616 91246 583652
rect 91742 582120 91798 582176
rect 91742 580760 91798 580816
rect 91742 579400 91798 579456
rect 91098 576680 91154 576736
rect 91098 575320 91154 575376
rect 91098 573960 91154 574016
rect 91190 572600 91246 572656
rect 91098 571396 91154 571432
rect 91098 571376 91100 571396
rect 91100 571376 91152 571396
rect 91152 571376 91154 571396
rect 91098 570016 91154 570072
rect 91098 568656 91154 568712
rect 91466 567296 91522 567352
rect 91374 565836 91376 565856
rect 91376 565836 91428 565856
rect 91428 565836 91430 565856
rect 91374 565800 91430 565836
rect 91374 564460 91430 564496
rect 91374 564440 91376 564460
rect 91376 564440 91428 564460
rect 91428 564440 91430 564460
rect 91374 563100 91430 563136
rect 91374 563080 91376 563100
rect 91376 563080 91428 563100
rect 91428 563080 91430 563100
rect 91098 561448 91154 561504
rect 91190 558728 91246 558784
rect 91098 556008 91154 556064
rect 91098 554784 91154 554840
rect 91098 554648 91154 554704
rect 91098 552100 91100 552120
rect 91100 552100 91152 552120
rect 91152 552100 91154 552120
rect 91098 552064 91154 552100
rect 91098 550724 91154 550760
rect 91098 550704 91100 550724
rect 91100 550704 91152 550724
rect 91152 550704 91154 550724
rect 91098 549344 91154 549400
rect 91098 547848 91154 547904
rect 91098 545148 91154 545184
rect 91098 545128 91100 545148
rect 91100 545128 91152 545148
rect 91152 545128 91154 545148
rect 91098 542428 91154 542464
rect 91098 542408 91100 542428
rect 91100 542408 91152 542428
rect 91152 542408 91154 542428
rect 91098 541184 91154 541240
rect 91098 539708 91154 539744
rect 91098 539688 91100 539708
rect 91100 539688 91152 539708
rect 91152 539688 91154 539708
rect 91282 557368 91338 557424
rect 92110 553288 92166 553344
rect 91374 547984 91430 548040
rect 91282 546488 91338 546544
rect 90454 535472 90510 535528
rect 91558 546508 91614 546544
rect 91558 546488 91560 546508
rect 91560 546488 91612 546508
rect 91612 546488 91614 546508
rect 92386 542272 92442 542328
rect 90454 459584 90510 459640
rect 91558 450472 91614 450528
rect 90362 444896 90418 444952
rect 92386 449112 92442 449168
rect 96618 592048 96674 592104
rect 95882 590824 95938 590880
rect 95146 547848 95202 547904
rect 94594 464344 94650 464400
rect 95882 469784 95938 469840
rect 95146 460128 95202 460184
rect 93030 447072 93086 447128
rect 93030 444624 93086 444680
rect 94502 444624 94558 444680
rect 97262 590960 97318 591016
rect 97906 543768 97962 543824
rect 97998 531392 98054 531448
rect 97906 471144 97962 471200
rect 154118 702480 154174 702536
rect 98642 451288 98698 451344
rect 96618 445712 96674 445768
rect 97630 445712 97686 445768
rect 101494 479440 101550 479496
rect 101586 456048 101642 456104
rect 104254 468424 104310 468480
rect 106186 554784 106242 554840
rect 104162 457000 104218 457056
rect 102138 445712 102194 445768
rect 111062 589464 111118 589520
rect 108394 464344 108450 464400
rect 108302 447752 108358 447808
rect 109498 444488 109554 444544
rect 111522 444488 111578 444544
rect 112534 458768 112590 458824
rect 119342 585656 119398 585712
rect 116122 446392 116178 446448
rect 113178 445712 113234 445768
rect 114374 445712 114430 445768
rect 115202 445712 115258 445768
rect 114374 444488 114430 444544
rect 117594 445712 117650 445768
rect 118606 445712 118662 445768
rect 120078 444624 120134 444680
rect 120630 417016 120686 417072
rect 85670 391040 85726 391096
rect 92754 391040 92810 391096
rect 69938 390360 69994 390416
rect 67730 378800 67786 378856
rect 69662 363704 69718 363760
rect 67546 299784 67602 299840
rect 67362 289992 67418 290048
rect 66810 286728 66866 286784
rect 66902 285640 66958 285696
rect 66258 284552 66314 284608
rect 66810 282376 66866 282432
rect 66810 279112 66866 279168
rect 66902 278024 66958 278080
rect 66350 276120 66406 276176
rect 66810 273944 66866 274000
rect 66718 272856 66774 272912
rect 66810 271804 66812 271824
rect 66812 271804 66864 271824
rect 66864 271804 66866 271824
rect 66810 271768 66866 271804
rect 66810 268504 66866 268560
rect 67546 283464 67602 283520
rect 67454 281288 67510 281344
rect 67178 280220 67234 280256
rect 67178 280200 67180 280220
rect 67180 280200 67232 280220
rect 67232 280200 67234 280220
rect 66994 277208 67050 277264
rect 67178 266328 67234 266384
rect 66902 265240 66958 265296
rect 66442 264152 66498 264208
rect 66902 263064 66958 263120
rect 66534 261976 66590 262032
rect 66350 260908 66406 260944
rect 66350 260888 66352 260908
rect 66352 260888 66404 260908
rect 66404 260888 66406 260908
rect 66258 258068 66260 258088
rect 66260 258068 66312 258088
rect 66312 258068 66314 258088
rect 66258 258032 66314 258068
rect 66810 257624 66866 257680
rect 66626 254360 66682 254416
rect 66810 253272 66866 253328
rect 66810 251096 66866 251152
rect 66810 246744 66866 246800
rect 66810 244568 66866 244624
rect 66810 243480 66866 243536
rect 66166 216552 66222 216608
rect 64510 212472 64566 212528
rect 62762 197920 62818 197976
rect 61934 190304 61990 190360
rect 66074 129240 66130 129296
rect 65522 128016 65578 128072
rect 64970 126248 65026 126304
rect 64786 125568 64842 125624
rect 64970 125568 65026 125624
rect 65982 122576 66038 122632
rect 66166 125160 66222 125216
rect 66166 82728 66222 82784
rect 64786 81368 64842 81424
rect 62026 77152 62082 77208
rect 64786 65592 64842 65648
rect 67362 256536 67418 256592
rect 67270 252184 67326 252240
rect 67270 235728 67326 235784
rect 67730 324536 67786 324592
rect 69386 329432 69442 329488
rect 71870 390632 71926 390688
rect 73342 389000 73398 389056
rect 74538 388320 74594 388376
rect 79506 388728 79562 388784
rect 77850 388320 77906 388376
rect 73158 371864 73214 371920
rect 73066 345072 73122 345128
rect 76562 373224 76618 373280
rect 75826 364928 75882 364984
rect 75734 360168 75790 360224
rect 75182 331200 75238 331256
rect 75826 331200 75882 331256
rect 77482 329432 77538 329488
rect 79874 352688 79930 352744
rect 83922 384920 83978 384976
rect 85670 390768 85726 390824
rect 79966 331764 80022 331800
rect 79966 331744 79968 331764
rect 79968 331744 80020 331764
rect 80020 331744 80022 331764
rect 81438 342352 81494 342408
rect 83830 335960 83886 336016
rect 86222 351056 86278 351112
rect 86958 367240 87014 367296
rect 86314 349696 86370 349752
rect 89810 390360 89866 390416
rect 91282 390360 91338 390416
rect 90362 389000 90418 389056
rect 89626 370504 89682 370560
rect 89534 357992 89590 358048
rect 87602 353912 87658 353968
rect 91006 386416 91062 386472
rect 92478 388628 92480 388648
rect 92480 388628 92532 388648
rect 92532 388628 92534 388648
rect 92478 388592 92534 388628
rect 102138 390496 102194 390552
rect 94226 390360 94282 390416
rect 93766 388592 93822 388648
rect 91098 365744 91154 365800
rect 92294 377304 92350 377360
rect 93122 367512 93178 367568
rect 92294 365744 92350 365800
rect 92386 345752 92442 345808
rect 97354 390360 97410 390416
rect 96158 389000 96214 389056
rect 95238 388456 95294 388512
rect 95146 379480 95202 379536
rect 95146 343712 95202 343768
rect 96342 338680 96398 338736
rect 98826 390360 98882 390416
rect 100758 390224 100814 390280
rect 99286 385600 99342 385656
rect 99286 371320 99342 371376
rect 99194 355428 99250 355464
rect 99194 355408 99196 355428
rect 99196 355408 99248 355428
rect 99248 355408 99250 355428
rect 99194 349696 99250 349752
rect 97814 341536 97870 341592
rect 94226 331200 94282 331256
rect 94870 331200 94926 331256
rect 97814 335688 97870 335744
rect 102230 389272 102286 389328
rect 104990 390360 105046 390416
rect 106554 390360 106610 390416
rect 100758 360168 100814 360224
rect 101126 360168 101182 360224
rect 99378 353504 99434 353560
rect 100666 352552 100722 352608
rect 100574 345616 100630 345672
rect 100758 340040 100814 340096
rect 108026 390360 108082 390416
rect 107474 388456 107530 388512
rect 103426 360848 103482 360904
rect 101402 331744 101458 331800
rect 104162 337320 104218 337376
rect 103242 331744 103298 331800
rect 106922 351872 106978 351928
rect 107474 351872 107530 351928
rect 104990 349016 105046 349072
rect 109498 390360 109554 390416
rect 108394 389408 108450 389464
rect 108762 361664 108818 361720
rect 112902 389000 112958 389056
rect 106922 335960 106978 336016
rect 110234 339632 110290 339688
rect 115938 390360 115994 390416
rect 118790 390360 118846 390416
rect 116122 389000 116178 389056
rect 117134 389000 117190 389056
rect 117594 389000 117650 389056
rect 118606 389000 118662 389056
rect 120446 388456 120502 388512
rect 118974 386960 119030 387016
rect 116582 377984 116638 378040
rect 117134 377984 117190 378040
rect 116582 376760 116638 376816
rect 114558 372680 114614 372736
rect 111062 357584 111118 357640
rect 111062 352688 111118 352744
rect 111614 342216 111670 342272
rect 114374 350512 114430 350568
rect 114650 339904 114706 339960
rect 119986 375264 120042 375320
rect 118882 349152 118938 349208
rect 119894 346432 119950 346488
rect 116582 338816 116638 338872
rect 117042 334056 117098 334112
rect 121642 440000 121698 440056
rect 121642 428440 121698 428496
rect 121550 417424 121606 417480
rect 122746 428440 122802 428496
rect 122102 397296 122158 397352
rect 121550 394848 121606 394904
rect 121458 392536 121514 392592
rect 121550 382880 121606 382936
rect 123022 447752 123078 447808
rect 123022 435240 123078 435296
rect 123022 425992 123078 426048
rect 122930 421912 122986 421968
rect 122930 415148 122932 415168
rect 122932 415148 122984 415168
rect 122984 415148 122986 415168
rect 122930 415112 122986 415148
rect 122102 368464 122158 368520
rect 122746 368464 122802 368520
rect 120722 353912 120778 353968
rect 124862 538736 124918 538792
rect 123114 424088 123170 424144
rect 123482 424088 123538 424144
rect 124126 444216 124182 444272
rect 124126 442040 124182 442096
rect 124126 437824 124182 437880
rect 124126 433200 124182 433256
rect 124034 431024 124090 431080
rect 124126 412700 124128 412720
rect 124128 412700 124180 412720
rect 124180 412700 124182 412720
rect 124126 412664 124182 412700
rect 123574 411304 123630 411360
rect 124126 408312 124182 408368
rect 124126 406172 124128 406192
rect 124128 406172 124180 406192
rect 124180 406172 124182 406192
rect 124126 406136 124182 406172
rect 123850 403688 123906 403744
rect 123942 401512 123998 401568
rect 124126 399336 124182 399392
rect 123758 397296 123814 397352
rect 126886 549344 126942 549400
rect 124310 420860 124312 420880
rect 124312 420860 124364 420880
rect 124364 420860 124366 420880
rect 124310 420824 124366 420860
rect 124310 419600 124366 419656
rect 124218 384920 124274 384976
rect 124402 382472 124458 382528
rect 124126 364384 124182 364440
rect 124034 356668 124036 356688
rect 124036 356668 124088 356688
rect 124088 356668 124090 356688
rect 124034 356632 124090 356668
rect 122194 356224 122250 356280
rect 125506 360168 125562 360224
rect 124954 351056 125010 351112
rect 124954 338272 125010 338328
rect 124678 331336 124734 331392
rect 125598 348880 125654 348936
rect 126794 348880 126850 348936
rect 125506 331336 125562 331392
rect 124954 329840 125010 329896
rect 126334 340176 126390 340232
rect 126886 340176 126942 340232
rect 127806 342488 127862 342544
rect 133142 536560 133198 536616
rect 130474 370640 130530 370696
rect 130382 369008 130438 369064
rect 131026 367376 131082 367432
rect 130382 350648 130438 350704
rect 131026 350648 131082 350704
rect 129002 343848 129058 343904
rect 129646 343848 129702 343904
rect 130750 332424 130806 332480
rect 129002 331744 129058 331800
rect 133786 361664 133842 361720
rect 133694 347792 133750 347848
rect 132498 333240 132554 333296
rect 137926 546488 137982 546544
rect 137282 391312 137338 391368
rect 134522 344256 134578 344312
rect 133970 336912 134026 336968
rect 137374 369008 137430 369064
rect 137190 340856 137246 340912
rect 134890 335552 134946 335608
rect 134522 332424 134578 332480
rect 134246 331336 134302 331392
rect 135718 331744 135774 331800
rect 136454 329976 136510 330032
rect 141422 513304 141478 513360
rect 142066 513304 142122 513360
rect 140778 446392 140834 446448
rect 141422 444896 141478 444952
rect 137926 340856 137982 340912
rect 140042 346976 140098 347032
rect 139398 339632 139454 339688
rect 140042 334600 140098 334656
rect 142894 536968 142950 537024
rect 142894 447072 142950 447128
rect 142986 380160 143042 380216
rect 143354 363568 143410 363624
rect 143446 340176 143502 340232
rect 141882 334192 141938 334248
rect 144550 332152 144606 332208
rect 146114 357992 146170 358048
rect 148414 535336 148470 535392
rect 148966 535336 149022 535392
rect 147586 363024 147642 363080
rect 147586 360848 147642 360904
rect 145562 332152 145618 332208
rect 144826 331744 144882 331800
rect 145286 331200 145342 331256
rect 147678 353504 147734 353560
rect 147770 350784 147826 350840
rect 148322 350784 148378 350840
rect 147678 349696 147734 349752
rect 148506 378120 148562 378176
rect 151082 369144 151138 369200
rect 151726 360168 151782 360224
rect 149426 356088 149482 356144
rect 149426 350376 149482 350432
rect 150346 346976 150402 347032
rect 148414 335960 148470 336016
rect 149702 331336 149758 331392
rect 150254 331336 150310 331392
rect 150438 331200 150494 331256
rect 160834 559000 160890 559056
rect 155222 456864 155278 456920
rect 153842 451288 153898 451344
rect 153934 372580 153936 372600
rect 153936 372580 153988 372600
rect 153988 372580 153990 372600
rect 153934 372544 153990 372580
rect 152462 359216 152518 359272
rect 153106 359216 153162 359272
rect 151818 358944 151874 359000
rect 152646 358944 152702 359000
rect 153106 358808 153162 358864
rect 152462 334600 152518 334656
rect 153014 332832 153070 332888
rect 152646 331200 152702 331256
rect 154210 338136 154266 338192
rect 154762 336912 154818 336968
rect 155314 389272 155370 389328
rect 155222 338000 155278 338056
rect 160742 535744 160798 535800
rect 156602 386416 156658 386472
rect 156510 344936 156566 344992
rect 156510 340040 156566 340096
rect 157246 338000 157302 338056
rect 156786 337320 156842 337376
rect 157338 331472 157394 331528
rect 156970 329840 157026 329896
rect 155958 329740 155960 329760
rect 155960 329740 156012 329760
rect 156012 329740 156014 329760
rect 155958 329704 156014 329740
rect 156694 329568 156750 329624
rect 152646 329160 152702 329216
rect 67822 308488 67878 308544
rect 67730 270680 67786 270736
rect 67638 269592 67694 269648
rect 67546 259800 67602 259856
rect 67638 245656 67694 245712
rect 67362 224848 67418 224904
rect 67730 238448 67786 238504
rect 156878 327664 156934 327720
rect 156786 327256 156842 327312
rect 157430 329024 157486 329080
rect 157338 310392 157394 310448
rect 80978 241984 81034 242040
rect 69662 241848 69718 241904
rect 68374 239536 68430 239592
rect 71686 238720 71742 238776
rect 72422 240080 72478 240136
rect 69662 206896 69718 206952
rect 72698 240080 72754 240136
rect 73802 241440 73858 241496
rect 77022 239400 77078 239456
rect 76562 238720 76618 238776
rect 74630 234504 74686 234560
rect 76562 223352 76618 223408
rect 75182 220768 75238 220824
rect 74538 220496 74594 220552
rect 73802 210296 73858 210352
rect 154670 241984 154726 242040
rect 81254 224712 81310 224768
rect 81346 209480 81402 209536
rect 83646 239536 83702 239592
rect 83462 208256 83518 208312
rect 82910 206760 82966 206816
rect 78678 199960 78734 200016
rect 72422 196560 72478 196616
rect 85670 224984 85726 225040
rect 86866 226072 86922 226128
rect 86866 224984 86922 225040
rect 86222 220632 86278 220688
rect 89534 221992 89590 222048
rect 86866 200640 86922 200696
rect 91006 227432 91062 227488
rect 89810 226344 89866 226400
rect 91006 226344 91062 226400
rect 85578 192480 85634 192536
rect 91190 233008 91246 233064
rect 93858 241440 93914 241496
rect 92570 238176 92626 238232
rect 92478 206624 92534 206680
rect 91006 202272 91062 202328
rect 94916 241440 94972 241496
rect 95238 212336 95294 212392
rect 96526 212336 96582 212392
rect 93950 209616 94006 209672
rect 95146 209616 95202 209672
rect 93766 206624 93822 206680
rect 90914 186904 90970 186960
rect 99286 215872 99342 215928
rect 100666 217640 100722 217696
rect 97906 199824 97962 199880
rect 96526 190984 96582 191040
rect 95146 188400 95202 188456
rect 101954 237224 102010 237280
rect 101402 236000 101458 236056
rect 101954 236000 102010 236056
rect 101402 226208 101458 226264
rect 102230 237224 102286 237280
rect 103610 234368 103666 234424
rect 102046 210840 102102 210896
rect 104806 195200 104862 195256
rect 110694 239808 110750 239864
rect 107750 235184 107806 235240
rect 110326 230288 110382 230344
rect 111890 239400 111946 239456
rect 111798 215056 111854 215112
rect 112994 215056 113050 215112
rect 115846 239400 115902 239456
rect 115202 225936 115258 225992
rect 117134 213696 117190 213752
rect 113086 204992 113142 205048
rect 117226 200776 117282 200832
rect 119986 219000 120042 219056
rect 121366 202816 121422 202872
rect 128358 219136 128414 219192
rect 130106 240896 130162 240952
rect 129830 234368 129886 234424
rect 133142 223488 133198 223544
rect 133694 223216 133750 223272
rect 131026 210976 131082 211032
rect 133142 207984 133198 208040
rect 135442 232872 135498 232928
rect 136546 228792 136602 228848
rect 135166 224304 135222 224360
rect 137282 237088 137338 237144
rect 129646 205536 129702 205592
rect 138018 227568 138074 227624
rect 140778 235184 140834 235240
rect 140778 234232 140834 234288
rect 139582 231648 139638 231704
rect 139490 227296 139546 227352
rect 138018 221856 138074 221912
rect 141422 213560 141478 213616
rect 122746 198056 122802 198112
rect 107566 194384 107622 194440
rect 129002 193840 129058 193896
rect 100666 187040 100722 187096
rect 93766 185544 93822 185600
rect 98458 180784 98514 180840
rect 97446 179424 97502 179480
rect 98458 177520 98514 177576
rect 97446 176840 97502 176896
rect 101954 183640 102010 183696
rect 103334 182144 103390 182200
rect 101954 177520 102010 177576
rect 105726 180920 105782 180976
rect 107014 179560 107070 179616
rect 105726 177520 105782 177576
rect 112258 182280 112314 182336
rect 108946 177520 109002 177576
rect 110326 177520 110382 177576
rect 114466 177520 114522 177576
rect 115846 177520 115902 177576
rect 117226 177520 117282 177576
rect 112258 177384 112314 177440
rect 123482 177520 123538 177576
rect 107014 176976 107070 177032
rect 119802 176976 119858 177032
rect 100666 176704 100722 176760
rect 102046 176704 102102 176760
rect 103334 176704 103390 176760
rect 125046 176704 125102 176760
rect 128174 176704 128230 176760
rect 142250 235864 142306 235920
rect 146114 227568 146170 227624
rect 147494 231512 147550 231568
rect 146206 223488 146262 223544
rect 143446 219000 143502 219056
rect 143354 217776 143410 217832
rect 150070 241168 150126 241224
rect 151726 241168 151782 241224
rect 150622 235592 150678 235648
rect 148966 204176 149022 204232
rect 152002 240080 152058 240136
rect 153106 240080 153162 240136
rect 152738 237360 152794 237416
rect 152370 235748 152426 235784
rect 152370 235728 152372 235748
rect 152372 235728 152424 235748
rect 152424 235728 152426 235748
rect 152922 235728 152978 235784
rect 152462 219000 152518 219056
rect 153382 238584 153438 238640
rect 153382 235864 153438 235920
rect 153566 235864 153622 235920
rect 153106 204856 153162 204912
rect 151726 202136 151782 202192
rect 155222 239944 155278 240000
rect 156694 241984 156750 242040
rect 155682 240080 155738 240136
rect 155774 239944 155830 240000
rect 155498 234504 155554 234560
rect 155682 234524 155738 234560
rect 155682 234504 155684 234524
rect 155684 234504 155736 234524
rect 155736 234504 155738 234524
rect 155958 235184 156014 235240
rect 155314 231648 155370 231704
rect 155774 231648 155830 231704
rect 155222 223352 155278 223408
rect 154486 195336 154542 195392
rect 142066 194520 142122 194576
rect 158074 385600 158130 385656
rect 159454 389408 159510 389464
rect 159362 374584 159418 374640
rect 158166 324400 158222 324456
rect 159362 369144 159418 369200
rect 158810 339632 158866 339688
rect 160098 378664 160154 378720
rect 159454 342080 159510 342136
rect 159362 338000 159418 338056
rect 158810 335960 158866 336016
rect 158902 335416 158958 335472
rect 158902 327528 158958 327584
rect 158902 326440 158958 326496
rect 158994 326304 159050 326360
rect 158718 324264 158774 324320
rect 158718 322088 158774 322144
rect 158718 321000 158774 321056
rect 158718 318824 158774 318880
rect 158718 317736 158774 317792
rect 158902 323176 158958 323232
rect 158810 316648 158866 316704
rect 159362 319368 159418 319424
rect 158718 315560 158774 315616
rect 158718 314472 158774 314528
rect 158718 313384 158774 313440
rect 158166 309848 158222 309904
rect 158718 306856 158774 306912
rect 158810 305768 158866 305824
rect 158718 304680 158774 304736
rect 158074 291760 158130 291816
rect 158074 287680 158130 287736
rect 157982 255176 158038 255232
rect 157338 233008 157394 233064
rect 157338 224712 157394 224768
rect 158902 300056 158958 300112
rect 158718 297064 158774 297120
rect 158718 294888 158774 294944
rect 158810 293800 158866 293856
rect 158718 292984 158774 293040
rect 158718 291896 158774 291952
rect 158718 290808 158774 290864
rect 158810 289720 158866 289776
rect 159270 288632 159326 288688
rect 158718 287544 158774 287600
rect 158810 286456 158866 286512
rect 158718 285368 158774 285424
rect 158718 284316 158720 284336
rect 158720 284316 158772 284336
rect 158772 284316 158774 284336
rect 158718 284280 158774 284316
rect 158718 282104 158774 282160
rect 158718 281016 158774 281072
rect 158718 279928 158774 279984
rect 158718 278860 158774 278896
rect 158718 278840 158720 278860
rect 158720 278840 158772 278860
rect 158772 278840 158774 278860
rect 158718 276664 158774 276720
rect 158718 275576 158774 275632
rect 158718 274488 158774 274544
rect 158810 273400 158866 273456
rect 158718 271224 158774 271280
rect 158718 269068 158774 269104
rect 158718 269048 158720 269068
rect 158720 269048 158772 269068
rect 158772 269048 158774 269068
rect 158258 267960 158314 268016
rect 158718 265784 158774 265840
rect 158718 262520 158774 262576
rect 158994 261432 159050 261488
rect 158810 258168 158866 258224
rect 158718 257080 158774 257136
rect 158718 256264 158774 256320
rect 158534 255176 158590 255232
rect 158166 242120 158222 242176
rect 158718 253000 158774 253056
rect 158718 250824 158774 250880
rect 158810 249736 158866 249792
rect 158902 248648 158958 248704
rect 158718 244316 158774 244352
rect 158718 244296 158720 244316
rect 158720 244296 158772 244316
rect 158772 244296 158774 244316
rect 158718 243208 158774 243264
rect 158718 233144 158774 233200
rect 159546 311208 159602 311264
rect 160006 307944 160062 308000
rect 160190 329568 160246 329624
rect 160190 326440 160246 326496
rect 160742 316648 160798 316704
rect 159546 305632 159602 305688
rect 159914 299240 159970 299296
rect 159914 296112 159970 296168
rect 160006 295976 160062 296032
rect 159454 283192 159510 283248
rect 159178 232756 159234 232792
rect 159178 232736 159180 232756
rect 159180 232736 159232 232756
rect 159232 232736 159234 232756
rect 159362 232736 159418 232792
rect 157982 199824 158038 199880
rect 159638 271768 159694 271824
rect 159638 270136 159694 270192
rect 160098 260752 160154 260808
rect 159730 249056 159786 249112
rect 159546 247560 159602 247616
rect 160006 244840 160062 244896
rect 160006 224168 160062 224224
rect 160190 241032 160246 241088
rect 162122 370640 162178 370696
rect 160834 296792 160890 296848
rect 160834 251776 160890 251832
rect 160742 206624 160798 206680
rect 160098 202816 160154 202872
rect 161570 240896 161626 240952
rect 160926 226072 160982 226128
rect 162766 344256 162822 344312
rect 162858 342080 162914 342136
rect 162766 260616 162822 260672
rect 162950 327664 163006 327720
rect 162950 288496 163006 288552
rect 164974 339496 165030 339552
rect 165158 337320 165214 337376
rect 165158 324944 165214 325000
rect 165066 323584 165122 323640
rect 164974 322088 165030 322144
rect 164882 313248 164938 313304
rect 165434 313248 165490 313304
rect 164882 303592 164938 303648
rect 163502 262112 163558 262168
rect 163502 254496 163558 254552
rect 162490 234232 162546 234288
rect 162214 233688 162270 233744
rect 162766 233688 162822 233744
rect 162122 210976 162178 211032
rect 162766 233280 162822 233336
rect 163778 261432 163834 261488
rect 164146 254088 164202 254144
rect 163686 250416 163742 250472
rect 163686 234504 163742 234560
rect 163594 230288 163650 230344
rect 173806 557504 173862 557560
rect 169022 526360 169078 526416
rect 166262 363704 166318 363760
rect 165894 332696 165950 332752
rect 167182 388320 167238 388376
rect 165526 303592 165582 303648
rect 167642 343712 167698 343768
rect 166354 298696 166410 298752
rect 165066 262112 165122 262168
rect 165066 242800 165122 242856
rect 165526 253136 165582 253192
rect 164882 228928 164938 228984
rect 163502 223216 163558 223272
rect 162766 210976 162822 211032
rect 162766 210704 162822 210760
rect 162214 205536 162270 205592
rect 158074 199416 158130 199472
rect 156786 196832 156842 196888
rect 156602 193840 156658 193896
rect 133142 178608 133198 178664
rect 166354 276120 166410 276176
rect 166446 266328 166502 266384
rect 168102 328344 168158 328400
rect 166906 266328 166962 266384
rect 166814 255448 166870 255504
rect 166722 237360 166778 237416
rect 163502 187176 163558 187232
rect 160742 178744 160798 178800
rect 133786 177520 133842 177576
rect 134798 177520 134854 177576
rect 148230 177520 148286 177576
rect 130750 176724 130806 176760
rect 130750 176704 130752 176724
rect 130752 176704 130804 176724
rect 130804 176704 130806 176724
rect 132406 176704 132462 176760
rect 136086 176740 136088 176760
rect 136088 176740 136140 176760
rect 136140 176740 136142 176760
rect 136086 176704 136142 176740
rect 158994 176740 158996 176760
rect 158996 176740 159048 176760
rect 159048 176740 159050 176760
rect 158994 176704 159050 176740
rect 129462 175616 129518 175672
rect 164974 176976 165030 177032
rect 164882 175208 164938 175264
rect 165158 175616 165214 175672
rect 67638 123528 67694 123584
rect 67454 120808 67510 120864
rect 67362 100680 67418 100736
rect 67546 102312 67602 102368
rect 67546 94968 67602 95024
rect 166354 183640 166410 183696
rect 168102 269728 168158 269784
rect 167826 249192 167882 249248
rect 167918 242800 167974 242856
rect 167918 241576 167974 241632
rect 167734 237360 167790 237416
rect 167642 231512 167698 231568
rect 166998 220496 167054 220552
rect 167918 237088 167974 237144
rect 168286 242800 168342 242856
rect 169114 337456 169170 337512
rect 170494 356768 170550 356824
rect 170402 336776 170458 336832
rect 169666 302368 169722 302424
rect 170402 284280 170458 284336
rect 169206 280472 169262 280528
rect 168470 241984 168526 242040
rect 168378 237360 168434 237416
rect 169666 247016 169722 247072
rect 167826 199416 167882 199472
rect 167642 199280 167698 199336
rect 166906 182008 166962 182064
rect 167642 178200 167698 178256
rect 166538 175344 166594 175400
rect 169022 192616 169078 192672
rect 169022 186904 169078 186960
rect 167918 175480 167974 175536
rect 167826 171536 167882 171592
rect 166262 106800 166318 106856
rect 164974 101360 165030 101416
rect 113178 94696 113234 94752
rect 130750 94696 130806 94752
rect 74814 92384 74870 92440
rect 88062 92112 88118 92168
rect 86866 91296 86922 91352
rect 85486 91160 85542 91216
rect 86774 91160 86830 91216
rect 86774 84088 86830 84144
rect 91650 91976 91706 92032
rect 89074 91160 89130 91216
rect 91006 91160 91062 91216
rect 88062 90344 88118 90400
rect 89718 86808 89774 86864
rect 89074 85448 89130 85504
rect 86866 76472 86922 76528
rect 77206 64232 77262 64288
rect 75826 61376 75882 61432
rect 79966 62736 80022 62792
rect 78586 58520 78642 58576
rect 77390 3304 77446 3360
rect 82726 59880 82782 59936
rect 87602 75248 87658 75304
rect 95054 91296 95110 91352
rect 93674 91160 93730 91216
rect 91650 89528 91706 89584
rect 95146 91160 95202 91216
rect 96526 91160 96582 91216
rect 96526 83952 96582 84008
rect 162858 94424 162914 94480
rect 119710 93336 119766 93392
rect 123022 93336 123078 93392
rect 103426 93200 103482 93256
rect 97354 92384 97410 92440
rect 100114 92384 100170 92440
rect 103150 92384 103206 92440
rect 98734 91296 98790 91352
rect 97814 91160 97870 91216
rect 99286 91160 99342 91216
rect 98734 86672 98790 86728
rect 97814 80008 97870 80064
rect 93766 69672 93822 69728
rect 95146 68176 95202 68232
rect 100574 91160 100630 91216
rect 102046 91160 102102 91216
rect 100574 85176 100630 85232
rect 108578 92384 108634 92440
rect 116766 92384 116822 92440
rect 124126 92384 124182 92440
rect 134430 92420 134432 92440
rect 134432 92420 134484 92440
rect 134484 92420 134486 92440
rect 134430 92384 134486 92420
rect 151358 92384 151414 92440
rect 104254 91160 104310 91216
rect 104806 91160 104862 91216
rect 105542 91160 105598 91216
rect 106186 91160 106242 91216
rect 107474 91160 107530 91216
rect 108486 91160 108542 91216
rect 104254 88168 104310 88224
rect 105542 85312 105598 85368
rect 106186 82592 106242 82648
rect 106186 82048 106242 82104
rect 98642 18536 98698 18592
rect 103426 24112 103482 24168
rect 107566 77968 107622 78024
rect 110142 91704 110198 91760
rect 111706 91296 111762 91352
rect 114374 91296 114430 91352
rect 115478 91296 115534 91352
rect 115754 91296 115810 91352
rect 110326 91160 110382 91216
rect 111614 91160 111670 91216
rect 110142 89664 110198 89720
rect 112994 91160 113050 91216
rect 114466 91160 114522 91216
rect 113086 80824 113142 80880
rect 115478 87896 115534 87952
rect 115846 91160 115902 91216
rect 115294 74432 115350 74488
rect 121182 91704 121238 91760
rect 117134 91160 117190 91216
rect 118606 91160 118662 91216
rect 119986 91160 120042 91216
rect 117226 76608 117282 76664
rect 116582 67496 116638 67552
rect 121366 91160 121422 91216
rect 121826 91160 121882 91216
rect 122746 91160 122802 91216
rect 124034 91160 124090 91216
rect 122102 66816 122158 66872
rect 136454 91704 136510 91760
rect 126702 91452 126758 91488
rect 126702 91432 126704 91452
rect 126704 91432 126756 91452
rect 126756 91432 126758 91452
rect 125506 91296 125562 91352
rect 126702 91296 126758 91352
rect 125414 91160 125470 91216
rect 126794 91160 126850 91216
rect 128266 91160 128322 91216
rect 125506 68312 125562 68368
rect 129646 91160 129702 91216
rect 132406 91160 132462 91216
rect 151542 91296 151598 91352
rect 136454 89392 136510 89448
rect 133786 86536 133842 86592
rect 151726 91160 151782 91216
rect 152462 91160 152518 91216
rect 153198 90888 153254 90944
rect 161938 90344 161994 90400
rect 161938 88032 161994 88088
rect 162858 90888 162914 90944
rect 162122 89392 162178 89448
rect 162030 85176 162086 85232
rect 165526 94968 165582 95024
rect 164974 87896 165030 87952
rect 170586 294480 170642 294536
rect 170586 268368 170642 268424
rect 170494 253952 170550 254008
rect 172242 455388 172298 455424
rect 172242 455368 172244 455388
rect 172244 455368 172296 455388
rect 172296 455368 172298 455388
rect 171782 450064 171838 450120
rect 172518 373224 172574 373280
rect 171874 349696 171930 349752
rect 171782 306448 171838 306504
rect 171230 275168 171286 275224
rect 171046 253952 171102 254008
rect 171138 247016 171194 247072
rect 170954 240896 171010 240952
rect 177394 549480 177450 549536
rect 175094 532480 175150 532536
rect 175002 384240 175058 384296
rect 175002 383696 175058 383752
rect 174542 353368 174598 353424
rect 173806 353232 173862 353288
rect 173806 352552 173862 352608
rect 173346 350784 173402 350840
rect 172610 314608 172666 314664
rect 173162 285776 173218 285832
rect 172518 275848 172574 275904
rect 172334 250416 172390 250472
rect 171874 244976 171930 245032
rect 172334 244840 172390 244896
rect 171690 242936 171746 242992
rect 171138 227296 171194 227352
rect 172334 243480 172390 243536
rect 172058 227296 172114 227352
rect 170402 184184 170458 184240
rect 169114 180784 169170 180840
rect 169390 177248 169446 177304
rect 169206 176840 169262 176896
rect 171874 210296 171930 210352
rect 171874 200912 171930 200968
rect 173254 279656 173310 279712
rect 173438 273264 173494 273320
rect 175002 318824 175058 318880
rect 174634 305768 174690 305824
rect 174542 262928 174598 262984
rect 173438 229744 173494 229800
rect 172426 217232 172482 217288
rect 171874 198056 171930 198112
rect 172058 198056 172114 198112
rect 171782 173848 171838 173904
rect 173254 200640 173310 200696
rect 174818 257216 174874 257272
rect 174818 249192 174874 249248
rect 174542 186224 174598 186280
rect 173346 179560 173402 179616
rect 169022 131688 169078 131744
rect 167826 111696 167882 111752
rect 167826 110064 167882 110120
rect 167734 108704 167790 108760
rect 166538 86672 166594 86728
rect 167826 89528 167882 89584
rect 169298 93472 169354 93528
rect 169298 89120 169354 89176
rect 169206 86536 169262 86592
rect 169022 74432 169078 74488
rect 141422 44784 141478 44840
rect 135258 18536 135314 18592
rect 133142 15816 133198 15872
rect 132958 3440 133014 3496
rect 144826 39208 144882 39264
rect 170586 105168 170642 105224
rect 174542 119312 174598 119368
rect 173438 100000 173494 100056
rect 173438 84088 173494 84144
rect 180154 545264 180210 545320
rect 178774 537104 178830 537160
rect 177394 391176 177450 391232
rect 176014 345072 176070 345128
rect 176658 345888 176714 345944
rect 176658 345616 176714 345672
rect 177946 373224 178002 373280
rect 177854 345888 177910 345944
rect 177486 338272 177542 338328
rect 177302 311072 177358 311128
rect 177486 310528 177542 310584
rect 177854 310528 177910 310584
rect 176934 309032 176990 309088
rect 176934 308352 176990 308408
rect 176566 272448 176622 272504
rect 176566 271904 176622 271960
rect 176014 227296 176070 227352
rect 175186 210840 175242 210896
rect 177486 269728 177542 269784
rect 177302 254496 177358 254552
rect 177302 234368 177358 234424
rect 176658 234232 176714 234288
rect 177946 308352 178002 308408
rect 177854 264968 177910 265024
rect 178682 346976 178738 347032
rect 178682 345616 178738 345672
rect 178038 295024 178094 295080
rect 178682 273264 178738 273320
rect 177946 234232 178002 234288
rect 177946 224304 178002 224360
rect 177394 223352 177450 223408
rect 178038 223624 178094 223680
rect 178866 278704 178922 278760
rect 180246 352552 180302 352608
rect 180154 317328 180210 317384
rect 180338 347792 180394 347848
rect 180338 304952 180394 305008
rect 180706 304952 180762 305008
rect 180246 259392 180302 259448
rect 180246 257896 180302 257952
rect 178958 241848 179014 241904
rect 179326 241848 179382 241904
rect 179418 239400 179474 239456
rect 178958 238448 179014 238504
rect 179418 238448 179474 238504
rect 178866 232872 178922 232928
rect 180062 225936 180118 225992
rect 178774 210840 178830 210896
rect 178682 203496 178738 203552
rect 177394 178064 177450 178120
rect 180062 210296 180118 210352
rect 180062 204992 180118 205048
rect 177394 90480 177450 90536
rect 177302 87488 177358 87544
rect 178682 92112 178738 92168
rect 177394 82728 177450 82784
rect 177302 35128 177358 35184
rect 176566 30232 176622 30288
rect 175094 19216 175150 19272
rect 180154 202408 180210 202464
rect 181442 246472 181498 246528
rect 181718 335688 181774 335744
rect 180338 182144 180394 182200
rect 180246 178608 180302 178664
rect 182914 368328 182970 368384
rect 182454 249872 182510 249928
rect 182454 249056 182510 249112
rect 182086 234368 182142 234424
rect 182086 233280 182142 233336
rect 182822 233008 182878 233064
rect 182086 230424 182142 230480
rect 181534 183504 181590 183560
rect 181534 180920 181590 180976
rect 183006 258032 183062 258088
rect 188526 560360 188582 560416
rect 186226 553424 186282 553480
rect 184846 541048 184902 541104
rect 184386 287816 184442 287872
rect 184294 267824 184350 267880
rect 183466 249872 183522 249928
rect 183098 243072 183154 243128
rect 183374 243072 183430 243128
rect 184294 233144 184350 233200
rect 183466 228248 183522 228304
rect 183466 226072 183522 226128
rect 184202 207576 184258 207632
rect 180338 83952 180394 84008
rect 181626 88168 181682 88224
rect 180154 44784 180210 44840
rect 181718 85448 181774 85504
rect 182914 91024 182970 91080
rect 180062 10240 180118 10296
rect 185582 382472 185638 382528
rect 185582 339632 185638 339688
rect 185582 315288 185638 315344
rect 184846 313112 184902 313168
rect 185582 312568 185638 312624
rect 184754 273264 184810 273320
rect 184754 244840 184810 244896
rect 184294 201048 184350 201104
rect 184294 187176 184350 187232
rect 185674 293936 185730 293992
rect 185766 273264 185822 273320
rect 186226 273264 186282 273320
rect 187146 369008 187202 369064
rect 188342 534928 188398 534984
rect 187698 378256 187754 378312
rect 187606 350376 187662 350432
rect 187606 349968 187662 350024
rect 188986 378256 189042 378312
rect 189170 380976 189226 381032
rect 189170 375128 189226 375184
rect 189078 360304 189134 360360
rect 188526 349968 188582 350024
rect 187606 302368 187662 302424
rect 187606 283056 187662 283112
rect 187514 281424 187570 281480
rect 186318 261432 186374 261488
rect 185582 230288 185638 230344
rect 186134 214648 186190 214704
rect 185582 208936 185638 208992
rect 184386 182280 184442 182336
rect 184294 123392 184350 123448
rect 187422 233144 187478 233200
rect 188434 273264 188490 273320
rect 187514 222808 187570 222864
rect 185674 179424 185730 179480
rect 186962 179968 187018 180024
rect 186962 94560 187018 94616
rect 186962 88984 187018 89040
rect 185674 82592 185730 82648
rect 185582 20576 185638 20632
rect 187146 101360 187202 101416
rect 188342 246472 188398 246528
rect 188434 231784 188490 231840
rect 188434 211792 188490 211848
rect 188434 202272 188490 202328
rect 189078 256944 189134 257000
rect 188618 231784 188674 231840
rect 189814 382336 189870 382392
rect 191654 552064 191710 552120
rect 191102 356224 191158 356280
rect 189906 342488 189962 342544
rect 189906 331880 189962 331936
rect 189814 290536 189870 290592
rect 192574 545400 192630 545456
rect 192574 518064 192630 518120
rect 192758 378120 192814 378176
rect 192574 353504 192630 353560
rect 192482 345888 192538 345944
rect 191654 338680 191710 338736
rect 191194 292576 191250 292632
rect 190458 264832 190514 264888
rect 190274 256944 190330 257000
rect 191746 284824 191802 284880
rect 191470 247016 191526 247072
rect 190458 240896 190514 240952
rect 190366 240760 190422 240816
rect 190274 229880 190330 229936
rect 189814 221856 189870 221912
rect 189722 133864 189778 133920
rect 191746 267824 191802 267880
rect 191654 262928 191710 262984
rect 191562 241440 191618 241496
rect 190366 175752 190422 175808
rect 188434 44784 188490 44840
rect 188342 6704 188398 6760
rect 186962 6160 187018 6216
rect 191654 221448 191710 221504
rect 191838 245676 191894 245712
rect 191838 245656 191840 245676
rect 191840 245656 191892 245676
rect 191892 245656 191894 245676
rect 191930 200776 191986 200832
rect 191746 185680 191802 185736
rect 192666 241712 192722 241768
rect 192666 241576 192722 241632
rect 192666 234504 192722 234560
rect 192482 178880 192538 178936
rect 191194 131688 191250 131744
rect 193862 292576 193918 292632
rect 195334 545128 195390 545184
rect 195242 542408 195298 542464
rect 195794 446392 195850 446448
rect 195334 379480 195390 379536
rect 195242 375944 195298 376000
rect 194506 375264 194562 375320
rect 195334 372544 195390 372600
rect 195426 371864 195482 371920
rect 195334 368464 195390 368520
rect 194874 361800 194930 361856
rect 194046 356632 194102 356688
rect 194874 356632 194930 356688
rect 193954 287816 194010 287872
rect 194230 287408 194286 287464
rect 194506 272312 194562 272368
rect 195150 265512 195206 265568
rect 195150 264968 195206 265024
rect 194414 253136 194470 253192
rect 194322 241440 194378 241496
rect 194230 240760 194286 240816
rect 194046 240624 194102 240680
rect 193954 236544 194010 236600
rect 193862 227432 193918 227488
rect 194414 229744 194470 229800
rect 194414 228384 194470 228440
rect 193862 212472 193918 212528
rect 193126 199416 193182 199472
rect 195518 348336 195574 348392
rect 195426 260888 195482 260944
rect 195334 257624 195390 257680
rect 195242 245656 195298 245712
rect 195242 231240 195298 231296
rect 194506 181328 194562 181384
rect 193862 117952 193918 118008
rect 192666 109656 192722 109712
rect 192574 103808 192630 103864
rect 192574 81368 192630 81424
rect 195886 377576 195942 377632
rect 196806 543904 196862 543960
rect 197358 534520 197414 534576
rect 197358 532208 197414 532264
rect 197358 529760 197414 529816
rect 197358 527312 197414 527368
rect 197358 524728 197414 524784
rect 197358 522280 197414 522336
rect 197358 517384 197414 517440
rect 197358 514936 197414 514992
rect 198002 512488 198058 512544
rect 197358 510176 197414 510232
rect 197358 507592 197414 507648
rect 197358 497800 197414 497856
rect 197358 495508 197414 495544
rect 197358 495488 197360 495508
rect 197360 495488 197412 495508
rect 197412 495488 197414 495508
rect 197358 492904 197414 492960
rect 197358 488144 197414 488200
rect 197358 485560 197414 485616
rect 197358 480664 197414 480720
rect 197358 478216 197414 478272
rect 197358 475768 197414 475824
rect 197358 473356 197360 473376
rect 197360 473356 197412 473376
rect 197412 473356 197414 473376
rect 197358 473320 197414 473356
rect 197266 470872 197322 470928
rect 197174 382472 197230 382528
rect 196714 353912 196770 353968
rect 195978 267144 196034 267200
rect 197358 468424 197414 468480
rect 197358 465976 197414 466032
rect 197358 463256 197414 463312
rect 197358 460808 197414 460864
rect 197358 458360 197414 458416
rect 197358 448588 197414 448624
rect 197358 448568 197360 448588
rect 197360 448568 197412 448588
rect 197412 448568 197414 448588
rect 197358 446120 197414 446176
rect 197358 443808 197414 443864
rect 197726 441396 197728 441416
rect 197728 441396 197780 441416
rect 197780 441396 197782 441416
rect 197726 441360 197782 441396
rect 197358 438932 197414 438968
rect 197358 438912 197360 438932
rect 197360 438912 197412 438932
rect 197412 438912 197414 438932
rect 197358 436328 197414 436384
rect 197358 431432 197414 431488
rect 197358 428984 197414 429040
rect 197358 426536 197414 426592
rect 197358 424088 197414 424144
rect 197358 419192 197414 419248
rect 197358 416780 197360 416800
rect 197360 416780 197412 416800
rect 197412 416780 197414 416800
rect 197358 416744 197414 416780
rect 197358 414296 197414 414352
rect 197358 411848 197414 411904
rect 197358 409536 197414 409592
rect 197358 406952 197414 407008
rect 197358 399608 197414 399664
rect 197358 397160 197414 397216
rect 197358 394732 197414 394768
rect 197358 394712 197360 394732
rect 197360 394712 197412 394732
rect 197412 394712 197414 394732
rect 197358 387368 197414 387424
rect 197358 380024 197414 380080
rect 198278 500384 198334 500440
rect 207662 556144 207718 556200
rect 198830 553968 198886 554024
rect 198646 529760 198702 529816
rect 198738 505144 198794 505200
rect 198554 455912 198610 455968
rect 198462 419600 198518 419656
rect 198462 392264 198518 392320
rect 198002 346568 198058 346624
rect 197358 345092 197414 345128
rect 197358 345072 197360 345092
rect 197360 345072 197412 345092
rect 197412 345072 197414 345092
rect 197266 309712 197322 309768
rect 197174 287272 197230 287328
rect 197358 282376 197414 282432
rect 197358 280220 197414 280256
rect 197358 280200 197360 280220
rect 197360 280200 197412 280220
rect 197412 280200 197414 280220
rect 197358 279404 197414 279440
rect 197358 279384 197360 279404
rect 197360 279384 197412 279404
rect 197412 279384 197414 279404
rect 197358 278604 197360 278624
rect 197360 278604 197412 278624
rect 197412 278604 197414 278624
rect 197358 278568 197414 278604
rect 198370 278024 198426 278080
rect 197358 276664 197414 276720
rect 197266 275848 197322 275904
rect 197358 275032 197414 275088
rect 197450 274488 197506 274544
rect 197358 272856 197414 272912
rect 197358 271496 197414 271552
rect 197358 269320 197414 269376
rect 197450 268776 197506 268832
rect 197358 267960 197414 268016
rect 197358 266600 197414 266656
rect 197450 264424 197506 264480
rect 197358 263628 197414 263664
rect 197358 263608 197360 263628
rect 197360 263608 197412 263628
rect 197412 263608 197414 263628
rect 198002 262268 198058 262304
rect 198002 262248 198004 262268
rect 198004 262248 198056 262268
rect 198056 262248 198058 262268
rect 197358 261432 197414 261488
rect 197358 260072 197414 260128
rect 197358 259256 197414 259312
rect 197358 258712 197414 258768
rect 197358 257352 197414 257408
rect 196622 240488 196678 240544
rect 196622 236680 196678 236736
rect 195610 188536 195666 188592
rect 195242 3984 195298 4040
rect 197174 237904 197230 237960
rect 197174 237360 197230 237416
rect 196714 211112 196770 211168
rect 197358 256536 197414 256592
rect 197358 254360 197414 254416
rect 197358 253544 197414 253600
rect 197358 253000 197414 253056
rect 197358 251660 197414 251696
rect 197358 251640 197360 251660
rect 197360 251640 197412 251660
rect 197412 251640 197414 251660
rect 197450 250824 197506 250880
rect 197358 250008 197414 250064
rect 197358 249464 197414 249520
rect 197818 248684 197820 248704
rect 197820 248684 197872 248704
rect 197872 248684 197874 248704
rect 197818 248648 197874 248684
rect 198646 453464 198702 453520
rect 198830 463256 198886 463312
rect 198830 433880 198886 433936
rect 201406 542680 201462 542736
rect 201314 536016 201370 536072
rect 199750 535880 199806 535936
rect 204074 538600 204130 538656
rect 202786 538464 202842 538520
rect 201406 535880 201462 535936
rect 204166 538228 204168 538248
rect 204168 538228 204220 538248
rect 204220 538228 204222 538248
rect 204166 538192 204222 538228
rect 200394 535472 200450 535528
rect 202050 535472 202106 535528
rect 201406 535336 201462 535392
rect 206282 545400 206338 545456
rect 207018 542272 207074 542328
rect 207662 542272 207718 542328
rect 207018 541184 207074 541240
rect 206282 536832 206338 536888
rect 208674 536016 208730 536072
rect 216678 557504 216734 557560
rect 218702 542680 218758 542736
rect 222474 538464 222530 538520
rect 225326 546624 225382 546680
rect 230478 545264 230534 545320
rect 255962 589328 256018 589384
rect 235262 553424 235318 553480
rect 233882 537104 233938 537160
rect 247038 554784 247094 554840
rect 243542 543904 243598 543960
rect 248510 545128 248566 545184
rect 253938 542544 253994 542600
rect 263598 560224 263654 560280
rect 264242 560224 264298 560280
rect 263598 559000 263654 559056
rect 255962 541184 256018 541240
rect 257342 541184 257398 541240
rect 255594 538328 255650 538384
rect 262218 550704 262274 550760
rect 266358 538736 266414 538792
rect 265530 538192 265586 538248
rect 303618 564440 303674 564496
rect 273994 538736 274050 538792
rect 278042 547848 278098 547904
rect 285126 552064 285182 552120
rect 290094 549480 290150 549536
rect 300030 546488 300086 546544
rect 307114 539688 307170 539744
rect 331218 553968 331274 554024
rect 316590 546488 316646 546544
rect 320178 541320 320234 541376
rect 323674 540096 323730 540152
rect 339958 549344 340014 549400
rect 337106 538192 337162 538248
rect 341522 540232 341578 540288
rect 348238 541048 348294 541104
rect 345386 539552 345442 539608
rect 356242 560360 356298 560416
rect 349986 539588 349988 539608
rect 349988 539588 350040 539608
rect 350040 539588 350042 539608
rect 349986 539552 350042 539588
rect 350354 538328 350410 538384
rect 353942 543768 353998 543824
rect 353666 536968 353722 537024
rect 356150 542408 356206 542464
rect 313370 535744 313426 535800
rect 308402 535608 308458 535664
rect 342258 535608 342314 535664
rect 302330 535472 302386 535528
rect 221094 535336 221150 535392
rect 354678 535336 354734 535392
rect 199750 533296 199806 533352
rect 199658 378120 199714 378176
rect 199658 377440 199714 377496
rect 199474 376488 199530 376544
rect 199382 320864 199438 320920
rect 356242 522960 356298 523016
rect 356242 496032 356298 496088
rect 356242 492632 356298 492688
rect 357622 540232 357678 540288
rect 358818 538328 358874 538384
rect 357898 532072 357954 532128
rect 358726 532072 358782 532128
rect 358726 529624 358782 529680
rect 358726 527196 358782 527232
rect 358726 527176 358728 527196
rect 358728 527176 358780 527196
rect 358780 527176 358782 527196
rect 358726 524728 358782 524784
rect 358726 522280 358782 522336
rect 357622 519832 357678 519888
rect 358726 519832 358782 519888
rect 358726 517384 358782 517440
rect 358082 514936 358138 514992
rect 357438 512624 357494 512680
rect 356702 507592 356758 507648
rect 356334 490320 356390 490376
rect 199842 376080 199898 376136
rect 201406 377440 201462 377496
rect 199474 314608 199530 314664
rect 200118 314744 200174 314800
rect 199658 314608 199714 314664
rect 199658 313928 199714 313984
rect 198554 262792 198610 262848
rect 199934 293256 199990 293312
rect 199290 287136 199346 287192
rect 199382 284416 199438 284472
rect 199290 282920 199346 282976
rect 198646 262248 198702 262304
rect 199934 281560 199990 281616
rect 201406 364928 201462 364984
rect 202234 377576 202290 377632
rect 200762 314744 200818 314800
rect 200210 301416 200266 301472
rect 201406 301452 201408 301472
rect 201408 301452 201460 301472
rect 201460 301452 201462 301472
rect 201406 301416 201462 301452
rect 200854 300736 200910 300792
rect 200762 299376 200818 299432
rect 200394 286320 200450 286376
rect 203522 367376 203578 367432
rect 202786 361800 202842 361856
rect 202234 343712 202290 343768
rect 203522 331744 203578 331800
rect 203522 329024 203578 329080
rect 202786 317464 202842 317520
rect 202142 304816 202198 304872
rect 201590 294480 201646 294536
rect 201130 285640 201186 285696
rect 201682 291896 201738 291952
rect 201498 289176 201554 289232
rect 201498 284824 201554 284880
rect 202234 287272 202290 287328
rect 202878 300736 202934 300792
rect 202878 291896 202934 291952
rect 205638 356768 205694 356824
rect 205178 325080 205234 325136
rect 204442 299376 204498 299432
rect 204994 299412 204996 299432
rect 204996 299412 205048 299432
rect 205048 299412 205050 299432
rect 204994 299376 205050 299412
rect 203522 291080 203578 291136
rect 204166 291080 204222 291136
rect 204166 289856 204222 289912
rect 203706 285776 203762 285832
rect 204718 288088 204774 288144
rect 204258 287136 204314 287192
rect 204718 285912 204774 285968
rect 208490 376080 208546 376136
rect 207662 344256 207718 344312
rect 206466 340856 206522 340912
rect 206374 337456 206430 337512
rect 206282 323720 206338 323776
rect 206466 319368 206522 319424
rect 206374 311888 206430 311944
rect 206926 311888 206982 311944
rect 205546 285640 205602 285696
rect 207662 311208 207718 311264
rect 209134 349016 209190 349072
rect 209686 349016 209742 349072
rect 209134 348336 209190 348392
rect 208490 311072 208546 311128
rect 208490 307808 208546 307864
rect 206834 285640 206890 285696
rect 207570 285640 207626 285696
rect 209134 298152 209190 298208
rect 209410 298152 209466 298208
rect 211802 375944 211858 376000
rect 209778 297472 209834 297528
rect 211802 302504 211858 302560
rect 214562 374040 214618 374096
rect 211894 290400 211950 290456
rect 211802 288088 211858 288144
rect 211986 285640 212042 285696
rect 214654 316648 214710 316704
rect 215114 316648 215170 316704
rect 214562 312432 214618 312488
rect 213918 310392 213974 310448
rect 215114 310392 215170 310448
rect 218702 369144 218758 369200
rect 216126 363024 216182 363080
rect 216034 358808 216090 358864
rect 214010 285640 214066 285696
rect 214746 285640 214802 285696
rect 214010 284960 214066 285016
rect 216126 340040 216182 340096
rect 216034 325080 216090 325136
rect 216034 320728 216090 320784
rect 215942 285776 215998 285832
rect 218058 304816 218114 304872
rect 219346 321544 219402 321600
rect 221462 374040 221518 374096
rect 221462 355272 221518 355328
rect 222842 365744 222898 365800
rect 222198 349696 222254 349752
rect 219438 314064 219494 314120
rect 218242 301008 218298 301064
rect 218702 301008 218758 301064
rect 218058 297064 218114 297120
rect 218058 295024 218114 295080
rect 218058 289312 218114 289368
rect 216678 287680 216734 287736
rect 217690 287272 217746 287328
rect 216218 285640 216274 285696
rect 217322 284416 217378 284472
rect 218058 285776 218114 285832
rect 219714 300736 219770 300792
rect 218702 300056 218758 300112
rect 219714 299648 219770 299704
rect 218702 295160 218758 295216
rect 220174 300736 220230 300792
rect 220726 292576 220782 292632
rect 220726 290536 220782 290592
rect 220082 285776 220138 285832
rect 222934 338136 222990 338192
rect 223026 304136 223082 304192
rect 223026 295296 223082 295352
rect 221646 289856 221702 289912
rect 221462 285640 221518 285696
rect 222842 288496 222898 288552
rect 222842 286320 222898 286376
rect 224314 344256 224370 344312
rect 225602 343712 225658 343768
rect 214470 283872 214526 283928
rect 216402 283872 216458 283928
rect 218794 283872 218850 283928
rect 224314 284416 224370 284472
rect 225050 285912 225106 285968
rect 225694 322088 225750 322144
rect 225694 299512 225750 299568
rect 225970 298696 226026 298752
rect 225602 285640 225658 285696
rect 227718 348472 227774 348528
rect 226982 340720 227038 340776
rect 226338 297336 226394 297392
rect 226522 285640 226578 285696
rect 227442 299512 227498 299568
rect 228454 353368 228510 353424
rect 228914 296928 228970 296984
rect 228362 295160 228418 295216
rect 223762 283872 223818 283928
rect 227994 283872 228050 283928
rect 229742 332560 229798 332616
rect 233882 375944 233938 376000
rect 233882 375128 233938 375184
rect 232502 356632 232558 356688
rect 231122 341400 231178 341456
rect 230478 331064 230534 331120
rect 231214 331064 231270 331120
rect 231122 309712 231178 309768
rect 231674 311208 231730 311264
rect 231674 309168 231730 309224
rect 231214 306584 231270 306640
rect 231122 293256 231178 293312
rect 230386 292032 230442 292088
rect 229742 287136 229798 287192
rect 229466 283872 229522 283928
rect 232226 307672 232282 307728
rect 232226 306448 232282 306504
rect 233882 319504 233938 319560
rect 232594 307672 232650 307728
rect 232594 296792 232650 296848
rect 232502 289720 232558 289776
rect 232594 287816 232650 287872
rect 232778 285912 232834 285968
rect 236642 348336 236698 348392
rect 235262 337456 235318 337512
rect 236642 329976 236698 330032
rect 235262 311072 235318 311128
rect 235538 311072 235594 311128
rect 234710 286320 234766 286376
rect 235998 289040 236054 289096
rect 236642 289720 236698 289776
rect 242898 371320 242954 371376
rect 243634 371320 243690 371376
rect 238942 334192 238998 334248
rect 238666 327256 238722 327312
rect 238114 324944 238170 325000
rect 237378 287272 237434 287328
rect 236642 285640 236698 285696
rect 238114 284416 238170 284472
rect 239126 331880 239182 331936
rect 241978 326440 242034 326496
rect 239954 292576 240010 292632
rect 239218 289312 239274 289368
rect 239218 287680 239274 287736
rect 241426 293936 241482 293992
rect 240966 289720 241022 289776
rect 243542 344256 243598 344312
rect 242254 323584 242310 323640
rect 242162 295296 242218 295352
rect 242806 293936 242862 293992
rect 242806 289584 242862 289640
rect 242806 289176 242862 289232
rect 242898 288360 242954 288416
rect 242898 287136 242954 287192
rect 245014 363568 245070 363624
rect 243634 341536 243690 341592
rect 244738 326304 244794 326360
rect 244738 322768 244794 322824
rect 244738 321680 244794 321736
rect 243634 308488 243690 308544
rect 243818 289584 243874 289640
rect 243542 288360 243598 288416
rect 244002 287272 244058 287328
rect 244094 284960 244150 285016
rect 244002 284824 244058 284880
rect 244002 284280 244058 284336
rect 231490 283872 231546 283928
rect 236366 283872 236422 283928
rect 236734 283872 236790 283928
rect 200026 280200 200082 280256
rect 244094 284008 244150 284064
rect 247038 375264 247094 375320
rect 246302 351872 246358 351928
rect 244370 282376 244426 282432
rect 244278 278024 244334 278080
rect 199934 276664 199990 276720
rect 199842 270136 199898 270192
rect 197358 247832 197414 247888
rect 197726 245112 197782 245168
rect 198646 245112 198702 245168
rect 198554 244296 198610 244352
rect 197358 243752 197414 243808
rect 197358 242120 197414 242176
rect 199750 241848 199806 241904
rect 198830 241576 198886 241632
rect 199566 240624 199622 240680
rect 198738 240352 198794 240408
rect 199658 240488 199714 240544
rect 199750 240080 199806 240136
rect 198002 214648 198058 214704
rect 197266 182960 197322 183016
rect 196714 177112 196770 177168
rect 198738 224984 198794 225040
rect 198830 204312 198886 204368
rect 198830 204040 198886 204096
rect 200026 273672 200082 273728
rect 244278 270172 244280 270192
rect 244280 270172 244332 270192
rect 244332 270172 244334 270192
rect 244278 270136 244334 270172
rect 244002 254632 244058 254688
rect 200210 240080 200266 240136
rect 201038 240080 201094 240136
rect 200578 239944 200634 240000
rect 200210 237360 200266 237416
rect 201406 239944 201462 240000
rect 201406 237224 201462 237280
rect 202050 237904 202106 237960
rect 201590 234232 201646 234288
rect 201498 233824 201554 233880
rect 201498 229880 201554 229936
rect 201590 210296 201646 210352
rect 201590 206352 201646 206408
rect 202234 233824 202290 233880
rect 202602 240080 202658 240136
rect 202786 237260 202788 237280
rect 202788 237260 202840 237280
rect 202840 237260 202842 237280
rect 202786 237224 202842 237260
rect 202418 234232 202474 234288
rect 202878 231104 202934 231160
rect 203522 236952 203578 237008
rect 202418 196832 202474 196888
rect 202234 196696 202290 196752
rect 201406 187176 201462 187232
rect 196806 93608 196862 93664
rect 196622 3848 196678 3904
rect 199474 127200 199530 127256
rect 199382 124752 199438 124808
rect 198094 85312 198150 85368
rect 198646 104760 198702 104816
rect 198186 77152 198242 77208
rect 199474 80008 199530 80064
rect 200946 89664 201002 89720
rect 202418 189760 202474 189816
rect 202234 90344 202290 90400
rect 202418 93880 202474 93936
rect 204166 228384 204222 228440
rect 205822 238584 205878 238640
rect 205638 235220 205640 235240
rect 205640 235220 205692 235240
rect 205692 235220 205694 235240
rect 205638 235184 205694 235220
rect 204442 227296 204498 227352
rect 204442 226344 204498 226400
rect 204166 225936 204222 225992
rect 203614 210296 203670 210352
rect 204718 206896 204774 206952
rect 204902 193160 204958 193216
rect 203614 175072 203670 175128
rect 205086 200912 205142 200968
rect 205638 213696 205694 213752
rect 206282 209480 206338 209536
rect 205086 186904 205142 186960
rect 205638 186224 205694 186280
rect 205178 93744 205234 93800
rect 207938 240080 207994 240136
rect 208306 240080 208362 240136
rect 208306 238176 208362 238232
rect 207662 237088 207718 237144
rect 207570 228384 207626 228440
rect 208398 237224 208454 237280
rect 209686 229064 209742 229120
rect 209042 228928 209098 228984
rect 208490 219000 208546 219056
rect 208490 214920 208546 214976
rect 207110 206760 207166 206816
rect 207110 205672 207166 205728
rect 207662 205672 207718 205728
rect 210698 240080 210754 240136
rect 210698 237360 210754 237416
rect 211250 235456 211306 235512
rect 209778 220632 209834 220688
rect 210422 220632 210478 220688
rect 209686 215056 209742 215112
rect 209042 200776 209098 200832
rect 209042 178880 209098 178936
rect 206374 135496 206430 135552
rect 206374 94424 206430 94480
rect 206466 93744 206522 93800
rect 206282 55120 206338 55176
rect 209226 178744 209282 178800
rect 209226 124752 209282 124808
rect 209318 117952 209374 118008
rect 211894 236000 211950 236056
rect 210606 220088 210662 220144
rect 210422 206216 210478 206272
rect 210422 201048 210478 201104
rect 210422 177384 210478 177440
rect 209318 92384 209374 92440
rect 209134 92248 209190 92304
rect 210606 98640 210662 98696
rect 210514 91568 210570 91624
rect 204902 22616 204958 22672
rect 212446 235456 212502 235512
rect 212722 207848 212778 207904
rect 212722 207032 212778 207088
rect 214194 231784 214250 231840
rect 215114 239944 215170 240000
rect 214562 213696 214618 213752
rect 213274 212472 213330 212528
rect 213274 207032 213330 207088
rect 214470 205572 214472 205592
rect 214472 205572 214524 205592
rect 214524 205572 214526 205592
rect 214470 205536 214526 205572
rect 215298 235728 215354 235784
rect 215298 235184 215354 235240
rect 215298 231240 215354 231296
rect 215298 213832 215354 213888
rect 215298 212608 215354 212664
rect 216678 237360 216734 237416
rect 216586 235184 216642 235240
rect 216034 219408 216090 219464
rect 215942 213968 215998 214024
rect 215850 193840 215906 193896
rect 214562 180648 214618 180704
rect 211894 180104 211950 180160
rect 213918 175616 213974 175672
rect 213918 174936 213974 174992
rect 214010 174256 214066 174312
rect 213918 173576 213974 173632
rect 214010 172896 214066 172952
rect 213918 172216 213974 172272
rect 214838 177248 214894 177304
rect 214102 171536 214158 171592
rect 213918 171012 213974 171048
rect 213918 170992 213920 171012
rect 213920 170992 213972 171012
rect 213972 170992 213974 171012
rect 214010 170312 214066 170368
rect 213918 169652 213974 169688
rect 213918 169632 213920 169652
rect 213920 169632 213972 169652
rect 213972 169632 213974 169652
rect 214010 168952 214066 169008
rect 213918 168308 213920 168328
rect 213920 168308 213972 168328
rect 213972 168308 213974 168328
rect 213918 168272 213974 168308
rect 214010 167592 214066 167648
rect 213918 166948 213920 166968
rect 213920 166948 213972 166968
rect 213972 166948 213974 166968
rect 213918 166912 213974 166948
rect 214010 166368 214066 166424
rect 213918 165008 213974 165064
rect 214010 164328 214066 164384
rect 214562 175228 214618 175264
rect 214562 175208 214564 175228
rect 214564 175208 214616 175228
rect 214616 175208 214618 175228
rect 214562 175072 214618 175128
rect 216034 213560 216090 213616
rect 217506 240080 217562 240136
rect 218426 240080 218482 240136
rect 217506 237360 217562 237416
rect 218150 237360 218206 237416
rect 217322 210432 217378 210488
rect 216678 207984 216734 208040
rect 216678 207032 216734 207088
rect 217322 207032 217378 207088
rect 218978 239808 219034 239864
rect 219346 239808 219402 239864
rect 218426 237360 218482 237416
rect 218242 216416 218298 216472
rect 219530 237224 219586 237280
rect 219438 237088 219494 237144
rect 221002 238448 221058 238504
rect 220818 238312 220874 238368
rect 221002 237360 221058 237416
rect 220358 236544 220414 236600
rect 220082 234640 220138 234696
rect 220174 226344 220230 226400
rect 215942 177248 215998 177304
rect 215390 173848 215446 173904
rect 214838 165688 214894 165744
rect 214470 163648 214526 163704
rect 213918 162968 213974 163024
rect 213918 162288 213974 162344
rect 214010 161744 214066 161800
rect 213918 161064 213974 161120
rect 214010 160384 214066 160440
rect 213918 159704 213974 159760
rect 214010 159024 214066 159080
rect 213918 158344 213974 158400
rect 213918 157120 213974 157176
rect 214010 156440 214066 156496
rect 213918 155760 213974 155816
rect 214010 155080 214066 155136
rect 214010 154400 214066 154456
rect 213918 153720 213974 153776
rect 213918 153040 213974 153096
rect 213366 151816 213422 151872
rect 214470 152496 214526 152552
rect 213274 147192 213330 147248
rect 213182 139848 213238 139904
rect 211986 136584 212042 136640
rect 211986 119312 212042 119368
rect 211894 90480 211950 90536
rect 213918 150476 213974 150512
rect 213918 150456 213920 150476
rect 213920 150456 213972 150476
rect 213972 150456 213974 150476
rect 214010 149776 214066 149832
rect 213918 149096 213974 149152
rect 213918 147872 213974 147928
rect 213918 146512 213974 146568
rect 214010 145832 214066 145888
rect 213918 145152 213974 145208
rect 213918 143792 213974 143848
rect 214010 143248 214066 143304
rect 213918 142568 213974 142624
rect 214838 157664 214894 157720
rect 214654 151136 214710 151192
rect 214562 148416 214618 148472
rect 213918 141888 213974 141944
rect 213918 140528 213974 140584
rect 214010 139168 214066 139224
rect 213918 138624 213974 138680
rect 213918 137264 213974 137320
rect 215942 144472 215998 144528
rect 214562 141208 214618 141264
rect 214102 137944 214158 138000
rect 213918 134544 213974 134600
rect 214010 133320 214066 133376
rect 213918 132640 213974 132696
rect 213918 131960 213974 132016
rect 213918 130600 213974 130656
rect 214010 129920 214066 129976
rect 214010 129240 214066 129296
rect 213918 128696 213974 128752
rect 213918 128016 213974 128072
rect 213918 126656 213974 126712
rect 214010 125296 214066 125352
rect 213918 124616 213974 124672
rect 213918 124072 213974 124128
rect 213458 123392 213514 123448
rect 213274 118768 213330 118824
rect 213366 106120 213422 106176
rect 211986 88032 212042 88088
rect 211802 87624 211858 87680
rect 214010 122712 214066 122768
rect 213918 122032 213974 122088
rect 214010 121352 214066 121408
rect 213918 120672 213974 120728
rect 214010 119992 214066 120048
rect 213918 119448 213974 119504
rect 214010 118088 214066 118144
rect 213918 117408 213974 117464
rect 214010 116728 214066 116784
rect 213918 116048 213974 116104
rect 214010 115368 214066 115424
rect 213918 114824 213974 114880
rect 214010 114144 214066 114200
rect 213918 113464 213974 113520
rect 214010 112784 214066 112840
rect 213918 112104 213974 112160
rect 214010 111424 214066 111480
rect 213918 110744 213974 110800
rect 214010 110200 214066 110256
rect 213918 109520 213974 109576
rect 214010 108840 214066 108896
rect 213918 108160 213974 108216
rect 214010 107480 214066 107536
rect 213918 106800 213974 106856
rect 213918 104916 213974 104952
rect 213918 104896 213920 104916
rect 213920 104896 213972 104916
rect 213972 104896 213974 104916
rect 214838 135224 214894 135280
rect 214654 131280 214710 131336
rect 213918 103556 213974 103592
rect 213918 103536 213920 103556
rect 213920 103536 213972 103556
rect 213972 103536 213974 103556
rect 214010 102856 214066 102912
rect 213918 102196 213974 102232
rect 213918 102176 213920 102196
rect 213920 102176 213972 102196
rect 213972 102176 213974 102196
rect 213918 101496 213974 101552
rect 214562 100952 214618 101008
rect 213918 100272 213974 100328
rect 214470 99592 214526 99648
rect 214010 98912 214066 98968
rect 213918 98232 213974 98288
rect 213918 97552 213974 97608
rect 215298 100000 215354 100056
rect 216034 125976 216090 126032
rect 215942 98640 215998 98696
rect 214746 96872 214802 96928
rect 214562 89120 214618 89176
rect 214838 96328 214894 96384
rect 214838 86808 214894 86864
rect 216126 106664 216182 106720
rect 220358 227568 220414 227624
rect 221462 237360 221518 237416
rect 221462 212608 221518 212664
rect 220174 190304 220230 190360
rect 223394 238584 223450 238640
rect 223762 236000 223818 236056
rect 222106 214512 222162 214568
rect 221922 209480 221978 209536
rect 224222 234640 224278 234696
rect 223486 189896 223542 189952
rect 225050 238448 225106 238504
rect 225142 237360 225198 237416
rect 225786 240080 225842 240136
rect 225786 237360 225842 237416
rect 226982 238312 227038 238368
rect 226154 234368 226210 234424
rect 225234 213152 225290 213208
rect 224958 183504 225014 183560
rect 225878 183640 225934 183696
rect 225602 182824 225658 182880
rect 221462 178880 221518 178936
rect 226246 182280 226302 182336
rect 227074 233280 227130 233336
rect 227074 226344 227130 226400
rect 227534 237360 227590 237416
rect 226982 181464 227038 181520
rect 226338 178880 226394 178936
rect 227074 178880 227130 178936
rect 226338 176840 226394 176896
rect 227626 233280 227682 233336
rect 227718 233144 227774 233200
rect 228178 232872 228234 232928
rect 227718 205672 227774 205728
rect 227718 182144 227774 182200
rect 227718 178608 227774 178664
rect 230570 240080 230626 240136
rect 229834 236544 229890 236600
rect 229650 236000 229706 236056
rect 229650 232736 229706 232792
rect 230570 231648 230626 231704
rect 228638 183504 228694 183560
rect 229374 180104 229430 180160
rect 228362 179016 228418 179072
rect 227810 176568 227866 176624
rect 227810 176024 227866 176080
rect 221186 175888 221242 175944
rect 224222 175888 224278 175944
rect 229190 174020 229192 174040
rect 229192 174020 229244 174040
rect 229244 174020 229246 174040
rect 229190 173984 229246 174020
rect 229098 173712 229154 173768
rect 230386 179696 230442 179752
rect 229742 176704 229798 176760
rect 229282 170856 229338 170912
rect 229190 164328 229246 164384
rect 229742 170312 229798 170368
rect 229374 155760 229430 155816
rect 231858 239400 231914 239456
rect 231490 228928 231546 228984
rect 231122 217912 231178 217968
rect 230570 178608 230626 178664
rect 230662 176568 230718 176624
rect 230570 174664 230626 174720
rect 230570 174392 230626 174448
rect 229834 162016 229890 162072
rect 230754 173340 230756 173360
rect 230756 173340 230808 173360
rect 230808 173340 230810 173360
rect 230754 173304 230810 173340
rect 230754 170448 230810 170504
rect 230662 160928 230718 160984
rect 230754 158616 230810 158672
rect 230570 158072 230626 158128
rect 231766 171808 231822 171864
rect 231582 171400 231638 171456
rect 231766 169904 231822 169960
rect 231214 168952 231270 169008
rect 231766 168544 231822 168600
rect 231398 168000 231454 168056
rect 231766 167592 231822 167648
rect 232594 240080 232650 240136
rect 232778 238312 232834 238368
rect 232594 228384 232650 228440
rect 232502 224984 232558 225040
rect 231950 216008 232006 216064
rect 231766 166676 231768 166696
rect 231768 166676 231820 166696
rect 231820 166676 231822 166696
rect 231766 166640 231822 166676
rect 231122 166096 231178 166152
rect 231490 164736 231546 164792
rect 231766 163784 231822 163840
rect 231674 162832 231730 162888
rect 230938 161880 230994 161936
rect 231766 159568 231822 159624
rect 231122 159024 231178 159080
rect 230846 157664 230902 157720
rect 229834 152496 229890 152552
rect 229742 146240 229798 146296
rect 229650 144064 229706 144120
rect 229650 141616 229706 141672
rect 229098 140664 229154 140720
rect 229742 136856 229798 136912
rect 229742 133592 229798 133648
rect 229742 123256 229798 123312
rect 229098 96736 229154 96792
rect 225050 95920 225106 95976
rect 226430 95920 226486 95976
rect 229006 95920 229062 95976
rect 229006 95512 229062 95568
rect 228546 95240 228602 95296
rect 220818 94696 220874 94752
rect 224222 94560 224278 94616
rect 225602 94560 225658 94616
rect 218794 93064 218850 93120
rect 217322 89120 217378 89176
rect 221462 91704 221518 91760
rect 220174 83408 220230 83464
rect 221462 53080 221518 53136
rect 196806 3304 196862 3360
rect 184202 2624 184258 2680
rect 222934 84904 222990 84960
rect 226430 87488 226486 87544
rect 228362 79600 228418 79656
rect 228546 79464 228602 79520
rect 229926 131416 229982 131472
rect 230570 153720 230626 153776
rect 230570 151952 230626 152008
rect 230662 151000 230718 151056
rect 230570 149096 230626 149152
rect 231674 157936 231730 157992
rect 231306 155216 231362 155272
rect 232778 226208 232834 226264
rect 232502 199416 232558 199472
rect 232042 173984 232098 174040
rect 231674 154264 231730 154320
rect 231766 153856 231822 153912
rect 231582 153312 231638 153368
rect 233238 178064 233294 178120
rect 234066 238720 234122 238776
rect 233514 215192 233570 215248
rect 235354 227568 235410 227624
rect 237930 240080 237986 240136
rect 236826 239944 236882 240000
rect 234986 216552 235042 216608
rect 235906 216552 235962 216608
rect 235262 214648 235318 214704
rect 234434 208392 234490 208448
rect 232686 157800 232742 157856
rect 231122 149640 231178 149696
rect 230754 148144 230810 148200
rect 230570 147736 230626 147792
rect 230754 147192 230810 147248
rect 230662 144880 230718 144936
rect 230386 142976 230442 143032
rect 230570 136312 230626 136368
rect 231306 149096 231362 149152
rect 231766 146784 231822 146840
rect 231674 145696 231730 145752
rect 231306 145288 231362 145344
rect 231214 135904 231270 135960
rect 231306 135360 231362 135416
rect 231122 130600 231178 130656
rect 231030 129784 231086 129840
rect 231674 144336 231730 144392
rect 231766 143928 231822 143984
rect 231766 143420 231768 143440
rect 231768 143420 231820 143440
rect 231820 143420 231822 143440
rect 231766 143384 231822 143420
rect 231766 138216 231822 138272
rect 231766 137808 231822 137864
rect 231766 134952 231822 135008
rect 231490 134000 231546 134056
rect 231490 133048 231546 133104
rect 231398 132504 231454 132560
rect 231766 131552 231822 131608
rect 231398 131144 231454 131200
rect 231766 130192 231822 130248
rect 231306 129240 231362 129296
rect 230754 128832 230810 128888
rect 231674 128288 231730 128344
rect 231674 128016 231730 128072
rect 230662 127880 230718 127936
rect 231214 126792 231270 126848
rect 230570 125976 230626 126032
rect 230754 124480 230810 124536
rect 230018 123528 230074 123584
rect 231030 122168 231086 122224
rect 230662 118904 230718 118960
rect 230570 117408 230626 117464
rect 230846 117000 230902 117056
rect 231306 126384 231362 126440
rect 231490 125024 231546 125080
rect 231306 124752 231362 124808
rect 231214 121624 231270 121680
rect 231214 120536 231270 120592
rect 231122 114552 231178 114608
rect 230662 113600 230718 113656
rect 231030 112648 231086 112704
rect 231122 112104 231178 112160
rect 230570 111288 230626 111344
rect 230938 107072 230994 107128
rect 230754 104624 230810 104680
rect 230478 100816 230534 100872
rect 230570 99456 230626 99512
rect 230754 98912 230810 98968
rect 230754 98504 230810 98560
rect 231030 97960 231086 98016
rect 230478 96192 230534 96248
rect 229926 93064 229982 93120
rect 231766 127336 231822 127392
rect 231674 124072 231730 124128
rect 231766 122576 231822 122632
rect 231766 120672 231822 120728
rect 231490 120264 231546 120320
rect 231674 119992 231730 120048
rect 231766 119720 231822 119776
rect 231674 119312 231730 119368
rect 231398 116320 231454 116376
rect 231306 111696 231362 111752
rect 231766 116456 231822 116512
rect 231674 116048 231730 116104
rect 231490 115096 231546 115152
rect 231490 114180 231492 114200
rect 231492 114180 231544 114200
rect 231544 114180 231546 114200
rect 231490 114144 231546 114180
rect 231674 113192 231730 113248
rect 231766 112240 231822 112296
rect 231674 111016 231730 111072
rect 231766 110744 231822 110800
rect 231674 109792 231730 109848
rect 231490 107888 231546 107944
rect 231582 106528 231638 106584
rect 231398 105576 231454 105632
rect 231582 105168 231638 105224
rect 231490 103672 231546 103728
rect 231766 109384 231822 109440
rect 231766 108432 231822 108488
rect 231766 104216 231822 104272
rect 231214 103264 231270 103320
rect 231398 102720 231454 102776
rect 231674 102720 231730 102776
rect 231490 101768 231546 101824
rect 231214 101224 231270 101280
rect 231766 102312 231822 102368
rect 231766 101360 231822 101416
rect 231766 100408 231822 100464
rect 231674 99864 231730 99920
rect 234710 169496 234766 169552
rect 234618 168544 234674 168600
rect 234618 165144 234674 165200
rect 233882 155216 233938 155272
rect 233790 145832 233846 145888
rect 232778 116592 232834 116648
rect 232594 105440 232650 105496
rect 231398 98640 231454 98696
rect 231398 97552 231454 97608
rect 231306 96600 231362 96656
rect 231306 82728 231362 82784
rect 235262 135768 235318 135824
rect 234158 123392 234214 123448
rect 234066 122032 234122 122088
rect 233882 105576 233938 105632
rect 235538 166232 235594 166288
rect 236090 168408 236146 168464
rect 235538 157936 235594 157992
rect 235446 126792 235502 126848
rect 236826 168408 236882 168464
rect 238850 232872 238906 232928
rect 239402 232872 239458 232928
rect 239402 231920 239458 231976
rect 238298 231240 238354 231296
rect 238114 223488 238170 223544
rect 239402 220768 239458 220824
rect 238758 210296 238814 210352
rect 240322 235592 240378 235648
rect 240690 235320 240746 235376
rect 240690 230424 240746 230480
rect 240782 227432 240838 227488
rect 240046 223352 240102 223408
rect 238850 208256 238906 208312
rect 238758 207712 238814 207768
rect 238022 174528 238078 174584
rect 237378 166232 237434 166288
rect 238022 164464 238078 164520
rect 235354 104624 235410 104680
rect 235446 82048 235502 82104
rect 238390 167592 238446 167648
rect 238114 154808 238170 154864
rect 238022 128016 238078 128072
rect 237010 125432 237066 125488
rect 236734 84904 236790 84960
rect 236642 76608 236698 76664
rect 239034 176024 239090 176080
rect 238942 170312 238998 170368
rect 239034 163376 239090 163432
rect 239402 139440 239458 139496
rect 238206 117952 238262 118008
rect 238114 103944 238170 104000
rect 239494 118768 239550 118824
rect 241702 237496 241758 237552
rect 240966 210976 241022 211032
rect 241058 179560 241114 179616
rect 240874 146920 240930 146976
rect 242162 239264 242218 239320
rect 241794 237360 241850 237416
rect 242162 238448 242218 238504
rect 244094 241304 244150 241360
rect 243634 238584 243690 238640
rect 241702 174256 241758 174312
rect 240874 128696 240930 128752
rect 239862 115504 239918 115560
rect 239678 115096 239734 115152
rect 243634 233008 243690 233064
rect 242806 225936 242862 225992
rect 242254 219136 242310 219192
rect 242254 172896 242310 172952
rect 242438 150048 242494 150104
rect 242346 146648 242402 146704
rect 242254 133456 242310 133512
rect 242162 117544 242218 117600
rect 241518 95648 241574 95704
rect 241150 83408 241206 83464
rect 242254 110744 242310 110800
rect 244462 270952 244518 271008
rect 248510 345480 248566 345536
rect 247682 335552 247738 335608
rect 247222 334056 247278 334112
rect 245750 289720 245806 289776
rect 245750 288496 245806 288552
rect 245658 276664 245714 276720
rect 246946 283736 247002 283792
rect 246854 283212 246910 283248
rect 246854 283192 246856 283212
rect 246856 283192 246908 283212
rect 246908 283192 246910 283212
rect 245934 281560 245990 281616
rect 245934 281016 245990 281072
rect 245934 278840 245990 278896
rect 246302 278024 246358 278080
rect 245934 277480 245990 277536
rect 245934 275884 245936 275904
rect 245936 275884 245988 275904
rect 245988 275884 245990 275904
rect 245934 275848 245990 275884
rect 245750 275304 245806 275360
rect 245658 274488 245714 274544
rect 245842 273672 245898 273728
rect 245750 273128 245806 273184
rect 245934 272312 245990 272368
rect 245934 271496 245990 271552
rect 245842 269592 245898 269648
rect 245750 266600 245806 266656
rect 245658 265820 245660 265840
rect 245660 265820 245712 265840
rect 245712 265820 245714 265840
rect 245658 265784 245714 265820
rect 246026 264424 246082 264480
rect 245842 263880 245898 263936
rect 244554 258168 244610 258224
rect 245934 262268 245990 262304
rect 245934 262248 245936 262268
rect 245936 262248 245988 262268
rect 245988 262248 245990 262268
rect 245750 261704 245806 261760
rect 246026 261432 246082 261488
rect 245842 260924 245844 260944
rect 245844 260924 245896 260944
rect 245896 260924 245898 260944
rect 245842 260888 245898 260924
rect 246394 259528 246450 259584
rect 245750 258712 245806 258768
rect 245750 257352 245806 257408
rect 245658 256536 245714 256592
rect 245750 255992 245806 256048
rect 245842 254360 245898 254416
rect 245934 253836 245990 253872
rect 245934 253816 245936 253836
rect 245936 253816 245988 253836
rect 245988 253816 245990 253836
rect 246026 253000 246082 253056
rect 245934 252184 245990 252240
rect 245934 251640 245990 251696
rect 245934 250824 245990 250880
rect 245842 250280 245898 250336
rect 244462 248648 244518 248704
rect 245658 248104 245714 248160
rect 245934 247288 245990 247344
rect 245842 246472 245898 246528
rect 245934 245928 245990 245984
rect 245658 245112 245714 245168
rect 244370 226072 244426 226128
rect 244370 225256 244426 225312
rect 244370 225120 244426 225176
rect 244370 219272 244426 219328
rect 246302 244568 246358 244624
rect 245842 243752 245898 243808
rect 245750 241576 245806 241632
rect 245934 239264 245990 239320
rect 246394 242392 246450 242448
rect 246946 240760 247002 240816
rect 247314 287816 247370 287872
rect 247314 260072 247370 260128
rect 246302 223352 246358 223408
rect 244370 179968 244426 180024
rect 244278 172760 244334 172816
rect 242990 148688 243046 148744
rect 243542 138080 243598 138136
rect 242346 104760 242402 104816
rect 242530 104080 242586 104136
rect 242346 100000 242402 100056
rect 242346 75248 242402 75304
rect 243910 153176 243966 153232
rect 243910 124752 243966 124808
rect 245198 145560 245254 145616
rect 244922 113328 244978 113384
rect 242898 26832 242954 26888
rect 245842 181328 245898 181384
rect 245750 140120 245806 140176
rect 245934 174528 245990 174584
rect 247038 167048 247094 167104
rect 245934 144064 245990 144120
rect 245290 135904 245346 135960
rect 246302 121624 246358 121680
rect 245198 107480 245254 107536
rect 246670 132776 246726 132832
rect 246578 108024 246634 108080
rect 242898 7520 242954 7576
rect 246210 3848 246266 3904
rect 246670 105576 246726 105632
rect 246578 76472 246634 76528
rect 246486 64232 246542 64288
rect 247866 141344 247922 141400
rect 249706 279384 249762 279440
rect 248602 221992 248658 222048
rect 249706 213696 249762 213752
rect 249246 174256 249302 174312
rect 249062 159024 249118 159080
rect 248510 156712 248566 156768
rect 248418 145696 248474 145752
rect 247774 100816 247830 100872
rect 247682 57160 247738 57216
rect 249062 118632 249118 118688
rect 247774 48864 247830 48920
rect 249982 297064 250038 297120
rect 253202 364928 253258 364984
rect 252650 332832 252706 332888
rect 250442 202408 250498 202464
rect 250442 165960 250498 166016
rect 249890 162424 249946 162480
rect 250534 150864 250590 150920
rect 249154 65456 249210 65512
rect 249798 50904 249854 50960
rect 249154 46144 249210 46200
rect 249982 13776 250038 13832
rect 251362 252456 251418 252512
rect 251270 249736 251326 249792
rect 252374 249736 252430 249792
rect 251270 248920 251326 248976
rect 251914 215872 251970 215928
rect 251914 215192 251970 215248
rect 251270 210704 251326 210760
rect 254582 338680 254638 338736
rect 253938 318824 253994 318880
rect 252742 261432 252798 261488
rect 254214 308488 254270 308544
rect 253202 269184 253258 269240
rect 253202 211792 253258 211848
rect 252650 183640 252706 183696
rect 251822 168544 251878 168600
rect 251178 159976 251234 160032
rect 250534 111016 250590 111072
rect 251914 154808 251970 154864
rect 250718 105576 250774 105632
rect 250718 87624 250774 87680
rect 256146 310392 256202 310448
rect 255962 310256 256018 310312
rect 255962 298152 256018 298208
rect 255410 291760 255466 291816
rect 255318 267824 255374 267880
rect 255410 266192 255466 266248
rect 255410 265512 255466 265568
rect 254122 231784 254178 231840
rect 254122 231104 254178 231160
rect 254030 217776 254086 217832
rect 255410 245676 255466 245712
rect 255410 245656 255412 245676
rect 255412 245656 255464 245676
rect 255464 245656 255466 245676
rect 256146 291760 256202 291816
rect 258078 367648 258134 367704
rect 256790 310392 256846 310448
rect 257342 310256 257398 310312
rect 256790 303728 256846 303784
rect 256698 240216 256754 240272
rect 253938 178608 253994 178664
rect 252742 172352 252798 172408
rect 253478 171536 253534 171592
rect 253202 132912 253258 132968
rect 254582 152904 254638 152960
rect 253478 132368 253534 132424
rect 253294 107752 253350 107808
rect 251822 51720 251878 51776
rect 253478 75112 253534 75168
rect 254766 151816 254822 151872
rect 254674 114552 254730 114608
rect 254582 68312 254638 68368
rect 255962 142704 256018 142760
rect 256146 142704 256202 142760
rect 254766 110336 254822 110392
rect 254766 91704 254822 91760
rect 255962 65592 256018 65648
rect 256238 116456 256294 116512
rect 259550 328480 259606 328536
rect 259550 285912 259606 285968
rect 260746 242956 260802 242992
rect 260746 242936 260748 242956
rect 260748 242936 260800 242956
rect 260800 242936 260802 242956
rect 260102 239944 260158 240000
rect 259550 222128 259606 222184
rect 259366 210976 259422 211032
rect 260746 222128 260802 222184
rect 260102 209616 260158 209672
rect 257434 163104 257490 163160
rect 258906 161880 258962 161936
rect 257526 149640 257582 149696
rect 257526 108976 257582 109032
rect 257618 101360 257674 101416
rect 257526 77832 257582 77888
rect 257434 64096 257490 64152
rect 254674 50224 254730 50280
rect 251822 33768 251878 33824
rect 250534 15136 250590 15192
rect 250534 13776 250590 13832
rect 255962 25608 256018 25664
rect 254582 24112 254638 24168
rect 253478 15816 253534 15872
rect 253478 15272 253534 15328
rect 254582 15272 254638 15328
rect 253202 11736 253258 11792
rect 257066 3984 257122 4040
rect 257342 3984 257398 4040
rect 260102 170176 260158 170232
rect 258906 121352 258962 121408
rect 260102 117816 260158 117872
rect 259274 115096 259330 115152
rect 258998 105440 259054 105496
rect 258906 73752 258962 73808
rect 259458 53896 259514 53952
rect 255870 3440 255926 3496
rect 256606 3440 256662 3496
rect 260194 69672 260250 69728
rect 262218 293120 262274 293176
rect 260930 237224 260986 237280
rect 262310 266328 262366 266384
rect 262770 266192 262826 266248
rect 262862 241304 262918 241360
rect 262310 226888 262366 226944
rect 265070 349152 265126 349208
rect 263690 347656 263746 347712
rect 264242 347656 264298 347712
rect 264242 346432 264298 346488
rect 263690 301008 263746 301064
rect 263598 212472 263654 212528
rect 264334 269728 264390 269784
rect 263598 204176 263654 204232
rect 263598 203496 263654 203552
rect 266358 296112 266414 296168
rect 264978 192480 265034 192536
rect 264334 179968 264390 180024
rect 269762 351192 269818 351248
rect 267830 209480 267886 209536
rect 269854 231240 269910 231296
rect 272706 376760 272762 376816
rect 270590 331744 270646 331800
rect 271142 284008 271198 284064
rect 270590 216552 270646 216608
rect 273258 313928 273314 313984
rect 272522 302368 272578 302424
rect 273258 286340 273314 286376
rect 273258 286320 273260 286340
rect 273260 286320 273312 286340
rect 273312 286320 273314 286340
rect 274086 309168 274142 309224
rect 273994 285776 274050 285832
rect 271878 227568 271934 227624
rect 271878 226888 271934 226944
rect 271786 216552 271842 216608
rect 271786 215872 271842 215928
rect 271142 182960 271198 183016
rect 272062 182144 272118 182200
rect 272062 181328 272118 181384
rect 274086 225528 274142 225584
rect 275374 296928 275430 296984
rect 281446 376624 281502 376680
rect 275374 178744 275430 178800
rect 273994 178608 274050 178664
rect 278042 304952 278098 305008
rect 277398 280744 277454 280800
rect 276846 219408 276902 219464
rect 276754 207576 276810 207632
rect 281446 375264 281502 375320
rect 279422 374040 279478 374096
rect 281446 374040 281502 374096
rect 278226 314744 278282 314800
rect 278134 287680 278190 287736
rect 283378 367104 283434 367160
rect 283562 367104 283618 367160
rect 283378 366288 283434 366344
rect 279422 304136 279478 304192
rect 278778 289040 278834 289096
rect 280342 280200 280398 280256
rect 279422 193840 279478 193896
rect 278778 177112 278834 177168
rect 278042 176704 278098 176760
rect 264978 175616 265034 175672
rect 265070 175208 265126 175264
rect 264978 173984 265034 174040
rect 265714 174800 265770 174856
rect 265070 173576 265126 173632
rect 264978 172624 265034 172680
rect 265070 172216 265126 172272
rect 264978 171400 265034 171456
rect 264978 170992 265034 171048
rect 264242 170040 264298 170096
rect 262862 166912 262918 166968
rect 261482 119312 261538 119368
rect 260746 93608 260802 93664
rect 260378 55120 260434 55176
rect 260378 53896 260434 53952
rect 260102 10240 260158 10296
rect 262770 137536 262826 137592
rect 262770 137128 262826 137184
rect 262678 136312 262734 136368
rect 262678 135768 262734 135824
rect 262770 133184 262826 133240
rect 262770 132776 262826 132832
rect 263138 145560 263194 145616
rect 262862 126928 262918 126984
rect 262862 120672 262918 120728
rect 262954 120264 263010 120320
rect 261666 98640 261722 98696
rect 261850 88984 261906 89040
rect 261574 69536 261630 69592
rect 262954 106392 263010 106448
rect 264978 169632 265034 169688
rect 265070 168816 265126 168872
rect 264978 167864 265034 167920
rect 265070 167456 265126 167512
rect 279330 173712 279386 173768
rect 279330 172216 279386 172272
rect 282182 316648 282238 316704
rect 282182 291896 282238 291952
rect 279422 169088 279478 169144
rect 280250 187176 280306 187232
rect 280066 176432 280122 176488
rect 279882 176024 279938 176080
rect 279606 175752 279662 175808
rect 279606 174256 279662 174312
rect 279514 166776 279570 166832
rect 264978 166232 265034 166288
rect 265622 165824 265678 165880
rect 265070 165280 265126 165336
rect 264978 164872 265034 164928
rect 265254 164056 265310 164112
rect 265070 163648 265126 163704
rect 264978 162868 264980 162888
rect 264980 162868 265032 162888
rect 265032 162868 265034 162888
rect 264978 162832 265034 162868
rect 265070 162288 265126 162344
rect 264978 161508 264980 161528
rect 264980 161508 265032 161528
rect 265032 161508 265034 161528
rect 264978 161472 265034 161508
rect 265070 161064 265126 161120
rect 264978 160656 265034 160712
rect 265070 159704 265126 159760
rect 264978 158888 265034 158944
rect 265070 158480 265126 158536
rect 264978 157664 265034 157720
rect 265070 156712 265126 156768
rect 264978 156304 265034 156360
rect 265162 155896 265218 155952
rect 264978 154536 265034 154592
rect 264978 153720 265034 153776
rect 264978 152904 265034 152960
rect 264334 152496 264390 152552
rect 264978 151136 265034 151192
rect 265070 150728 265126 150784
rect 264978 149912 265034 149968
rect 265070 149640 265126 149696
rect 265162 149504 265218 149560
rect 265070 148960 265126 149016
rect 264978 147756 265034 147792
rect 264978 147736 264980 147756
rect 264980 147736 265032 147756
rect 265032 147736 265034 147756
rect 265070 147328 265126 147384
rect 264978 146396 265034 146432
rect 264978 146376 264980 146396
rect 264980 146376 265032 146396
rect 265032 146376 265034 146396
rect 265070 145968 265126 146024
rect 264978 145152 265034 145208
rect 265162 145696 265218 145752
rect 265070 144744 265126 144800
rect 264978 144336 265034 144392
rect 265162 143792 265218 143848
rect 264610 142568 264666 142624
rect 264334 139168 264390 139224
rect 263138 120808 263194 120864
rect 264242 108704 264298 108760
rect 262954 57160 263010 57216
rect 264978 142180 265034 142216
rect 264978 142160 264980 142180
rect 264980 142160 265032 142180
rect 265032 142160 265034 142180
rect 280250 164872 280306 164928
rect 265806 157120 265862 157176
rect 265990 154128 266046 154184
rect 265714 148552 265770 148608
rect 265162 141344 265218 141400
rect 264978 140820 265034 140856
rect 264978 140800 264980 140820
rect 264980 140800 265032 140820
rect 265032 140800 265034 140820
rect 264978 139984 265034 140040
rect 264978 138624 265034 138680
rect 264978 136992 265034 137048
rect 264978 136176 265034 136232
rect 265070 135632 265126 135688
rect 264978 132640 265034 132696
rect 264426 108568 264482 108624
rect 264334 105168 264390 105224
rect 265070 131824 265126 131880
rect 264978 131416 265034 131472
rect 264978 129648 265034 129704
rect 265622 128424 265678 128480
rect 264978 127880 265034 127936
rect 265070 127084 265126 127120
rect 265070 127064 265072 127084
rect 265072 127064 265124 127084
rect 265124 127064 265126 127084
rect 264978 126248 265034 126304
rect 265070 125296 265126 125352
rect 264978 124480 265034 124536
rect 264978 124072 265034 124128
rect 265070 123664 265126 123720
rect 264978 121896 265034 121952
rect 265070 121080 265126 121136
rect 264978 119720 265034 119776
rect 264978 118496 265034 118552
rect 265070 117136 265126 117192
rect 264978 116320 265034 116376
rect 265070 115504 265126 115560
rect 264978 115096 265034 115152
rect 264978 113736 265034 113792
rect 265254 112512 265310 112568
rect 264978 111968 265034 112024
rect 265070 111560 265126 111616
rect 264978 111152 265034 111208
rect 265070 109928 265126 109984
rect 264978 109520 265034 109576
rect 264978 106936 265034 106992
rect 264978 105984 265034 106040
rect 265070 105576 265126 105632
rect 264978 103808 265034 103864
rect 264978 103400 265034 103456
rect 264518 102720 264574 102776
rect 264886 102584 264942 102640
rect 264978 101768 265034 101824
rect 265070 101224 265126 101280
rect 265070 100000 265126 100056
rect 264978 99592 265034 99648
rect 264978 98640 265034 98696
rect 265070 97824 265126 97880
rect 264978 97008 265034 97064
rect 264886 94560 264942 94616
rect 265806 143384 265862 143440
rect 265714 125840 265770 125896
rect 265898 141752 265954 141808
rect 280342 161064 280398 161120
rect 279330 144744 279386 144800
rect 266082 141208 266138 141264
rect 267002 134408 267058 134464
rect 265898 123392 265954 123448
rect 266266 108976 266322 109032
rect 265806 98232 265862 98288
rect 265806 79328 265862 79384
rect 265714 66816 265770 66872
rect 279330 133320 279386 133376
rect 267094 122848 267150 122904
rect 280158 121352 280214 121408
rect 279330 120128 279386 120184
rect 267646 115912 267702 115968
rect 267186 100408 267242 100464
rect 267738 110336 267794 110392
rect 267186 72528 267242 72584
rect 267094 68176 267150 68232
rect 267002 58520 267058 58576
rect 267830 95512 267886 95568
rect 267738 19216 267794 19272
rect 268382 19216 268438 19272
rect 261758 11600 261814 11656
rect 260102 3576 260158 3632
rect 260654 3576 260710 3632
rect 266358 3304 266414 3360
rect 270498 94560 270554 94616
rect 271878 94424 271934 94480
rect 275926 92248 275982 92304
rect 273994 62736 274050 62792
rect 273258 30232 273314 30288
rect 273902 30232 273958 30288
rect 279330 104216 279386 104272
rect 278042 86128 278098 86184
rect 281446 172896 281502 172952
rect 282366 306584 282422 306640
rect 283194 299648 283250 299704
rect 282274 270544 282330 270600
rect 282918 179424 282974 179480
rect 281814 175480 281870 175536
rect 282826 174664 282882 174720
rect 282734 174256 282790 174312
rect 282826 173984 282882 174040
rect 281814 170856 281870 170912
rect 282826 169360 282882 169416
rect 282826 167864 282882 167920
rect 282734 167048 282790 167104
rect 282826 165552 282882 165608
rect 281814 164092 281816 164112
rect 281816 164092 281868 164112
rect 281868 164092 281870 164112
rect 281814 164056 281870 164092
rect 282182 163240 282238 163296
rect 282826 162560 282882 162616
rect 282274 161744 282330 161800
rect 282642 160248 282698 160304
rect 282826 159432 282882 159488
rect 282734 158752 282790 158808
rect 282090 157936 282146 157992
rect 281722 151816 281778 151872
rect 281906 149640 281962 149696
rect 281722 138932 281724 138952
rect 281724 138932 281776 138952
rect 281776 138932 281778 138952
rect 281722 138896 281778 138932
rect 282550 155660 282552 155680
rect 282552 155660 282604 155680
rect 282604 155660 282606 155680
rect 282550 155624 282606 155660
rect 282826 154128 282882 154184
rect 282366 153448 282422 153504
rect 282826 152632 282882 152688
rect 282734 151136 282790 151192
rect 282826 150340 282882 150376
rect 282826 150320 282828 150340
rect 282828 150320 282880 150340
rect 282880 150320 282882 150340
rect 282734 148824 282790 148880
rect 282826 148008 282882 148064
rect 282826 147328 282882 147384
rect 282734 146512 282790 146568
rect 282826 145832 282882 145888
rect 282550 145016 282606 145072
rect 282458 143520 282514 143576
rect 282826 142704 282882 142760
rect 282826 142060 282828 142080
rect 282828 142060 282880 142080
rect 282880 142060 282882 142080
rect 282826 142024 282882 142060
rect 282734 141208 282790 141264
rect 282826 140392 282882 140448
rect 282642 138216 282698 138272
rect 282826 137400 282882 137456
rect 282182 136584 282238 136640
rect 282826 135904 282882 135960
rect 282826 135088 282882 135144
rect 282458 134408 282514 134464
rect 285586 367104 285642 367160
rect 284298 199960 284354 200016
rect 284298 199416 284354 199472
rect 283562 179968 283618 180024
rect 281630 128968 281686 129024
rect 281538 126792 281594 126848
rect 280434 119176 280490 119232
rect 281630 124480 281686 124536
rect 282826 131280 282882 131336
rect 282274 130600 282330 130656
rect 282642 129784 282698 129840
rect 282826 128288 282882 128344
rect 282826 127472 282882 127528
rect 282826 125976 282882 126032
rect 282182 125160 282238 125216
rect 282090 123664 282146 123720
rect 282642 122984 282698 123040
rect 282826 122168 282882 122224
rect 282826 119856 282882 119912
rect 281722 115368 281778 115424
rect 282826 118360 282882 118416
rect 282826 117544 282882 117600
rect 282826 116864 282882 116920
rect 282274 116048 282330 116104
rect 282458 114552 282514 114608
rect 282274 113736 282330 113792
rect 282826 113092 282828 113112
rect 282828 113092 282880 113112
rect 282880 113092 282882 113112
rect 282826 113056 282882 113092
rect 282826 112240 282882 112296
rect 282274 110744 282330 110800
rect 282826 109248 282882 109304
rect 282182 108432 282238 108488
rect 282366 107752 282422 107808
rect 281630 106936 281686 106992
rect 281814 106120 281870 106176
rect 281722 103164 281724 103184
rect 281724 103164 281776 103184
rect 281776 103164 281778 103184
rect 281722 103128 281778 103164
rect 281722 100816 281778 100872
rect 281906 103944 281962 104000
rect 287058 367512 287114 367568
rect 287058 327120 287114 327176
rect 285586 207576 285642 207632
rect 285034 192616 285090 192672
rect 284574 176432 284630 176488
rect 289726 322768 289782 322824
rect 288530 289856 288586 289912
rect 288438 194384 288494 194440
rect 288714 202136 288770 202192
rect 288714 201492 288716 201512
rect 288716 201492 288768 201512
rect 288768 201492 288770 201512
rect 288714 201456 288770 201492
rect 288714 178744 288770 178800
rect 291842 341536 291898 341592
rect 291198 298696 291254 298752
rect 291290 288496 291346 288552
rect 290002 177384 290058 177440
rect 291382 178608 291438 178664
rect 291290 153720 291346 153776
rect 291106 117136 291162 117192
rect 282826 102312 282882 102368
rect 282826 99320 282882 99376
rect 281998 98504 282054 98560
rect 282826 97824 282882 97880
rect 282734 97008 282790 97064
rect 282826 96328 282882 96384
rect 281630 91024 281686 91080
rect 281630 90344 281686 90400
rect 277490 22616 277546 22672
rect 278686 2624 278742 2680
rect 288346 60424 288402 60480
rect 284390 20576 284446 20632
rect 284942 20576 284998 20632
rect 287794 5616 287850 5672
rect 288346 5616 288402 5672
rect 289082 6704 289138 6760
rect 292486 213832 292542 213888
rect 293222 213832 293278 213888
rect 297362 331200 297418 331256
rect 298006 331220 298062 331256
rect 298006 331200 298008 331220
rect 298008 331200 298060 331220
rect 298060 331200 298062 331220
rect 295338 294480 295394 294536
rect 295246 238312 295302 238368
rect 292670 99320 292726 99376
rect 293222 99320 293278 99376
rect 294234 179968 294290 180024
rect 295982 184320 296038 184376
rect 295338 33088 295394 33144
rect 290186 3440 290242 3496
rect 294878 3440 294934 3496
rect 295890 13640 295946 13696
rect 296074 44784 296130 44840
rect 296074 33088 296130 33144
rect 297362 231920 297418 231976
rect 296902 196696 296958 196752
rect 299570 261296 299626 261352
rect 299478 208120 299534 208176
rect 299478 207576 299534 207632
rect 299386 147736 299442 147792
rect 298742 101360 298798 101416
rect 298098 86944 298154 87000
rect 297362 72392 297418 72448
rect 297362 8200 297418 8256
rect 295982 3848 296038 3904
rect 299754 207712 299810 207768
rect 300122 203632 300178 203688
rect 300122 33768 300178 33824
rect 299662 13116 299718 13152
rect 299662 13096 299664 13116
rect 299664 13096 299716 13116
rect 299716 13096 299718 13116
rect 302882 299512 302938 299568
rect 307758 369008 307814 369064
rect 304998 342216 305054 342272
rect 305642 342216 305698 342272
rect 304998 306448 305054 306504
rect 303618 291080 303674 291136
rect 303618 266328 303674 266384
rect 303618 140820 303674 140856
rect 303618 140800 303620 140820
rect 303620 140800 303672 140820
rect 303672 140800 303674 140820
rect 302882 64096 302938 64152
rect 302974 35128 303030 35184
rect 302974 34584 303030 34640
rect 302882 23296 302938 23352
rect 303526 23296 303582 23352
rect 300122 3848 300178 3904
rect 300766 3440 300822 3496
rect 304262 291080 304318 291136
rect 304262 290400 304318 290456
rect 304446 266328 304502 266384
rect 305090 238720 305146 238776
rect 304998 156032 305054 156088
rect 304262 34584 304318 34640
rect 306470 214512 306526 214568
rect 309046 260072 309102 260128
rect 309046 259392 309102 259448
rect 307114 223624 307170 223680
rect 309874 259392 309930 259448
rect 313278 337320 313334 337376
rect 314658 292576 314714 292632
rect 315118 292576 315174 292632
rect 313462 231104 313518 231160
rect 319626 376624 319682 376680
rect 315302 213152 315358 213208
rect 316682 228248 316738 228304
rect 314014 84768 314070 84824
rect 313922 82764 313924 82784
rect 313924 82764 313976 82784
rect 313976 82764 313978 82784
rect 313922 82728 313978 82764
rect 310518 17856 310574 17912
rect 314014 9560 314070 9616
rect 320178 361664 320234 361720
rect 320822 361664 320878 361720
rect 319442 351192 319498 351248
rect 317418 313248 317474 313304
rect 317326 215056 317382 215112
rect 316774 195336 316830 195392
rect 318798 307808 318854 307864
rect 318154 302232 318210 302288
rect 318246 211112 318302 211168
rect 318062 195200 318118 195256
rect 319442 73752 319498 73808
rect 322294 357992 322350 358048
rect 320914 185680 320970 185736
rect 324686 358128 324742 358184
rect 325606 358128 325662 358184
rect 324686 357448 324742 357504
rect 324318 345616 324374 345672
rect 323030 321544 323086 321600
rect 322202 139440 322258 139496
rect 318522 3304 318578 3360
rect 323674 221448 323730 221504
rect 326342 352552 326398 352608
rect 324962 191120 325018 191176
rect 328458 358128 328514 358184
rect 327078 228928 327134 228984
rect 322202 3712 322258 3768
rect 325054 37848 325110 37904
rect 331862 371864 331918 371920
rect 329102 140800 329158 140856
rect 326342 3984 326398 4040
rect 329102 3304 329158 3360
rect 331954 235320 332010 235376
rect 341154 374584 341210 374640
rect 338026 360984 338082 361040
rect 337382 360168 337438 360224
rect 338026 360168 338082 360224
rect 336094 236000 336150 236056
rect 335358 137672 335414 137728
rect 338118 335416 338174 335472
rect 344282 319368 344338 319424
rect 342994 235184 343050 235240
rect 340970 3440 341026 3496
rect 347042 340040 347098 340096
rect 351182 377304 351238 377360
rect 355322 377576 355378 377632
rect 353942 366288 353998 366344
rect 353298 360032 353354 360088
rect 349802 315288 349858 315344
rect 344282 3440 344338 3496
rect 352562 284960 352618 285016
rect 351182 196560 351238 196616
rect 349802 94424 349858 94480
rect 346950 3304 347006 3360
rect 352654 138624 352710 138680
rect 356242 423680 356298 423736
rect 356334 382336 356390 382392
rect 356334 377576 356390 377632
rect 357162 495488 357218 495544
rect 358726 510040 358782 510096
rect 358726 505164 358782 505200
rect 358726 505144 358728 505164
rect 358728 505144 358780 505164
rect 358780 505144 358782 505164
rect 358726 502696 358782 502752
rect 358634 493040 358690 493096
rect 358726 487736 358782 487792
rect 358082 487192 358138 487248
rect 358082 485288 358138 485344
rect 357898 470620 357954 470656
rect 357898 470600 357900 470620
rect 357900 470600 357952 470620
rect 357952 470600 357954 470620
rect 357438 458360 357494 458416
rect 357530 438912 357586 438968
rect 357438 373224 357494 373280
rect 357898 436328 357954 436384
rect 358726 482840 358782 482896
rect 358726 480392 358782 480448
rect 358726 477944 358782 478000
rect 358542 473048 358598 473104
rect 358726 465704 358782 465760
rect 358450 460808 358506 460864
rect 358726 455912 358782 455968
rect 358726 453464 358782 453520
rect 358726 451016 358782 451072
rect 358726 448704 358782 448760
rect 358726 446120 358782 446176
rect 358726 443672 358782 443728
rect 358726 441224 358782 441280
rect 358726 438932 358782 438968
rect 358726 438912 358728 438932
rect 358728 438912 358780 438932
rect 358780 438912 358782 438932
rect 358726 433880 358782 433936
rect 358726 431432 358782 431488
rect 358726 428984 358782 429040
rect 358726 426536 358782 426592
rect 358726 421640 358782 421696
rect 358726 419192 358782 419248
rect 358726 416780 358728 416800
rect 358728 416780 358780 416800
rect 358780 416780 358782 416800
rect 358726 416744 358782 416780
rect 358726 414296 358782 414352
rect 358726 411848 358782 411904
rect 358726 409400 358782 409456
rect 358726 406952 358782 407008
rect 358726 404232 358782 404288
rect 358726 401784 358782 401840
rect 358634 399336 358690 399392
rect 358726 394440 358782 394496
rect 357622 391992 357678 392048
rect 357714 389544 357770 389600
rect 358726 387096 358782 387152
rect 358726 384648 358782 384704
rect 358634 379752 358690 379808
rect 358082 375128 358138 375184
rect 357530 362208 357586 362264
rect 356150 311072 356206 311128
rect 356794 311072 356850 311128
rect 355322 233144 355378 233200
rect 356794 204856 356850 204912
rect 356702 142432 356758 142488
rect 352562 65456 352618 65512
rect 358910 497800 358966 497856
rect 359002 463256 359058 463312
rect 359094 396888 359150 396944
rect 359462 308352 359518 308408
rect 362958 538192 363014 538248
rect 361854 377304 361910 377360
rect 361762 364928 361818 364984
rect 361486 245656 361542 245712
rect 352562 3984 352618 4040
rect 351642 3848 351698 3904
rect 363234 370640 363290 370696
rect 364338 269728 364394 269784
rect 365994 375944 366050 376000
rect 365902 372544 365958 372600
rect 363694 226888 363750 226944
rect 361486 96464 361542 96520
rect 367374 341400 367430 341456
rect 367742 284824 367798 284880
rect 368662 393372 368718 393408
rect 368662 393352 368664 393372
rect 368664 393352 368716 393372
rect 368716 393352 368718 393372
rect 368662 370504 368718 370560
rect 368570 366288 368626 366344
rect 371422 371864 371478 371920
rect 367742 101224 367798 101280
rect 371974 229064 372030 229120
rect 374642 328752 374698 328808
rect 374734 208936 374790 208992
rect 380990 541184 381046 541240
rect 380898 535608 380954 535664
rect 378874 374584 378930 374640
rect 378138 351056 378194 351112
rect 378782 266192 378838 266248
rect 376758 134408 376814 134464
rect 377402 102720 377458 102776
rect 380990 246200 381046 246256
rect 380898 194520 380954 194576
rect 385130 372680 385186 372736
rect 385682 372680 385738 372736
rect 380898 139304 380954 139360
rect 380898 138624 380954 138680
rect 382922 104080 382978 104136
rect 376022 3848 376078 3904
rect 359462 3304 359518 3360
rect 385682 99592 385738 99648
rect 387062 99456 387118 99512
rect 389822 317464 389878 317520
rect 389178 293936 389234 293992
rect 388442 99184 388498 99240
rect 391202 198056 391258 198112
rect 392674 310528 392730 310584
rect 392582 99728 392638 99784
rect 582654 697176 582710 697232
rect 582562 683848 582618 683904
rect 582378 670656 582434 670712
rect 580354 554784 580410 554840
rect 579894 537784 579950 537840
rect 397458 188264 397514 188320
rect 395986 145560 396042 145616
rect 396722 142296 396778 142352
rect 395526 142160 395582 142216
rect 395434 134408 395490 134464
rect 395434 132640 395490 132696
rect 394054 97688 394110 97744
rect 393962 95104 394018 95160
rect 393318 94424 393374 94480
rect 393318 88168 393374 88224
rect 397366 115776 397422 115832
rect 397550 139340 397552 139360
rect 397552 139340 397604 139360
rect 397604 139340 397606 139360
rect 397550 139304 397606 139340
rect 397918 137264 397974 137320
rect 397642 136176 397698 136232
rect 397550 135360 397606 135416
rect 397642 134680 397698 134736
rect 397550 133456 397606 133512
rect 398470 131688 398526 131744
rect 398654 129648 398710 129704
rect 397550 128968 397606 129024
rect 397550 128152 397606 128208
rect 397550 127064 397606 127120
rect 397550 126268 397606 126304
rect 397550 126248 397552 126268
rect 397552 126248 397604 126268
rect 397604 126248 397606 126268
rect 397550 125160 397606 125216
rect 397642 124344 397698 124400
rect 397550 123256 397606 123312
rect 397550 122304 397606 122360
rect 400770 142160 400826 142216
rect 401690 180784 401746 180840
rect 405738 206352 405794 206408
rect 404358 184184 404414 184240
rect 398838 130872 398894 130928
rect 398194 121352 398250 121408
rect 398746 120536 398802 120592
rect 397550 119720 397606 119776
rect 397550 118532 397552 118552
rect 397552 118532 397604 118552
rect 397604 118532 397606 118552
rect 397550 118496 397606 118532
rect 397642 117816 397698 117872
rect 397550 116728 397606 116784
rect 397550 114824 397606 114880
rect 397550 114008 397606 114064
rect 397642 113056 397698 113112
rect 397734 111968 397790 112024
rect 397458 111288 397514 111344
rect 397550 110200 397606 110256
rect 397458 109248 397514 109304
rect 397458 108160 397514 108216
rect 397550 107480 397606 107536
rect 397458 106664 397514 106720
rect 397458 105576 397514 105632
rect 397458 104796 397460 104816
rect 397460 104796 397512 104816
rect 397512 104796 397514 104816
rect 397458 104760 397514 104796
rect 397642 104080 397698 104136
rect 397458 102856 397514 102912
rect 397458 101632 397514 101688
rect 397550 100816 397606 100872
rect 397458 99320 397514 99376
rect 405830 185544 405886 185600
rect 405922 145560 405978 145616
rect 406290 142432 406346 142488
rect 407210 224168 407266 224224
rect 409878 143384 409934 143440
rect 412638 220088 412694 220144
rect 411994 199280 412050 199336
rect 411442 145560 411498 145616
rect 410890 143384 410946 143440
rect 418802 367104 418858 367160
rect 416778 233280 416834 233336
rect 419906 139576 419962 139632
rect 418710 139440 418766 139496
rect 425702 200776 425758 200832
rect 420918 143384 420974 143440
rect 422114 143384 422170 143440
rect 426438 197920 426494 197976
rect 580354 524456 580410 524512
rect 580262 484608 580318 484664
rect 580262 471416 580318 471472
rect 580354 378392 580410 378448
rect 580262 377984 580318 378040
rect 429198 222808 429254 222864
rect 428462 206216 428518 206272
rect 430578 181328 430634 181384
rect 427818 142296 427874 142352
rect 426530 140800 426586 140856
rect 434718 224984 434774 225040
rect 431958 142160 432014 142216
rect 432970 142160 433026 142216
rect 433982 139984 434038 140040
rect 442998 287136 443054 287192
rect 436190 204312 436246 204368
rect 435362 140800 435418 140856
rect 440238 200640 440294 200696
rect 420550 139712 420606 139768
rect 420550 139440 420606 139496
rect 426898 139440 426954 139496
rect 428738 139440 428794 139496
rect 429474 139440 429530 139496
rect 434994 139440 435050 139496
rect 439042 139440 439098 139496
rect 399850 137672 399906 137728
rect 439962 131960 440018 132016
rect 441710 179696 441766 179752
rect 440330 177248 440386 177304
rect 441618 160656 441674 160712
rect 440514 140800 440570 140856
rect 440422 139984 440478 140040
rect 440422 128696 440478 128752
rect 440422 125840 440478 125896
rect 440330 109112 440386 109168
rect 440238 106392 440294 106448
rect 401414 100680 401470 100736
rect 399482 39208 399538 39264
rect 421654 100680 421710 100736
rect 425058 100680 425114 100736
rect 428646 100680 428702 100736
rect 404450 99728 404506 99784
rect 404542 99592 404598 99648
rect 405554 99592 405610 99648
rect 407578 99320 407634 99376
rect 408590 93744 408646 93800
rect 410062 95240 410118 95296
rect 416410 96464 416466 96520
rect 422114 99456 422170 99512
rect 425886 99456 425942 99512
rect 425426 92384 425482 92440
rect 427818 97688 427874 97744
rect 429658 99184 429714 99240
rect 429842 95784 429898 95840
rect 432602 96872 432658 96928
rect 430670 88168 430726 88224
rect 437202 95104 437258 95160
rect 438490 96872 438546 96928
rect 441710 140800 441766 140856
rect 442170 138216 442226 138272
rect 441986 130600 442042 130656
rect 442906 137128 442962 137184
rect 442906 136176 442962 136232
rect 442906 135088 442962 135144
rect 442906 133220 442908 133240
rect 442908 133220 442960 133240
rect 442960 133220 442962 133240
rect 442906 133184 442962 133220
rect 444470 189760 444526 189816
rect 443182 134408 443238 134464
rect 442906 132404 442908 132424
rect 442908 132404 442960 132424
rect 442960 132404 442962 132424
rect 442906 132368 442962 132404
rect 442906 129648 442962 129704
rect 442906 127744 442962 127800
rect 442906 126656 442962 126712
rect 442906 124108 442908 124128
rect 442908 124108 442960 124128
rect 442960 124108 442962 124128
rect 442906 124072 442962 124108
rect 442814 123256 442870 123312
rect 442998 122032 443054 122088
rect 442906 121352 442962 121408
rect 442630 120264 442686 120320
rect 442906 119448 442962 119504
rect 441710 118632 441766 118688
rect 440514 117544 440570 117600
rect 441710 116592 441766 116648
rect 440514 114688 440570 114744
rect 441618 101632 441674 101688
rect 442906 115504 442962 115560
rect 442354 113736 442410 113792
rect 442170 111696 442226 111752
rect 442354 111016 442410 111072
rect 441802 110064 441858 110120
rect 442906 108160 442962 108216
rect 442538 107208 442594 107264
rect 441986 104352 442042 104408
rect 442906 103536 442962 103592
rect 442722 102584 442778 102640
rect 443090 71712 443146 71768
rect 448518 229744 448574 229800
rect 447322 138624 447378 138680
rect 449898 203496 449954 203552
rect 448610 189624 448666 189680
rect 451278 190984 451334 191040
rect 582470 644000 582526 644056
rect 582470 551248 582526 551304
rect 582470 511264 582526 511320
rect 582562 458088 582618 458144
rect 582470 431568 582526 431624
rect 582378 375264 582434 375320
rect 582378 365064 582434 365120
rect 580170 272176 580226 272232
rect 580906 179152 580962 179208
rect 582470 165824 582526 165880
rect 580170 139304 580226 139360
rect 580170 125976 580226 126032
rect 582930 630808 582986 630864
rect 582746 617480 582802 617536
rect 582838 577632 582894 577688
rect 582746 541592 582802 541648
rect 582746 535472 582802 535528
rect 582654 404912 582710 404968
rect 583022 590960 583078 591016
rect 583114 564304 583170 564360
rect 583114 556144 583170 556200
rect 583758 556144 583814 556200
rect 583114 536832 583170 536888
rect 583114 458088 583170 458144
rect 583022 418240 583078 418296
rect 582930 404912 582986 404968
rect 582838 376624 582894 376680
rect 582930 351872 582986 351928
rect 582838 325216 582894 325272
rect 582746 298696 582802 298752
rect 582838 234640 582894 234696
rect 582746 152632 582802 152688
rect 582654 145560 582710 145616
rect 580170 99456 580226 99512
rect 582470 95240 582526 95296
rect 582378 86128 582434 86184
rect 582378 72936 582434 72992
rect 452658 8200 452714 8256
rect 582654 59608 582710 59664
rect 582746 33088 582802 33144
rect 582562 19760 582618 19816
rect 582470 6568 582526 6624
rect 583666 334600 583722 334656
rect 583022 312024 583078 312080
rect 583022 266192 583078 266248
rect 583022 258848 583078 258904
rect 583114 245520 583170 245576
rect 583298 232328 583354 232384
rect 583114 211112 583170 211168
rect 583114 192480 583170 192536
rect 583022 112784 583078 112840
rect 583206 186904 583262 186960
rect 582930 46280 582986 46336
rect 583390 219000 583446 219056
rect 583574 211112 583630 211168
rect 583482 205400 583538 205456
<< metal3 >>
rect 69606 702476 69612 702540
rect 69676 702538 69682 702540
rect 154113 702538 154179 702541
rect 69676 702536 154179 702538
rect 69676 702480 154118 702536
rect 154174 702480 154179 702536
rect 69676 702478 154179 702480
rect 69676 702476 69682 702478
rect 154113 702475 154179 702478
rect -960 697220 480 697460
rect 582649 697234 582715 697237
rect 583520 697234 584960 697324
rect 582649 697232 584960 697234
rect 582649 697176 582654 697232
rect 582710 697176 584960 697232
rect 582649 697174 584960 697176
rect 582649 697171 582715 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 3417 684314 3483 684317
rect -960 684312 3483 684314
rect -960 684256 3422 684312
rect 3478 684256 3483 684312
rect -960 684254 3483 684256
rect -960 684164 480 684254
rect 3417 684251 3483 684254
rect 582557 683906 582623 683909
rect 583520 683906 584960 683996
rect 582557 683904 584960 683906
rect 582557 683848 582562 683904
rect 582618 683848 584960 683904
rect 582557 683846 584960 683848
rect 582557 683843 582623 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3509 671258 3575 671261
rect -960 671256 3575 671258
rect -960 671200 3514 671256
rect 3570 671200 3575 671256
rect -960 671198 3575 671200
rect -960 671108 480 671198
rect 3509 671195 3575 671198
rect 582373 670714 582439 670717
rect 583520 670714 584960 670804
rect 582373 670712 584960 670714
rect 582373 670656 582378 670712
rect 582434 670656 584960 670712
rect 582373 670654 584960 670656
rect 582373 670651 582439 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 3417 658202 3483 658205
rect -960 658200 3483 658202
rect -960 658144 3422 658200
rect 3478 658144 3483 658200
rect -960 658142 3483 658144
rect -960 658052 480 658142
rect 3417 658139 3483 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 582465 644058 582531 644061
rect 583520 644058 584960 644148
rect 582465 644056 584960 644058
rect 582465 644000 582470 644056
rect 582526 644000 584960 644056
rect 582465 643998 584960 644000
rect 582465 643995 582531 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 3509 632090 3575 632093
rect -960 632088 3575 632090
rect -960 632032 3514 632088
rect 3570 632032 3575 632088
rect -960 632030 3575 632032
rect -960 631940 480 632030
rect 3509 632027 3575 632030
rect 582925 630866 582991 630869
rect 583520 630866 584960 630956
rect 582925 630864 584960 630866
rect 582925 630808 582930 630864
rect 582986 630808 584960 630864
rect 582925 630806 584960 630808
rect 582925 630803 582991 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 3509 619170 3575 619173
rect -960 619168 3575 619170
rect -960 619112 3514 619168
rect 3570 619112 3575 619168
rect -960 619110 3575 619112
rect -960 619020 480 619110
rect 3509 619107 3575 619110
rect 582741 617538 582807 617541
rect 583520 617538 584960 617628
rect 582741 617536 584960 617538
rect 582741 617480 582746 617536
rect 582802 617480 584960 617536
rect 582741 617478 584960 617480
rect 582741 617475 582807 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 3509 606114 3575 606117
rect -960 606112 3575 606114
rect -960 606056 3514 606112
rect 3570 606056 3575 606112
rect -960 606054 3575 606056
rect -960 605964 480 606054
rect 3509 606051 3575 606054
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 74901 592106 74967 592109
rect 96613 592106 96679 592109
rect 74901 592104 96679 592106
rect 74901 592048 74906 592104
rect 74962 592048 96618 592104
rect 96674 592048 96679 592104
rect 74901 592046 96679 592048
rect 74901 592043 74967 592046
rect 96613 592043 96679 592046
rect 77661 591018 77727 591021
rect 97257 591018 97323 591021
rect 77661 591016 97323 591018
rect 77661 590960 77666 591016
rect 77722 590960 97262 591016
rect 97318 590960 97323 591016
rect 77661 590958 97323 590960
rect 77661 590955 77727 590958
rect 97257 590955 97323 590958
rect 583017 591018 583083 591021
rect 583520 591018 584960 591108
rect 583017 591016 584960 591018
rect 583017 590960 583022 591016
rect 583078 590960 584960 591016
rect 583017 590958 584960 590960
rect 583017 590955 583083 590958
rect 82261 590882 82327 590885
rect 95877 590882 95943 590885
rect 82261 590880 95943 590882
rect 82261 590824 82266 590880
rect 82322 590824 95882 590880
rect 95938 590824 95943 590880
rect 583520 590868 584960 590958
rect 82261 590822 95943 590824
rect 82261 590819 82327 590822
rect 95877 590819 95943 590822
rect 66110 590684 66116 590748
rect 66180 590746 66186 590748
rect 70301 590746 70367 590749
rect 71129 590746 71195 590749
rect 66180 590744 71195 590746
rect 66180 590688 70306 590744
rect 70362 590688 71134 590744
rect 71190 590688 71195 590744
rect 66180 590686 71195 590688
rect 66180 590684 66186 590686
rect 70301 590683 70367 590686
rect 71129 590683 71195 590686
rect 70301 589930 70367 589933
rect 90357 589930 90423 589933
rect 70301 589928 90423 589930
rect 70301 589872 70306 589928
rect 70362 589872 90362 589928
rect 90418 589872 90423 589928
rect 70301 589870 90423 589872
rect 70301 589867 70367 589870
rect 90357 589867 90423 589870
rect 83181 589522 83247 589525
rect 111057 589522 111123 589525
rect 83181 589520 111123 589522
rect 83181 589464 83186 589520
rect 83242 589464 111062 589520
rect 111118 589464 111123 589520
rect 83181 589462 111123 589464
rect 83181 589459 83247 589462
rect 111057 589459 111123 589462
rect 81341 589386 81407 589389
rect 93761 589386 93827 589389
rect 255957 589386 256023 589389
rect 81341 589384 256023 589386
rect 81341 589328 81346 589384
rect 81402 589328 93766 589384
rect 93822 589328 255962 589384
rect 256018 589328 256023 589384
rect 81341 589326 256023 589328
rect 81341 589323 81407 589326
rect 93761 589323 93827 589326
rect 255957 589323 256023 589326
rect 72417 588706 72483 588709
rect 93117 588706 93183 588709
rect 72417 588704 93183 588706
rect 72417 588648 72422 588704
rect 72478 588648 93122 588704
rect 93178 588648 93183 588704
rect 72417 588646 93183 588648
rect 72417 588643 72483 588646
rect 93117 588643 93183 588646
rect 88057 588570 88123 588573
rect 88190 588570 88196 588572
rect 88057 588568 88196 588570
rect 88057 588512 88062 588568
rect 88118 588512 88196 588568
rect 88057 588510 88196 588512
rect 88057 588507 88123 588510
rect 88190 588508 88196 588510
rect 88260 588508 88266 588572
rect 66805 588434 66871 588437
rect 66805 588432 68908 588434
rect 66805 588376 66810 588432
rect 66866 588376 68908 588432
rect 66805 588374 68908 588376
rect 66805 588371 66871 588374
rect 91737 587618 91803 587621
rect 88596 587616 91803 587618
rect 88596 587560 91742 587616
rect 91798 587560 91803 587616
rect 88596 587558 91803 587560
rect 91737 587555 91803 587558
rect 66253 586530 66319 586533
rect 66253 586528 66362 586530
rect 66253 586472 66258 586528
rect 66314 586472 66362 586528
rect 66253 586467 66362 586472
rect 66302 586394 66362 586467
rect 68878 586394 68938 587044
rect 66302 586334 68938 586394
rect 89713 586258 89779 586261
rect 88596 586256 89779 586258
rect 88596 586200 89718 586256
rect 89774 586200 89779 586256
rect 88596 586198 89779 586200
rect 89713 586195 89779 586198
rect 66805 585714 66871 585717
rect 66805 585712 68908 585714
rect 66805 585656 66810 585712
rect 66866 585656 68908 585712
rect 66805 585654 68908 585656
rect 66805 585651 66871 585654
rect 88190 585652 88196 585716
rect 88260 585714 88266 585716
rect 119337 585714 119403 585717
rect 88260 585712 119403 585714
rect 88260 585656 119342 585712
rect 119398 585656 119403 585712
rect 88260 585654 119403 585656
rect 88260 585652 88266 585654
rect 119337 585651 119403 585654
rect 91369 584898 91435 584901
rect 88596 584896 91435 584898
rect 88596 584840 91374 584896
rect 91430 584840 91435 584896
rect 88596 584838 91435 584840
rect 91369 584835 91435 584838
rect 67725 584354 67791 584357
rect 67725 584352 68908 584354
rect 67725 584296 67730 584352
rect 67786 584296 68908 584352
rect 67725 584294 68908 584296
rect 67725 584291 67791 584294
rect 91185 583674 91251 583677
rect 88596 583672 91251 583674
rect 88596 583616 91190 583672
rect 91246 583616 91251 583672
rect 88596 583614 91251 583616
rect 91185 583611 91251 583614
rect 66805 582994 66871 582997
rect 66805 582992 68908 582994
rect 66805 582936 66810 582992
rect 66866 582936 68908 582992
rect 66805 582934 68908 582936
rect 66805 582931 66871 582934
rect 69422 582252 69428 582316
rect 69492 582252 69498 582316
rect 66713 581770 66779 581773
rect 69430 581770 69490 582252
rect 91737 582178 91803 582181
rect 88596 582176 91803 582178
rect 88596 582120 91742 582176
rect 91798 582120 91803 582176
rect 88596 582118 91803 582120
rect 91737 582115 91803 582118
rect 66713 581768 69490 581770
rect 66713 581712 66718 581768
rect 66774 581740 69490 581768
rect 66774 581712 69460 581740
rect 66713 581710 69460 581712
rect 66713 581707 66779 581710
rect 91737 580818 91803 580821
rect 88596 580816 91803 580818
rect 88596 580760 91742 580816
rect 91798 580760 91803 580816
rect 88596 580758 91803 580760
rect 91737 580755 91803 580758
rect 66805 580274 66871 580277
rect 66805 580272 68908 580274
rect 66805 580216 66810 580272
rect 66866 580216 68908 580272
rect 66805 580214 68908 580216
rect 66805 580211 66871 580214
rect -960 580002 480 580092
rect 3417 580002 3483 580005
rect -960 580000 3483 580002
rect -960 579944 3422 580000
rect 3478 579944 3483 580000
rect -960 579942 3483 579944
rect -960 579852 480 579942
rect 3417 579939 3483 579942
rect 91737 579458 91803 579461
rect 88596 579456 91803 579458
rect 88596 579400 91742 579456
rect 91798 579400 91803 579456
rect 88596 579398 91803 579400
rect 91737 579395 91803 579398
rect 67817 578914 67883 578917
rect 67817 578912 68908 578914
rect 67817 578856 67822 578912
rect 67878 578856 68908 578912
rect 67817 578854 68908 578856
rect 67817 578851 67883 578854
rect 91134 578098 91140 578100
rect 88596 578038 91140 578098
rect 91134 578036 91140 578038
rect 91204 578036 91210 578100
rect 582833 577690 582899 577693
rect 583520 577690 584960 577780
rect 582833 577688 584960 577690
rect 582833 577632 582838 577688
rect 582894 577632 584960 577688
rect 582833 577630 584960 577632
rect 582833 577627 582899 577630
rect 67541 577554 67607 577557
rect 67541 577552 68908 577554
rect 67541 577496 67546 577552
rect 67602 577496 68908 577552
rect 583520 577540 584960 577630
rect 67541 577494 68908 577496
rect 67541 577491 67607 577494
rect 91093 576738 91159 576741
rect 88596 576736 91159 576738
rect 88596 576680 91098 576736
rect 91154 576680 91159 576736
rect 88596 576678 91159 576680
rect 91093 576675 91159 576678
rect 67449 576194 67515 576197
rect 67449 576192 68908 576194
rect 67449 576136 67454 576192
rect 67510 576136 68908 576192
rect 67449 576134 68908 576136
rect 67449 576131 67515 576134
rect 91093 575378 91159 575381
rect 88596 575376 91159 575378
rect 88596 575320 91098 575376
rect 91154 575320 91159 575376
rect 88596 575318 91159 575320
rect 91093 575315 91159 575318
rect 67357 574970 67423 574973
rect 67357 574968 68908 574970
rect 67357 574912 67362 574968
rect 67418 574912 68908 574968
rect 67357 574910 68908 574912
rect 67357 574907 67423 574910
rect 91093 574018 91159 574021
rect 88596 574016 91159 574018
rect 88596 573960 91098 574016
rect 91154 573960 91159 574016
rect 88596 573958 91159 573960
rect 91093 573955 91159 573958
rect 65977 573474 66043 573477
rect 65977 573472 68908 573474
rect 65977 573416 65982 573472
rect 66038 573416 68908 573472
rect 65977 573414 68908 573416
rect 65977 573411 66043 573414
rect 91185 572658 91251 572661
rect 88596 572656 91251 572658
rect 88596 572600 91190 572656
rect 91246 572600 91251 572656
rect 88596 572598 91251 572600
rect 91185 572595 91251 572598
rect 66805 572114 66871 572117
rect 66805 572112 68908 572114
rect 66805 572056 66810 572112
rect 66866 572056 68908 572112
rect 66805 572054 68908 572056
rect 66805 572051 66871 572054
rect 91093 571434 91159 571437
rect 88596 571432 91159 571434
rect 88596 571376 91098 571432
rect 91154 571376 91159 571432
rect 88596 571374 91159 571376
rect 91093 571371 91159 571374
rect 67357 570754 67423 570757
rect 67357 570752 68908 570754
rect 67357 570696 67362 570752
rect 67418 570696 68908 570752
rect 67357 570694 68908 570696
rect 67357 570691 67423 570694
rect 91093 570074 91159 570077
rect 88596 570072 91159 570074
rect 88596 570016 91098 570072
rect 91154 570016 91159 570072
rect 88596 570014 91159 570016
rect 91093 570011 91159 570014
rect 66805 569394 66871 569397
rect 66805 569392 68908 569394
rect 66805 569336 66810 569392
rect 66866 569336 68908 569392
rect 66805 569334 68908 569336
rect 66805 569331 66871 569334
rect 91093 568714 91159 568717
rect 88596 568712 91159 568714
rect 88596 568656 91098 568712
rect 91154 568656 91159 568712
rect 88596 568654 91159 568656
rect 91093 568651 91159 568654
rect 66805 568034 66871 568037
rect 66805 568032 68908 568034
rect 66805 567976 66810 568032
rect 66866 567976 68908 568032
rect 66805 567974 68908 567976
rect 66805 567971 66871 567974
rect 89805 567354 89871 567357
rect 91461 567354 91527 567357
rect 88596 567352 91527 567354
rect 88596 567296 89810 567352
rect 89866 567296 91466 567352
rect 91522 567296 91527 567352
rect 88596 567294 91527 567296
rect 89805 567291 89871 567294
rect 91461 567291 91527 567294
rect -960 566946 480 567036
rect 3417 566946 3483 566949
rect -960 566944 3483 566946
rect -960 566888 3422 566944
rect 3478 566888 3483 566944
rect -960 566886 3483 566888
rect -960 566796 480 566886
rect 3417 566883 3483 566886
rect 67633 566674 67699 566677
rect 67633 566672 68908 566674
rect 67633 566616 67638 566672
rect 67694 566616 68908 566672
rect 67633 566614 68908 566616
rect 67633 566611 67699 566614
rect 91369 565858 91435 565861
rect 88596 565856 91435 565858
rect 88596 565800 91374 565856
rect 91430 565800 91435 565856
rect 88596 565798 91435 565800
rect 91369 565795 91435 565798
rect 66805 565042 66871 565045
rect 66805 565040 68908 565042
rect 66805 564984 66810 565040
rect 66866 564984 68908 565040
rect 66805 564982 68908 564984
rect 66805 564979 66871 564982
rect 91369 564498 91435 564501
rect 88596 564496 91435 564498
rect 88596 564440 91374 564496
rect 91430 564440 91435 564496
rect 88596 564438 91435 564440
rect 91369 564435 91435 564438
rect 178534 564436 178540 564500
rect 178604 564498 178610 564500
rect 303613 564498 303679 564501
rect 178604 564496 303679 564498
rect 178604 564440 303618 564496
rect 303674 564440 303679 564496
rect 178604 564438 303679 564440
rect 178604 564436 178610 564438
rect 303613 564435 303679 564438
rect 583109 564362 583175 564365
rect 583520 564362 584960 564452
rect 583109 564360 584960 564362
rect 583109 564304 583114 564360
rect 583170 564304 584960 564360
rect 583109 564302 584960 564304
rect 583109 564299 583175 564302
rect 583520 564212 584960 564302
rect 66805 563682 66871 563685
rect 66805 563680 68908 563682
rect 66805 563624 66810 563680
rect 66866 563624 68908 563680
rect 66805 563622 68908 563624
rect 66805 563619 66871 563622
rect 91369 563138 91435 563141
rect 88596 563136 91435 563138
rect 88596 563080 91374 563136
rect 91430 563080 91435 563136
rect 88596 563078 91435 563080
rect 91369 563075 91435 563078
rect 66805 562322 66871 562325
rect 66805 562320 68908 562322
rect 66805 562264 66810 562320
rect 66866 562264 68908 562320
rect 66805 562262 68908 562264
rect 66805 562259 66871 562262
rect 91093 561506 91159 561509
rect 88596 561504 91159 561506
rect 88596 561448 91098 561504
rect 91154 561448 91159 561504
rect 88596 561446 91159 561448
rect 91093 561443 91159 561446
rect 66805 560962 66871 560965
rect 66805 560960 68908 560962
rect 66805 560904 66810 560960
rect 66866 560904 68908 560960
rect 66805 560902 68908 560904
rect 66805 560899 66871 560902
rect 188521 560418 188587 560421
rect 356237 560418 356303 560421
rect 188521 560416 356303 560418
rect 188521 560360 188526 560416
rect 188582 560360 356242 560416
rect 356298 560360 356303 560416
rect 188521 560358 356303 560360
rect 188521 560355 188587 560358
rect 356237 560355 356303 560358
rect 263593 560282 263659 560285
rect 264237 560282 264303 560285
rect 263593 560280 264303 560282
rect 263593 560224 263598 560280
rect 263654 560224 264242 560280
rect 264298 560224 264303 560280
rect 263593 560222 264303 560224
rect 263593 560219 263659 560222
rect 264237 560219 264303 560222
rect 88885 560146 88951 560149
rect 89621 560146 89687 560149
rect 88596 560144 89687 560146
rect 88596 560088 88890 560144
rect 88946 560088 89626 560144
rect 89682 560088 89687 560144
rect 88596 560086 89687 560088
rect 88885 560083 88951 560086
rect 89621 560083 89687 560086
rect 66069 559602 66135 559605
rect 66069 559600 68908 559602
rect 66069 559544 66074 559600
rect 66130 559544 68908 559600
rect 66069 559542 68908 559544
rect 66069 559539 66135 559542
rect 160829 559058 160895 559061
rect 263593 559058 263659 559061
rect 160829 559056 263659 559058
rect 160829 559000 160834 559056
rect 160890 559000 263598 559056
rect 263654 559000 263659 559056
rect 160829 558998 263659 559000
rect 160829 558995 160895 558998
rect 263593 558995 263659 558998
rect 91185 558786 91251 558789
rect 88596 558784 91251 558786
rect 88596 558728 91190 558784
rect 91246 558728 91251 558784
rect 88596 558726 91251 558728
rect 91185 558723 91251 558726
rect 66253 558378 66319 558381
rect 66253 558376 68908 558378
rect 66253 558320 66258 558376
rect 66314 558320 68908 558376
rect 66253 558318 68908 558320
rect 66253 558315 66319 558318
rect 173801 557562 173867 557565
rect 216673 557562 216739 557565
rect 173801 557560 216739 557562
rect 173801 557504 173806 557560
rect 173862 557504 216678 557560
rect 216734 557504 216739 557560
rect 173801 557502 216739 557504
rect 173801 557499 173867 557502
rect 216673 557499 216739 557502
rect 91277 557426 91343 557429
rect 88596 557424 91343 557426
rect 88596 557368 91282 557424
rect 91338 557368 91343 557424
rect 88596 557366 91343 557368
rect 91277 557363 91343 557366
rect 67398 556820 67404 556884
rect 67468 556882 67474 556884
rect 67468 556822 68908 556882
rect 67468 556820 67474 556822
rect 207657 556202 207723 556205
rect 583109 556202 583175 556205
rect 583753 556202 583819 556205
rect 207657 556200 583819 556202
rect 207657 556144 207662 556200
rect 207718 556144 583114 556200
rect 583170 556144 583758 556200
rect 583814 556144 583819 556200
rect 207657 556142 583819 556144
rect 207657 556139 207723 556142
rect 583109 556139 583175 556142
rect 583753 556139 583819 556142
rect 91093 556066 91159 556069
rect 88596 556064 91159 556066
rect 88596 556008 91098 556064
rect 91154 556008 91159 556064
rect 88596 556006 91159 556008
rect 91093 556003 91159 556006
rect 66805 555522 66871 555525
rect 66805 555520 68908 555522
rect 66805 555464 66810 555520
rect 66866 555464 68908 555520
rect 66805 555462 68908 555464
rect 66805 555459 66871 555462
rect 91093 554842 91159 554845
rect 106181 554842 106247 554845
rect 247033 554842 247099 554845
rect 580349 554842 580415 554845
rect 91093 554840 580415 554842
rect 91093 554784 91098 554840
rect 91154 554784 106186 554840
rect 106242 554784 247038 554840
rect 247094 554784 580354 554840
rect 580410 554784 580415 554840
rect 91093 554782 580415 554784
rect 91093 554779 91159 554782
rect 106181 554779 106247 554782
rect 247033 554779 247099 554782
rect 580349 554779 580415 554782
rect 91093 554706 91159 554709
rect 88596 554704 91159 554706
rect 88596 554648 91098 554704
rect 91154 554648 91159 554704
rect 88596 554646 91159 554648
rect 91093 554643 91159 554646
rect 66437 554162 66503 554165
rect 66437 554160 68908 554162
rect 66437 554104 66442 554160
rect 66498 554104 68908 554160
rect 66437 554102 68908 554104
rect 66437 554099 66503 554102
rect 198825 554026 198891 554029
rect 331213 554026 331279 554029
rect 198825 554024 331279 554026
rect -960 553890 480 553980
rect 198825 553968 198830 554024
rect 198886 553968 331218 554024
rect 331274 553968 331279 554024
rect 198825 553966 331279 553968
rect 198825 553963 198891 553966
rect 331213 553963 331279 553966
rect 3325 553890 3391 553893
rect -960 553888 3391 553890
rect -960 553832 3330 553888
rect 3386 553832 3391 553888
rect -960 553830 3391 553832
rect -960 553740 480 553830
rect 3325 553827 3391 553830
rect 186221 553482 186287 553485
rect 235257 553482 235323 553485
rect 186221 553480 235323 553482
rect 186221 553424 186226 553480
rect 186282 553424 235262 553480
rect 235318 553424 235323 553480
rect 186221 553422 235323 553424
rect 186221 553419 186287 553422
rect 235257 553419 235323 553422
rect 92105 553346 92171 553349
rect 88596 553344 92171 553346
rect 88596 553288 92110 553344
rect 92166 553288 92171 553344
rect 88596 553286 92171 553288
rect 92105 553283 92171 553286
rect 67449 552802 67515 552805
rect 67449 552800 68908 552802
rect 67449 552744 67454 552800
rect 67510 552744 68908 552800
rect 67449 552742 68908 552744
rect 67449 552739 67515 552742
rect 91093 552122 91159 552125
rect 88596 552120 91159 552122
rect 88596 552064 91098 552120
rect 91154 552064 91159 552120
rect 88596 552062 91159 552064
rect 91093 552059 91159 552062
rect 191649 552122 191715 552125
rect 285121 552122 285187 552125
rect 191649 552120 285187 552122
rect 191649 552064 191654 552120
rect 191710 552064 285126 552120
rect 285182 552064 285187 552120
rect 191649 552062 285187 552064
rect 191649 552059 191715 552062
rect 285121 552059 285187 552062
rect 66662 551380 66668 551444
rect 66732 551442 66738 551444
rect 66732 551382 68908 551442
rect 66732 551380 66738 551382
rect 198590 551244 198596 551308
rect 198660 551306 198666 551308
rect 582465 551306 582531 551309
rect 198660 551304 582531 551306
rect 198660 551248 582470 551304
rect 582526 551248 582531 551304
rect 198660 551246 582531 551248
rect 198660 551244 198666 551246
rect 582465 551243 582531 551246
rect 583520 551020 584960 551260
rect 91093 550762 91159 550765
rect 88596 550760 91159 550762
rect 88596 550704 91098 550760
rect 91154 550704 91159 550760
rect 88596 550702 91159 550704
rect 91093 550699 91159 550702
rect 184790 550700 184796 550764
rect 184860 550762 184866 550764
rect 262213 550762 262279 550765
rect 184860 550760 262279 550762
rect 184860 550704 262218 550760
rect 262274 550704 262279 550760
rect 184860 550702 262279 550704
rect 184860 550700 184866 550702
rect 262213 550699 262279 550702
rect 66805 550082 66871 550085
rect 66805 550080 68908 550082
rect 66805 550024 66810 550080
rect 66866 550024 68908 550080
rect 66805 550022 68908 550024
rect 66805 550019 66871 550022
rect 177389 549538 177455 549541
rect 290089 549538 290155 549541
rect 177389 549536 290155 549538
rect 177389 549480 177394 549536
rect 177450 549480 290094 549536
rect 290150 549480 290155 549536
rect 177389 549478 290155 549480
rect 177389 549475 177455 549478
rect 290089 549475 290155 549478
rect 91093 549402 91159 549405
rect 88596 549400 91159 549402
rect 88596 549344 91098 549400
rect 91154 549344 91159 549400
rect 88596 549342 91159 549344
rect 91093 549339 91159 549342
rect 126881 549402 126947 549405
rect 339953 549402 340019 549405
rect 126881 549400 340019 549402
rect 126881 549344 126886 549400
rect 126942 549344 339958 549400
rect 340014 549344 340019 549400
rect 126881 549342 340019 549344
rect 126881 549339 126947 549342
rect 339953 549339 340019 549342
rect 66805 548722 66871 548725
rect 66805 548720 68908 548722
rect 66805 548664 66810 548720
rect 66866 548664 68908 548720
rect 66805 548662 68908 548664
rect 66805 548659 66871 548662
rect 91369 548042 91435 548045
rect 88596 548040 91435 548042
rect 88596 547984 91374 548040
rect 91430 547984 91435 548040
rect 88596 547982 91435 547984
rect 91369 547979 91435 547982
rect 91093 547906 91159 547909
rect 95141 547906 95207 547909
rect 278037 547906 278103 547909
rect 91093 547904 278103 547906
rect 91093 547848 91098 547904
rect 91154 547848 95146 547904
rect 95202 547848 278042 547904
rect 278098 547848 278103 547904
rect 91093 547846 278103 547848
rect 91093 547843 91159 547846
rect 95141 547843 95207 547846
rect 278037 547843 278103 547846
rect 66897 547362 66963 547365
rect 66897 547360 68908 547362
rect 66897 547304 66902 547360
rect 66958 547304 68908 547360
rect 66897 547302 68908 547304
rect 66897 547299 66963 547302
rect 170254 546620 170260 546684
rect 170324 546682 170330 546684
rect 225321 546682 225387 546685
rect 170324 546680 225387 546682
rect 170324 546624 225326 546680
rect 225382 546624 225387 546680
rect 170324 546622 225387 546624
rect 170324 546620 170330 546622
rect 225321 546619 225387 546622
rect 91277 546546 91343 546549
rect 91553 546546 91619 546549
rect 88596 546544 91619 546546
rect 88596 546488 91282 546544
rect 91338 546488 91558 546544
rect 91614 546488 91619 546544
rect 88596 546486 91619 546488
rect 91277 546483 91343 546486
rect 91553 546483 91619 546486
rect 137921 546546 137987 546549
rect 300025 546546 300091 546549
rect 137921 546544 300091 546546
rect 137921 546488 137926 546544
rect 137982 546488 300030 546544
rect 300086 546488 300091 546544
rect 137921 546486 300091 546488
rect 137921 546483 137987 546486
rect 300025 546483 300091 546486
rect 316585 546546 316651 546549
rect 358854 546546 358860 546548
rect 316585 546544 358860 546546
rect 316585 546488 316590 546544
rect 316646 546488 358860 546544
rect 316585 546486 358860 546488
rect 316585 546483 316651 546486
rect 358854 546484 358860 546486
rect 358924 546484 358930 546548
rect 66897 546002 66963 546005
rect 66897 546000 68908 546002
rect 66897 545944 66902 546000
rect 66958 545944 68908 546000
rect 66897 545942 68908 545944
rect 66897 545939 66963 545942
rect 192569 545458 192635 545461
rect 206277 545458 206343 545461
rect 192569 545456 206343 545458
rect 192569 545400 192574 545456
rect 192630 545400 206282 545456
rect 206338 545400 206343 545456
rect 192569 545398 206343 545400
rect 192569 545395 192635 545398
rect 206277 545395 206343 545398
rect 180149 545322 180215 545325
rect 230473 545322 230539 545325
rect 180149 545320 230539 545322
rect 180149 545264 180154 545320
rect 180210 545264 230478 545320
rect 230534 545264 230539 545320
rect 180149 545262 230539 545264
rect 180149 545259 180215 545262
rect 230473 545259 230539 545262
rect 91093 545186 91159 545189
rect 88596 545184 91159 545186
rect 88596 545128 91098 545184
rect 91154 545128 91159 545184
rect 88596 545126 91159 545128
rect 91093 545123 91159 545126
rect 195329 545186 195395 545189
rect 248505 545186 248571 545189
rect 195329 545184 248571 545186
rect 195329 545128 195334 545184
rect 195390 545128 248510 545184
rect 248566 545128 248571 545184
rect 195329 545126 248571 545128
rect 195329 545123 195395 545126
rect 248505 545123 248571 545126
rect 66897 544642 66963 544645
rect 66897 544640 68908 544642
rect 66897 544584 66902 544640
rect 66958 544584 68908 544640
rect 66897 544582 68908 544584
rect 66897 544579 66963 544582
rect 196801 543962 196867 543965
rect 243537 543962 243603 543965
rect 196801 543960 243603 543962
rect 196801 543904 196806 543960
rect 196862 543904 243542 543960
rect 243598 543904 243603 543960
rect 196801 543902 243603 543904
rect 196801 543899 196867 543902
rect 243537 543899 243603 543902
rect 97901 543826 97967 543829
rect 353937 543826 354003 543829
rect 88596 543824 354003 543826
rect 88596 543768 97906 543824
rect 97962 543768 353942 543824
rect 353998 543768 354003 543824
rect 88596 543766 354003 543768
rect 97901 543763 97967 543766
rect 353937 543763 354003 543766
rect 66897 543282 66963 543285
rect 66897 543280 68908 543282
rect 66897 543224 66902 543280
rect 66958 543224 68908 543280
rect 66897 543222 68908 543224
rect 66897 543219 66963 543222
rect 201401 542738 201467 542741
rect 218697 542738 218763 542741
rect 201401 542736 218763 542738
rect 201401 542680 201406 542736
rect 201462 542680 218702 542736
rect 218758 542680 218763 542736
rect 201401 542678 218763 542680
rect 201401 542675 201467 542678
rect 218697 542675 218763 542678
rect 197854 542540 197860 542604
rect 197924 542602 197930 542604
rect 253933 542602 253999 542605
rect 197924 542600 253999 542602
rect 197924 542544 253938 542600
rect 253994 542544 253999 542600
rect 197924 542542 253999 542544
rect 197924 542540 197930 542542
rect 253933 542539 253999 542542
rect 91093 542466 91159 542469
rect 88596 542464 91159 542466
rect 88596 542408 91098 542464
rect 91154 542408 91159 542464
rect 88596 542406 91159 542408
rect 91093 542403 91159 542406
rect 195237 542466 195303 542469
rect 356145 542466 356211 542469
rect 195237 542464 356211 542466
rect 195237 542408 195242 542464
rect 195298 542408 356150 542464
rect 356206 542408 356211 542464
rect 195237 542406 356211 542408
rect 195237 542403 195303 542406
rect 356145 542403 356211 542406
rect 65977 542330 66043 542333
rect 69422 542330 69428 542332
rect 65977 542328 69428 542330
rect 65977 542272 65982 542328
rect 66038 542272 69428 542328
rect 65977 542270 69428 542272
rect 65977 542267 66043 542270
rect 69422 542268 69428 542270
rect 69492 542268 69498 542332
rect 91134 542268 91140 542332
rect 91204 542330 91210 542332
rect 92381 542330 92447 542333
rect 91204 542328 92447 542330
rect 91204 542272 92386 542328
rect 92442 542272 92447 542328
rect 91204 542270 92447 542272
rect 91204 542268 91210 542270
rect 92381 542267 92447 542270
rect 207013 542330 207079 542333
rect 207657 542330 207723 542333
rect 207013 542328 207723 542330
rect 207013 542272 207018 542328
rect 207074 542272 207662 542328
rect 207718 542272 207723 542328
rect 207013 542270 207723 542272
rect 207013 542267 207079 542270
rect 207657 542267 207723 542270
rect 66989 541922 67055 541925
rect 66989 541920 68908 541922
rect 66989 541864 66994 541920
rect 67050 541864 68908 541920
rect 66989 541862 68908 541864
rect 66989 541859 67055 541862
rect 582741 541650 582807 541653
rect 383610 541648 582807 541650
rect 383610 541592 582746 541648
rect 582802 541592 582807 541648
rect 383610 541590 582807 541592
rect 320173 541378 320239 541381
rect 353334 541378 353340 541380
rect 320173 541376 353340 541378
rect 320173 541320 320178 541376
rect 320234 541320 353340 541376
rect 320173 541318 353340 541320
rect 320173 541315 320239 541318
rect 353334 541316 353340 541318
rect 353404 541316 353410 541380
rect 91093 541242 91159 541245
rect 88596 541240 91159 541242
rect 88596 541184 91098 541240
rect 91154 541184 91159 541240
rect 88596 541182 91159 541184
rect 91093 541179 91159 541182
rect 199326 541180 199332 541244
rect 199396 541242 199402 541244
rect 207013 541242 207079 541245
rect 199396 541240 207079 541242
rect 199396 541184 207018 541240
rect 207074 541184 207079 541240
rect 199396 541182 207079 541184
rect 199396 541180 199402 541182
rect 207013 541179 207079 541182
rect 255957 541242 256023 541245
rect 257337 541242 257403 541245
rect 380985 541242 381051 541245
rect 383610 541242 383670 541590
rect 582741 541587 582807 541590
rect 255957 541240 383670 541242
rect 255957 541184 255962 541240
rect 256018 541184 257342 541240
rect 257398 541184 380990 541240
rect 381046 541184 383670 541240
rect 255957 541182 383670 541184
rect 255957 541179 256023 541182
rect 257337 541179 257403 541182
rect 380985 541179 381051 541182
rect 184841 541106 184907 541109
rect 348233 541106 348299 541109
rect 184841 541104 348299 541106
rect 184841 541048 184846 541104
rect 184902 541048 348238 541104
rect 348294 541048 348299 541104
rect 184841 541046 348299 541048
rect 184841 541043 184907 541046
rect 348233 541043 348299 541046
rect -960 540684 480 540924
rect 67541 539610 67607 539613
rect 69430 539610 69490 540532
rect 341517 540290 341583 540293
rect 357617 540290 357683 540293
rect 341517 540288 357683 540290
rect 341517 540232 341522 540288
rect 341578 540232 357622 540288
rect 357678 540232 357683 540288
rect 341517 540230 357683 540232
rect 341517 540227 341583 540230
rect 357617 540227 357683 540230
rect 88793 540154 88859 540157
rect 323669 540154 323735 540157
rect 88793 540152 323735 540154
rect 88793 540096 88798 540152
rect 88854 540096 323674 540152
rect 323730 540096 323735 540152
rect 88793 540094 323735 540096
rect 88793 540091 88859 540094
rect 323669 540091 323735 540094
rect 91093 539746 91159 539749
rect 88596 539744 91159 539746
rect 88596 539688 91098 539744
rect 91154 539688 91159 539744
rect 88596 539686 91159 539688
rect 91093 539683 91159 539686
rect 185342 539684 185348 539748
rect 185412 539746 185418 539748
rect 307109 539746 307175 539749
rect 185412 539744 307175 539746
rect 185412 539688 307114 539744
rect 307170 539688 307175 539744
rect 185412 539686 307175 539688
rect 185412 539684 185418 539686
rect 307109 539683 307175 539686
rect 345381 539610 345447 539613
rect 349981 539610 350047 539613
rect 67541 539608 74550 539610
rect 67541 539552 67546 539608
rect 67602 539552 74550 539608
rect 67541 539550 74550 539552
rect 67541 539547 67607 539550
rect 74490 538794 74550 539550
rect 345381 539608 350047 539610
rect 345381 539552 345386 539608
rect 345442 539552 349986 539608
rect 350042 539552 350047 539608
rect 345381 539550 350047 539552
rect 345381 539547 345447 539550
rect 349981 539547 350047 539550
rect 124857 538794 124923 538797
rect 74490 538792 124923 538794
rect 74490 538736 124862 538792
rect 124918 538736 124923 538792
rect 74490 538734 124923 538736
rect 124857 538731 124923 538734
rect 266353 538794 266419 538797
rect 273989 538794 274055 538797
rect 266353 538792 274055 538794
rect 266353 538736 266358 538792
rect 266414 538736 273994 538792
rect 274050 538736 274055 538792
rect 266353 538734 274055 538736
rect 266353 538731 266419 538734
rect 273989 538731 274055 538734
rect 196566 538596 196572 538660
rect 196636 538658 196642 538660
rect 204069 538658 204135 538661
rect 196636 538656 204135 538658
rect 196636 538600 204074 538656
rect 204130 538600 204135 538656
rect 196636 538598 204135 538600
rect 196636 538596 196642 538598
rect 204069 538595 204135 538598
rect 202781 538522 202847 538525
rect 222469 538522 222535 538525
rect 202781 538520 222535 538522
rect 202781 538464 202786 538520
rect 202842 538464 222474 538520
rect 222530 538464 222535 538520
rect 202781 538462 222535 538464
rect 202781 538459 202847 538462
rect 222469 538459 222535 538462
rect 194358 538324 194364 538388
rect 194428 538386 194434 538388
rect 255589 538386 255655 538389
rect 194428 538384 255655 538386
rect 194428 538328 255594 538384
rect 255650 538328 255655 538384
rect 194428 538326 255655 538328
rect 194428 538324 194434 538326
rect 255589 538323 255655 538326
rect 350349 538386 350415 538389
rect 358813 538386 358879 538389
rect 350349 538384 358879 538386
rect 350349 538328 350354 538384
rect 350410 538328 358818 538384
rect 358874 538328 358879 538384
rect 350349 538326 358879 538328
rect 350349 538323 350415 538326
rect 358813 538323 358879 538326
rect 204161 538250 204227 538253
rect 265525 538250 265591 538253
rect 204161 538248 265591 538250
rect 204161 538192 204166 538248
rect 204222 538192 265530 538248
rect 265586 538192 265591 538248
rect 204161 538190 265591 538192
rect 204161 538187 204227 538190
rect 265525 538187 265591 538190
rect 337101 538250 337167 538253
rect 362953 538250 363019 538253
rect 337101 538248 363019 538250
rect 337101 538192 337106 538248
rect 337162 538192 362958 538248
rect 363014 538192 363019 538248
rect 337101 538190 363019 538192
rect 337101 538187 337167 538190
rect 362953 538187 363019 538190
rect 579889 537842 579955 537845
rect 583520 537842 584960 537932
rect 579889 537840 584960 537842
rect 579889 537784 579894 537840
rect 579950 537784 584960 537840
rect 579889 537782 584960 537784
rect 579889 537779 579955 537782
rect 583520 537692 584960 537782
rect 67081 537434 67147 537437
rect 67398 537434 67404 537436
rect 67081 537432 67404 537434
rect 67081 537376 67086 537432
rect 67142 537376 67404 537432
rect 67081 537374 67404 537376
rect 67081 537371 67147 537374
rect 67398 537372 67404 537374
rect 67468 537372 67474 537436
rect 178769 537162 178835 537165
rect 233877 537162 233943 537165
rect 178769 537160 233943 537162
rect 178769 537104 178774 537160
rect 178830 537104 233882 537160
rect 233938 537104 233943 537160
rect 178769 537102 233943 537104
rect 178769 537099 178835 537102
rect 233877 537099 233943 537102
rect 142889 537026 142955 537029
rect 353661 537026 353727 537029
rect 142889 537024 353727 537026
rect 142889 536968 142894 537024
rect 142950 536968 353666 537024
rect 353722 536968 353727 537024
rect 142889 536966 353727 536968
rect 142889 536963 142955 536966
rect 353661 536963 353727 536966
rect 206277 536890 206343 536893
rect 583109 536890 583175 536893
rect 206277 536888 583175 536890
rect 206277 536832 206282 536888
rect 206338 536832 583114 536888
rect 583170 536832 583175 536888
rect 206277 536830 583175 536832
rect 206277 536827 206343 536830
rect 583109 536827 583175 536830
rect 66161 536754 66227 536757
rect 76741 536754 76807 536757
rect 66161 536752 76807 536754
rect 66161 536696 66166 536752
rect 66222 536696 76746 536752
rect 76802 536696 76807 536752
rect 66161 536694 76807 536696
rect 66161 536691 66227 536694
rect 76741 536691 76807 536694
rect 75177 536618 75243 536621
rect 133137 536618 133203 536621
rect 75177 536616 133203 536618
rect 75177 536560 75182 536616
rect 75238 536560 133142 536616
rect 133198 536560 133203 536616
rect 75177 536558 133203 536560
rect 75177 536555 75243 536558
rect 133137 536555 133203 536558
rect 14457 536074 14523 536077
rect 45461 536074 45527 536077
rect 73153 536074 73219 536077
rect 14457 536072 73219 536074
rect 14457 536016 14462 536072
rect 14518 536016 45466 536072
rect 45522 536016 73158 536072
rect 73214 536016 73219 536072
rect 14457 536014 73219 536016
rect 14457 536011 14523 536014
rect 45461 536011 45527 536014
rect 73153 536011 73219 536014
rect 201309 536074 201375 536077
rect 208669 536074 208735 536077
rect 201309 536072 208735 536074
rect 201309 536016 201314 536072
rect 201370 536016 208674 536072
rect 208730 536016 208735 536072
rect 201309 536014 208735 536016
rect 201309 536011 201375 536014
rect 208669 536011 208735 536014
rect 199745 535938 199811 535941
rect 201401 535938 201467 535941
rect 199745 535936 201467 535938
rect 199745 535880 199750 535936
rect 199806 535880 201406 535936
rect 201462 535880 201467 535936
rect 199745 535878 201467 535880
rect 199745 535875 199811 535878
rect 201401 535875 201467 535878
rect 160737 535802 160803 535805
rect 313365 535802 313431 535805
rect 160737 535800 313431 535802
rect 160737 535744 160742 535800
rect 160798 535744 313370 535800
rect 313426 535744 313431 535800
rect 160737 535742 313431 535744
rect 160737 535739 160803 535742
rect 313365 535739 313431 535742
rect 80053 535666 80119 535669
rect 308397 535666 308463 535669
rect 80053 535664 308463 535666
rect 80053 535608 80058 535664
rect 80114 535608 308402 535664
rect 308458 535608 308463 535664
rect 80053 535606 308463 535608
rect 80053 535603 80119 535606
rect 308397 535603 308463 535606
rect 342253 535666 342319 535669
rect 380893 535666 380959 535669
rect 342253 535664 380959 535666
rect 342253 535608 342258 535664
rect 342314 535608 380898 535664
rect 380954 535608 380959 535664
rect 342253 535606 380959 535608
rect 342253 535603 342319 535606
rect 380893 535603 380959 535606
rect 69565 535532 69631 535533
rect 69565 535530 69612 535532
rect 69520 535528 69612 535530
rect 69520 535472 69570 535528
rect 69520 535470 69612 535472
rect 69565 535468 69612 535470
rect 69676 535468 69682 535532
rect 70485 535530 70551 535533
rect 72325 535532 72391 535533
rect 71630 535530 71636 535532
rect 70485 535528 71636 535530
rect 70485 535472 70490 535528
rect 70546 535472 71636 535528
rect 70485 535470 71636 535472
rect 69565 535467 69631 535468
rect 70485 535467 70551 535470
rect 71630 535468 71636 535470
rect 71700 535468 71706 535532
rect 72325 535530 72372 535532
rect 72280 535528 72372 535530
rect 72280 535472 72330 535528
rect 72280 535470 72372 535472
rect 72325 535468 72372 535470
rect 72436 535468 72442 535532
rect 84285 535530 84351 535533
rect 90449 535530 90515 535533
rect 84285 535528 90515 535530
rect 84285 535472 84290 535528
rect 84346 535472 90454 535528
rect 90510 535472 90515 535528
rect 84285 535470 90515 535472
rect 72325 535467 72391 535468
rect 84285 535467 84351 535470
rect 90449 535467 90515 535470
rect 199510 535468 199516 535532
rect 199580 535530 199586 535532
rect 200389 535530 200455 535533
rect 199580 535528 200455 535530
rect 199580 535472 200394 535528
rect 200450 535472 200455 535528
rect 199580 535470 200455 535472
rect 199580 535468 199586 535470
rect 200389 535467 200455 535470
rect 200614 535468 200620 535532
rect 200684 535530 200690 535532
rect 202045 535530 202111 535533
rect 200684 535528 202111 535530
rect 200684 535472 202050 535528
rect 202106 535472 202111 535528
rect 200684 535470 202111 535472
rect 200684 535468 200690 535470
rect 202045 535467 202111 535470
rect 302325 535530 302391 535533
rect 582741 535530 582807 535533
rect 302325 535528 582807 535530
rect 302325 535472 302330 535528
rect 302386 535472 582746 535528
rect 582802 535472 582807 535528
rect 302325 535470 582807 535472
rect 302325 535467 302391 535470
rect 582741 535467 582807 535470
rect 148409 535394 148475 535397
rect 148961 535394 149027 535397
rect 201401 535394 201467 535397
rect 221089 535394 221155 535397
rect 148409 535392 201467 535394
rect 148409 535336 148414 535392
rect 148470 535336 148966 535392
rect 149022 535336 201406 535392
rect 201462 535336 201467 535392
rect 148409 535334 201467 535336
rect 148409 535331 148475 535334
rect 148961 535331 149027 535334
rect 201401 535331 201467 535334
rect 209730 535392 221155 535394
rect 209730 535336 221094 535392
rect 221150 535336 221155 535392
rect 209730 535334 221155 535336
rect 188337 534986 188403 534989
rect 209730 534986 209790 535334
rect 221089 535331 221155 535334
rect 354673 535394 354739 535397
rect 354673 535392 355610 535394
rect 354673 535336 354678 535392
rect 354734 535336 355610 535392
rect 354673 535334 355610 535336
rect 354673 535331 354739 535334
rect 188337 534984 209790 534986
rect 188337 534928 188342 534984
rect 188398 534928 209790 534984
rect 188337 534926 209790 534928
rect 188337 534923 188403 534926
rect 355550 534684 355610 535334
rect 197353 534578 197419 534581
rect 197353 534576 200100 534578
rect 197353 534520 197358 534576
rect 197414 534520 200100 534576
rect 197353 534518 200100 534520
rect 197353 534515 197419 534518
rect 53741 533354 53807 533357
rect 199745 533354 199811 533357
rect 53741 533352 199811 533354
rect 53741 533296 53746 533352
rect 53802 533296 199750 533352
rect 199806 533296 199811 533352
rect 53741 533294 199811 533296
rect 53741 533291 53807 533294
rect 199745 533291 199811 533294
rect 175089 532538 175155 532541
rect 200062 532538 200068 532540
rect 175089 532536 200068 532538
rect 175089 532480 175094 532536
rect 175150 532480 200068 532536
rect 175089 532478 200068 532480
rect 175089 532475 175155 532478
rect 200062 532476 200068 532478
rect 200132 532476 200138 532540
rect 197353 532266 197419 532269
rect 197353 532264 200100 532266
rect 197353 532208 197358 532264
rect 197414 532208 200100 532264
rect 197353 532206 200100 532208
rect 197353 532203 197419 532206
rect 357893 532130 357959 532133
rect 358721 532130 358787 532133
rect 356132 532128 358787 532130
rect 356132 532072 357898 532128
rect 357954 532072 358726 532128
rect 358782 532072 358787 532128
rect 356132 532070 358787 532072
rect 357893 532067 357959 532070
rect 358721 532067 358787 532070
rect 97993 531452 98059 531453
rect 97942 531450 97948 531452
rect 97902 531390 97948 531450
rect 98012 531448 98059 531452
rect 98054 531392 98059 531448
rect 97942 531388 97948 531390
rect 98012 531388 98059 531392
rect 97993 531387 98059 531388
rect 197353 529818 197419 529821
rect 198641 529818 198707 529821
rect 197353 529816 200100 529818
rect 197353 529760 197358 529816
rect 197414 529760 198646 529816
rect 198702 529760 200100 529816
rect 197353 529758 200100 529760
rect 197353 529755 197419 529758
rect 198641 529755 198707 529758
rect 358721 529682 358787 529685
rect 356132 529680 358787 529682
rect 356132 529624 358726 529680
rect 358782 529624 358787 529680
rect 356132 529622 358787 529624
rect 358721 529619 358787 529622
rect -960 527914 480 528004
rect 3417 527914 3483 527917
rect -960 527912 3483 527914
rect -960 527856 3422 527912
rect 3478 527856 3483 527912
rect -960 527854 3483 527856
rect -960 527764 480 527854
rect 3417 527851 3483 527854
rect 197353 527370 197419 527373
rect 197353 527368 200100 527370
rect 197353 527312 197358 527368
rect 197414 527312 200100 527368
rect 197353 527310 200100 527312
rect 197353 527307 197419 527310
rect 358721 527234 358787 527237
rect 356132 527232 358787 527234
rect 356132 527176 358726 527232
rect 358782 527176 358787 527232
rect 356132 527174 358787 527176
rect 358721 527171 358787 527174
rect 169017 526418 169083 526421
rect 197854 526418 197860 526420
rect 169017 526416 197860 526418
rect 169017 526360 169022 526416
rect 169078 526360 197860 526416
rect 169017 526358 197860 526360
rect 169017 526355 169083 526358
rect 197854 526356 197860 526358
rect 197924 526356 197930 526420
rect 197353 524786 197419 524789
rect 358721 524786 358787 524789
rect 197353 524784 200100 524786
rect 197353 524728 197358 524784
rect 197414 524728 200100 524784
rect 197353 524726 200100 524728
rect 356132 524784 358787 524786
rect 356132 524728 358726 524784
rect 358782 524728 358787 524784
rect 356132 524726 358787 524728
rect 197353 524723 197419 524726
rect 358721 524723 358787 524726
rect 580349 524514 580415 524517
rect 583520 524514 584960 524604
rect 580349 524512 584960 524514
rect 580349 524456 580354 524512
rect 580410 524456 584960 524512
rect 580349 524454 584960 524456
rect 580349 524451 580415 524454
rect 583520 524364 584960 524454
rect 168966 523636 168972 523700
rect 169036 523698 169042 523700
rect 199510 523698 199516 523700
rect 169036 523638 199516 523698
rect 169036 523636 169042 523638
rect 199510 523636 199516 523638
rect 199580 523636 199586 523700
rect 66662 522956 66668 523020
rect 66732 523018 66738 523020
rect 67081 523018 67147 523021
rect 356237 523018 356303 523021
rect 66732 523016 67147 523018
rect 66732 522960 67086 523016
rect 67142 522960 67147 523016
rect 66732 522958 67147 522960
rect 66732 522956 66738 522958
rect 67081 522955 67147 522958
rect 356102 523016 356303 523018
rect 356102 522960 356242 523016
rect 356298 522960 356303 523016
rect 356102 522958 356303 522960
rect 66478 522820 66484 522884
rect 66548 522882 66554 522884
rect 66897 522882 66963 522885
rect 66548 522880 66963 522882
rect 66548 522824 66902 522880
rect 66958 522824 66963 522880
rect 66548 522822 66963 522824
rect 66548 522820 66554 522822
rect 66897 522819 66963 522822
rect 197353 522338 197419 522341
rect 356102 522338 356162 522958
rect 356237 522955 356303 522958
rect 358721 522338 358787 522341
rect 197353 522336 200100 522338
rect 197353 522280 197358 522336
rect 197414 522280 200100 522336
rect 356102 522336 358787 522338
rect 356102 522308 358726 522336
rect 197353 522278 200100 522280
rect 356132 522280 358726 522308
rect 358782 522280 358787 522336
rect 356132 522278 358787 522280
rect 197353 522275 197419 522278
rect 358721 522275 358787 522278
rect 357617 519890 357683 519893
rect 358721 519890 358787 519893
rect 356132 519888 358787 519890
rect 161974 518876 161980 518940
rect 162044 518938 162050 518940
rect 200070 518938 200130 519860
rect 356132 519832 357622 519888
rect 357678 519832 358726 519888
rect 358782 519832 358787 519888
rect 356132 519830 358787 519832
rect 357617 519827 357683 519830
rect 358721 519827 358787 519830
rect 162044 518878 200130 518938
rect 162044 518876 162050 518878
rect 50981 518122 51047 518125
rect 191782 518122 191788 518124
rect 50981 518120 191788 518122
rect 50981 518064 50986 518120
rect 51042 518064 191788 518120
rect 50981 518062 191788 518064
rect 50981 518059 51047 518062
rect 191782 518060 191788 518062
rect 191852 518122 191858 518124
rect 192569 518122 192635 518125
rect 191852 518120 192635 518122
rect 191852 518064 192574 518120
rect 192630 518064 192635 518120
rect 191852 518062 192635 518064
rect 191852 518060 191858 518062
rect 192569 518059 192635 518062
rect 50797 517578 50863 517581
rect 50981 517578 51047 517581
rect 50797 517576 51047 517578
rect 50797 517520 50802 517576
rect 50858 517520 50986 517576
rect 51042 517520 51047 517576
rect 50797 517518 51047 517520
rect 50797 517515 50863 517518
rect 50981 517515 51047 517518
rect 197353 517442 197419 517445
rect 358721 517442 358787 517445
rect 197353 517440 200100 517442
rect 197353 517384 197358 517440
rect 197414 517384 200100 517440
rect 197353 517382 200100 517384
rect 356132 517440 358787 517442
rect 356132 517384 358726 517440
rect 358782 517384 358787 517440
rect 356132 517382 358787 517384
rect 197353 517379 197419 517382
rect 358721 517379 358787 517382
rect 197353 514994 197419 514997
rect 358077 514994 358143 514997
rect 197353 514992 200100 514994
rect -960 514858 480 514948
rect 197353 514936 197358 514992
rect 197414 514936 200100 514992
rect 197353 514934 200100 514936
rect 356132 514992 358143 514994
rect 356132 514936 358082 514992
rect 358138 514936 358143 514992
rect 356132 514934 358143 514936
rect 197353 514931 197419 514934
rect 358077 514931 358143 514934
rect 3509 514858 3575 514861
rect -960 514856 3575 514858
rect -960 514800 3514 514856
rect 3570 514800 3575 514856
rect -960 514798 3575 514800
rect -960 514708 480 514798
rect 3509 514795 3575 514798
rect 141417 513362 141483 513365
rect 142061 513362 142127 513365
rect 199326 513362 199332 513364
rect 141417 513360 199332 513362
rect 141417 513304 141422 513360
rect 141478 513304 142066 513360
rect 142122 513304 199332 513360
rect 141417 513302 199332 513304
rect 141417 513299 141483 513302
rect 142061 513299 142127 513302
rect 199326 513300 199332 513302
rect 199396 513300 199402 513364
rect 357433 512682 357499 512685
rect 356132 512680 357499 512682
rect 356132 512624 357438 512680
rect 357494 512624 357499 512680
rect 356132 512622 357499 512624
rect 357433 512619 357499 512622
rect 197997 512546 198063 512549
rect 197997 512544 200100 512546
rect 197997 512488 198002 512544
rect 198058 512488 200100 512544
rect 197997 512486 200100 512488
rect 197997 512483 198063 512486
rect 582465 511322 582531 511325
rect 583520 511322 584960 511412
rect 582465 511320 584960 511322
rect 582465 511264 582470 511320
rect 582526 511264 584960 511320
rect 582465 511262 584960 511264
rect 582465 511259 582531 511262
rect 583520 511172 584960 511262
rect 197353 510234 197419 510237
rect 197353 510232 200100 510234
rect 197353 510176 197358 510232
rect 197414 510176 200100 510232
rect 197353 510174 200100 510176
rect 197353 510171 197419 510174
rect 358721 510098 358787 510101
rect 356132 510096 358787 510098
rect 356132 510040 358726 510096
rect 358782 510040 358787 510096
rect 356132 510038 358787 510040
rect 358721 510035 358787 510038
rect 197353 507650 197419 507653
rect 356697 507650 356763 507653
rect 197353 507648 200100 507650
rect 197353 507592 197358 507648
rect 197414 507592 200100 507648
rect 197353 507590 200100 507592
rect 356132 507648 356763 507650
rect 356132 507592 356702 507648
rect 356758 507592 356763 507648
rect 356132 507590 356763 507592
rect 197353 507587 197419 507590
rect 356697 507587 356763 507590
rect 198733 505202 198799 505205
rect 358721 505202 358787 505205
rect 198733 505200 200100 505202
rect 198733 505144 198738 505200
rect 198794 505144 200100 505200
rect 198733 505142 200100 505144
rect 356132 505200 358787 505202
rect 356132 505144 358726 505200
rect 358782 505144 358787 505200
rect 356132 505142 358787 505144
rect 198733 505139 198799 505142
rect 358721 505139 358787 505142
rect 358721 502754 358787 502757
rect 356132 502752 358787 502754
rect 188838 502420 188844 502484
rect 188908 502482 188914 502484
rect 200070 502482 200130 502724
rect 356132 502696 358726 502752
rect 358782 502696 358787 502752
rect 356132 502694 358787 502696
rect 358721 502691 358787 502694
rect 188908 502422 200130 502482
rect 188908 502420 188914 502422
rect -960 501802 480 501892
rect 3509 501802 3575 501805
rect -960 501800 3575 501802
rect -960 501744 3514 501800
rect 3570 501744 3575 501800
rect -960 501742 3575 501744
rect -960 501652 480 501742
rect 3509 501739 3575 501742
rect 198273 500442 198339 500445
rect 198590 500442 198596 500444
rect 198273 500440 198596 500442
rect 198273 500384 198278 500440
rect 198334 500384 198596 500440
rect 198273 500382 198596 500384
rect 198273 500379 198339 500382
rect 198590 500380 198596 500382
rect 198660 500442 198666 500444
rect 198660 500382 200100 500442
rect 198660 500380 198666 500382
rect 356102 499900 356162 500276
rect 356094 499836 356100 499900
rect 356164 499836 356170 499900
rect 197353 497858 197419 497861
rect 358905 497858 358971 497861
rect 197353 497856 200100 497858
rect 197353 497800 197358 497856
rect 197414 497800 200100 497856
rect 197353 497798 200100 497800
rect 356132 497856 358971 497858
rect 356132 497800 358910 497856
rect 358966 497800 358971 497856
rect 583520 497844 584960 498084
rect 356132 497798 358971 497800
rect 197353 497795 197419 497798
rect 358905 497795 358971 497798
rect 356237 496090 356303 496093
rect 356102 496088 356303 496090
rect 356102 496032 356242 496088
rect 356298 496032 356303 496088
rect 356102 496030 356303 496032
rect 197353 495546 197419 495549
rect 356102 495546 356162 496030
rect 356237 496027 356303 496030
rect 357157 495546 357223 495549
rect 197353 495544 200100 495546
rect 197353 495488 197358 495544
rect 197414 495488 200100 495544
rect 356102 495544 357223 495546
rect 356102 495516 357162 495544
rect 197353 495486 200100 495488
rect 356132 495488 357162 495516
rect 357218 495488 357223 495544
rect 356132 495486 357223 495488
rect 197353 495483 197419 495486
rect 357157 495483 357223 495486
rect 358629 493098 358695 493101
rect 356132 493096 358695 493098
rect 356132 493068 358634 493096
rect 356102 493040 358634 493068
rect 358690 493040 358695 493096
rect 356102 493038 358695 493040
rect 197353 492962 197419 492965
rect 197353 492960 200100 492962
rect 197353 492904 197358 492960
rect 197414 492904 200100 492960
rect 197353 492902 200100 492904
rect 197353 492899 197419 492902
rect 356102 492690 356162 493038
rect 358629 493035 358695 493038
rect 356237 492690 356303 492693
rect 356102 492688 356303 492690
rect 356102 492632 356242 492688
rect 356298 492632 356303 492688
rect 356102 492630 356303 492632
rect 356237 492627 356303 492630
rect 195094 490452 195100 490516
rect 195164 490514 195170 490516
rect 195164 490454 200100 490514
rect 195164 490452 195170 490454
rect 356329 490378 356395 490381
rect 356132 490376 356395 490378
rect 356132 490320 356334 490376
rect 356390 490320 356395 490376
rect 356132 490318 356395 490320
rect 356329 490315 356395 490318
rect -960 488596 480 488836
rect 197353 488202 197419 488205
rect 197353 488200 200100 488202
rect 197353 488144 197358 488200
rect 197414 488144 200100 488200
rect 197353 488142 200100 488144
rect 197353 488139 197419 488142
rect 358721 487794 358787 487797
rect 356132 487792 358787 487794
rect 356132 487736 358726 487792
rect 358782 487736 358787 487792
rect 356132 487734 358787 487736
rect 358721 487731 358787 487734
rect 358077 487250 358143 487253
rect 361614 487250 361620 487252
rect 358077 487248 361620 487250
rect 358077 487192 358082 487248
rect 358138 487192 361620 487248
rect 358077 487190 361620 487192
rect 358077 487187 358143 487190
rect 361614 487188 361620 487190
rect 361684 487188 361690 487252
rect 197353 485618 197419 485621
rect 197353 485616 200100 485618
rect 197353 485560 197358 485616
rect 197414 485560 200100 485616
rect 197353 485558 200100 485560
rect 197353 485555 197419 485558
rect 358077 485346 358143 485349
rect 356132 485344 358143 485346
rect 356132 485288 358082 485344
rect 358138 485288 358143 485344
rect 356132 485286 358143 485288
rect 358077 485283 358143 485286
rect 580257 484666 580323 484669
rect 583520 484666 584960 484756
rect 580257 484664 584960 484666
rect 580257 484608 580262 484664
rect 580318 484608 584960 484664
rect 580257 484606 584960 484608
rect 580257 484603 580323 484606
rect 583520 484516 584960 484606
rect 198406 483108 198412 483172
rect 198476 483170 198482 483172
rect 198476 483110 200100 483170
rect 198476 483108 198482 483110
rect 358721 482898 358787 482901
rect 356132 482896 358787 482898
rect 356132 482840 358726 482896
rect 358782 482840 358787 482896
rect 356132 482838 358787 482840
rect 358721 482835 358787 482838
rect 197353 480722 197419 480725
rect 197353 480720 200100 480722
rect 197353 480664 197358 480720
rect 197414 480664 200100 480720
rect 197353 480662 200100 480664
rect 197353 480659 197419 480662
rect 358721 480450 358787 480453
rect 356132 480448 358787 480450
rect 356132 480392 358726 480448
rect 358782 480392 358787 480448
rect 356132 480390 358787 480392
rect 358721 480387 358787 480390
rect 101489 479498 101555 479501
rect 122598 479498 122604 479500
rect 101489 479496 122604 479498
rect 101489 479440 101494 479496
rect 101550 479440 122604 479496
rect 101489 479438 122604 479440
rect 101489 479435 101555 479438
rect 122598 479436 122604 479438
rect 122668 479436 122674 479500
rect 197353 478274 197419 478277
rect 197353 478272 200100 478274
rect 197353 478216 197358 478272
rect 197414 478216 200100 478272
rect 197353 478214 200100 478216
rect 197353 478211 197419 478214
rect 358721 478002 358787 478005
rect 356132 478000 358787 478002
rect 356132 477944 358726 478000
rect 358782 477944 358787 478000
rect 356132 477942 358787 477944
rect 358721 477939 358787 477942
rect 197353 475826 197419 475829
rect 197353 475824 200100 475826
rect -960 475690 480 475780
rect 197353 475768 197358 475824
rect 197414 475768 200100 475824
rect 197353 475766 200100 475768
rect 197353 475763 197419 475766
rect 3325 475690 3391 475693
rect -960 475688 3391 475690
rect -960 475632 3330 475688
rect 3386 475632 3391 475688
rect -960 475630 3391 475632
rect -960 475540 480 475630
rect 3325 475627 3391 475630
rect 356646 475554 356652 475556
rect 356132 475494 356652 475554
rect 356646 475492 356652 475494
rect 356716 475492 356722 475556
rect 197353 473378 197419 473381
rect 197353 473376 200100 473378
rect 197353 473320 197358 473376
rect 197414 473320 200100 473376
rect 197353 473318 200100 473320
rect 197353 473315 197419 473318
rect 358537 473106 358603 473109
rect 356132 473104 358603 473106
rect 356132 473048 358542 473104
rect 358598 473048 358603 473104
rect 356132 473046 358603 473048
rect 358537 473043 358603 473046
rect 580257 471474 580323 471477
rect 583520 471474 584960 471564
rect 580257 471472 584960 471474
rect 580257 471416 580262 471472
rect 580318 471416 584960 471472
rect 580257 471414 584960 471416
rect 580257 471411 580323 471414
rect 583520 471324 584960 471414
rect 97901 471202 97967 471205
rect 106406 471202 106412 471204
rect 97901 471200 106412 471202
rect 97901 471144 97906 471200
rect 97962 471144 106412 471200
rect 97901 471142 106412 471144
rect 97901 471139 97967 471142
rect 106406 471140 106412 471142
rect 106476 471140 106482 471204
rect 197261 470930 197327 470933
rect 197261 470928 200100 470930
rect 197261 470872 197266 470928
rect 197322 470872 200100 470928
rect 197261 470870 200100 470872
rect 197261 470867 197327 470870
rect 357893 470658 357959 470661
rect 356132 470656 357959 470658
rect 356132 470600 357898 470656
rect 357954 470600 357959 470656
rect 356132 470598 357959 470600
rect 357893 470595 357959 470598
rect 95877 469842 95943 469845
rect 104934 469842 104940 469844
rect 95877 469840 104940 469842
rect 95877 469784 95882 469840
rect 95938 469784 104940 469840
rect 95877 469782 104940 469784
rect 95877 469779 95943 469782
rect 104934 469780 104940 469782
rect 105004 469780 105010 469844
rect 104249 468482 104315 468485
rect 115974 468482 115980 468484
rect 104249 468480 115980 468482
rect 104249 468424 104254 468480
rect 104310 468424 115980 468480
rect 104249 468422 115980 468424
rect 104249 468419 104315 468422
rect 115974 468420 115980 468422
rect 116044 468420 116050 468484
rect 197353 468482 197419 468485
rect 197353 468480 200100 468482
rect 197353 468424 197358 468480
rect 197414 468424 200100 468480
rect 197353 468422 200100 468424
rect 197353 468419 197419 468422
rect 356102 467938 356162 468180
rect 356278 467938 356284 467940
rect 356102 467878 356284 467938
rect 356278 467876 356284 467878
rect 356348 467876 356354 467940
rect 197353 466034 197419 466037
rect 197353 466032 200100 466034
rect 197353 465976 197358 466032
rect 197414 465976 200100 466032
rect 197353 465974 200100 465976
rect 197353 465971 197419 465974
rect 86217 465762 86283 465765
rect 91134 465762 91140 465764
rect 86217 465760 91140 465762
rect 86217 465704 86222 465760
rect 86278 465704 91140 465760
rect 86217 465702 91140 465704
rect 86217 465699 86283 465702
rect 91134 465700 91140 465702
rect 91204 465700 91210 465764
rect 358721 465762 358787 465765
rect 356132 465760 358787 465762
rect 356132 465704 358726 465760
rect 358782 465704 358787 465760
rect 356132 465702 358787 465704
rect 358721 465699 358787 465702
rect 81433 464402 81499 464405
rect 89662 464402 89668 464404
rect 81433 464400 89668 464402
rect 81433 464344 81438 464400
rect 81494 464344 89668 464400
rect 81433 464342 89668 464344
rect 81433 464339 81499 464342
rect 89662 464340 89668 464342
rect 89732 464340 89738 464404
rect 94589 464402 94655 464405
rect 107694 464402 107700 464404
rect 94589 464400 107700 464402
rect 94589 464344 94594 464400
rect 94650 464344 107700 464400
rect 94589 464342 107700 464344
rect 94589 464339 94655 464342
rect 107694 464340 107700 464342
rect 107764 464340 107770 464404
rect 108389 464402 108455 464405
rect 117998 464402 118004 464404
rect 108389 464400 118004 464402
rect 108389 464344 108394 464400
rect 108450 464344 118004 464400
rect 108389 464342 118004 464344
rect 108389 464339 108455 464342
rect 117998 464340 118004 464342
rect 118068 464340 118074 464404
rect 197353 463314 197419 463317
rect 198825 463314 198891 463317
rect 358997 463314 359063 463317
rect 197353 463312 200100 463314
rect 197353 463256 197358 463312
rect 197414 463256 198830 463312
rect 198886 463256 200100 463312
rect 197353 463254 200100 463256
rect 356132 463312 359063 463314
rect 356132 463256 359002 463312
rect 359058 463256 359063 463312
rect 356132 463254 359063 463256
rect 197353 463251 197419 463254
rect 198825 463251 198891 463254
rect 358997 463251 359063 463254
rect 82813 462906 82879 462909
rect 92606 462906 92612 462908
rect 82813 462904 92612 462906
rect 82813 462848 82818 462904
rect 82874 462848 92612 462904
rect 82813 462846 92612 462848
rect 82813 462843 82879 462846
rect 92606 462844 92612 462846
rect 92676 462844 92682 462908
rect -960 462634 480 462724
rect 3509 462634 3575 462637
rect -960 462632 3575 462634
rect -960 462576 3514 462632
rect 3570 462576 3575 462632
rect -960 462574 3575 462576
rect -960 462484 480 462574
rect 3509 462571 3575 462574
rect 197353 460866 197419 460869
rect 358445 460866 358511 460869
rect 197353 460864 200100 460866
rect 197353 460808 197358 460864
rect 197414 460808 200100 460864
rect 197353 460806 200100 460808
rect 356132 460864 358511 460866
rect 356132 460808 358450 460864
rect 358506 460808 358511 460864
rect 356132 460806 358511 460808
rect 197353 460803 197419 460806
rect 358445 460803 358511 460806
rect 95141 460186 95207 460189
rect 111742 460186 111748 460188
rect 95141 460184 111748 460186
rect 95141 460128 95146 460184
rect 95202 460128 111748 460184
rect 95141 460126 111748 460128
rect 95141 460123 95207 460126
rect 111742 460124 111748 460126
rect 111812 460124 111818 460188
rect 90449 459642 90515 459645
rect 93894 459642 93900 459644
rect 90449 459640 93900 459642
rect 90449 459584 90454 459640
rect 90510 459584 93900 459640
rect 90449 459582 93900 459584
rect 90449 459579 90515 459582
rect 93894 459580 93900 459582
rect 93964 459580 93970 459644
rect 112529 458826 112595 458829
rect 118734 458826 118740 458828
rect 112529 458824 118740 458826
rect 112529 458768 112534 458824
rect 112590 458768 118740 458824
rect 112529 458766 118740 458768
rect 112529 458763 112595 458766
rect 118734 458764 118740 458766
rect 118804 458764 118810 458828
rect 197353 458418 197419 458421
rect 198774 458418 198780 458420
rect 197353 458416 198780 458418
rect 197353 458360 197358 458416
rect 197414 458360 198780 458416
rect 197353 458358 198780 458360
rect 197353 458355 197419 458358
rect 198774 458356 198780 458358
rect 198844 458418 198850 458420
rect 357433 458418 357499 458421
rect 198844 458358 200100 458418
rect 356132 458416 357499 458418
rect 356132 458360 357438 458416
rect 357494 458360 357499 458416
rect 356132 458358 357499 458360
rect 198844 458356 198850 458358
rect 357433 458355 357499 458358
rect 582557 458146 582623 458149
rect 583109 458146 583175 458149
rect 583520 458146 584960 458236
rect 582557 458144 584960 458146
rect 582557 458088 582562 458144
rect 582618 458088 583114 458144
rect 583170 458088 584960 458144
rect 582557 458086 584960 458088
rect 582557 458083 582623 458086
rect 583109 458083 583175 458086
rect 583520 457996 584960 458086
rect 88333 457466 88399 457469
rect 100702 457466 100708 457468
rect 88333 457464 100708 457466
rect 88333 457408 88338 457464
rect 88394 457408 100708 457464
rect 88333 457406 100708 457408
rect 88333 457403 88399 457406
rect 100702 457404 100708 457406
rect 100772 457404 100778 457468
rect 104157 457058 104223 457061
rect 108982 457058 108988 457060
rect 104157 457056 108988 457058
rect 104157 457000 104162 457056
rect 104218 457000 108988 457056
rect 104157 456998 108988 457000
rect 104157 456995 104223 456998
rect 108982 456996 108988 456998
rect 109052 456996 109058 457060
rect 69013 456922 69079 456925
rect 69790 456922 69796 456924
rect 69013 456920 69796 456922
rect 69013 456864 69018 456920
rect 69074 456864 69796 456920
rect 69013 456862 69796 456864
rect 69013 456859 69079 456862
rect 69790 456860 69796 456862
rect 69860 456922 69866 456924
rect 155217 456922 155283 456925
rect 69860 456920 155283 456922
rect 69860 456864 155222 456920
rect 155278 456864 155283 456920
rect 69860 456862 155283 456864
rect 69860 456860 69866 456862
rect 155217 456859 155283 456862
rect 87137 456106 87203 456109
rect 98126 456106 98132 456108
rect 87137 456104 98132 456106
rect 87137 456048 87142 456104
rect 87198 456048 98132 456104
rect 87137 456046 98132 456048
rect 87137 456043 87203 456046
rect 98126 456044 98132 456046
rect 98196 456044 98202 456108
rect 101581 456106 101647 456109
rect 102174 456106 102180 456108
rect 101581 456104 102180 456106
rect 101581 456048 101586 456104
rect 101642 456048 102180 456104
rect 101581 456046 102180 456048
rect 101581 456043 101647 456046
rect 102174 456044 102180 456046
rect 102244 456044 102250 456108
rect 198549 455970 198615 455973
rect 358721 455970 358787 455973
rect 198549 455968 200100 455970
rect 198549 455912 198554 455968
rect 198610 455912 200100 455968
rect 198549 455910 200100 455912
rect 356132 455968 358787 455970
rect 356132 455912 358726 455968
rect 358782 455912 358787 455968
rect 356132 455910 358787 455912
rect 198549 455907 198615 455910
rect 358721 455907 358787 455910
rect 82813 455426 82879 455429
rect 172237 455426 172303 455429
rect 82813 455424 172303 455426
rect 82813 455368 82818 455424
rect 82874 455368 172242 455424
rect 172298 455368 172303 455424
rect 82813 455366 172303 455368
rect 82813 455363 82879 455366
rect 172237 455363 172303 455366
rect 198641 453522 198707 453525
rect 358721 453522 358787 453525
rect 198641 453520 200100 453522
rect 198641 453464 198646 453520
rect 198702 453464 200100 453520
rect 198641 453462 200100 453464
rect 356132 453520 358787 453522
rect 356132 453464 358726 453520
rect 358782 453464 358787 453520
rect 356132 453462 358787 453464
rect 198641 453459 198707 453462
rect 358721 453459 358787 453462
rect 61837 453250 61903 453253
rect 75177 453250 75243 453253
rect 61837 453248 75243 453250
rect 61837 453192 61842 453248
rect 61898 453192 75182 453248
rect 75238 453192 75243 453248
rect 61837 453190 75243 453192
rect 61837 453187 61903 453190
rect 75177 453187 75243 453190
rect 86861 453250 86927 453253
rect 96654 453250 96660 453252
rect 86861 453248 96660 453250
rect 86861 453192 86866 453248
rect 86922 453192 96660 453248
rect 86861 453190 96660 453192
rect 86861 453187 86927 453190
rect 96654 453188 96660 453190
rect 96724 453188 96730 453252
rect 98637 451346 98703 451349
rect 153837 451346 153903 451349
rect 98637 451344 153903 451346
rect 98637 451288 98642 451344
rect 98698 451288 153842 451344
rect 153898 451288 153903 451344
rect 98637 451286 153903 451288
rect 98637 451283 98703 451286
rect 153837 451283 153903 451286
rect 358721 451074 358787 451077
rect 356132 451072 358787 451074
rect 66110 450468 66116 450532
rect 66180 450530 66186 450532
rect 91553 450530 91619 450533
rect 66180 450528 93870 450530
rect 66180 450472 91558 450528
rect 91614 450472 93870 450528
rect 66180 450470 93870 450472
rect 66180 450468 66186 450470
rect 91553 450467 91619 450470
rect 93810 450122 93870 450470
rect 171777 450122 171843 450125
rect 93810 450120 171843 450122
rect 93810 450064 171782 450120
rect 171838 450064 171843 450120
rect 93810 450062 171843 450064
rect 171777 450059 171843 450062
rect 160686 449924 160692 449988
rect 160756 449986 160762 449988
rect 200070 449986 200130 451044
rect 356132 451016 358726 451072
rect 358782 451016 358787 451072
rect 356132 451014 358787 451016
rect 358721 451011 358787 451014
rect 160756 449926 200130 449986
rect 160756 449924 160762 449926
rect -960 449578 480 449668
rect 3141 449578 3207 449581
rect -960 449576 3207 449578
rect -960 449520 3146 449576
rect 3202 449520 3207 449576
rect -960 449518 3207 449520
rect -960 449428 480 449518
rect 3141 449515 3207 449518
rect 92381 449170 92447 449173
rect 120206 449170 120212 449172
rect 92381 449168 120212 449170
rect 92381 449112 92386 449168
rect 92442 449112 120212 449168
rect 92381 449110 120212 449112
rect 92381 449107 92447 449110
rect 120206 449108 120212 449110
rect 120276 449108 120282 449172
rect 358721 448762 358787 448765
rect 356132 448760 358787 448762
rect 356132 448704 358726 448760
rect 358782 448704 358787 448760
rect 356132 448702 358787 448704
rect 358721 448699 358787 448702
rect 72693 448628 72759 448629
rect 72693 448624 72740 448628
rect 72804 448626 72810 448628
rect 197353 448626 197419 448629
rect 72693 448568 72698 448624
rect 72693 448564 72740 448568
rect 72804 448566 72850 448626
rect 197353 448624 200100 448626
rect 197353 448568 197358 448624
rect 197414 448568 200100 448624
rect 197353 448566 200100 448568
rect 72804 448564 72810 448566
rect 72693 448563 72759 448564
rect 197353 448563 197419 448566
rect 50797 447810 50863 447813
rect 80881 447810 80947 447813
rect 50797 447808 80947 447810
rect 50797 447752 50802 447808
rect 50858 447752 80886 447808
rect 80942 447752 80947 447808
rect 50797 447750 80947 447752
rect 50797 447747 50863 447750
rect 80881 447747 80947 447750
rect 84193 447810 84259 447813
rect 95182 447810 95188 447812
rect 84193 447808 95188 447810
rect 84193 447752 84198 447808
rect 84254 447752 95188 447808
rect 84193 447750 95188 447752
rect 84193 447747 84259 447750
rect 95182 447748 95188 447750
rect 95252 447748 95258 447812
rect 108297 447810 108363 447813
rect 123017 447810 123083 447813
rect 108297 447808 123083 447810
rect 108297 447752 108302 447808
rect 108358 447752 123022 447808
rect 123078 447752 123083 447808
rect 108297 447750 123083 447752
rect 108297 447747 108363 447750
rect 123017 447747 123083 447750
rect 93025 447130 93091 447133
rect 142889 447130 142955 447133
rect 93025 447128 142955 447130
rect 93025 447072 93030 447128
rect 93086 447072 142894 447128
rect 142950 447072 142955 447128
rect 93025 447070 142955 447072
rect 93025 447067 93091 447070
rect 142889 447067 142955 447070
rect 116117 446450 116183 446453
rect 140773 446450 140839 446453
rect 116117 446448 140839 446450
rect 116117 446392 116122 446448
rect 116178 446392 140778 446448
rect 140834 446392 140839 446448
rect 116117 446390 140839 446392
rect 116117 446387 116183 446390
rect 140773 446387 140839 446390
rect 194542 446388 194548 446452
rect 194612 446450 194618 446452
rect 195789 446450 195855 446453
rect 194612 446448 195855 446450
rect 194612 446392 195794 446448
rect 195850 446392 195855 446448
rect 194612 446390 195855 446392
rect 194612 446388 194618 446390
rect 195789 446387 195855 446390
rect 197353 446178 197419 446181
rect 358721 446178 358787 446181
rect 197353 446176 200100 446178
rect 197353 446120 197358 446176
rect 197414 446120 200100 446176
rect 197353 446118 200100 446120
rect 356132 446176 358787 446178
rect 356132 446120 358726 446176
rect 358782 446120 358787 446176
rect 356132 446118 358787 446120
rect 197353 446115 197419 446118
rect 358721 446115 358787 446118
rect 60641 445770 60707 445773
rect 85573 445770 85639 445773
rect 60641 445768 85639 445770
rect 60641 445712 60646 445768
rect 60702 445712 85578 445768
rect 85634 445712 85639 445768
rect 60641 445710 85639 445712
rect 60641 445707 60707 445710
rect 85573 445707 85639 445710
rect 96470 445708 96476 445772
rect 96540 445770 96546 445772
rect 96613 445770 96679 445773
rect 97625 445770 97691 445773
rect 96540 445768 97691 445770
rect 96540 445712 96618 445768
rect 96674 445712 97630 445768
rect 97686 445712 97691 445768
rect 96540 445710 97691 445712
rect 96540 445708 96546 445710
rect 96613 445707 96679 445710
rect 97625 445707 97691 445710
rect 100518 445708 100524 445772
rect 100588 445770 100594 445772
rect 102133 445770 102199 445773
rect 100588 445768 102199 445770
rect 100588 445712 102138 445768
rect 102194 445712 102199 445768
rect 100588 445710 102199 445712
rect 100588 445708 100594 445710
rect 102133 445707 102199 445710
rect 113173 445770 113239 445773
rect 114369 445770 114435 445773
rect 113173 445768 114435 445770
rect 113173 445712 113178 445768
rect 113234 445712 114374 445768
rect 114430 445712 114435 445768
rect 113173 445710 114435 445712
rect 113173 445707 113239 445710
rect 114369 445707 114435 445710
rect 115197 445770 115263 445773
rect 115790 445770 115796 445772
rect 115197 445768 115796 445770
rect 115197 445712 115202 445768
rect 115258 445712 115796 445768
rect 115197 445710 115796 445712
rect 115197 445707 115263 445710
rect 115790 445708 115796 445710
rect 115860 445708 115866 445772
rect 117589 445770 117655 445773
rect 118601 445772 118667 445773
rect 118550 445770 118556 445772
rect 117589 445768 118556 445770
rect 118620 445768 118667 445772
rect 117589 445712 117594 445768
rect 117650 445712 118556 445768
rect 118662 445712 118667 445768
rect 117589 445710 118556 445712
rect 117589 445707 117655 445710
rect 118550 445708 118556 445710
rect 118620 445708 118667 445712
rect 118601 445707 118667 445708
rect 90357 444954 90423 444957
rect 141417 444954 141483 444957
rect 90357 444952 141483 444954
rect 90357 444896 90362 444952
rect 90418 444896 141422 444952
rect 141478 444896 141483 444952
rect 90357 444894 141483 444896
rect 90357 444891 90423 444894
rect 141417 444891 141483 444894
rect 115790 444756 115796 444820
rect 115860 444818 115866 444820
rect 124254 444818 124260 444820
rect 115860 444758 124260 444818
rect 115860 444756 115866 444758
rect 124254 444756 124260 444758
rect 124324 444756 124330 444820
rect 52269 444682 52335 444685
rect 93025 444682 93091 444685
rect 94497 444684 94563 444685
rect 94446 444682 94452 444684
rect 52269 444680 93091 444682
rect 52269 444624 52274 444680
rect 52330 444624 93030 444680
rect 93086 444624 93091 444680
rect 52269 444622 93091 444624
rect 94406 444622 94452 444682
rect 94516 444680 94563 444684
rect 120073 444682 120139 444685
rect 94558 444624 94563 444680
rect 52269 444619 52335 444622
rect 93025 444619 93091 444622
rect 94446 444620 94452 444622
rect 94516 444620 94563 444624
rect 94497 444619 94563 444620
rect 103470 444680 120139 444682
rect 103470 444624 120078 444680
rect 120134 444624 120139 444680
rect 583520 444668 584960 444908
rect 103470 444622 120139 444624
rect 87045 444546 87111 444549
rect 103470 444546 103530 444622
rect 120073 444619 120139 444622
rect 87045 444544 103530 444546
rect 87045 444488 87050 444544
rect 87106 444488 103530 444544
rect 87045 444486 103530 444488
rect 87045 444483 87111 444486
rect 108798 444484 108804 444548
rect 108868 444546 108874 444548
rect 109493 444546 109559 444549
rect 108868 444544 109559 444546
rect 108868 444488 109498 444544
rect 109554 444488 109559 444544
rect 108868 444486 109559 444488
rect 108868 444484 108874 444486
rect 109493 444483 109559 444486
rect 111517 444548 111583 444549
rect 114369 444548 114435 444549
rect 111517 444544 111564 444548
rect 111628 444546 111634 444548
rect 114318 444546 114324 444548
rect 111517 444488 111522 444544
rect 111517 444484 111564 444488
rect 111628 444486 111674 444546
rect 114278 444486 114324 444546
rect 114388 444544 114435 444548
rect 114430 444488 114435 444544
rect 111628 444484 111634 444486
rect 114318 444484 114324 444486
rect 114388 444484 114435 444488
rect 111517 444483 111583 444484
rect 114369 444483 114435 444484
rect 124121 444274 124187 444277
rect 120612 444272 124187 444274
rect 120612 444216 124126 444272
rect 124182 444216 124187 444272
rect 120612 444214 124187 444216
rect 124121 444211 124187 444214
rect 197353 443866 197419 443869
rect 197353 443864 200100 443866
rect 197353 443808 197358 443864
rect 197414 443808 200100 443864
rect 197353 443806 200100 443808
rect 197353 443803 197419 443806
rect 358721 443730 358787 443733
rect 356132 443728 358787 443730
rect 356132 443672 358726 443728
rect 358782 443672 358787 443728
rect 356132 443670 358787 443672
rect 358721 443667 358787 443670
rect 67357 442234 67423 442237
rect 67766 442234 67772 442236
rect 67357 442232 67772 442234
rect 67357 442176 67362 442232
rect 67418 442176 67772 442232
rect 67357 442174 67772 442176
rect 67357 442171 67423 442174
rect 67766 442172 67772 442174
rect 67836 442234 67842 442236
rect 67836 442174 68908 442234
rect 67836 442172 67842 442174
rect 124121 442098 124187 442101
rect 120612 442096 124187 442098
rect 120612 442040 124126 442096
rect 124182 442040 124187 442096
rect 120612 442038 124187 442040
rect 124121 442035 124187 442038
rect 197721 441418 197787 441421
rect 197721 441416 200100 441418
rect 197721 441360 197726 441416
rect 197782 441360 200100 441416
rect 197721 441358 200100 441360
rect 197721 441355 197787 441358
rect 358721 441282 358787 441285
rect 356132 441280 358787 441282
rect 356132 441224 358726 441280
rect 358782 441224 358787 441280
rect 356132 441222 358787 441224
rect 358721 441219 358787 441222
rect 121637 440058 121703 440061
rect 120612 440056 121703 440058
rect 120612 440000 121642 440056
rect 121698 440000 121703 440056
rect 120612 439998 121703 440000
rect 121637 439995 121703 439998
rect 66345 439922 66411 439925
rect 66345 439920 68908 439922
rect 66345 439864 66350 439920
rect 66406 439864 68908 439920
rect 66345 439862 68908 439864
rect 66345 439859 66411 439862
rect 197353 438970 197419 438973
rect 357525 438970 357591 438973
rect 358721 438970 358787 438973
rect 197353 438968 200100 438970
rect 197353 438912 197358 438968
rect 197414 438912 200100 438968
rect 197353 438910 200100 438912
rect 356132 438968 358787 438970
rect 356132 438912 357530 438968
rect 357586 438912 358726 438968
rect 358782 438912 358787 438968
rect 356132 438910 358787 438912
rect 197353 438907 197419 438910
rect 357525 438907 357591 438910
rect 358721 438907 358787 438910
rect 124121 437882 124187 437885
rect 120612 437880 124187 437882
rect 120612 437824 124126 437880
rect 124182 437824 124187 437880
rect 120612 437822 124187 437824
rect 124121 437819 124187 437822
rect 66805 437746 66871 437749
rect 66805 437744 68908 437746
rect 66805 437688 66810 437744
rect 66866 437688 68908 437744
rect 66805 437686 68908 437688
rect 66805 437683 66871 437686
rect -960 436508 480 436748
rect 197353 436386 197419 436389
rect 357893 436386 357959 436389
rect 197353 436384 200100 436386
rect 197353 436328 197358 436384
rect 197414 436328 200100 436384
rect 197353 436326 200100 436328
rect 356132 436384 357959 436386
rect 356132 436328 357898 436384
rect 357954 436328 357959 436384
rect 356132 436326 357959 436328
rect 197353 436323 197419 436326
rect 357893 436323 357959 436326
rect 66253 435434 66319 435437
rect 66253 435432 68908 435434
rect 66253 435376 66258 435432
rect 66314 435376 68908 435432
rect 66253 435374 68908 435376
rect 66253 435371 66319 435374
rect 121678 435298 121684 435300
rect 120612 435238 121684 435298
rect 121678 435236 121684 435238
rect 121748 435298 121754 435300
rect 123017 435298 123083 435301
rect 121748 435296 123083 435298
rect 121748 435240 123022 435296
rect 123078 435240 123083 435296
rect 121748 435238 123083 435240
rect 121748 435236 121754 435238
rect 123017 435235 123083 435238
rect 198825 433938 198891 433941
rect 358721 433938 358787 433941
rect 198825 433936 200100 433938
rect 198825 433880 198830 433936
rect 198886 433880 200100 433936
rect 198825 433878 200100 433880
rect 356132 433936 358787 433938
rect 356132 433880 358726 433936
rect 358782 433880 358787 433936
rect 356132 433878 358787 433880
rect 198825 433875 198891 433878
rect 358721 433875 358787 433878
rect 66253 433258 66319 433261
rect 124121 433258 124187 433261
rect 66253 433256 68908 433258
rect 66253 433200 66258 433256
rect 66314 433200 68908 433256
rect 66253 433198 68908 433200
rect 120612 433256 124187 433258
rect 120612 433200 124126 433256
rect 124182 433200 124187 433256
rect 120612 433198 124187 433200
rect 66253 433195 66319 433198
rect 124121 433195 124187 433198
rect 582465 431626 582531 431629
rect 583520 431626 584960 431716
rect 582465 431624 584960 431626
rect 582465 431568 582470 431624
rect 582526 431568 584960 431624
rect 582465 431566 584960 431568
rect 582465 431563 582531 431566
rect 197353 431490 197419 431493
rect 358721 431490 358787 431493
rect 197353 431488 200100 431490
rect 197353 431432 197358 431488
rect 197414 431432 200100 431488
rect 197353 431430 200100 431432
rect 356132 431488 358787 431490
rect 356132 431432 358726 431488
rect 358782 431432 358787 431488
rect 583520 431476 584960 431566
rect 356132 431430 358787 431432
rect 197353 431427 197419 431430
rect 358721 431427 358787 431430
rect 66529 431082 66595 431085
rect 124029 431082 124095 431085
rect 66529 431080 68908 431082
rect 66529 431024 66534 431080
rect 66590 431024 68908 431080
rect 120060 431080 124095 431082
rect 120060 431052 124034 431080
rect 66529 431022 68908 431024
rect 120030 431024 124034 431052
rect 124090 431024 124095 431080
rect 120030 431022 124095 431024
rect 66529 431019 66595 431022
rect 120030 430676 120090 431022
rect 124029 431019 124095 431022
rect 120022 430612 120028 430676
rect 120092 430612 120098 430676
rect 197353 429042 197419 429045
rect 358721 429042 358787 429045
rect 197353 429040 200100 429042
rect 197353 428984 197358 429040
rect 197414 428984 200100 429040
rect 197353 428982 200100 428984
rect 356132 429040 358787 429042
rect 356132 428984 358726 429040
rect 358782 428984 358787 429040
rect 356132 428982 358787 428984
rect 197353 428979 197419 428982
rect 358721 428979 358787 428982
rect 66805 428634 66871 428637
rect 66805 428632 68908 428634
rect 66805 428576 66810 428632
rect 66866 428576 68908 428632
rect 66805 428574 68908 428576
rect 66805 428571 66871 428574
rect 121637 428498 121703 428501
rect 122741 428498 122807 428501
rect 120612 428496 122807 428498
rect 120612 428440 121642 428496
rect 121698 428440 122746 428496
rect 122802 428440 122807 428496
rect 120612 428438 122807 428440
rect 121637 428435 121703 428438
rect 122741 428435 122807 428438
rect 197353 426594 197419 426597
rect 358721 426594 358787 426597
rect 197353 426592 200100 426594
rect 197353 426536 197358 426592
rect 197414 426536 200100 426592
rect 197353 426534 200100 426536
rect 356132 426592 358787 426594
rect 356132 426536 358726 426592
rect 358782 426536 358787 426592
rect 356132 426534 358787 426536
rect 197353 426531 197419 426534
rect 358721 426531 358787 426534
rect 66805 426322 66871 426325
rect 66805 426320 68908 426322
rect 66805 426264 66810 426320
rect 66866 426264 68908 426320
rect 66805 426262 68908 426264
rect 66805 426259 66871 426262
rect 120214 426052 120274 426292
rect 120206 425988 120212 426052
rect 120276 426050 120282 426052
rect 123017 426050 123083 426053
rect 120276 426048 123083 426050
rect 120276 425992 123022 426048
rect 123078 425992 123083 426048
rect 120276 425990 123083 425992
rect 120276 425988 120282 425990
rect 123017 425987 123083 425990
rect 66069 424282 66135 424285
rect 66069 424280 68908 424282
rect 66069 424224 66074 424280
rect 66130 424224 68908 424280
rect 66069 424222 68908 424224
rect 66069 424219 66135 424222
rect 123109 424146 123175 424149
rect 123477 424146 123543 424149
rect 120612 424144 123543 424146
rect 120612 424088 123114 424144
rect 123170 424088 123482 424144
rect 123538 424088 123543 424144
rect 120612 424086 123543 424088
rect 123109 424083 123175 424086
rect 123477 424083 123543 424086
rect 197353 424146 197419 424149
rect 197353 424144 200100 424146
rect 197353 424088 197358 424144
rect 197414 424088 200100 424144
rect 197353 424086 200100 424088
rect 197353 424083 197419 424086
rect 356102 423738 356162 424116
rect 356237 423738 356303 423741
rect 356102 423736 356303 423738
rect -960 423602 480 423692
rect 356102 423680 356242 423736
rect 356298 423680 356303 423736
rect 356102 423678 356303 423680
rect 356237 423675 356303 423678
rect 3141 423602 3207 423605
rect -960 423600 3207 423602
rect -960 423544 3146 423600
rect 3202 423544 3207 423600
rect -960 423542 3207 423544
rect -960 423452 480 423542
rect 3141 423539 3207 423542
rect 66621 421970 66687 421973
rect 122925 421970 122991 421973
rect 66621 421968 68908 421970
rect 66621 421912 66626 421968
rect 66682 421912 68908 421968
rect 66621 421910 68908 421912
rect 120612 421968 122991 421970
rect 120612 421912 122930 421968
rect 122986 421912 122991 421968
rect 120612 421910 122991 421912
rect 66621 421907 66687 421910
rect 122925 421907 122991 421910
rect 198590 421636 198596 421700
rect 198660 421698 198666 421700
rect 358721 421698 358787 421701
rect 198660 421638 200100 421698
rect 356132 421696 358787 421698
rect 356132 421640 358726 421696
rect 358782 421640 358787 421696
rect 356132 421638 358787 421640
rect 198660 421636 198666 421638
rect 358721 421635 358787 421638
rect 124305 420884 124371 420885
rect 124254 420882 124260 420884
rect 124214 420822 124260 420882
rect 124324 420880 124371 420884
rect 124366 420824 124371 420880
rect 124254 420820 124260 420822
rect 124324 420820 124371 420824
rect 124305 420819 124371 420820
rect 66662 419596 66668 419660
rect 66732 419658 66738 419660
rect 67725 419658 67791 419661
rect 124305 419658 124371 419661
rect 66732 419656 68908 419658
rect 66732 419600 67730 419656
rect 67786 419600 68908 419656
rect 66732 419598 68908 419600
rect 120612 419656 124371 419658
rect 120612 419600 124310 419656
rect 124366 419600 124371 419656
rect 120612 419598 124371 419600
rect 66732 419596 66738 419598
rect 67725 419595 67791 419598
rect 124305 419595 124371 419598
rect 198457 419658 198523 419661
rect 198958 419658 198964 419660
rect 198457 419656 198964 419658
rect 198457 419600 198462 419656
rect 198518 419600 198964 419656
rect 198457 419598 198964 419600
rect 198457 419595 198523 419598
rect 198958 419596 198964 419598
rect 199028 419596 199034 419660
rect 197353 419250 197419 419253
rect 358721 419250 358787 419253
rect 197353 419248 200100 419250
rect 197353 419192 197358 419248
rect 197414 419192 200100 419248
rect 197353 419190 200100 419192
rect 356132 419248 358787 419250
rect 356132 419192 358726 419248
rect 358782 419192 358787 419248
rect 356132 419190 358787 419192
rect 197353 419187 197419 419190
rect 358721 419187 358787 419190
rect 583017 418298 583083 418301
rect 583520 418298 584960 418388
rect 583017 418296 584960 418298
rect 583017 418240 583022 418296
rect 583078 418240 584960 418296
rect 583017 418238 584960 418240
rect 583017 418235 583083 418238
rect 583520 418148 584960 418238
rect 121545 417482 121611 417485
rect 120612 417480 121611 417482
rect 120612 417452 121550 417480
rect 120582 417424 121550 417452
rect 121606 417424 121611 417480
rect 120582 417422 121611 417424
rect 68878 416802 68938 417316
rect 120582 417077 120642 417422
rect 121545 417419 121611 417422
rect 120582 417072 120691 417077
rect 120582 417016 120630 417072
rect 120686 417016 120691 417072
rect 120582 417014 120691 417016
rect 120625 417011 120691 417014
rect 66854 416742 68938 416802
rect 197353 416802 197419 416805
rect 358721 416802 358787 416805
rect 197353 416800 200100 416802
rect 197353 416744 197358 416800
rect 197414 416744 200100 416800
rect 197353 416742 200100 416744
rect 356132 416800 358787 416802
rect 356132 416744 358726 416800
rect 358782 416744 358787 416800
rect 356132 416742 358787 416744
rect 56501 416666 56567 416669
rect 64597 416666 64663 416669
rect 66854 416666 66914 416742
rect 197353 416739 197419 416742
rect 358721 416739 358787 416742
rect 56501 416664 66914 416666
rect 56501 416608 56506 416664
rect 56562 416608 64602 416664
rect 64658 416608 66914 416664
rect 56501 416606 66914 416608
rect 56501 416603 56567 416606
rect 64597 416603 64663 416606
rect 52177 415442 52243 415445
rect 56501 415442 56567 415445
rect 52177 415440 56567 415442
rect 52177 415384 52182 415440
rect 52238 415384 56506 415440
rect 56562 415384 56567 415440
rect 52177 415382 56567 415384
rect 52177 415379 52243 415382
rect 56501 415379 56567 415382
rect 66805 415170 66871 415173
rect 122925 415170 122991 415173
rect 66805 415168 68908 415170
rect 66805 415112 66810 415168
rect 66866 415112 68908 415168
rect 66805 415110 68908 415112
rect 120612 415168 122991 415170
rect 120612 415112 122930 415168
rect 122986 415112 122991 415168
rect 120612 415110 122991 415112
rect 66805 415107 66871 415110
rect 122925 415107 122991 415110
rect 197353 414354 197419 414357
rect 358721 414354 358787 414357
rect 197353 414352 200100 414354
rect 197353 414296 197358 414352
rect 197414 414296 200100 414352
rect 197353 414294 200100 414296
rect 356132 414352 358787 414354
rect 356132 414296 358726 414352
rect 358782 414296 358787 414352
rect 356132 414294 358787 414296
rect 197353 414291 197419 414294
rect 358721 414291 358787 414294
rect 67449 412858 67515 412861
rect 67449 412856 68908 412858
rect 67449 412800 67454 412856
rect 67510 412800 68908 412856
rect 67449 412798 68908 412800
rect 67449 412795 67515 412798
rect 124121 412722 124187 412725
rect 120612 412720 124187 412722
rect 120612 412664 124126 412720
rect 124182 412664 124187 412720
rect 120612 412662 124187 412664
rect 124121 412659 124187 412662
rect 197353 411906 197419 411909
rect 358721 411906 358787 411909
rect 197353 411904 200100 411906
rect 197353 411848 197358 411904
rect 197414 411848 200100 411904
rect 197353 411846 200100 411848
rect 356132 411904 358787 411906
rect 356132 411848 358726 411904
rect 358782 411848 358787 411904
rect 356132 411846 358787 411848
rect 197353 411843 197419 411846
rect 358721 411843 358787 411846
rect 123569 411362 123635 411365
rect 154614 411362 154620 411364
rect 122790 411360 154620 411362
rect 122790 411304 123574 411360
rect 123630 411304 154620 411360
rect 122790 411302 154620 411304
rect 122790 411226 122850 411302
rect 123569 411299 123635 411302
rect 154614 411300 154620 411302
rect 154684 411300 154690 411364
rect 120582 411166 122850 411226
rect 66713 410682 66779 410685
rect 66713 410680 68908 410682
rect -960 410546 480 410636
rect 66713 410624 66718 410680
rect 66774 410624 68908 410680
rect 120582 410652 120642 411166
rect 66713 410622 68908 410624
rect 66713 410619 66779 410622
rect 3417 410546 3483 410549
rect -960 410544 3483 410546
rect -960 410488 3422 410544
rect 3478 410488 3483 410544
rect -960 410486 3483 410488
rect -960 410396 480 410486
rect 3417 410483 3483 410486
rect 197353 409594 197419 409597
rect 197353 409592 200100 409594
rect 197353 409536 197358 409592
rect 197414 409536 200100 409592
rect 197353 409534 200100 409536
rect 197353 409531 197419 409534
rect 358721 409458 358787 409461
rect 356132 409456 358787 409458
rect 356132 409400 358726 409456
rect 358782 409400 358787 409456
rect 356132 409398 358787 409400
rect 358721 409395 358787 409398
rect 124121 408370 124187 408373
rect 120612 408368 124187 408370
rect 69246 407828 69306 408340
rect 120612 408312 124126 408368
rect 124182 408312 124187 408368
rect 120612 408310 124187 408312
rect 124121 408307 124187 408310
rect 69238 407764 69244 407828
rect 69308 407764 69314 407828
rect 60549 407146 60615 407149
rect 69238 407146 69244 407148
rect 60549 407144 69244 407146
rect 60549 407088 60554 407144
rect 60610 407088 69244 407144
rect 60549 407086 69244 407088
rect 60549 407083 60615 407086
rect 69238 407084 69244 407086
rect 69308 407084 69314 407148
rect 197353 407010 197419 407013
rect 358721 407010 358787 407013
rect 197353 407008 200100 407010
rect 197353 406952 197358 407008
rect 197414 406952 200100 407008
rect 197353 406950 200100 406952
rect 356132 407008 358787 407010
rect 356132 406952 358726 407008
rect 358782 406952 358787 407008
rect 356132 406950 358787 406952
rect 197353 406947 197419 406950
rect 358721 406947 358787 406950
rect 66345 406194 66411 406197
rect 124121 406194 124187 406197
rect 66345 406192 68908 406194
rect 66345 406136 66350 406192
rect 66406 406136 68908 406192
rect 66345 406134 68908 406136
rect 120612 406192 124187 406194
rect 120612 406136 124126 406192
rect 124182 406136 124187 406192
rect 120612 406134 124187 406136
rect 66345 406131 66411 406134
rect 124121 406131 124187 406134
rect 582649 404970 582715 404973
rect 582925 404970 582991 404973
rect 583520 404970 584960 405060
rect 582649 404968 584960 404970
rect 582649 404912 582654 404968
rect 582710 404912 582930 404968
rect 582986 404912 584960 404968
rect 582649 404910 584960 404912
rect 582649 404907 582715 404910
rect 582925 404907 582991 404910
rect 583520 404820 584960 404910
rect 186814 404500 186820 404564
rect 186884 404562 186890 404564
rect 186884 404502 200100 404562
rect 186884 404500 186890 404502
rect 358721 404290 358787 404293
rect 356132 404288 358787 404290
rect 356132 404232 358726 404288
rect 358782 404232 358787 404288
rect 356132 404230 358787 404232
rect 358721 404227 358787 404230
rect 66345 403746 66411 403749
rect 122598 403746 122604 403748
rect 66345 403744 68908 403746
rect 66345 403688 66350 403744
rect 66406 403688 68908 403744
rect 66345 403686 68908 403688
rect 120612 403686 122604 403746
rect 66345 403683 66411 403686
rect 122598 403684 122604 403686
rect 122668 403746 122674 403748
rect 123845 403746 123911 403749
rect 122668 403744 123911 403746
rect 122668 403688 123850 403744
rect 123906 403688 123911 403744
rect 122668 403686 123911 403688
rect 122668 403684 122674 403686
rect 123845 403683 123911 403686
rect 177430 401644 177436 401708
rect 177500 401706 177506 401708
rect 200070 401706 200130 402084
rect 358721 401842 358787 401845
rect 356132 401840 358787 401842
rect 356132 401784 358726 401840
rect 358782 401784 358787 401840
rect 356132 401782 358787 401784
rect 358721 401779 358787 401782
rect 177500 401646 200130 401706
rect 177500 401644 177506 401646
rect 66345 401570 66411 401573
rect 123937 401570 124003 401573
rect 66345 401568 68908 401570
rect 66345 401512 66350 401568
rect 66406 401512 68908 401568
rect 66345 401510 68908 401512
rect 120612 401568 124003 401570
rect 120612 401512 123942 401568
rect 123998 401512 124003 401568
rect 120612 401510 124003 401512
rect 66345 401507 66411 401510
rect 123937 401507 124003 401510
rect 197353 399666 197419 399669
rect 197353 399664 200100 399666
rect 197353 399608 197358 399664
rect 197414 399608 200100 399664
rect 197353 399606 200100 399608
rect 197353 399603 197419 399606
rect 66345 399394 66411 399397
rect 124121 399394 124187 399397
rect 358629 399394 358695 399397
rect 66345 399392 68908 399394
rect 66345 399336 66350 399392
rect 66406 399336 68908 399392
rect 66345 399334 68908 399336
rect 120612 399392 124187 399394
rect 120612 399336 124126 399392
rect 124182 399336 124187 399392
rect 120612 399334 124187 399336
rect 356132 399392 358695 399394
rect 356132 399336 358634 399392
rect 358690 399336 358695 399392
rect 356132 399334 358695 399336
rect 66345 399331 66411 399334
rect 124121 399331 124187 399334
rect 358629 399331 358695 399334
rect -960 397490 480 397580
rect 2773 397490 2839 397493
rect -960 397488 2839 397490
rect -960 397432 2778 397488
rect 2834 397432 2839 397488
rect -960 397430 2839 397432
rect -960 397340 480 397430
rect 2773 397427 2839 397430
rect 122097 397354 122163 397357
rect 123753 397354 123819 397357
rect 120582 397352 123819 397354
rect 120582 397296 122102 397352
rect 122158 397296 123758 397352
rect 123814 397296 123819 397352
rect 120582 397294 123819 397296
rect 120582 397052 120642 397294
rect 122097 397291 122163 397294
rect 123753 397291 123819 397294
rect 197353 397218 197419 397221
rect 197353 397216 200100 397218
rect 197353 397160 197358 397216
rect 197414 397160 200100 397216
rect 197353 397158 200100 397160
rect 197353 397155 197419 397158
rect 66989 396946 67055 396949
rect 67357 396946 67423 396949
rect 359089 396946 359155 396949
rect 66989 396944 68908 396946
rect 66989 396888 66994 396944
rect 67050 396888 67362 396944
rect 67418 396888 68908 396944
rect 66989 396886 68908 396888
rect 356132 396944 359155 396946
rect 356132 396888 359094 396944
rect 359150 396888 359155 396944
rect 356132 396886 359155 396888
rect 66989 396883 67055 396886
rect 67357 396883 67423 396886
rect 359089 396883 359155 396886
rect 67265 395994 67331 395997
rect 67541 395994 67607 395997
rect 67265 395992 67607 395994
rect 67265 395936 67270 395992
rect 67326 395936 67546 395992
rect 67602 395936 67607 395992
rect 67265 395934 67607 395936
rect 67265 395931 67331 395934
rect 67541 395931 67607 395934
rect 67541 394906 67607 394909
rect 121545 394906 121611 394909
rect 67541 394904 68908 394906
rect 67541 394848 67546 394904
rect 67602 394848 68908 394904
rect 67541 394846 68908 394848
rect 120612 394904 121611 394906
rect 120612 394848 121550 394904
rect 121606 394848 121611 394904
rect 120612 394846 121611 394848
rect 67541 394843 67607 394846
rect 121545 394843 121611 394846
rect 197353 394770 197419 394773
rect 197353 394768 200100 394770
rect 197353 394712 197358 394768
rect 197414 394712 200100 394768
rect 197353 394710 200100 394712
rect 197353 394707 197419 394710
rect 358721 394498 358787 394501
rect 356132 394496 358787 394498
rect 356132 394440 358726 394496
rect 358782 394440 358787 394496
rect 356132 394438 358787 394440
rect 358721 394435 358787 394438
rect 368657 393410 368723 393413
rect 400254 393410 400260 393412
rect 368657 393408 400260 393410
rect 368657 393352 368662 393408
rect 368718 393352 400260 393408
rect 368657 393350 400260 393352
rect 368657 393347 368723 393350
rect 400254 393348 400260 393350
rect 400324 393348 400330 393412
rect 66805 392594 66871 392597
rect 121453 392594 121519 392597
rect 66805 392592 68908 392594
rect 66805 392536 66810 392592
rect 66866 392536 68908 392592
rect 66805 392534 68908 392536
rect 120612 392592 121519 392594
rect 120612 392536 121458 392592
rect 121514 392536 121519 392592
rect 120612 392534 121519 392536
rect 66805 392531 66871 392534
rect 121453 392531 121519 392534
rect 198457 392322 198523 392325
rect 180750 392320 200100 392322
rect 180750 392264 198462 392320
rect 198518 392264 200100 392320
rect 180750 392262 200100 392264
rect 119470 392124 119476 392188
rect 119540 392186 119546 392188
rect 180750 392186 180810 392262
rect 198457 392259 198523 392262
rect 119540 392126 180810 392186
rect 119540 392124 119546 392126
rect 357617 392050 357683 392053
rect 356132 392048 357683 392050
rect 356132 391992 357622 392048
rect 357678 391992 357683 392048
rect 356132 391990 357683 391992
rect 357617 391987 357683 391990
rect 583520 391628 584960 391868
rect 64689 391370 64755 391373
rect 137277 391370 137343 391373
rect 64689 391368 70410 391370
rect 64689 391312 64694 391368
rect 64750 391312 70410 391368
rect 64689 391310 70410 391312
rect 64689 391307 64755 391310
rect 70350 391098 70410 391310
rect 89670 391368 137343 391370
rect 89670 391312 137282 391368
rect 137338 391312 137343 391368
rect 89670 391310 137343 391312
rect 71814 391172 71820 391236
rect 71884 391234 71890 391236
rect 71884 391174 84946 391234
rect 71884 391172 71890 391174
rect 70350 391038 80070 391098
rect 80010 390826 80070 391038
rect 84886 390962 84946 391174
rect 85665 391098 85731 391101
rect 89670 391098 89730 391310
rect 137277 391307 137343 391310
rect 177389 391234 177455 391237
rect 93810 391232 177455 391234
rect 93810 391176 177394 391232
rect 177450 391176 177455 391232
rect 93810 391174 177455 391176
rect 85665 391096 89730 391098
rect 85665 391040 85670 391096
rect 85726 391040 89730 391096
rect 85665 391038 89730 391040
rect 85665 391035 85731 391038
rect 92606 391036 92612 391100
rect 92676 391098 92682 391100
rect 92749 391098 92815 391101
rect 92676 391096 92815 391098
rect 92676 391040 92754 391096
rect 92810 391040 92815 391096
rect 92676 391038 92815 391040
rect 92676 391036 92682 391038
rect 92749 391035 92815 391038
rect 93810 390962 93870 391174
rect 177389 391171 177455 391174
rect 84886 390902 93870 390962
rect 85665 390826 85731 390829
rect 80010 390824 85731 390826
rect 80010 390768 85670 390824
rect 85726 390768 85731 390824
rect 80010 390766 85731 390768
rect 85665 390763 85731 390766
rect 71865 390692 71931 390693
rect 71814 390628 71820 390692
rect 71884 390690 71931 390692
rect 71884 390688 71976 390690
rect 71926 390632 71976 390688
rect 71884 390630 71976 390632
rect 71884 390628 71931 390630
rect 71865 390627 71931 390628
rect 102133 390556 102199 390557
rect 102133 390554 102180 390556
rect 102088 390552 102180 390554
rect 102088 390496 102138 390552
rect 102088 390494 102180 390496
rect 102133 390492 102180 390494
rect 102244 390492 102250 390556
rect 102133 390491 102199 390492
rect 69606 390356 69612 390420
rect 69676 390418 69682 390420
rect 69933 390418 69999 390421
rect 69676 390416 69999 390418
rect 69676 390360 69938 390416
rect 69994 390360 69999 390416
rect 69676 390358 69999 390360
rect 69676 390356 69682 390358
rect 69933 390355 69999 390358
rect 89478 390356 89484 390420
rect 89548 390418 89554 390420
rect 89805 390418 89871 390421
rect 89548 390416 89871 390418
rect 89548 390360 89810 390416
rect 89866 390360 89871 390416
rect 89548 390358 89871 390360
rect 89548 390356 89554 390358
rect 89805 390355 89871 390358
rect 91134 390356 91140 390420
rect 91204 390418 91210 390420
rect 91277 390418 91343 390421
rect 91204 390416 91343 390418
rect 91204 390360 91282 390416
rect 91338 390360 91343 390416
rect 91204 390358 91343 390360
rect 91204 390356 91210 390358
rect 91277 390355 91343 390358
rect 93894 390356 93900 390420
rect 93964 390418 93970 390420
rect 94221 390418 94287 390421
rect 93964 390416 94287 390418
rect 93964 390360 94226 390416
rect 94282 390360 94287 390416
rect 93964 390358 94287 390360
rect 93964 390356 93970 390358
rect 94221 390355 94287 390358
rect 96654 390356 96660 390420
rect 96724 390418 96730 390420
rect 97349 390418 97415 390421
rect 96724 390416 97415 390418
rect 96724 390360 97354 390416
rect 97410 390360 97415 390416
rect 96724 390358 97415 390360
rect 96724 390356 96730 390358
rect 97349 390355 97415 390358
rect 98126 390356 98132 390420
rect 98196 390418 98202 390420
rect 98821 390418 98887 390421
rect 104985 390420 105051 390421
rect 104934 390418 104940 390420
rect 98196 390416 98887 390418
rect 98196 390360 98826 390416
rect 98882 390360 98887 390416
rect 98196 390358 98887 390360
rect 104894 390358 104940 390418
rect 105004 390416 105051 390420
rect 105046 390360 105051 390416
rect 98196 390356 98202 390358
rect 98821 390355 98887 390358
rect 104934 390356 104940 390358
rect 105004 390356 105051 390360
rect 106406 390356 106412 390420
rect 106476 390418 106482 390420
rect 106549 390418 106615 390421
rect 106476 390416 106615 390418
rect 106476 390360 106554 390416
rect 106610 390360 106615 390416
rect 106476 390358 106615 390360
rect 106476 390356 106482 390358
rect 104985 390355 105051 390356
rect 106549 390355 106615 390358
rect 107694 390356 107700 390420
rect 107764 390418 107770 390420
rect 108021 390418 108087 390421
rect 107764 390416 108087 390418
rect 107764 390360 108026 390416
rect 108082 390360 108087 390416
rect 107764 390358 108087 390360
rect 107764 390356 107770 390358
rect 108021 390355 108087 390358
rect 108982 390356 108988 390420
rect 109052 390418 109058 390420
rect 109493 390418 109559 390421
rect 109052 390416 109559 390418
rect 109052 390360 109498 390416
rect 109554 390360 109559 390416
rect 109052 390358 109559 390360
rect 109052 390356 109058 390358
rect 109493 390355 109559 390358
rect 115933 390420 115999 390421
rect 118785 390420 118851 390421
rect 115933 390416 115980 390420
rect 116044 390418 116050 390420
rect 118734 390418 118740 390420
rect 115933 390360 115938 390416
rect 115933 390356 115980 390360
rect 116044 390358 116090 390418
rect 118694 390358 118740 390418
rect 118804 390416 118851 390420
rect 118846 390360 118851 390416
rect 116044 390356 116050 390358
rect 118734 390356 118740 390358
rect 118804 390356 118851 390360
rect 115933 390355 115999 390356
rect 118785 390355 118851 390356
rect 100753 390284 100819 390285
rect 100702 390282 100708 390284
rect 100662 390222 100708 390282
rect 100772 390280 100819 390284
rect 100814 390224 100819 390280
rect 100702 390220 100708 390222
rect 100772 390220 100819 390224
rect 100753 390219 100819 390220
rect 108389 389466 108455 389469
rect 159449 389466 159515 389469
rect 108389 389464 159515 389466
rect 108389 389408 108394 389464
rect 108450 389408 159454 389464
rect 159510 389408 159515 389464
rect 108389 389406 159515 389408
rect 108389 389403 108455 389406
rect 159449 389403 159515 389406
rect 102225 389330 102291 389333
rect 155309 389330 155375 389333
rect 102225 389328 155375 389330
rect 102225 389272 102230 389328
rect 102286 389272 155314 389328
rect 155370 389272 155375 389328
rect 102225 389270 155375 389272
rect 102225 389267 102291 389270
rect 155309 389267 155375 389270
rect 64597 389194 64663 389197
rect 200070 389194 200130 389844
rect 357709 389602 357775 389605
rect 356132 389600 357775 389602
rect 356132 389544 357714 389600
rect 357770 389544 357775 389600
rect 356132 389542 357775 389544
rect 357709 389539 357775 389542
rect 64597 389192 200130 389194
rect 64597 389136 64602 389192
rect 64658 389136 200130 389192
rect 64597 389134 200130 389136
rect 64597 389131 64663 389134
rect 73337 389058 73403 389061
rect 90357 389058 90423 389061
rect 73337 389056 90423 389058
rect 73337 389000 73342 389056
rect 73398 389000 90362 389056
rect 90418 389000 90423 389056
rect 73337 388998 90423 389000
rect 73337 388995 73403 388998
rect 90357 388995 90423 388998
rect 95182 388996 95188 389060
rect 95252 389058 95258 389060
rect 96153 389058 96219 389061
rect 95252 389056 96219 389058
rect 95252 389000 96158 389056
rect 96214 389000 96219 389056
rect 95252 388998 96219 389000
rect 95252 388996 95258 388998
rect 96153 388995 96219 388998
rect 111742 388996 111748 389060
rect 111812 389058 111818 389060
rect 112897 389058 112963 389061
rect 111812 389056 112963 389058
rect 111812 389000 112902 389056
rect 112958 389000 112963 389056
rect 111812 388998 112963 389000
rect 111812 388996 111818 388998
rect 112897 388995 112963 388998
rect 116117 389058 116183 389061
rect 117129 389058 117195 389061
rect 116117 389056 117195 389058
rect 116117 389000 116122 389056
rect 116178 389000 117134 389056
rect 117190 389000 117195 389056
rect 116117 388998 117195 389000
rect 116117 388995 116183 388998
rect 117129 388995 117195 388998
rect 117589 389058 117655 389061
rect 117998 389058 118004 389060
rect 117589 389056 118004 389058
rect 117589 389000 117594 389056
rect 117650 389000 118004 389056
rect 117589 388998 118004 389000
rect 117589 388995 117655 388998
rect 117998 388996 118004 388998
rect 118068 389058 118074 389060
rect 118601 389058 118667 389061
rect 118068 389056 118667 389058
rect 118068 389000 118606 389056
rect 118662 389000 118667 389056
rect 118068 388998 118667 389000
rect 118068 388996 118074 388998
rect 118601 388995 118667 388998
rect 61837 388786 61903 388789
rect 79501 388786 79567 388789
rect 61837 388784 79567 388786
rect 61837 388728 61842 388784
rect 61898 388728 79506 388784
rect 79562 388728 79567 388784
rect 61837 388726 79567 388728
rect 61837 388723 61903 388726
rect 79501 388723 79567 388726
rect 92473 388650 92539 388653
rect 93761 388650 93827 388653
rect 97942 388650 97948 388652
rect 92473 388648 97948 388650
rect 92473 388592 92478 388648
rect 92534 388592 93766 388648
rect 93822 388592 97948 388648
rect 92473 388590 97948 388592
rect 92473 388587 92539 388590
rect 93761 388587 93827 388590
rect 97942 388588 97948 388590
rect 98012 388588 98018 388652
rect 95233 388514 95299 388517
rect 96470 388514 96476 388516
rect 95233 388512 96476 388514
rect 95233 388456 95238 388512
rect 95294 388456 96476 388512
rect 95233 388454 96476 388456
rect 95233 388451 95299 388454
rect 96470 388452 96476 388454
rect 96540 388452 96546 388516
rect 107469 388514 107535 388517
rect 120441 388514 120507 388517
rect 107469 388512 120507 388514
rect 107469 388456 107474 388512
rect 107530 388456 120446 388512
rect 120502 388456 120507 388512
rect 107469 388454 120507 388456
rect 107469 388451 107535 388454
rect 120441 388451 120507 388454
rect 61837 388378 61903 388381
rect 72366 388378 72372 388380
rect 61837 388376 72372 388378
rect 61837 388320 61842 388376
rect 61898 388320 72372 388376
rect 61837 388318 72372 388320
rect 61837 388315 61903 388318
rect 72366 388316 72372 388318
rect 72436 388378 72442 388380
rect 74533 388378 74599 388381
rect 72436 388376 74599 388378
rect 72436 388320 74538 388376
rect 74594 388320 74599 388376
rect 72436 388318 74599 388320
rect 72436 388316 72442 388318
rect 74533 388315 74599 388318
rect 77845 388378 77911 388381
rect 167177 388378 167243 388381
rect 77845 388376 167243 388378
rect 77845 388320 77850 388376
rect 77906 388320 167182 388376
rect 167238 388320 167243 388376
rect 77845 388318 167243 388320
rect 77845 388315 77911 388318
rect 167177 388315 167243 388318
rect 197353 387426 197419 387429
rect 197353 387424 200100 387426
rect 197353 387368 197358 387424
rect 197414 387368 200100 387424
rect 197353 387366 200100 387368
rect 197353 387363 197419 387366
rect 358721 387154 358787 387157
rect 356132 387152 358787 387154
rect 356132 387096 358726 387152
rect 358782 387096 358787 387152
rect 356132 387094 358787 387096
rect 358721 387091 358787 387094
rect 7557 387018 7623 387021
rect 118969 387018 119035 387021
rect 7557 387016 119035 387018
rect 7557 386960 7562 387016
rect 7618 386960 118974 387016
rect 119030 386960 119035 387016
rect 7557 386958 119035 386960
rect 7557 386955 7623 386958
rect 118969 386955 119035 386958
rect 91001 386474 91067 386477
rect 156597 386474 156663 386477
rect 91001 386472 156663 386474
rect 91001 386416 91006 386472
rect 91062 386416 156602 386472
rect 156658 386416 156663 386472
rect 91001 386414 156663 386416
rect 91001 386411 91067 386414
rect 156597 386411 156663 386414
rect 4797 385658 4863 385661
rect 95182 385658 95188 385660
rect 4797 385656 95188 385658
rect 4797 385600 4802 385656
rect 4858 385600 95188 385656
rect 4797 385598 95188 385600
rect 4797 385595 4863 385598
rect 95182 385596 95188 385598
rect 95252 385596 95258 385660
rect 99281 385658 99347 385661
rect 158069 385658 158135 385661
rect 99281 385656 158135 385658
rect 99281 385600 99286 385656
rect 99342 385600 158074 385656
rect 158130 385600 158135 385656
rect 99281 385598 158135 385600
rect 99281 385595 99347 385598
rect 158069 385595 158135 385598
rect 83917 384980 83983 384981
rect 83917 384978 83964 384980
rect 83836 384976 83964 384978
rect 84028 384978 84034 384980
rect 124213 384978 124279 384981
rect 84028 384976 124279 384978
rect 83836 384920 83922 384976
rect 84028 384920 124218 384976
rect 124274 384920 124279 384976
rect 83836 384918 83964 384920
rect 83917 384916 83964 384918
rect 84028 384918 124279 384920
rect 84028 384916 84034 384918
rect 83917 384915 83983 384916
rect 124213 384915 124279 384918
rect 197302 384916 197308 384980
rect 197372 384978 197378 384980
rect 197372 384918 200100 384978
rect 197372 384916 197378 384918
rect 358721 384706 358787 384709
rect 356132 384704 358787 384706
rect 356132 384648 358726 384704
rect 358782 384648 358787 384704
rect 356132 384646 358787 384648
rect 358721 384643 358787 384646
rect -960 384284 480 384524
rect 61929 384298 61995 384301
rect 174997 384298 175063 384301
rect 61929 384296 175063 384298
rect 61929 384240 61934 384296
rect 61990 384240 175002 384296
rect 175058 384240 175063 384296
rect 61929 384238 175063 384240
rect 61929 384235 61995 384238
rect 174997 384235 175063 384238
rect 174997 383754 175063 383757
rect 197302 383754 197308 383756
rect 174997 383752 197308 383754
rect 174997 383696 175002 383752
rect 175058 383696 197308 383752
rect 174997 383694 197308 383696
rect 174997 383691 175063 383694
rect 197302 383692 197308 383694
rect 197372 383692 197378 383756
rect 57697 382938 57763 382941
rect 121545 382938 121611 382941
rect 57697 382936 121611 382938
rect 57697 382880 57702 382936
rect 57758 382880 121550 382936
rect 121606 382880 121611 382936
rect 57697 382878 121611 382880
rect 57697 382875 57763 382878
rect 121545 382875 121611 382878
rect 124397 382530 124463 382533
rect 185577 382530 185643 382533
rect 124397 382528 185643 382530
rect 124397 382472 124402 382528
rect 124458 382472 185582 382528
rect 185638 382472 185643 382528
rect 124397 382470 185643 382472
rect 124397 382467 124463 382470
rect 185577 382467 185643 382470
rect 197169 382530 197235 382533
rect 197169 382528 200100 382530
rect 197169 382472 197174 382528
rect 197230 382472 200100 382528
rect 197169 382470 200100 382472
rect 197169 382467 197235 382470
rect 60549 382394 60615 382397
rect 189809 382394 189875 382397
rect 356329 382394 356395 382397
rect 60549 382392 189875 382394
rect 60549 382336 60554 382392
rect 60610 382336 189814 382392
rect 189870 382336 189875 382392
rect 60549 382334 189875 382336
rect 356132 382392 356395 382394
rect 356132 382336 356334 382392
rect 356390 382336 356395 382392
rect 356132 382334 356395 382336
rect 60549 382331 60615 382334
rect 189809 382331 189875 382334
rect 356329 382331 356395 382334
rect 65517 381034 65583 381037
rect 66069 381034 66135 381037
rect 189165 381034 189231 381037
rect 65517 381032 189231 381034
rect 65517 380976 65522 381032
rect 65578 380976 66074 381032
rect 66130 380976 189170 381032
rect 189226 380976 189231 381032
rect 65517 380974 189231 380976
rect 65517 380971 65583 380974
rect 66069 380971 66135 380974
rect 189165 380971 189231 380974
rect 142981 380218 143047 380221
rect 158662 380218 158668 380220
rect 142981 380216 158668 380218
rect 142981 380160 142986 380216
rect 143042 380160 158668 380216
rect 142981 380158 158668 380160
rect 142981 380155 143047 380158
rect 158662 380156 158668 380158
rect 158732 380156 158738 380220
rect 197353 380082 197419 380085
rect 197353 380080 200100 380082
rect 197353 380024 197358 380080
rect 197414 380024 200100 380080
rect 197353 380022 200100 380024
rect 197353 380019 197419 380022
rect 358629 379810 358695 379813
rect 356132 379808 358695 379810
rect 356132 379752 358634 379808
rect 358690 379752 358695 379808
rect 356132 379750 358695 379752
rect 358629 379747 358695 379750
rect 95141 379538 95207 379541
rect 195329 379538 195395 379541
rect 95141 379536 195395 379538
rect 95141 379480 95146 379536
rect 95202 379480 195334 379536
rect 195390 379480 195395 379536
rect 95141 379478 195395 379480
rect 95141 379475 95207 379478
rect 195329 379475 195395 379478
rect 67725 378858 67791 378861
rect 124806 378858 124812 378860
rect 67725 378856 124812 378858
rect 67725 378800 67730 378856
rect 67786 378800 124812 378856
rect 67725 378798 124812 378800
rect 67725 378795 67791 378798
rect 124806 378796 124812 378798
rect 124876 378796 124882 378860
rect 53649 378722 53715 378725
rect 160093 378722 160159 378725
rect 53649 378720 160159 378722
rect 53649 378664 53654 378720
rect 53710 378664 160098 378720
rect 160154 378664 160159 378720
rect 53649 378662 160159 378664
rect 53649 378659 53715 378662
rect 160093 378659 160159 378662
rect 580349 378450 580415 378453
rect 583520 378450 584960 378540
rect 580349 378448 584960 378450
rect 580349 378392 580354 378448
rect 580410 378392 584960 378448
rect 580349 378390 584960 378392
rect 580349 378387 580415 378390
rect 187693 378314 187759 378317
rect 188981 378314 189047 378317
rect 200614 378314 200620 378316
rect 187693 378312 200620 378314
rect 187693 378256 187698 378312
rect 187754 378256 188986 378312
rect 189042 378256 200620 378312
rect 187693 378254 200620 378256
rect 187693 378251 187759 378254
rect 188981 378251 189047 378254
rect 200614 378252 200620 378254
rect 200684 378252 200690 378316
rect 583520 378300 584960 378390
rect 148501 378178 148567 378181
rect 192753 378178 192819 378181
rect 148501 378176 192819 378178
rect 148501 378120 148506 378176
rect 148562 378120 192758 378176
rect 192814 378120 192819 378176
rect 148501 378118 192819 378120
rect 148501 378115 148567 378118
rect 192753 378115 192819 378118
rect 194358 378116 194364 378180
rect 194428 378178 194434 378180
rect 199653 378178 199719 378181
rect 194428 378176 199719 378178
rect 194428 378120 199658 378176
rect 199714 378120 199719 378176
rect 194428 378118 199719 378120
rect 194428 378116 194434 378118
rect 199653 378115 199719 378118
rect 116577 378042 116643 378045
rect 117129 378042 117195 378045
rect 116577 378040 117195 378042
rect 116577 377984 116582 378040
rect 116638 377984 117134 378040
rect 117190 377984 117195 378040
rect 116577 377982 117195 377984
rect 116577 377979 116643 377982
rect 117129 377979 117195 377982
rect 197302 377980 197308 378044
rect 197372 378042 197378 378044
rect 580257 378042 580323 378045
rect 197372 378040 580323 378042
rect 197372 377984 580262 378040
rect 580318 377984 580323 378040
rect 197372 377982 580323 377984
rect 197372 377980 197378 377982
rect 580257 377979 580323 377982
rect 195881 377634 195947 377637
rect 202229 377634 202295 377637
rect 195881 377632 202295 377634
rect 195881 377576 195886 377632
rect 195942 377576 202234 377632
rect 202290 377576 202295 377632
rect 195881 377574 202295 377576
rect 195881 377571 195947 377574
rect 202229 377571 202295 377574
rect 355317 377634 355383 377637
rect 356329 377634 356395 377637
rect 355317 377632 356395 377634
rect 355317 377576 355322 377632
rect 355378 377576 356334 377632
rect 356390 377576 356395 377632
rect 355317 377574 356395 377576
rect 355317 377571 355383 377574
rect 356329 377571 356395 377574
rect 199653 377498 199719 377501
rect 201401 377498 201467 377501
rect 199653 377496 201467 377498
rect 199653 377440 199658 377496
rect 199714 377440 201406 377496
rect 201462 377440 201467 377496
rect 199653 377438 201467 377440
rect 199653 377435 199719 377438
rect 201401 377435 201467 377438
rect 92289 377362 92355 377365
rect 120022 377362 120028 377364
rect 92289 377360 120028 377362
rect 92289 377304 92294 377360
rect 92350 377304 120028 377360
rect 92289 377302 120028 377304
rect 92289 377299 92355 377302
rect 120022 377300 120028 377302
rect 120092 377300 120098 377364
rect 351177 377362 351243 377365
rect 361849 377362 361915 377365
rect 351177 377360 361915 377362
rect 351177 377304 351182 377360
rect 351238 377304 361854 377360
rect 361910 377304 361915 377360
rect 351177 377302 361915 377304
rect 351177 377299 351243 377302
rect 361849 377299 361915 377302
rect 116577 376818 116643 376821
rect 272701 376818 272767 376821
rect 116577 376816 272767 376818
rect 116577 376760 116582 376816
rect 116638 376760 272706 376816
rect 272762 376760 272767 376816
rect 116577 376758 272767 376760
rect 116577 376755 116643 376758
rect 272701 376755 272767 376758
rect 65885 376682 65951 376685
rect 281441 376682 281507 376685
rect 65885 376680 281507 376682
rect 65885 376624 65890 376680
rect 65946 376624 281446 376680
rect 281502 376624 281507 376680
rect 65885 376622 281507 376624
rect 65885 376619 65951 376622
rect 281441 376619 281507 376622
rect 319621 376682 319687 376685
rect 582833 376682 582899 376685
rect 319621 376680 582899 376682
rect 319621 376624 319626 376680
rect 319682 376624 582838 376680
rect 582894 376624 582899 376680
rect 319621 376622 582899 376624
rect 319621 376619 319687 376622
rect 582833 376619 582899 376622
rect 198958 376484 198964 376548
rect 199028 376546 199034 376548
rect 199469 376546 199535 376549
rect 199028 376544 199535 376546
rect 199028 376488 199474 376544
rect 199530 376488 199535 376544
rect 199028 376486 199535 376488
rect 199028 376484 199034 376486
rect 199469 376483 199535 376486
rect 199837 376138 199903 376141
rect 208485 376138 208551 376141
rect 199837 376136 208551 376138
rect 199837 376080 199842 376136
rect 199898 376080 208490 376136
rect 208546 376080 208551 376136
rect 199837 376078 208551 376080
rect 199837 376075 199903 376078
rect 208485 376075 208551 376078
rect 195237 376002 195303 376005
rect 211797 376002 211863 376005
rect 195237 376000 211863 376002
rect 195237 375944 195242 376000
rect 195298 375944 211802 376000
rect 211858 375944 211863 376000
rect 195237 375942 211863 375944
rect 195237 375939 195303 375942
rect 211797 375939 211863 375942
rect 233877 376002 233943 376005
rect 365989 376002 366055 376005
rect 233877 376000 366055 376002
rect 233877 375944 233882 376000
rect 233938 375944 365994 376000
rect 366050 375944 366055 376000
rect 233877 375942 366055 375944
rect 233877 375939 233943 375942
rect 365989 375939 366055 375942
rect 114318 375260 114324 375324
rect 114388 375322 114394 375324
rect 119981 375322 120047 375325
rect 114388 375320 120047 375322
rect 114388 375264 119986 375320
rect 120042 375264 120047 375320
rect 114388 375262 120047 375264
rect 114388 375260 114394 375262
rect 119981 375259 120047 375262
rect 194501 375322 194567 375325
rect 247033 375322 247099 375325
rect 194501 375320 247099 375322
rect 194501 375264 194506 375320
rect 194562 375264 247038 375320
rect 247094 375264 247099 375320
rect 194501 375262 247099 375264
rect 194501 375259 194567 375262
rect 247033 375259 247099 375262
rect 281441 375322 281507 375325
rect 582373 375322 582439 375325
rect 281441 375320 582439 375322
rect 281441 375264 281446 375320
rect 281502 375264 582378 375320
rect 582434 375264 582439 375320
rect 281441 375262 582439 375264
rect 281441 375259 281507 375262
rect 582373 375259 582439 375262
rect 189165 375186 189231 375189
rect 233877 375186 233943 375189
rect 189165 375184 233943 375186
rect 189165 375128 189170 375184
rect 189226 375128 233882 375184
rect 233938 375128 233943 375184
rect 189165 375126 233943 375128
rect 189165 375123 189231 375126
rect 233877 375123 233943 375126
rect 358077 375186 358143 375189
rect 358854 375186 358860 375188
rect 358077 375184 358860 375186
rect 358077 375128 358082 375184
rect 358138 375128 358860 375184
rect 358077 375126 358860 375128
rect 358077 375123 358143 375126
rect 358854 375124 358860 375126
rect 358924 375124 358930 375188
rect 159357 374642 159423 374645
rect 166390 374642 166396 374644
rect 159357 374640 166396 374642
rect 159357 374584 159362 374640
rect 159418 374584 166396 374640
rect 159357 374582 166396 374584
rect 159357 374579 159423 374582
rect 166390 374580 166396 374582
rect 166460 374580 166466 374644
rect 341149 374642 341215 374645
rect 378869 374642 378935 374645
rect 341149 374640 378935 374642
rect 341149 374584 341154 374640
rect 341210 374584 378874 374640
rect 378930 374584 378935 374640
rect 341149 374582 378935 374584
rect 341149 374579 341215 374582
rect 378869 374579 378935 374582
rect 62021 374098 62087 374101
rect 214557 374098 214623 374101
rect 62021 374096 214623 374098
rect 62021 374040 62026 374096
rect 62082 374040 214562 374096
rect 214618 374040 214623 374096
rect 62021 374038 214623 374040
rect 62021 374035 62087 374038
rect 214557 374035 214623 374038
rect 221457 374098 221523 374101
rect 253054 374098 253060 374100
rect 221457 374096 253060 374098
rect 221457 374040 221462 374096
rect 221518 374040 253060 374096
rect 221457 374038 253060 374040
rect 221457 374035 221523 374038
rect 253054 374036 253060 374038
rect 253124 374036 253130 374100
rect 279417 374098 279483 374101
rect 281441 374098 281507 374101
rect 279417 374096 281507 374098
rect 279417 374040 279422 374096
rect 279478 374040 281446 374096
rect 281502 374040 281507 374096
rect 279417 374038 281507 374040
rect 279417 374035 279483 374038
rect 281441 374035 281507 374038
rect 76557 373282 76623 373285
rect 172513 373282 172579 373285
rect 76557 373280 172579 373282
rect 76557 373224 76562 373280
rect 76618 373224 172518 373280
rect 172574 373224 172579 373280
rect 76557 373222 172579 373224
rect 76557 373219 76623 373222
rect 172513 373219 172579 373222
rect 177941 373282 178007 373285
rect 357433 373282 357499 373285
rect 177941 373280 357499 373282
rect 177941 373224 177946 373280
rect 178002 373224 357438 373280
rect 357494 373224 357499 373280
rect 177941 373222 357499 373224
rect 177941 373219 178007 373222
rect 357433 373219 357499 373222
rect 114553 372738 114619 372741
rect 385125 372738 385191 372741
rect 385677 372738 385743 372741
rect 114553 372736 385743 372738
rect 114553 372680 114558 372736
rect 114614 372680 385130 372736
rect 385186 372680 385682 372736
rect 385738 372680 385743 372736
rect 114553 372678 385743 372680
rect 114553 372675 114619 372678
rect 385125 372675 385191 372678
rect 385677 372675 385743 372678
rect 18597 372602 18663 372605
rect 153929 372602 153995 372605
rect 18597 372600 153995 372602
rect 18597 372544 18602 372600
rect 18658 372544 153934 372600
rect 153990 372544 153995 372600
rect 18597 372542 153995 372544
rect 18597 372539 18663 372542
rect 153929 372539 153995 372542
rect 195329 372602 195395 372605
rect 365897 372602 365963 372605
rect 195329 372600 365963 372602
rect 195329 372544 195334 372600
rect 195390 372544 365902 372600
rect 365958 372544 365963 372600
rect 195329 372542 365963 372544
rect 195329 372539 195395 372542
rect 365897 372539 365963 372542
rect 73153 371922 73219 371925
rect 119470 371922 119476 371924
rect 73153 371920 119476 371922
rect 73153 371864 73158 371920
rect 73214 371864 119476 371920
rect 73153 371862 119476 371864
rect 73153 371859 73219 371862
rect 119470 371860 119476 371862
rect 119540 371860 119546 371924
rect 195421 371922 195487 371925
rect 331857 371922 331923 371925
rect 371417 371922 371483 371925
rect 195421 371920 371483 371922
rect 195421 371864 195426 371920
rect 195482 371864 331862 371920
rect 331918 371864 371422 371920
rect 371478 371864 371483 371920
rect 195421 371862 371483 371864
rect 195421 371859 195487 371862
rect 331857 371859 331923 371862
rect 371417 371859 371483 371862
rect -960 371378 480 371468
rect 3233 371378 3299 371381
rect -960 371376 3299 371378
rect -960 371320 3238 371376
rect 3294 371320 3299 371376
rect -960 371318 3299 371320
rect -960 371228 480 371318
rect 3233 371315 3299 371318
rect 18597 371378 18663 371381
rect 19241 371378 19307 371381
rect 18597 371376 19307 371378
rect 18597 371320 18602 371376
rect 18658 371320 19246 371376
rect 19302 371320 19307 371376
rect 18597 371318 19307 371320
rect 18597 371315 18663 371318
rect 19241 371315 19307 371318
rect 99281 371378 99347 371381
rect 242893 371378 242959 371381
rect 243629 371378 243695 371381
rect 99281 371376 243695 371378
rect 99281 371320 99286 371376
rect 99342 371320 242898 371376
rect 242954 371320 243634 371376
rect 243690 371320 243695 371376
rect 99281 371318 243695 371320
rect 99281 371315 99347 371318
rect 242893 371315 242959 371318
rect 243629 371315 243695 371318
rect 130469 370698 130535 370701
rect 162117 370698 162183 370701
rect 363229 370698 363295 370701
rect 130469 370696 363295 370698
rect 130469 370640 130474 370696
rect 130530 370640 162122 370696
rect 162178 370640 363234 370696
rect 363290 370640 363295 370696
rect 130469 370638 363295 370640
rect 130469 370635 130535 370638
rect 162117 370635 162183 370638
rect 363229 370635 363295 370638
rect 89621 370562 89687 370565
rect 368657 370562 368723 370565
rect 89621 370560 368723 370562
rect 89621 370504 89626 370560
rect 89682 370504 368662 370560
rect 368718 370504 368723 370560
rect 89621 370502 368723 370504
rect 89621 370499 89687 370502
rect 368657 370499 368723 370502
rect 151077 369202 151143 369205
rect 159357 369202 159423 369205
rect 151077 369200 159423 369202
rect 151077 369144 151082 369200
rect 151138 369144 159362 369200
rect 159418 369144 159423 369200
rect 151077 369142 159423 369144
rect 151077 369139 151143 369142
rect 159357 369139 159423 369142
rect 198774 369140 198780 369204
rect 198844 369202 198850 369204
rect 218697 369202 218763 369205
rect 198844 369200 218763 369202
rect 198844 369144 218702 369200
rect 218758 369144 218763 369200
rect 198844 369142 218763 369144
rect 198844 369140 198850 369142
rect 218697 369139 218763 369142
rect 63401 369066 63467 369069
rect 130377 369066 130443 369069
rect 63401 369064 130443 369066
rect 63401 369008 63406 369064
rect 63462 369008 130382 369064
rect 130438 369008 130443 369064
rect 63401 369006 130443 369008
rect 63401 369003 63467 369006
rect 130377 369003 130443 369006
rect 137369 369066 137435 369069
rect 154062 369066 154068 369068
rect 137369 369064 154068 369066
rect 137369 369008 137374 369064
rect 137430 369008 154068 369064
rect 137369 369006 154068 369008
rect 137369 369003 137435 369006
rect 154062 369004 154068 369006
rect 154132 369004 154138 369068
rect 187141 369066 187207 369069
rect 307753 369066 307819 369069
rect 187141 369064 307819 369066
rect 187141 369008 187146 369064
rect 187202 369008 307758 369064
rect 307814 369008 307819 369064
rect 187141 369006 307819 369008
rect 187141 369003 187207 369006
rect 307753 369003 307819 369006
rect 122097 368522 122163 368525
rect 122741 368522 122807 368525
rect 195329 368522 195395 368525
rect 122097 368520 195395 368522
rect 122097 368464 122102 368520
rect 122158 368464 122746 368520
rect 122802 368464 195334 368520
rect 195390 368464 195395 368520
rect 122097 368462 195395 368464
rect 122097 368459 122163 368462
rect 122741 368459 122807 368462
rect 195329 368459 195395 368462
rect 182909 368386 182975 368389
rect 186814 368386 186820 368388
rect 182909 368384 186820 368386
rect 182909 368328 182914 368384
rect 182970 368328 186820 368384
rect 182909 368326 186820 368328
rect 182909 368323 182975 368326
rect 186814 368324 186820 368326
rect 186884 368324 186890 368388
rect 69790 367644 69796 367708
rect 69860 367706 69866 367708
rect 69860 367646 84210 367706
rect 69860 367644 69866 367646
rect 84150 367298 84210 367646
rect 200614 367644 200620 367708
rect 200684 367706 200690 367708
rect 258073 367706 258139 367709
rect 200684 367704 258139 367706
rect 200684 367648 258078 367704
rect 258134 367648 258139 367704
rect 200684 367646 258139 367648
rect 200684 367644 200690 367646
rect 258073 367643 258139 367646
rect 93117 367570 93183 367573
rect 287053 367570 287119 367573
rect 287646 367570 287652 367572
rect 93117 367568 287652 367570
rect 93117 367512 93122 367568
rect 93178 367512 287058 367568
rect 287114 367512 287652 367568
rect 93117 367510 287652 367512
rect 93117 367507 93183 367510
rect 287053 367507 287119 367510
rect 287646 367508 287652 367510
rect 287716 367508 287722 367572
rect 131021 367434 131087 367437
rect 203517 367434 203583 367437
rect 131021 367432 203583 367434
rect 131021 367376 131026 367432
rect 131082 367376 203522 367432
rect 203578 367376 203583 367432
rect 131021 367374 203583 367376
rect 131021 367371 131087 367374
rect 203517 367371 203583 367374
rect 86953 367298 87019 367301
rect 166206 367298 166212 367300
rect 84150 367296 166212 367298
rect 84150 367240 86958 367296
rect 87014 367240 166212 367296
rect 84150 367238 166212 367240
rect 86953 367235 87019 367238
rect 166206 367236 166212 367238
rect 166276 367236 166282 367300
rect 283373 367162 283439 367165
rect 283557 367162 283623 367165
rect 285581 367162 285647 367165
rect 418797 367162 418863 367165
rect 283373 367160 418863 367162
rect 283373 367104 283378 367160
rect 283434 367104 283562 367160
rect 283618 367104 285586 367160
rect 285642 367104 418802 367160
rect 418858 367104 418863 367160
rect 283373 367102 418863 367104
rect 283373 367099 283439 367102
rect 283557 367099 283623 367102
rect 285581 367099 285647 367102
rect 418797 367099 418863 367102
rect 56501 366346 56567 366349
rect 283373 366346 283439 366349
rect 56501 366344 283439 366346
rect 56501 366288 56506 366344
rect 56562 366288 283378 366344
rect 283434 366288 283439 366344
rect 56501 366286 283439 366288
rect 56501 366283 56567 366286
rect 283373 366283 283439 366286
rect 353937 366346 354003 366349
rect 368565 366346 368631 366349
rect 353937 366344 368631 366346
rect 353937 366288 353942 366344
rect 353998 366288 368570 366344
rect 368626 366288 368631 366344
rect 353937 366286 368631 366288
rect 353937 366283 354003 366286
rect 368565 366283 368631 366286
rect 91093 365802 91159 365805
rect 92289 365802 92355 365805
rect 222837 365802 222903 365805
rect 91093 365800 222903 365802
rect 91093 365744 91098 365800
rect 91154 365744 92294 365800
rect 92350 365744 222842 365800
rect 222898 365744 222903 365800
rect 91093 365742 222903 365744
rect 91093 365739 91159 365742
rect 92289 365739 92355 365742
rect 222837 365739 222903 365742
rect 582373 365122 582439 365125
rect 583520 365122 584960 365212
rect 582373 365120 584960 365122
rect 582373 365064 582378 365120
rect 582434 365064 584960 365120
rect 582373 365062 584960 365064
rect 582373 365059 582439 365062
rect 75821 364986 75887 364989
rect 194542 364986 194548 364988
rect 75821 364984 194548 364986
rect 75821 364928 75826 364984
rect 75882 364928 194548 364984
rect 75821 364926 194548 364928
rect 75821 364923 75887 364926
rect 194542 364924 194548 364926
rect 194612 364924 194618 364988
rect 201401 364986 201467 364989
rect 253197 364986 253263 364989
rect 361757 364986 361823 364989
rect 201401 364984 253263 364986
rect 201401 364928 201406 364984
rect 201462 364928 253202 364984
rect 253258 364928 253263 364984
rect 201401 364926 253263 364928
rect 201401 364923 201467 364926
rect 253197 364923 253263 364926
rect 277350 364984 361823 364986
rect 277350 364928 361762 364984
rect 361818 364928 361823 364984
rect 583520 364972 584960 365062
rect 277350 364926 361823 364928
rect 124121 364442 124187 364445
rect 267590 364442 267596 364444
rect 124121 364440 267596 364442
rect 124121 364384 124126 364440
rect 124182 364384 267596 364440
rect 124121 364382 267596 364384
rect 124121 364379 124187 364382
rect 267590 364380 267596 364382
rect 267660 364442 267666 364444
rect 277350 364442 277410 364926
rect 361757 364923 361823 364926
rect 267660 364382 277410 364442
rect 267660 364380 267666 364382
rect 69657 363762 69723 363765
rect 166257 363762 166323 363765
rect 69657 363760 166323 363762
rect 69657 363704 69662 363760
rect 69718 363704 166262 363760
rect 166318 363704 166323 363760
rect 69657 363702 166323 363704
rect 69657 363699 69723 363702
rect 166257 363699 166323 363702
rect 143349 363626 143415 363629
rect 245009 363626 245075 363629
rect 143349 363624 245075 363626
rect 143349 363568 143354 363624
rect 143410 363568 245014 363624
rect 245070 363568 245075 363624
rect 143349 363566 245075 363568
rect 143349 363563 143415 363566
rect 245009 363563 245075 363566
rect 147581 363082 147647 363085
rect 216121 363082 216187 363085
rect 147581 363080 216187 363082
rect 147581 363024 147586 363080
rect 147642 363024 216126 363080
rect 216182 363024 216187 363080
rect 147581 363022 216187 363024
rect 147581 363019 147647 363022
rect 216121 363019 216187 363022
rect 64689 362266 64755 362269
rect 357525 362266 357591 362269
rect 64689 362264 357591 362266
rect 64689 362208 64694 362264
rect 64750 362208 357530 362264
rect 357586 362208 357591 362264
rect 64689 362206 357591 362208
rect 64689 362203 64755 362206
rect 357525 362203 357591 362206
rect 194869 361858 194935 361861
rect 113130 361856 194935 361858
rect 113130 361800 194874 361856
rect 194930 361800 194935 361856
rect 113130 361798 194935 361800
rect 108757 361724 108823 361725
rect 108757 361720 108804 361724
rect 108868 361722 108874 361724
rect 113130 361722 113190 361798
rect 194869 361795 194935 361798
rect 202781 361858 202847 361861
rect 203006 361858 203012 361860
rect 202781 361856 203012 361858
rect 202781 361800 202786 361856
rect 202842 361800 203012 361856
rect 202781 361798 203012 361800
rect 202781 361795 202847 361798
rect 203006 361796 203012 361798
rect 203076 361796 203082 361860
rect 108757 361664 108762 361720
rect 108757 361660 108804 361664
rect 108868 361662 113190 361722
rect 133781 361722 133847 361725
rect 320173 361722 320239 361725
rect 320817 361722 320883 361725
rect 133781 361720 320883 361722
rect 133781 361664 133786 361720
rect 133842 361664 320178 361720
rect 320234 361664 320822 361720
rect 320878 361664 320883 361720
rect 133781 361662 320883 361664
rect 108868 361660 108874 361662
rect 108757 361659 108823 361660
rect 133781 361659 133847 361662
rect 320173 361659 320239 361662
rect 320817 361659 320883 361662
rect 338021 361042 338087 361045
rect 354438 361042 354444 361044
rect 338021 361040 354444 361042
rect 338021 360984 338026 361040
rect 338082 360984 354444 361040
rect 338021 360982 354444 360984
rect 338021 360979 338087 360982
rect 354438 360980 354444 360982
rect 354508 360980 354514 361044
rect 103421 360906 103487 360909
rect 147581 360906 147647 360909
rect 356278 360906 356284 360908
rect 103421 360904 147647 360906
rect 103421 360848 103426 360904
rect 103482 360848 147586 360904
rect 147642 360848 147647 360904
rect 103421 360846 147647 360848
rect 103421 360843 103487 360846
rect 147581 360843 147647 360846
rect 190410 360846 356284 360906
rect 189073 360362 189139 360365
rect 190410 360362 190470 360846
rect 356278 360844 356284 360846
rect 356348 360844 356354 360908
rect 132450 360360 190470 360362
rect 132450 360304 189078 360360
rect 189134 360304 190470 360360
rect 132450 360302 190470 360304
rect 75729 360226 75795 360229
rect 100753 360226 100819 360229
rect 101121 360226 101187 360229
rect 75729 360224 101187 360226
rect 75729 360168 75734 360224
rect 75790 360168 100758 360224
rect 100814 360168 101126 360224
rect 101182 360168 101187 360224
rect 75729 360166 101187 360168
rect 75729 360163 75795 360166
rect 100753 360163 100819 360166
rect 101121 360163 101187 360166
rect 124806 360164 124812 360228
rect 124876 360226 124882 360228
rect 125501 360226 125567 360229
rect 132450 360226 132510 360302
rect 189073 360299 189139 360302
rect 124876 360224 132510 360226
rect 124876 360168 125506 360224
rect 125562 360168 132510 360224
rect 124876 360166 132510 360168
rect 151721 360226 151787 360229
rect 337377 360226 337443 360229
rect 338021 360226 338087 360229
rect 151721 360224 338087 360226
rect 151721 360168 151726 360224
rect 151782 360168 337382 360224
rect 337438 360168 338026 360224
rect 338082 360168 338087 360224
rect 151721 360166 338087 360168
rect 124876 360164 124882 360166
rect 125501 360163 125567 360166
rect 151721 360163 151787 360166
rect 337377 360163 337443 360166
rect 338021 360163 338087 360166
rect 166390 360028 166396 360092
rect 166460 360090 166466 360092
rect 353293 360090 353359 360093
rect 166460 360088 353359 360090
rect 166460 360032 353298 360088
rect 353354 360032 353359 360088
rect 166460 360030 353359 360032
rect 166460 360028 166466 360030
rect 353293 360027 353359 360030
rect 81014 359348 81020 359412
rect 81084 359410 81090 359412
rect 356094 359410 356100 359412
rect 81084 359350 356100 359410
rect 81084 359348 81090 359350
rect 356094 359348 356100 359350
rect 356164 359348 356170 359412
rect 152457 359274 152523 359277
rect 153101 359274 153167 359277
rect 152457 359272 153167 359274
rect 152457 359216 152462 359272
rect 152518 359216 153106 359272
rect 153162 359216 153167 359272
rect 152457 359214 153167 359216
rect 152457 359211 152523 359214
rect 153101 359211 153167 359214
rect 3325 359002 3391 359005
rect 151813 359002 151879 359005
rect 152641 359002 152707 359005
rect 3325 359000 152707 359002
rect 3325 358944 3330 359000
rect 3386 358944 151818 359000
rect 151874 358944 152646 359000
rect 152702 358944 152707 359000
rect 3325 358942 152707 358944
rect 3325 358939 3391 358942
rect 151813 358939 151879 358942
rect 152641 358939 152707 358942
rect 153101 358866 153167 358869
rect 216029 358866 216095 358869
rect 153101 358864 216095 358866
rect 153101 358808 153106 358864
rect 153162 358808 216034 358864
rect 216090 358808 216095 358864
rect 153101 358806 216095 358808
rect 153101 358803 153167 358806
rect 216029 358803 216095 358806
rect -960 358458 480 358548
rect 3417 358458 3483 358461
rect -960 358456 3483 358458
rect -960 358400 3422 358456
rect 3478 358400 3483 358456
rect -960 358398 3483 358400
rect -960 358308 480 358398
rect 3417 358395 3483 358398
rect 324681 358186 324747 358189
rect 325601 358186 325667 358189
rect 328453 358186 328519 358189
rect 324681 358184 328519 358186
rect 324681 358128 324686 358184
rect 324742 358128 325606 358184
rect 325662 358128 328458 358184
rect 328514 358128 328519 358184
rect 324681 358126 328519 358128
rect 324681 358123 324747 358126
rect 325601 358123 325667 358126
rect 328453 358123 328519 358126
rect 89529 358050 89595 358053
rect 146109 358050 146175 358053
rect 89529 358048 146175 358050
rect 89529 357992 89534 358048
rect 89590 357992 146114 358048
rect 146170 357992 146175 358048
rect 89529 357990 146175 357992
rect 89529 357987 89595 357990
rect 146109 357987 146175 357990
rect 322289 358050 322355 358053
rect 353334 358050 353340 358052
rect 322289 358048 353340 358050
rect 322289 357992 322294 358048
rect 322350 357992 353340 358048
rect 322289 357990 353340 357992
rect 322289 357987 322355 357990
rect 353334 357988 353340 357990
rect 353404 357988 353410 358052
rect 111057 357642 111123 357645
rect 111558 357642 111564 357644
rect 111057 357640 111564 357642
rect 111057 357584 111062 357640
rect 111118 357584 111564 357640
rect 111057 357582 111564 357584
rect 111057 357579 111123 357582
rect 111558 357580 111564 357582
rect 111628 357642 111634 357644
rect 191230 357642 191236 357644
rect 111628 357582 191236 357642
rect 111628 357580 111634 357582
rect 191230 357580 191236 357582
rect 191300 357580 191306 357644
rect 65977 357506 66043 357509
rect 324681 357506 324747 357509
rect 65977 357504 324747 357506
rect 65977 357448 65982 357504
rect 66038 357448 324686 357504
rect 324742 357448 324747 357504
rect 65977 357446 324747 357448
rect 65977 357443 66043 357446
rect 324681 357443 324747 357446
rect 170489 356826 170555 356829
rect 205633 356826 205699 356829
rect 170489 356824 205699 356826
rect 170489 356768 170494 356824
rect 170550 356768 205638 356824
rect 205694 356768 205699 356824
rect 170489 356766 205699 356768
rect 170489 356763 170555 356766
rect 205633 356763 205699 356766
rect 124029 356690 124095 356693
rect 194041 356690 194107 356693
rect 124029 356688 194107 356690
rect 124029 356632 124034 356688
rect 124090 356632 194046 356688
rect 194102 356632 194107 356688
rect 124029 356630 194107 356632
rect 124029 356627 124095 356630
rect 194041 356627 194107 356630
rect 194869 356690 194935 356693
rect 232497 356690 232563 356693
rect 194869 356688 232563 356690
rect 194869 356632 194874 356688
rect 194930 356632 232502 356688
rect 232558 356632 232563 356688
rect 194869 356630 232563 356632
rect 194869 356627 194935 356630
rect 232497 356627 232563 356630
rect 122189 356282 122255 356285
rect 191097 356282 191163 356285
rect 122189 356280 191163 356282
rect 122189 356224 122194 356280
rect 122250 356224 191102 356280
rect 191158 356224 191163 356280
rect 122189 356222 191163 356224
rect 122189 356219 122255 356222
rect 191097 356219 191163 356222
rect 69606 356084 69612 356148
rect 69676 356146 69682 356148
rect 149421 356146 149487 356149
rect 69676 356144 149487 356146
rect 69676 356088 149426 356144
rect 149482 356088 149487 356144
rect 69676 356086 149487 356088
rect 69676 356084 69682 356086
rect 149421 356083 149487 356086
rect 99189 355466 99255 355469
rect 251214 355466 251220 355468
rect 99189 355464 251220 355466
rect 99189 355408 99194 355464
rect 99250 355408 251220 355464
rect 99189 355406 251220 355408
rect 99189 355403 99255 355406
rect 251214 355404 251220 355406
rect 251284 355404 251290 355468
rect 59169 355330 59235 355333
rect 221457 355330 221523 355333
rect 59169 355328 221523 355330
rect 59169 355272 59174 355328
rect 59230 355272 221462 355328
rect 221518 355272 221523 355328
rect 59169 355270 221523 355272
rect 59169 355267 59235 355270
rect 221457 355267 221523 355270
rect 87597 353970 87663 353973
rect 120717 353970 120783 353973
rect 196709 353970 196775 353973
rect 87597 353968 196775 353970
rect 87597 353912 87602 353968
rect 87658 353912 120722 353968
rect 120778 353912 196714 353968
rect 196770 353912 196775 353968
rect 87597 353910 196775 353912
rect 87597 353907 87663 353910
rect 120717 353907 120783 353910
rect 196709 353907 196775 353910
rect 99373 353562 99439 353565
rect 100518 353562 100524 353564
rect 99373 353560 100524 353562
rect 99373 353504 99378 353560
rect 99434 353504 100524 353560
rect 99373 353502 100524 353504
rect 99373 353499 99439 353502
rect 100518 353500 100524 353502
rect 100588 353562 100594 353564
rect 147673 353562 147739 353565
rect 192569 353562 192635 353565
rect 100588 353502 103530 353562
rect 100588 353500 100594 353502
rect 103470 353426 103530 353502
rect 147673 353560 192635 353562
rect 147673 353504 147678 353560
rect 147734 353504 192574 353560
rect 192630 353504 192635 353560
rect 147673 353502 192635 353504
rect 147673 353499 147739 353502
rect 192569 353499 192635 353502
rect 174537 353426 174603 353429
rect 228449 353426 228515 353429
rect 103470 353424 174603 353426
rect 103470 353368 174542 353424
rect 174598 353368 174603 353424
rect 103470 353366 174603 353368
rect 174537 353363 174603 353366
rect 195286 353424 228515 353426
rect 195286 353368 228454 353424
rect 228510 353368 228515 353424
rect 195286 353366 228515 353368
rect 173801 353290 173867 353293
rect 195286 353290 195346 353366
rect 228449 353363 228515 353366
rect 173801 353288 195346 353290
rect 173801 353232 173806 353288
rect 173862 353232 195346 353288
rect 173801 353230 195346 353232
rect 173801 353227 173867 353230
rect 79869 352746 79935 352749
rect 111057 352746 111123 352749
rect 79869 352744 111123 352746
rect 79869 352688 79874 352744
rect 79930 352688 111062 352744
rect 111118 352688 111123 352744
rect 79869 352686 111123 352688
rect 79869 352683 79935 352686
rect 111057 352683 111123 352686
rect 100661 352610 100727 352613
rect 173801 352610 173867 352613
rect 100661 352608 173867 352610
rect 100661 352552 100666 352608
rect 100722 352552 173806 352608
rect 173862 352552 173867 352608
rect 100661 352550 173867 352552
rect 100661 352547 100727 352550
rect 173801 352547 173867 352550
rect 180241 352610 180307 352613
rect 326337 352610 326403 352613
rect 180241 352608 326403 352610
rect 180241 352552 180246 352608
rect 180302 352552 326342 352608
rect 326398 352552 326403 352608
rect 180241 352550 326403 352552
rect 180241 352547 180307 352550
rect 326337 352547 326403 352550
rect 106917 351930 106983 351933
rect 107469 351930 107535 351933
rect 246297 351930 246363 351933
rect 106917 351928 246363 351930
rect 106917 351872 106922 351928
rect 106978 351872 107474 351928
rect 107530 351872 246302 351928
rect 246358 351872 246363 351928
rect 106917 351870 246363 351872
rect 106917 351867 106983 351870
rect 107469 351867 107535 351870
rect 246297 351867 246363 351870
rect 582925 351930 582991 351933
rect 583520 351930 584960 352020
rect 582925 351928 584960 351930
rect 582925 351872 582930 351928
rect 582986 351872 584960 351928
rect 582925 351870 584960 351872
rect 582925 351867 582991 351870
rect 583520 351780 584960 351870
rect 269757 351250 269823 351253
rect 319437 351250 319503 351253
rect 258030 351248 319503 351250
rect 258030 351192 269762 351248
rect 269818 351192 319442 351248
rect 319498 351192 319503 351248
rect 258030 351190 319503 351192
rect 86217 351114 86283 351117
rect 124949 351114 125015 351117
rect 86217 351112 125015 351114
rect 86217 351056 86222 351112
rect 86278 351056 124954 351112
rect 125010 351056 125015 351112
rect 86217 351054 125015 351056
rect 86217 351051 86283 351054
rect 124949 351051 125015 351054
rect 147765 350842 147831 350845
rect 148317 350842 148383 350845
rect 173341 350842 173407 350845
rect 147765 350840 173407 350842
rect 147765 350784 147770 350840
rect 147826 350784 148322 350840
rect 148378 350784 173346 350840
rect 173402 350784 173407 350840
rect 147765 350782 173407 350784
rect 147765 350779 147831 350782
rect 148317 350779 148383 350782
rect 173341 350779 173407 350782
rect 130377 350706 130443 350709
rect 131021 350706 131087 350709
rect 258030 350706 258090 351190
rect 269757 351187 269823 351190
rect 319437 351187 319503 351190
rect 378133 351114 378199 351117
rect 130377 350704 258090 350706
rect 130377 350648 130382 350704
rect 130438 350648 131026 350704
rect 131082 350648 258090 350704
rect 130377 350646 258090 350648
rect 296670 351112 378199 351114
rect 296670 351056 378138 351112
rect 378194 351056 378199 351112
rect 296670 351054 378199 351056
rect 130377 350643 130443 350646
rect 131021 350643 131087 350646
rect 114369 350570 114435 350573
rect 295926 350570 295932 350572
rect 114369 350568 295932 350570
rect 114369 350512 114374 350568
rect 114430 350512 295932 350568
rect 114369 350510 295932 350512
rect 114369 350507 114435 350510
rect 295926 350508 295932 350510
rect 295996 350570 296002 350572
rect 296670 350570 296730 351054
rect 378133 351051 378199 351054
rect 295996 350510 296730 350570
rect 295996 350508 296002 350510
rect 149421 350434 149487 350437
rect 187601 350434 187667 350437
rect 149421 350432 187667 350434
rect 149421 350376 149426 350432
rect 149482 350376 187606 350432
rect 187662 350376 187667 350432
rect 149421 350374 187667 350376
rect 149421 350371 149487 350374
rect 187601 350371 187667 350374
rect 187601 350026 187667 350029
rect 188521 350026 188587 350029
rect 187601 350024 188587 350026
rect 187601 349968 187606 350024
rect 187662 349968 188526 350024
rect 188582 349968 188587 350024
rect 187601 349966 188587 349968
rect 187601 349963 187667 349966
rect 188521 349963 188587 349966
rect 67950 349692 67956 349756
rect 68020 349754 68026 349756
rect 86309 349754 86375 349757
rect 68020 349752 86375 349754
rect 68020 349696 86314 349752
rect 86370 349696 86375 349752
rect 68020 349694 86375 349696
rect 68020 349692 68026 349694
rect 86309 349691 86375 349694
rect 99189 349754 99255 349757
rect 147673 349754 147739 349757
rect 99189 349752 147739 349754
rect 99189 349696 99194 349752
rect 99250 349696 147678 349752
rect 147734 349696 147739 349752
rect 99189 349694 147739 349696
rect 99189 349691 99255 349694
rect 147673 349691 147739 349694
rect 171869 349754 171935 349757
rect 222193 349754 222259 349757
rect 171869 349752 222259 349754
rect 171869 349696 171874 349752
rect 171930 349696 222198 349752
rect 222254 349696 222259 349752
rect 171869 349694 222259 349696
rect 171869 349691 171935 349694
rect 222193 349691 222259 349694
rect 118550 349148 118556 349212
rect 118620 349210 118626 349212
rect 118877 349210 118943 349213
rect 265065 349210 265131 349213
rect 118620 349208 265131 349210
rect 118620 349152 118882 349208
rect 118938 349152 265070 349208
rect 265126 349152 265131 349208
rect 118620 349150 265131 349152
rect 118620 349148 118626 349150
rect 118877 349147 118943 349150
rect 265065 349147 265131 349150
rect 104985 349074 105051 349077
rect 121678 349074 121684 349076
rect 104985 349072 121684 349074
rect 104985 349016 104990 349072
rect 105046 349016 121684 349072
rect 104985 349014 121684 349016
rect 104985 349011 105051 349014
rect 121678 349012 121684 349014
rect 121748 349074 121754 349076
rect 209129 349074 209195 349077
rect 209681 349074 209747 349077
rect 121748 349072 209747 349074
rect 121748 349016 209134 349072
rect 209190 349016 209686 349072
rect 209742 349016 209747 349072
rect 121748 349014 209747 349016
rect 121748 349012 121754 349014
rect 209129 349011 209195 349014
rect 209681 349011 209747 349014
rect 67766 348876 67772 348940
rect 67836 348938 67842 348940
rect 125593 348938 125659 348941
rect 126789 348938 126855 348941
rect 67836 348936 126855 348938
rect 67836 348880 125598 348936
rect 125654 348880 126794 348936
rect 126850 348880 126855 348936
rect 67836 348878 126855 348880
rect 67836 348876 67842 348878
rect 125593 348875 125659 348878
rect 126789 348875 126855 348878
rect 208894 348468 208900 348532
rect 208964 348530 208970 348532
rect 227713 348530 227779 348533
rect 208964 348528 227779 348530
rect 208964 348472 227718 348528
rect 227774 348472 227779 348528
rect 208964 348470 227779 348472
rect 208964 348468 208970 348470
rect 227713 348467 227779 348470
rect 67357 348394 67423 348397
rect 195513 348394 195579 348397
rect 67357 348392 195579 348394
rect 67357 348336 67362 348392
rect 67418 348336 195518 348392
rect 195574 348336 195579 348392
rect 67357 348334 195579 348336
rect 67357 348331 67423 348334
rect 195513 348331 195579 348334
rect 209129 348394 209195 348397
rect 236637 348394 236703 348397
rect 209129 348392 236703 348394
rect 209129 348336 209134 348392
rect 209190 348336 236642 348392
rect 236698 348336 236703 348392
rect 209129 348334 236703 348336
rect 209129 348331 209195 348334
rect 236637 348331 236703 348334
rect 133689 347850 133755 347853
rect 180333 347850 180399 347853
rect 133689 347848 180399 347850
rect 133689 347792 133694 347848
rect 133750 347792 180338 347848
rect 180394 347792 180399 347848
rect 133689 347790 180399 347792
rect 133689 347787 133755 347790
rect 180333 347787 180399 347790
rect 263685 347714 263751 347717
rect 264237 347714 264303 347717
rect 263685 347712 264303 347714
rect 263685 347656 263690 347712
rect 263746 347656 264242 347712
rect 264298 347656 264303 347712
rect 263685 347654 264303 347656
rect 263685 347651 263751 347654
rect 264237 347651 264303 347654
rect 66662 346972 66668 347036
rect 66732 347034 66738 347036
rect 140037 347034 140103 347037
rect 66732 347032 140103 347034
rect 66732 346976 140042 347032
rect 140098 346976 140103 347032
rect 66732 346974 140103 346976
rect 66732 346972 66738 346974
rect 140037 346971 140103 346974
rect 150341 347034 150407 347037
rect 178677 347034 178743 347037
rect 150341 347032 178743 347034
rect 150341 346976 150346 347032
rect 150402 346976 178682 347032
rect 178738 346976 178743 347032
rect 150341 346974 178743 346976
rect 150341 346971 150407 346974
rect 178677 346971 178743 346974
rect 60457 346626 60523 346629
rect 197997 346626 198063 346629
rect 60457 346624 198063 346626
rect 60457 346568 60462 346624
rect 60518 346568 198002 346624
rect 198058 346568 198063 346624
rect 60457 346566 198063 346568
rect 60457 346563 60523 346566
rect 197997 346563 198063 346566
rect 119889 346490 119955 346493
rect 264237 346490 264303 346493
rect 119889 346488 264303 346490
rect 119889 346432 119894 346488
rect 119950 346432 264242 346488
rect 264298 346432 264303 346488
rect 119889 346430 264303 346432
rect 119889 346427 119955 346430
rect 264237 346427 264303 346430
rect 176653 345946 176719 345949
rect 177849 345946 177915 345949
rect 192477 345946 192543 345949
rect 176653 345944 192543 345946
rect 176653 345888 176658 345944
rect 176714 345888 177854 345944
rect 177910 345888 192482 345944
rect 192538 345888 192543 345944
rect 176653 345886 192543 345888
rect 176653 345883 176719 345886
rect 177849 345883 177915 345886
rect 192477 345883 192543 345886
rect 92381 345810 92447 345813
rect 94446 345810 94452 345812
rect 92381 345808 94452 345810
rect 92381 345752 92386 345808
rect 92442 345752 94452 345808
rect 92381 345750 94452 345752
rect 92381 345747 92447 345750
rect 94446 345748 94452 345750
rect 94516 345810 94522 345812
rect 186814 345810 186820 345812
rect 94516 345750 186820 345810
rect 94516 345748 94522 345750
rect 186814 345748 186820 345750
rect 186884 345748 186890 345812
rect 100569 345674 100635 345677
rect 176653 345674 176719 345677
rect 100569 345672 176719 345674
rect 100569 345616 100574 345672
rect 100630 345616 176658 345672
rect 176714 345616 176719 345672
rect 100569 345614 176719 345616
rect 100569 345611 100635 345614
rect 176653 345611 176719 345614
rect 178677 345674 178743 345677
rect 324313 345674 324379 345677
rect 178677 345672 324379 345674
rect 178677 345616 178682 345672
rect 178738 345616 324318 345672
rect 324374 345616 324379 345672
rect 178677 345614 324379 345616
rect 178677 345611 178743 345614
rect 324313 345611 324379 345614
rect 248505 345540 248571 345541
rect 248454 345538 248460 345540
rect -960 345402 480 345492
rect 248414 345478 248460 345538
rect 248524 345536 248571 345540
rect 248566 345480 248571 345536
rect 248454 345476 248460 345478
rect 248524 345476 248571 345480
rect 248505 345475 248571 345476
rect 3509 345402 3575 345405
rect -960 345400 3575 345402
rect -960 345344 3514 345400
rect 3570 345344 3575 345400
rect -960 345342 3575 345344
rect -960 345252 480 345342
rect 3509 345339 3575 345342
rect 73061 345130 73127 345133
rect 176009 345130 176075 345133
rect 73061 345128 176075 345130
rect 73061 345072 73066 345128
rect 73122 345072 176014 345128
rect 176070 345072 176075 345128
rect 73061 345070 176075 345072
rect 73061 345067 73127 345070
rect 176009 345067 176075 345070
rect 197353 345130 197419 345133
rect 198406 345130 198412 345132
rect 197353 345128 198412 345130
rect 197353 345072 197358 345128
rect 197414 345072 198412 345128
rect 197353 345070 198412 345072
rect 197353 345067 197419 345070
rect 198406 345068 198412 345070
rect 198476 345068 198482 345132
rect 156505 344994 156571 344997
rect 196566 344994 196572 344996
rect 156505 344992 196572 344994
rect 156505 344936 156510 344992
rect 156566 344936 196572 344992
rect 156505 344934 196572 344936
rect 156505 344931 156571 344934
rect 196566 344932 196572 344934
rect 196636 344932 196642 344996
rect 134517 344314 134583 344317
rect 162761 344314 162827 344317
rect 207657 344314 207723 344317
rect 134517 344312 207723 344314
rect 134517 344256 134522 344312
rect 134578 344256 162766 344312
rect 162822 344256 207662 344312
rect 207718 344256 207723 344312
rect 134517 344254 207723 344256
rect 134517 344251 134583 344254
rect 162761 344251 162827 344254
rect 207657 344251 207723 344254
rect 224309 344314 224375 344317
rect 243537 344314 243603 344317
rect 224309 344312 243603 344314
rect 224309 344256 224314 344312
rect 224370 344256 243542 344312
rect 243598 344256 243603 344312
rect 224309 344254 243603 344256
rect 224309 344251 224375 344254
rect 243537 344251 243603 344254
rect 128997 343906 129063 343909
rect 129641 343906 129707 343909
rect 156454 343906 156460 343908
rect 128997 343904 156460 343906
rect 128997 343848 129002 343904
rect 129058 343848 129646 343904
rect 129702 343848 156460 343904
rect 128997 343846 156460 343848
rect 128997 343843 129063 343846
rect 129641 343843 129707 343846
rect 156454 343844 156460 343846
rect 156524 343844 156530 343908
rect 95141 343770 95207 343773
rect 167637 343770 167703 343773
rect 95141 343768 167703 343770
rect 95141 343712 95146 343768
rect 95202 343712 167642 343768
rect 167698 343712 167703 343768
rect 95141 343710 167703 343712
rect 95141 343707 95207 343710
rect 167637 343707 167703 343710
rect 202229 343770 202295 343773
rect 225597 343770 225663 343773
rect 202229 343768 225663 343770
rect 202229 343712 202234 343768
rect 202290 343712 225602 343768
rect 225658 343712 225663 343768
rect 202229 343710 225663 343712
rect 202229 343707 202295 343710
rect 225597 343707 225663 343710
rect 64781 342954 64847 342957
rect 111742 342954 111748 342956
rect 64781 342952 111748 342954
rect 64781 342896 64786 342952
rect 64842 342896 111748 342952
rect 64781 342894 111748 342896
rect 64781 342891 64847 342894
rect 111742 342892 111748 342894
rect 111812 342892 111818 342956
rect 127801 342546 127867 342549
rect 189901 342546 189967 342549
rect 127801 342544 189967 342546
rect 127801 342488 127806 342544
rect 127862 342488 189906 342544
rect 189962 342488 189967 342544
rect 127801 342486 189967 342488
rect 127801 342483 127867 342486
rect 189901 342483 189967 342486
rect 81433 342410 81499 342413
rect 230422 342410 230428 342412
rect 81433 342408 230428 342410
rect 81433 342352 81438 342408
rect 81494 342352 230428 342408
rect 81433 342350 230428 342352
rect 81433 342347 81499 342350
rect 230422 342348 230428 342350
rect 230492 342348 230498 342412
rect 111609 342274 111675 342277
rect 304993 342274 305059 342277
rect 305637 342274 305703 342277
rect 111609 342272 305703 342274
rect 111609 342216 111614 342272
rect 111670 342216 304998 342272
rect 305054 342216 305642 342272
rect 305698 342216 305703 342272
rect 111609 342214 305703 342216
rect 111609 342211 111675 342214
rect 304993 342211 305059 342214
rect 305637 342211 305703 342214
rect 159449 342138 159515 342141
rect 162853 342138 162919 342141
rect 159449 342136 162919 342138
rect 159449 342080 159454 342136
rect 159510 342080 162858 342136
rect 162914 342080 162919 342136
rect 159449 342078 162919 342080
rect 159449 342075 159515 342078
rect 162853 342075 162919 342078
rect 97809 341594 97875 341597
rect 157742 341594 157748 341596
rect 97809 341592 157748 341594
rect 97809 341536 97814 341592
rect 97870 341536 157748 341592
rect 97809 341534 157748 341536
rect 97809 341531 97875 341534
rect 157742 341532 157748 341534
rect 157812 341532 157818 341596
rect 243629 341594 243695 341597
rect 291837 341594 291903 341597
rect 243629 341592 291903 341594
rect 243629 341536 243634 341592
rect 243690 341536 291842 341592
rect 291898 341536 291903 341592
rect 243629 341534 291903 341536
rect 243629 341531 243695 341534
rect 291837 341531 291903 341534
rect 67357 341458 67423 341461
rect 219934 341458 219940 341460
rect 67357 341456 219940 341458
rect 67357 341400 67362 341456
rect 67418 341400 219940 341456
rect 67357 341398 219940 341400
rect 67357 341395 67423 341398
rect 219934 341396 219940 341398
rect 220004 341396 220010 341460
rect 231117 341458 231183 341461
rect 367369 341458 367435 341461
rect 231117 341456 367435 341458
rect 231117 341400 231122 341456
rect 231178 341400 367374 341456
rect 367430 341400 367435 341456
rect 231117 341398 367435 341400
rect 231117 341395 231183 341398
rect 367369 341395 367435 341398
rect 137185 340914 137251 340917
rect 137921 340914 137987 340917
rect 206461 340914 206527 340917
rect 137185 340912 206527 340914
rect 137185 340856 137190 340912
rect 137246 340856 137926 340912
rect 137982 340856 206466 340912
rect 206522 340856 206527 340912
rect 137185 340854 206527 340856
rect 137185 340851 137251 340854
rect 137921 340851 137987 340854
rect 206461 340851 206527 340854
rect 157742 340716 157748 340780
rect 157812 340778 157818 340780
rect 158478 340778 158484 340780
rect 157812 340718 158484 340778
rect 157812 340716 157818 340718
rect 158478 340716 158484 340718
rect 158548 340778 158554 340780
rect 226977 340778 227043 340781
rect 158548 340776 227043 340778
rect 158548 340720 226982 340776
rect 227038 340720 227043 340776
rect 158548 340718 227043 340720
rect 158548 340716 158554 340718
rect 226977 340715 227043 340718
rect 126329 340234 126395 340237
rect 126881 340234 126947 340237
rect 143441 340234 143507 340237
rect 158846 340234 158852 340236
rect 126329 340232 132510 340234
rect 126329 340176 126334 340232
rect 126390 340176 126886 340232
rect 126942 340176 132510 340232
rect 126329 340174 132510 340176
rect 126329 340171 126395 340174
rect 126881 340171 126947 340174
rect 16481 340098 16547 340101
rect 56409 340098 56475 340101
rect 100753 340098 100819 340101
rect 16481 340096 100819 340098
rect 16481 340040 16486 340096
rect 16542 340040 56414 340096
rect 56470 340040 100758 340096
rect 100814 340040 100819 340096
rect 16481 340038 100819 340040
rect 132450 340098 132510 340174
rect 143441 340232 158852 340234
rect 143441 340176 143446 340232
rect 143502 340176 158852 340232
rect 143441 340174 158852 340176
rect 143441 340171 143507 340174
rect 158846 340172 158852 340174
rect 158916 340172 158922 340236
rect 156505 340098 156571 340101
rect 132450 340096 156571 340098
rect 132450 340040 156510 340096
rect 156566 340040 156571 340096
rect 132450 340038 156571 340040
rect 16481 340035 16547 340038
rect 56409 340035 56475 340038
rect 100753 340035 100819 340038
rect 156505 340035 156571 340038
rect 216121 340098 216187 340101
rect 347037 340098 347103 340101
rect 216121 340096 347103 340098
rect 216121 340040 216126 340096
rect 216182 340040 347042 340096
rect 347098 340040 347103 340096
rect 216121 340038 347103 340040
rect 216121 340035 216187 340038
rect 347037 340035 347103 340038
rect 114645 339962 114711 339965
rect 115790 339962 115796 339964
rect 114645 339960 115796 339962
rect 114645 339904 114650 339960
rect 114706 339904 115796 339960
rect 114645 339902 115796 339904
rect 114645 339899 114711 339902
rect 115790 339900 115796 339902
rect 115860 339900 115866 339964
rect 110229 339690 110295 339693
rect 139393 339690 139459 339693
rect 110229 339688 139459 339690
rect 110229 339632 110234 339688
rect 110290 339632 139398 339688
rect 139454 339632 139459 339688
rect 110229 339630 139459 339632
rect 110229 339627 110295 339630
rect 139393 339627 139459 339630
rect 158805 339690 158871 339693
rect 185577 339690 185643 339693
rect 158805 339688 185643 339690
rect 158805 339632 158810 339688
rect 158866 339632 185582 339688
rect 185638 339632 185643 339688
rect 158805 339630 185643 339632
rect 158805 339627 158871 339630
rect 185577 339627 185643 339630
rect 115790 339492 115796 339556
rect 115860 339554 115866 339556
rect 164969 339554 165035 339557
rect 115860 339552 165035 339554
rect 115860 339496 164974 339552
rect 165030 339496 165035 339552
rect 115860 339494 165035 339496
rect 115860 339492 115866 339494
rect 164969 339491 165035 339494
rect 67766 338812 67772 338876
rect 67836 338874 67842 338876
rect 116577 338874 116643 338877
rect 67836 338872 116643 338874
rect 67836 338816 116582 338872
rect 116638 338816 116643 338872
rect 67836 338814 116643 338816
rect 67836 338812 67842 338814
rect 116577 338811 116643 338814
rect 96337 338738 96403 338741
rect 191649 338738 191715 338741
rect 254577 338738 254643 338741
rect 96337 338736 254643 338738
rect 96337 338680 96342 338736
rect 96398 338680 191654 338736
rect 191710 338680 254582 338736
rect 254638 338680 254643 338736
rect 96337 338678 254643 338680
rect 96337 338675 96403 338678
rect 191649 338675 191715 338678
rect 254577 338675 254643 338678
rect 583520 338452 584960 338692
rect 124949 338330 125015 338333
rect 177481 338330 177547 338333
rect 124949 338328 177547 338330
rect 124949 338272 124954 338328
rect 125010 338272 177486 338328
rect 177542 338272 177547 338328
rect 124949 338270 177547 338272
rect 124949 338267 125015 338270
rect 177481 338267 177547 338270
rect 154205 338194 154271 338197
rect 222929 338194 222995 338197
rect 154205 338192 222995 338194
rect 154205 338136 154210 338192
rect 154266 338136 222934 338192
rect 222990 338136 222995 338192
rect 154205 338134 222995 338136
rect 154205 338131 154271 338134
rect 222929 338131 222995 338134
rect 155217 338058 155283 338061
rect 157241 338058 157307 338061
rect 155217 338056 157307 338058
rect 155217 338000 155222 338056
rect 155278 338000 157246 338056
rect 157302 338000 157307 338056
rect 155217 337998 157307 338000
rect 155217 337995 155283 337998
rect 157241 337995 157307 337998
rect 159357 338058 159423 338061
rect 160870 338058 160876 338060
rect 159357 338056 160876 338058
rect 159357 338000 159362 338056
rect 159418 338000 160876 338056
rect 159357 337998 160876 338000
rect 159357 337995 159423 337998
rect 160870 337996 160876 337998
rect 160940 337996 160946 338060
rect 169109 337514 169175 337517
rect 206369 337514 206435 337517
rect 169109 337512 206435 337514
rect 169109 337456 169114 337512
rect 169170 337456 206374 337512
rect 206430 337456 206435 337512
rect 169109 337454 206435 337456
rect 169109 337451 169175 337454
rect 206369 337451 206435 337454
rect 213126 337452 213132 337516
rect 213196 337514 213202 337516
rect 235257 337514 235323 337517
rect 213196 337512 235323 337514
rect 213196 337456 235262 337512
rect 235318 337456 235323 337512
rect 213196 337454 235323 337456
rect 213196 337452 213202 337454
rect 235257 337451 235323 337454
rect 66110 337316 66116 337380
rect 66180 337378 66186 337380
rect 104157 337378 104223 337381
rect 66180 337376 104223 337378
rect 66180 337320 104162 337376
rect 104218 337320 104223 337376
rect 66180 337318 104223 337320
rect 66180 337316 66186 337318
rect 104157 337315 104223 337318
rect 156781 337378 156847 337381
rect 165153 337378 165219 337381
rect 156781 337376 165219 337378
rect 156781 337320 156786 337376
rect 156842 337320 165158 337376
rect 165214 337320 165219 337376
rect 156781 337318 165219 337320
rect 156781 337315 156847 337318
rect 165153 337315 165219 337318
rect 169518 337316 169524 337380
rect 169588 337378 169594 337380
rect 313273 337378 313339 337381
rect 169588 337376 313339 337378
rect 169588 337320 313278 337376
rect 313334 337320 313339 337376
rect 169588 337318 313339 337320
rect 169588 337316 169594 337318
rect 313273 337315 313339 337318
rect 133965 336970 134031 336973
rect 154757 336970 154823 336973
rect 133965 336968 154823 336970
rect 133965 336912 133970 336968
rect 134026 336912 154762 336968
rect 154818 336912 154823 336968
rect 133965 336910 154823 336912
rect 133965 336907 134031 336910
rect 154757 336907 154823 336910
rect 64597 336834 64663 336837
rect 170397 336834 170463 336837
rect 64597 336832 170463 336834
rect 64597 336776 64602 336832
rect 64658 336776 170402 336832
rect 170458 336776 170463 336832
rect 64597 336774 170463 336776
rect 64597 336771 64663 336774
rect 170397 336771 170463 336774
rect 83825 336018 83891 336021
rect 106917 336018 106983 336021
rect 83825 336016 106983 336018
rect 83825 335960 83830 336016
rect 83886 335960 106922 336016
rect 106978 335960 106983 336016
rect 83825 335958 106983 335960
rect 83825 335955 83891 335958
rect 106917 335955 106983 335958
rect 148409 336018 148475 336021
rect 158805 336018 158871 336021
rect 148409 336016 158871 336018
rect 148409 335960 148414 336016
rect 148470 335960 158810 336016
rect 158866 335960 158871 336016
rect 148409 335958 158871 335960
rect 148409 335955 148475 335958
rect 158805 335955 158871 335958
rect 97809 335746 97875 335749
rect 181713 335746 181779 335749
rect 97809 335744 181779 335746
rect 97809 335688 97814 335744
rect 97870 335688 181718 335744
rect 181774 335688 181779 335744
rect 97809 335686 181779 335688
rect 97809 335683 97875 335686
rect 181713 335683 181779 335686
rect 134885 335610 134951 335613
rect 247677 335610 247743 335613
rect 134885 335608 247743 335610
rect 134885 335552 134890 335608
rect 134946 335552 247682 335608
rect 247738 335552 247743 335608
rect 134885 335550 247743 335552
rect 134885 335547 134951 335550
rect 247677 335547 247743 335550
rect 158897 335474 158963 335477
rect 338113 335474 338179 335477
rect 158897 335472 338179 335474
rect 158897 335416 158902 335472
rect 158958 335416 338118 335472
rect 338174 335416 338179 335472
rect 158897 335414 338179 335416
rect 158897 335411 158963 335414
rect 338113 335411 338179 335414
rect 63125 334658 63191 334661
rect 140037 334658 140103 334661
rect 63125 334656 140103 334658
rect 63125 334600 63130 334656
rect 63186 334600 140042 334656
rect 140098 334600 140103 334656
rect 63125 334598 140103 334600
rect 63125 334595 63191 334598
rect 140037 334595 140103 334598
rect 152457 334658 152523 334661
rect 583661 334658 583727 334661
rect 152457 334656 583727 334658
rect 152457 334600 152462 334656
rect 152518 334600 583666 334656
rect 583722 334600 583727 334656
rect 152457 334598 583727 334600
rect 152457 334595 152523 334598
rect 583661 334595 583727 334598
rect 141877 334250 141943 334253
rect 238937 334250 239003 334253
rect 141877 334248 239003 334250
rect 141877 334192 141882 334248
rect 141938 334192 238942 334248
rect 238998 334192 239003 334248
rect 141877 334190 239003 334192
rect 141877 334187 141943 334190
rect 238937 334187 239003 334190
rect 117037 334114 117103 334117
rect 247217 334114 247283 334117
rect 117037 334112 247283 334114
rect 117037 334056 117042 334112
rect 117098 334056 247222 334112
rect 247278 334056 247283 334112
rect 117037 334054 247283 334056
rect 117037 334051 117103 334054
rect 247217 334051 247283 334054
rect 132493 333298 132559 333301
rect 152590 333298 152596 333300
rect 132493 333296 152596 333298
rect 132493 333240 132498 333296
rect 132554 333240 152596 333296
rect 132493 333238 152596 333240
rect 132493 333235 132559 333238
rect 152590 333236 152596 333238
rect 152660 333236 152666 333300
rect 153009 332890 153075 332893
rect 252645 332890 252711 332893
rect 153009 332888 252711 332890
rect 153009 332832 153014 332888
rect 153070 332832 252650 332888
rect 252706 332832 252711 332888
rect 153009 332830 252711 332832
rect 153009 332827 153075 332830
rect 252645 332827 252711 332830
rect 65885 332754 65951 332757
rect 165889 332754 165955 332757
rect 65885 332752 165955 332754
rect 65885 332696 65890 332752
rect 65946 332696 165894 332752
rect 165950 332696 165955 332752
rect 65885 332694 165955 332696
rect 65885 332691 65951 332694
rect 165889 332691 165955 332694
rect 69790 332556 69796 332620
rect 69860 332618 69866 332620
rect 229737 332618 229803 332621
rect 69860 332616 229803 332618
rect 69860 332560 229742 332616
rect 229798 332560 229803 332616
rect 69860 332558 229803 332560
rect 69860 332556 69866 332558
rect 229737 332555 229803 332558
rect 130745 332482 130811 332485
rect 134517 332482 134583 332485
rect 130745 332480 134583 332482
rect -960 332196 480 332436
rect 130745 332424 130750 332480
rect 130806 332424 134522 332480
rect 134578 332424 134583 332480
rect 130745 332422 134583 332424
rect 130745 332419 130811 332422
rect 134517 332419 134583 332422
rect 144545 332210 144611 332213
rect 145557 332210 145623 332213
rect 144545 332208 145623 332210
rect 144545 332152 144550 332208
rect 144606 332152 145562 332208
rect 145618 332152 145623 332208
rect 144545 332150 145623 332152
rect 144545 332147 144611 332150
rect 145557 332147 145623 332150
rect 189901 331938 189967 331941
rect 239121 331938 239187 331941
rect 189901 331936 239187 331938
rect 189901 331880 189906 331936
rect 189962 331880 239126 331936
rect 239182 331880 239187 331936
rect 189901 331878 239187 331880
rect 189901 331875 189967 331878
rect 239121 331875 239187 331878
rect 60641 331802 60707 331805
rect 79961 331802 80027 331805
rect 60641 331800 80027 331802
rect 60641 331744 60646 331800
rect 60702 331744 79966 331800
rect 80022 331744 80027 331800
rect 60641 331742 80027 331744
rect 60641 331739 60707 331742
rect 79961 331739 80027 331742
rect 82670 331740 82676 331804
rect 82740 331802 82746 331804
rect 101397 331802 101463 331805
rect 82740 331800 101463 331802
rect 82740 331744 101402 331800
rect 101458 331744 101463 331800
rect 82740 331742 101463 331744
rect 82740 331740 82746 331742
rect 101397 331739 101463 331742
rect 103237 331802 103303 331805
rect 128997 331802 129063 331805
rect 103237 331800 129063 331802
rect 103237 331744 103242 331800
rect 103298 331744 129002 331800
rect 129058 331744 129063 331800
rect 103237 331742 129063 331744
rect 103237 331739 103303 331742
rect 128997 331739 129063 331742
rect 135713 331802 135779 331805
rect 144821 331802 144887 331805
rect 177246 331802 177252 331804
rect 135713 331800 177252 331802
rect 135713 331744 135718 331800
rect 135774 331744 144826 331800
rect 144882 331744 177252 331800
rect 135713 331742 177252 331744
rect 135713 331739 135779 331742
rect 144821 331739 144887 331742
rect 177246 331740 177252 331742
rect 177316 331740 177322 331804
rect 203517 331802 203583 331805
rect 270585 331802 270651 331805
rect 203517 331800 270651 331802
rect 203517 331744 203522 331800
rect 203578 331744 270590 331800
rect 270646 331744 270651 331800
rect 203517 331742 270651 331744
rect 203517 331739 203583 331742
rect 270585 331739 270651 331742
rect 157333 331530 157399 331533
rect 157742 331530 157748 331532
rect 157333 331528 157748 331530
rect 157333 331472 157338 331528
rect 157394 331472 157748 331528
rect 157333 331470 157748 331472
rect 157333 331467 157399 331470
rect 157742 331468 157748 331470
rect 157812 331468 157818 331532
rect 124673 331394 124739 331397
rect 125501 331394 125567 331397
rect 124673 331392 125567 331394
rect 124673 331336 124678 331392
rect 124734 331336 125506 331392
rect 125562 331336 125567 331392
rect 124673 331334 125567 331336
rect 124673 331331 124739 331334
rect 125501 331331 125567 331334
rect 134241 331394 134307 331397
rect 141918 331394 141924 331396
rect 134241 331392 141924 331394
rect 134241 331336 134246 331392
rect 134302 331336 141924 331392
rect 134241 331334 141924 331336
rect 134241 331331 134307 331334
rect 141918 331332 141924 331334
rect 141988 331332 141994 331396
rect 149697 331394 149763 331397
rect 150249 331394 150315 331397
rect 178718 331394 178724 331396
rect 149697 331392 178724 331394
rect 149697 331336 149702 331392
rect 149758 331336 150254 331392
rect 150310 331336 178724 331392
rect 149697 331334 178724 331336
rect 149697 331331 149763 331334
rect 150249 331331 150315 331334
rect 178718 331332 178724 331334
rect 178788 331332 178794 331396
rect 75177 331258 75243 331261
rect 75678 331258 75684 331260
rect 75177 331256 75684 331258
rect 75177 331200 75182 331256
rect 75238 331200 75684 331256
rect 75177 331198 75684 331200
rect 75177 331195 75243 331198
rect 75678 331196 75684 331198
rect 75748 331258 75754 331260
rect 75821 331258 75887 331261
rect 75748 331256 75887 331258
rect 75748 331200 75826 331256
rect 75882 331200 75887 331256
rect 75748 331198 75887 331200
rect 75748 331196 75754 331198
rect 75821 331195 75887 331198
rect 94221 331258 94287 331261
rect 94865 331258 94931 331261
rect 145281 331258 145347 331261
rect 150433 331258 150499 331261
rect 94221 331256 135178 331258
rect 94221 331200 94226 331256
rect 94282 331200 94870 331256
rect 94926 331200 135178 331256
rect 94221 331198 135178 331200
rect 94221 331195 94287 331198
rect 94865 331195 94931 331198
rect 135118 331122 135178 331198
rect 145281 331256 150499 331258
rect 145281 331200 145286 331256
rect 145342 331200 150438 331256
rect 150494 331200 150499 331256
rect 145281 331198 150499 331200
rect 145281 331195 145347 331198
rect 150433 331195 150499 331198
rect 152641 331258 152707 331261
rect 297357 331258 297423 331261
rect 298001 331258 298067 331261
rect 152641 331256 298067 331258
rect 152641 331200 152646 331256
rect 152702 331200 297362 331256
rect 297418 331200 298006 331256
rect 298062 331200 298067 331256
rect 152641 331198 298067 331200
rect 152641 331195 152707 331198
rect 297357 331195 297423 331198
rect 298001 331195 298067 331198
rect 230473 331122 230539 331125
rect 231209 331122 231275 331125
rect 135118 331120 231275 331122
rect 135118 331064 230478 331120
rect 230534 331064 231214 331120
rect 231270 331064 231275 331120
rect 135118 331062 231275 331064
rect 230473 331059 230539 331062
rect 231209 331059 231275 331062
rect 136449 330034 136515 330037
rect 236637 330034 236703 330037
rect 136449 330032 236703 330034
rect 136449 329976 136454 330032
rect 136510 329976 236642 330032
rect 236698 329976 236703 330032
rect 136449 329974 236703 329976
rect 136449 329971 136515 329974
rect 236637 329971 236703 329974
rect 35157 329898 35223 329901
rect 124949 329898 125015 329901
rect 35157 329896 125015 329898
rect 35157 329840 35162 329896
rect 35218 329840 124954 329896
rect 125010 329840 125015 329896
rect 35157 329838 125015 329840
rect 35157 329835 35223 329838
rect 124949 329835 125015 329838
rect 151854 329836 151860 329900
rect 151924 329898 151930 329900
rect 156965 329898 157031 329901
rect 151924 329896 157031 329898
rect 151924 329840 156970 329896
rect 157026 329840 157031 329896
rect 151924 329838 157031 329840
rect 151924 329836 151930 329838
rect 156965 329835 157031 329838
rect 155953 329762 156019 329765
rect 157190 329762 157196 329764
rect 155953 329760 157196 329762
rect 155953 329704 155958 329760
rect 156014 329704 157196 329760
rect 155953 329702 157196 329704
rect 155953 329699 156019 329702
rect 157190 329700 157196 329702
rect 157260 329700 157266 329764
rect 156689 329626 156755 329629
rect 160185 329626 160251 329629
rect 156689 329624 160251 329626
rect 156689 329568 156694 329624
rect 156750 329568 160190 329624
rect 160246 329568 160251 329624
rect 156689 329566 160251 329568
rect 156689 329563 156755 329566
rect 160185 329563 160251 329566
rect 69381 329490 69447 329493
rect 69381 329488 69490 329490
rect 69381 329432 69386 329488
rect 69442 329432 69490 329488
rect 69381 329427 69490 329432
rect 77150 329428 77156 329492
rect 77220 329490 77226 329492
rect 77477 329490 77543 329493
rect 77220 329488 77543 329490
rect 77220 329432 77482 329488
rect 77538 329432 77543 329488
rect 77220 329430 77543 329432
rect 77220 329428 77226 329430
rect 77477 329427 77543 329430
rect 69430 328916 69490 329427
rect 152641 329220 152707 329221
rect 142286 329156 142292 329220
rect 142356 329218 142362 329220
rect 151670 329218 151676 329220
rect 142356 329158 151676 329218
rect 142356 329156 142362 329158
rect 151670 329156 151676 329158
rect 151740 329156 151746 329220
rect 152590 329218 152596 329220
rect 152550 329158 152596 329218
rect 152660 329216 152707 329220
rect 152702 329160 152707 329216
rect 152590 329156 152596 329158
rect 152660 329156 152707 329160
rect 152641 329155 152707 329156
rect 157425 329082 157491 329085
rect 203517 329082 203583 329085
rect 157425 329080 203583 329082
rect 157425 329024 157430 329080
rect 157486 329024 203522 329080
rect 203578 329024 203583 329080
rect 157425 329022 203583 329024
rect 157425 329019 157491 329022
rect 203517 329019 203583 329022
rect 374637 328810 374703 328813
rect 156646 328808 374703 328810
rect 156646 328752 374642 328808
rect 374698 328752 374703 328808
rect 156646 328750 374703 328752
rect 156646 328644 156706 328750
rect 374637 328747 374703 328750
rect 259545 328540 259611 328541
rect 259494 328538 259500 328540
rect 259454 328478 259500 328538
rect 259564 328536 259611 328540
rect 259606 328480 259611 328536
rect 259494 328476 259500 328478
rect 259564 328476 259611 328480
rect 259545 328475 259611 328476
rect 69422 328340 69428 328404
rect 69492 328340 69498 328404
rect 166206 328340 166212 328404
rect 166276 328402 166282 328404
rect 168097 328402 168163 328405
rect 166276 328400 168163 328402
rect 166276 328344 168102 328400
rect 168158 328344 168163 328400
rect 166276 328342 168163 328344
rect 166276 328340 166282 328342
rect 69430 327828 69490 328340
rect 168097 328339 168163 328342
rect 156873 327722 156939 327725
rect 162945 327722 163011 327725
rect 156873 327720 163011 327722
rect 156873 327664 156878 327720
rect 156934 327664 162950 327720
rect 163006 327664 163011 327720
rect 156873 327662 163011 327664
rect 156873 327659 156939 327662
rect 162945 327659 163011 327662
rect 158897 327586 158963 327589
rect 156676 327584 158963 327586
rect 156676 327528 158902 327584
rect 158958 327528 158963 327584
rect 156676 327526 158963 327528
rect 158897 327523 158963 327526
rect 156781 327314 156847 327317
rect 238661 327314 238727 327317
rect 156781 327312 238727 327314
rect 156781 327256 156786 327312
rect 156842 327256 238666 327312
rect 238722 327256 238727 327312
rect 156781 327254 238727 327256
rect 156781 327251 156847 327254
rect 238661 327251 238727 327254
rect 198406 327116 198412 327180
rect 198476 327178 198482 327180
rect 287053 327178 287119 327181
rect 198476 327176 287119 327178
rect 198476 327120 287058 327176
rect 287114 327120 287119 327176
rect 198476 327118 287119 327120
rect 198476 327116 198482 327118
rect 287053 327115 287119 327118
rect 66897 326770 66963 326773
rect 66897 326768 68908 326770
rect 66897 326712 66902 326768
rect 66958 326712 68908 326768
rect 66897 326710 68908 326712
rect 66897 326707 66963 326710
rect 158897 326498 158963 326501
rect 156676 326496 158963 326498
rect 156676 326440 158902 326496
rect 158958 326440 158963 326496
rect 156676 326438 158963 326440
rect 158897 326435 158963 326438
rect 160185 326498 160251 326501
rect 241973 326498 242039 326501
rect 160185 326496 242039 326498
rect 160185 326440 160190 326496
rect 160246 326440 241978 326496
rect 242034 326440 242039 326496
rect 160185 326438 242039 326440
rect 160185 326435 160251 326438
rect 241973 326435 242039 326438
rect 158989 326362 159055 326365
rect 244733 326362 244799 326365
rect 158989 326360 244799 326362
rect 158989 326304 158994 326360
rect 159050 326304 244738 326360
rect 244794 326304 244799 326360
rect 158989 326302 244799 326304
rect 158989 326299 159055 326302
rect 244733 326299 244799 326302
rect 66110 325620 66116 325684
rect 66180 325682 66186 325684
rect 66180 325622 68908 325682
rect 66180 325620 66186 325622
rect 157742 325410 157748 325412
rect 156676 325350 157748 325410
rect 157742 325348 157748 325350
rect 157812 325348 157818 325412
rect 582833 325274 582899 325277
rect 583520 325274 584960 325364
rect 582833 325272 584960 325274
rect 582833 325216 582838 325272
rect 582894 325216 584960 325272
rect 582833 325214 584960 325216
rect 582833 325211 582899 325214
rect 205173 325138 205239 325141
rect 216029 325138 216095 325141
rect 205173 325136 216095 325138
rect 205173 325080 205178 325136
rect 205234 325080 216034 325136
rect 216090 325080 216095 325136
rect 583520 325124 584960 325214
rect 205173 325078 216095 325080
rect 205173 325075 205239 325078
rect 216029 325075 216095 325078
rect 165153 325002 165219 325005
rect 237414 325002 237420 325004
rect 165153 325000 237420 325002
rect 165153 324944 165158 325000
rect 165214 324944 237420 325000
rect 165153 324942 237420 324944
rect 165153 324939 165219 324942
rect 237414 324940 237420 324942
rect 237484 324940 237490 325004
rect 238109 325002 238175 325005
rect 255262 325002 255268 325004
rect 238109 325000 255268 325002
rect 238109 324944 238114 325000
rect 238170 324944 255268 325000
rect 238109 324942 255268 324944
rect 238109 324939 238175 324942
rect 255262 324940 255268 324942
rect 255332 324940 255338 325004
rect 67725 324594 67791 324597
rect 67725 324592 68908 324594
rect 67725 324536 67730 324592
rect 67786 324536 68908 324592
rect 67725 324534 68908 324536
rect 67725 324531 67791 324534
rect 157742 324396 157748 324460
rect 157812 324458 157818 324460
rect 158161 324458 158227 324461
rect 157812 324456 158227 324458
rect 157812 324400 158166 324456
rect 158222 324400 158227 324456
rect 157812 324398 158227 324400
rect 157812 324396 157818 324398
rect 158161 324395 158227 324398
rect 158713 324322 158779 324325
rect 156676 324320 158779 324322
rect 156676 324264 158718 324320
rect 158774 324264 158779 324320
rect 156676 324262 158779 324264
rect 158713 324259 158779 324262
rect 69422 323988 69428 324052
rect 69492 323988 69498 324052
rect 69430 323476 69490 323988
rect 206277 323778 206343 323781
rect 249742 323778 249748 323780
rect 206277 323776 249748 323778
rect 206277 323720 206282 323776
rect 206338 323720 249748 323776
rect 206277 323718 249748 323720
rect 206277 323715 206343 323718
rect 249742 323716 249748 323718
rect 249812 323716 249818 323780
rect 165061 323642 165127 323645
rect 242249 323642 242315 323645
rect 165061 323640 242315 323642
rect 165061 323584 165066 323640
rect 165122 323584 242254 323640
rect 242310 323584 242315 323640
rect 165061 323582 242315 323584
rect 165061 323579 165127 323582
rect 242249 323579 242315 323582
rect 158897 323234 158963 323237
rect 156676 323232 158963 323234
rect 156676 323176 158902 323232
rect 158958 323176 158963 323232
rect 156676 323174 158963 323176
rect 158897 323171 158963 323174
rect 244733 322826 244799 322829
rect 289721 322826 289787 322829
rect 244733 322824 289787 322826
rect 244733 322768 244738 322824
rect 244794 322768 289726 322824
rect 289782 322768 289787 322824
rect 244733 322766 289787 322768
rect 244733 322763 244799 322766
rect 289721 322763 289787 322766
rect 66253 322418 66319 322421
rect 66253 322416 68908 322418
rect 66253 322360 66258 322416
rect 66314 322360 68908 322416
rect 66253 322358 68908 322360
rect 66253 322355 66319 322358
rect 158713 322148 158779 322149
rect 158662 322146 158668 322148
rect 156676 322086 158668 322146
rect 158732 322144 158779 322148
rect 158774 322088 158779 322144
rect 158662 322084 158668 322086
rect 158732 322084 158779 322088
rect 158713 322083 158779 322084
rect 164969 322146 165035 322149
rect 225689 322146 225755 322149
rect 164969 322144 225755 322146
rect 164969 322088 164974 322144
rect 165030 322088 225694 322144
rect 225750 322088 225755 322144
rect 164969 322086 225755 322088
rect 164969 322083 165035 322086
rect 225689 322083 225755 322086
rect 244733 321740 244799 321741
rect 244733 321738 244780 321740
rect 244688 321736 244780 321738
rect 244688 321680 244738 321736
rect 244688 321678 244780 321680
rect 244733 321676 244780 321678
rect 244844 321676 244850 321740
rect 244733 321675 244799 321676
rect 219341 321602 219407 321605
rect 323025 321602 323091 321605
rect 219341 321600 323091 321602
rect 219341 321544 219346 321600
rect 219402 321544 323030 321600
rect 323086 321544 323091 321600
rect 219341 321542 323091 321544
rect 219341 321539 219407 321542
rect 323025 321539 323091 321542
rect 66805 321330 66871 321333
rect 66805 321328 68908 321330
rect 66805 321272 66810 321328
rect 66866 321272 68908 321328
rect 66805 321270 68908 321272
rect 66805 321267 66871 321270
rect 158713 321058 158779 321061
rect 156676 321056 158779 321058
rect 156676 321000 158718 321056
rect 158774 321000 158779 321056
rect 156676 320998 158779 321000
rect 158713 320995 158779 320998
rect 199377 320922 199443 320925
rect 227662 320922 227668 320924
rect 199377 320920 227668 320922
rect 199377 320864 199382 320920
rect 199438 320864 227668 320920
rect 199377 320862 227668 320864
rect 199377 320859 199443 320862
rect 227662 320860 227668 320862
rect 227732 320860 227738 320924
rect 157190 320724 157196 320788
rect 157260 320786 157266 320788
rect 216029 320786 216095 320789
rect 157260 320784 216095 320786
rect 157260 320728 216034 320784
rect 216090 320728 216095 320784
rect 157260 320726 216095 320728
rect 157260 320724 157266 320726
rect 216029 320723 216095 320726
rect 66897 320242 66963 320245
rect 66897 320240 68908 320242
rect 66897 320184 66902 320240
rect 66958 320184 68908 320240
rect 66897 320182 68908 320184
rect 66897 320179 66963 320182
rect 156646 319426 156706 319940
rect 210734 319500 210740 319564
rect 210804 319562 210810 319564
rect 233877 319562 233943 319565
rect 210804 319560 233943 319562
rect 210804 319504 233882 319560
rect 233938 319504 233943 319560
rect 210804 319502 233943 319504
rect 210804 319500 210810 319502
rect 233877 319499 233943 319502
rect 159357 319426 159423 319429
rect 166390 319426 166396 319428
rect 156646 319424 166396 319426
rect -960 319290 480 319380
rect 156646 319368 159362 319424
rect 159418 319368 166396 319424
rect 156646 319366 166396 319368
rect 159357 319363 159423 319366
rect 166390 319364 166396 319366
rect 166460 319364 166466 319428
rect 206461 319426 206527 319429
rect 344277 319426 344343 319429
rect 206461 319424 344343 319426
rect 206461 319368 206466 319424
rect 206522 319368 344282 319424
rect 344338 319368 344343 319424
rect 206461 319366 344343 319368
rect 206461 319363 206527 319366
rect 344277 319363 344343 319366
rect 4061 319290 4127 319293
rect -960 319288 4127 319290
rect -960 319232 4066 319288
rect 4122 319232 4127 319288
rect -960 319230 4127 319232
rect -960 319140 480 319230
rect 4061 319227 4127 319230
rect 66989 319154 67055 319157
rect 66989 319152 68908 319154
rect 66989 319096 66994 319152
rect 67050 319096 68908 319152
rect 66989 319094 68908 319096
rect 66989 319091 67055 319094
rect 158713 318882 158779 318885
rect 156676 318880 158779 318882
rect 156676 318824 158718 318880
rect 158774 318824 158779 318880
rect 156676 318822 158779 318824
rect 158713 318819 158779 318822
rect 174997 318882 175063 318885
rect 253933 318882 253999 318885
rect 174997 318880 253999 318882
rect 174997 318824 175002 318880
rect 175058 318824 253938 318880
rect 253994 318824 253999 318880
rect 174997 318822 253999 318824
rect 174997 318819 175063 318822
rect 253933 318819 253999 318822
rect 66805 318066 66871 318069
rect 66805 318064 68908 318066
rect 66805 318008 66810 318064
rect 66866 318008 68908 318064
rect 66805 318006 68908 318008
rect 66805 318003 66871 318006
rect 158713 317794 158779 317797
rect 156676 317792 158779 317794
rect 156676 317736 158718 317792
rect 158774 317736 158779 317792
rect 156676 317734 158779 317736
rect 158713 317731 158779 317734
rect 202781 317522 202847 317525
rect 389817 317522 389883 317525
rect 202781 317520 389883 317522
rect 202781 317464 202786 317520
rect 202842 317464 389822 317520
rect 389878 317464 389883 317520
rect 202781 317462 389883 317464
rect 202781 317459 202847 317462
rect 389817 317459 389883 317462
rect 173014 317324 173020 317388
rect 173084 317386 173090 317388
rect 180149 317386 180215 317389
rect 173084 317384 180215 317386
rect 173084 317328 180154 317384
rect 180210 317328 180215 317384
rect 173084 317326 180215 317328
rect 173084 317324 173090 317326
rect 180149 317323 180215 317326
rect 66805 316978 66871 316981
rect 66805 316976 68908 316978
rect 66805 316920 66810 316976
rect 66866 316920 68908 316976
rect 66805 316918 68908 316920
rect 66805 316915 66871 316918
rect 158805 316706 158871 316709
rect 156676 316704 158871 316706
rect 156676 316648 158810 316704
rect 158866 316648 158871 316704
rect 156676 316646 158871 316648
rect 158805 316643 158871 316646
rect 160737 316706 160803 316709
rect 168966 316706 168972 316708
rect 160737 316704 168972 316706
rect 160737 316648 160742 316704
rect 160798 316648 168972 316704
rect 160737 316646 168972 316648
rect 160737 316643 160803 316646
rect 168966 316644 168972 316646
rect 169036 316644 169042 316708
rect 187550 316644 187556 316708
rect 187620 316706 187626 316708
rect 214649 316706 214715 316709
rect 187620 316704 214715 316706
rect 187620 316648 214654 316704
rect 214710 316648 214715 316704
rect 187620 316646 214715 316648
rect 187620 316644 187626 316646
rect 214649 316643 214715 316646
rect 215109 316706 215175 316709
rect 282177 316706 282243 316709
rect 215109 316704 282243 316706
rect 215109 316648 215114 316704
rect 215170 316648 282182 316704
rect 282238 316648 282243 316704
rect 215109 316646 282243 316648
rect 215109 316643 215175 316646
rect 282177 316643 282243 316646
rect 66529 315890 66595 315893
rect 66529 315888 68908 315890
rect 66529 315832 66534 315888
rect 66590 315832 68908 315888
rect 66529 315830 68908 315832
rect 66529 315827 66595 315830
rect 158713 315618 158779 315621
rect 156676 315616 158779 315618
rect 156676 315560 158718 315616
rect 158774 315560 158779 315616
rect 156676 315558 158779 315560
rect 158713 315555 158779 315558
rect 185577 315346 185643 315349
rect 349797 315346 349863 315349
rect 185577 315344 349863 315346
rect 185577 315288 185582 315344
rect 185638 315288 349802 315344
rect 349858 315288 349863 315344
rect 185577 315286 349863 315288
rect 185577 315283 185643 315286
rect 349797 315283 349863 315286
rect 66621 314802 66687 314805
rect 200113 314802 200179 314805
rect 200757 314802 200823 314805
rect 278221 314802 278287 314805
rect 66621 314800 68908 314802
rect 66621 314744 66626 314800
rect 66682 314744 68908 314800
rect 66621 314742 68908 314744
rect 200113 314800 278287 314802
rect 200113 314744 200118 314800
rect 200174 314744 200762 314800
rect 200818 314744 278226 314800
rect 278282 314744 278287 314800
rect 200113 314742 278287 314744
rect 66621 314739 66687 314742
rect 200113 314739 200179 314742
rect 200757 314739 200823 314742
rect 278221 314739 278287 314742
rect 166206 314604 166212 314668
rect 166276 314666 166282 314668
rect 172605 314666 172671 314669
rect 199469 314666 199535 314669
rect 199653 314666 199719 314669
rect 166276 314664 199719 314666
rect 166276 314608 172610 314664
rect 172666 314608 199474 314664
rect 199530 314608 199658 314664
rect 199714 314608 199719 314664
rect 166276 314606 199719 314608
rect 166276 314604 166282 314606
rect 172605 314603 172671 314606
rect 199469 314603 199535 314606
rect 199653 314603 199719 314606
rect 158713 314530 158779 314533
rect 156676 314528 158779 314530
rect 156676 314472 158718 314528
rect 158774 314472 158779 314528
rect 156676 314470 158779 314472
rect 158713 314467 158779 314470
rect 206870 314060 206876 314124
rect 206940 314122 206946 314124
rect 219433 314122 219499 314125
rect 206940 314120 219499 314122
rect 206940 314064 219438 314120
rect 219494 314064 219499 314120
rect 206940 314062 219499 314064
rect 206940 314060 206946 314062
rect 219433 314059 219499 314062
rect 66897 313986 66963 313989
rect 199653 313986 199719 313989
rect 273253 313986 273319 313989
rect 66897 313984 68908 313986
rect 66897 313928 66902 313984
rect 66958 313928 68908 313984
rect 66897 313926 68908 313928
rect 199653 313984 273319 313986
rect 199653 313928 199658 313984
rect 199714 313928 273258 313984
rect 273314 313928 273319 313984
rect 199653 313926 273319 313928
rect 66897 313923 66963 313926
rect 199653 313923 199719 313926
rect 273253 313923 273319 313926
rect 158713 313442 158779 313445
rect 156676 313440 158779 313442
rect 156676 313384 158718 313440
rect 158774 313384 158779 313440
rect 156676 313382 158779 313384
rect 158713 313379 158779 313382
rect 164877 313306 164943 313309
rect 165429 313306 165495 313309
rect 317413 313306 317479 313309
rect 164877 313304 317479 313306
rect 164877 313248 164882 313304
rect 164938 313248 165434 313304
rect 165490 313248 317418 313304
rect 317474 313248 317479 313304
rect 164877 313246 317479 313248
rect 164877 313243 164943 313246
rect 165429 313243 165495 313246
rect 317413 313243 317479 313246
rect 184841 313170 184907 313173
rect 191046 313170 191052 313172
rect 161430 313168 191052 313170
rect 161430 313112 184846 313168
rect 184902 313112 191052 313168
rect 161430 313110 191052 313112
rect 161430 313034 161490 313110
rect 184841 313107 184907 313110
rect 191046 313108 191052 313110
rect 191116 313108 191122 313172
rect 156646 312974 161490 313034
rect 66897 312898 66963 312901
rect 66897 312896 68908 312898
rect 66897 312840 66902 312896
rect 66958 312840 68908 312896
rect 66897 312838 68908 312840
rect 66897 312835 66963 312838
rect 156646 312324 156706 312974
rect 156822 312564 156828 312628
rect 156892 312626 156898 312628
rect 185577 312626 185643 312629
rect 156892 312624 185643 312626
rect 156892 312568 185582 312624
rect 185638 312568 185643 312624
rect 156892 312566 185643 312568
rect 156892 312564 156898 312566
rect 185577 312563 185643 312566
rect 199326 312428 199332 312492
rect 199396 312490 199402 312492
rect 214557 312490 214623 312493
rect 199396 312488 214623 312490
rect 199396 312432 214562 312488
rect 214618 312432 214623 312488
rect 199396 312430 214623 312432
rect 199396 312428 199402 312430
rect 214557 312427 214623 312430
rect 583017 312082 583083 312085
rect 583520 312082 584960 312172
rect 583017 312080 584960 312082
rect 583017 312024 583022 312080
rect 583078 312024 584960 312080
rect 583017 312022 584960 312024
rect 583017 312019 583083 312022
rect 206369 311946 206435 311949
rect 206921 311946 206987 311949
rect 240726 311946 240732 311948
rect 206369 311944 240732 311946
rect 206369 311888 206374 311944
rect 206430 311888 206926 311944
rect 206982 311888 240732 311944
rect 206369 311886 240732 311888
rect 206369 311883 206435 311886
rect 206921 311883 206987 311886
rect 240726 311884 240732 311886
rect 240796 311884 240802 311948
rect 583520 311932 584960 312022
rect 66989 311810 67055 311813
rect 66989 311808 68908 311810
rect 66989 311752 66994 311808
rect 67050 311752 68908 311808
rect 66989 311750 68908 311752
rect 66989 311747 67055 311750
rect 159541 311266 159607 311269
rect 156676 311264 159607 311266
rect 156676 311208 159546 311264
rect 159602 311208 159607 311264
rect 156676 311206 159607 311208
rect 159541 311203 159607 311206
rect 207657 311266 207723 311269
rect 231669 311266 231735 311269
rect 207657 311264 231735 311266
rect 207657 311208 207662 311264
rect 207718 311208 231674 311264
rect 231730 311208 231735 311264
rect 207657 311206 231735 311208
rect 207657 311203 207723 311206
rect 231669 311203 231735 311206
rect 177297 311130 177363 311133
rect 208485 311130 208551 311133
rect 177297 311128 208551 311130
rect 177297 311072 177302 311128
rect 177358 311072 208490 311128
rect 208546 311072 208551 311128
rect 177297 311070 208551 311072
rect 177297 311067 177363 311070
rect 208485 311067 208551 311070
rect 235257 311130 235323 311133
rect 235533 311130 235599 311133
rect 356145 311130 356211 311133
rect 356789 311130 356855 311133
rect 235257 311128 356855 311130
rect 235257 311072 235262 311128
rect 235318 311072 235538 311128
rect 235594 311072 356150 311128
rect 356206 311072 356794 311128
rect 356850 311072 356855 311128
rect 235257 311070 356855 311072
rect 235257 311067 235323 311070
rect 235533 311067 235599 311070
rect 356145 311067 356211 311070
rect 356789 311067 356855 311070
rect 67081 310722 67147 310725
rect 67081 310720 68908 310722
rect 67081 310664 67086 310720
rect 67142 310664 68908 310720
rect 67081 310662 68908 310664
rect 67081 310659 67147 310662
rect 177481 310586 177547 310589
rect 177849 310586 177915 310589
rect 392669 310586 392735 310589
rect 177481 310584 392735 310586
rect 177481 310528 177486 310584
rect 177542 310528 177854 310584
rect 177910 310528 392674 310584
rect 392730 310528 392735 310584
rect 177481 310526 392735 310528
rect 177481 310523 177547 310526
rect 177849 310523 177915 310526
rect 392669 310523 392735 310526
rect 157190 310388 157196 310452
rect 157260 310450 157266 310452
rect 157333 310450 157399 310453
rect 213913 310450 213979 310453
rect 215109 310450 215175 310453
rect 157260 310448 215175 310450
rect 157260 310392 157338 310448
rect 157394 310392 213918 310448
rect 213974 310392 215114 310448
rect 215170 310392 215175 310448
rect 157260 310390 215175 310392
rect 157260 310388 157266 310390
rect 157333 310387 157399 310390
rect 213913 310387 213979 310390
rect 215109 310387 215175 310390
rect 256141 310450 256207 310453
rect 256785 310450 256851 310453
rect 256141 310448 256851 310450
rect 256141 310392 256146 310448
rect 256202 310392 256790 310448
rect 256846 310392 256851 310448
rect 256141 310390 256851 310392
rect 256141 310387 256207 310390
rect 256785 310387 256851 310390
rect 255957 310314 256023 310317
rect 257337 310314 257403 310317
rect 255957 310312 257403 310314
rect 255957 310256 255962 310312
rect 256018 310256 257342 310312
rect 257398 310256 257403 310312
rect 255957 310254 257403 310256
rect 255957 310251 256023 310254
rect 257337 310251 257403 310254
rect 156646 309770 156706 310148
rect 158161 309906 158227 309909
rect 173198 309906 173204 309908
rect 158161 309904 173204 309906
rect 158161 309848 158166 309904
rect 158222 309848 173204 309904
rect 158161 309846 173204 309848
rect 158161 309843 158227 309846
rect 173198 309844 173204 309846
rect 173268 309844 173274 309908
rect 158846 309770 158852 309772
rect 156646 309710 158852 309770
rect 158846 309708 158852 309710
rect 158916 309770 158922 309772
rect 188286 309770 188292 309772
rect 158916 309710 188292 309770
rect 158916 309708 158922 309710
rect 188286 309708 188292 309710
rect 188356 309708 188362 309772
rect 197261 309770 197327 309773
rect 231117 309770 231183 309773
rect 197261 309768 231183 309770
rect 197261 309712 197266 309768
rect 197322 309712 231122 309768
rect 231178 309712 231183 309768
rect 197261 309710 231183 309712
rect 197261 309707 197327 309710
rect 231117 309707 231183 309710
rect 66897 309634 66963 309637
rect 66897 309632 68908 309634
rect 66897 309576 66902 309632
rect 66958 309576 68908 309632
rect 66897 309574 68908 309576
rect 66897 309571 66963 309574
rect 231669 309226 231735 309229
rect 274081 309226 274147 309229
rect 231669 309224 274147 309226
rect 231669 309168 231674 309224
rect 231730 309168 274086 309224
rect 274142 309168 274147 309224
rect 231669 309166 274147 309168
rect 231669 309163 231735 309166
rect 274081 309163 274147 309166
rect 176929 309090 176995 309093
rect 156676 309088 176995 309090
rect 156676 309032 176934 309088
rect 176990 309032 176995 309088
rect 156676 309030 176995 309032
rect 176929 309027 176995 309030
rect 67817 308546 67883 308549
rect 243629 308546 243695 308549
rect 254209 308546 254275 308549
rect 67817 308544 68908 308546
rect 67817 308488 67822 308544
rect 67878 308488 68908 308544
rect 67817 308486 68908 308488
rect 243629 308544 254275 308546
rect 243629 308488 243634 308544
rect 243690 308488 254214 308544
rect 254270 308488 254275 308544
rect 243629 308486 254275 308488
rect 67817 308483 67883 308486
rect 243629 308483 243695 308486
rect 254209 308483 254275 308486
rect 176929 308410 176995 308413
rect 177941 308410 178007 308413
rect 359457 308410 359523 308413
rect 176929 308408 359523 308410
rect 176929 308352 176934 308408
rect 176990 308352 177946 308408
rect 178002 308352 359462 308408
rect 359518 308352 359523 308408
rect 176929 308350 359523 308352
rect 176929 308347 176995 308350
rect 177941 308347 178007 308350
rect 359457 308347 359523 308350
rect 160001 308002 160067 308005
rect 156676 308000 160067 308002
rect 156676 307944 160006 308000
rect 160062 307944 160067 308000
rect 156676 307942 160067 307944
rect 160001 307939 160067 307942
rect 208485 307866 208551 307869
rect 318793 307866 318859 307869
rect 208485 307864 318859 307866
rect 208485 307808 208490 307864
rect 208546 307808 318798 307864
rect 318854 307808 318859 307864
rect 208485 307806 318859 307808
rect 208485 307803 208551 307806
rect 318793 307803 318859 307806
rect 232221 307730 232287 307733
rect 232589 307730 232655 307733
rect 232221 307728 232655 307730
rect 232221 307672 232226 307728
rect 232282 307672 232594 307728
rect 232650 307672 232655 307728
rect 232221 307670 232655 307672
rect 232221 307667 232287 307670
rect 232589 307667 232655 307670
rect 66897 307458 66963 307461
rect 66897 307456 68908 307458
rect 66897 307400 66902 307456
rect 66958 307400 68908 307456
rect 66897 307398 68908 307400
rect 66897 307395 66963 307398
rect 158713 306914 158779 306917
rect 156676 306912 158779 306914
rect 156676 306856 158718 306912
rect 158774 306856 158779 306912
rect 156676 306854 158779 306856
rect 158713 306851 158779 306854
rect 231209 306642 231275 306645
rect 282361 306642 282427 306645
rect 231209 306640 282427 306642
rect 231209 306584 231214 306640
rect 231270 306584 282366 306640
rect 282422 306584 282427 306640
rect 231209 306582 282427 306584
rect 231209 306579 231275 306582
rect 282361 306579 282427 306582
rect 171777 306506 171843 306509
rect 231894 306506 231900 306508
rect 171777 306504 231900 306506
rect 171777 306448 171782 306504
rect 171838 306448 231900 306504
rect 171777 306446 231900 306448
rect 171777 306443 171843 306446
rect 231894 306444 231900 306446
rect 231964 306444 231970 306508
rect 232221 306506 232287 306509
rect 304993 306506 305059 306509
rect 232221 306504 305059 306506
rect 232221 306448 232226 306504
rect 232282 306448 304998 306504
rect 305054 306448 305059 306504
rect 232221 306446 305059 306448
rect 232221 306443 232287 306446
rect 304993 306443 305059 306446
rect 66897 306370 66963 306373
rect 66897 306368 68908 306370
rect -960 306234 480 306324
rect 66897 306312 66902 306368
rect 66958 306312 68908 306368
rect 66897 306310 68908 306312
rect 66897 306307 66963 306310
rect 3509 306234 3575 306237
rect -960 306232 3575 306234
rect -960 306176 3514 306232
rect 3570 306176 3575 306232
rect -960 306174 3575 306176
rect -960 306084 480 306174
rect 3509 306171 3575 306174
rect 158805 305826 158871 305829
rect 156676 305824 158871 305826
rect 156676 305768 158810 305824
rect 158866 305768 158871 305824
rect 156676 305766 158871 305768
rect 158805 305763 158871 305766
rect 159030 305764 159036 305828
rect 159100 305826 159106 305828
rect 174629 305826 174695 305829
rect 159100 305824 174695 305826
rect 159100 305768 174634 305824
rect 174690 305768 174695 305824
rect 159100 305766 174695 305768
rect 159100 305764 159106 305766
rect 174629 305763 174695 305766
rect 159541 305690 159607 305693
rect 220854 305690 220860 305692
rect 159541 305688 220860 305690
rect 159541 305632 159546 305688
rect 159602 305632 220860 305688
rect 159541 305630 220860 305632
rect 159541 305627 159607 305630
rect 220854 305628 220860 305630
rect 220924 305628 220930 305692
rect 65977 305282 66043 305285
rect 65977 305280 68908 305282
rect 65977 305224 65982 305280
rect 66038 305224 68908 305280
rect 65977 305222 68908 305224
rect 65977 305219 66043 305222
rect 180333 305010 180399 305013
rect 180701 305010 180767 305013
rect 278037 305010 278103 305013
rect 180333 305008 278103 305010
rect 180333 304952 180338 305008
rect 180394 304952 180706 305008
rect 180762 304952 278042 305008
rect 278098 304952 278103 305008
rect 180333 304950 278103 304952
rect 180333 304947 180399 304950
rect 180701 304947 180767 304950
rect 278037 304947 278103 304950
rect 202137 304874 202203 304877
rect 218053 304874 218119 304877
rect 202137 304872 218119 304874
rect 202137 304816 202142 304872
rect 202198 304816 218058 304872
rect 218114 304816 218119 304872
rect 202137 304814 218119 304816
rect 202137 304811 202203 304814
rect 218053 304811 218119 304814
rect 158713 304738 158779 304741
rect 156676 304736 158779 304738
rect 156676 304680 158718 304736
rect 158774 304680 158779 304736
rect 156676 304678 158779 304680
rect 158713 304675 158779 304678
rect 66621 304194 66687 304197
rect 169518 304194 169524 304196
rect 66621 304192 68908 304194
rect 66621 304136 66626 304192
rect 66682 304136 68908 304192
rect 66621 304134 68908 304136
rect 161430 304134 169524 304194
rect 66621 304131 66687 304134
rect 161430 303650 161490 304134
rect 169518 304132 169524 304134
rect 169588 304194 169594 304196
rect 182766 304194 182772 304196
rect 169588 304134 182772 304194
rect 169588 304132 169594 304134
rect 182766 304132 182772 304134
rect 182836 304132 182842 304196
rect 223021 304194 223087 304197
rect 279417 304194 279483 304197
rect 223021 304192 279483 304194
rect 223021 304136 223026 304192
rect 223082 304136 279422 304192
rect 279478 304136 279483 304192
rect 223021 304134 279483 304136
rect 223021 304131 223087 304134
rect 279417 304131 279483 304134
rect 256785 303786 256851 303789
rect 171090 303784 256851 303786
rect 171090 303728 256790 303784
rect 256846 303728 256851 303784
rect 171090 303726 256851 303728
rect 156676 303590 161490 303650
rect 164877 303650 164943 303653
rect 165521 303650 165587 303653
rect 171090 303650 171150 303726
rect 256785 303723 256851 303726
rect 164877 303648 171150 303650
rect 164877 303592 164882 303648
rect 164938 303592 165526 303648
rect 165582 303592 171150 303648
rect 164877 303590 171150 303592
rect 164877 303587 164943 303590
rect 165521 303587 165587 303590
rect 65885 303106 65951 303109
rect 65885 303104 68908 303106
rect 65885 303048 65890 303104
rect 65946 303048 68908 303104
rect 65885 303046 68908 303048
rect 65885 303043 65951 303046
rect 211797 302562 211863 302565
rect 248638 302562 248644 302564
rect 211797 302560 248644 302562
rect 156646 302290 156706 302532
rect 211797 302504 211802 302560
rect 211858 302504 248644 302560
rect 211797 302502 248644 302504
rect 211797 302499 211863 302502
rect 248638 302500 248644 302502
rect 248708 302500 248714 302564
rect 168414 302364 168420 302428
rect 168484 302426 168490 302428
rect 169661 302426 169727 302429
rect 168484 302424 169727 302426
rect 168484 302368 169666 302424
rect 169722 302368 169727 302424
rect 168484 302366 169727 302368
rect 168484 302364 168490 302366
rect 169661 302363 169727 302366
rect 187601 302426 187667 302429
rect 272517 302426 272583 302429
rect 187601 302424 272583 302426
rect 187601 302368 187606 302424
rect 187662 302368 272522 302424
rect 272578 302368 272583 302424
rect 187601 302366 272583 302368
rect 187601 302363 187667 302366
rect 272517 302363 272583 302366
rect 318149 302290 318215 302293
rect 156646 302288 318215 302290
rect 156646 302232 318154 302288
rect 318210 302232 318215 302288
rect 156646 302230 318215 302232
rect 318149 302227 318215 302230
rect 66897 302018 66963 302021
rect 66897 302016 68908 302018
rect 66897 301960 66902 302016
rect 66958 301960 68908 302016
rect 66897 301958 68908 301960
rect 66897 301955 66963 301958
rect 66713 300930 66779 300933
rect 156646 300930 156706 301444
rect 197118 301412 197124 301476
rect 197188 301474 197194 301476
rect 200205 301474 200271 301477
rect 201401 301474 201467 301477
rect 197188 301472 201467 301474
rect 197188 301416 200210 301472
rect 200266 301416 201406 301472
rect 201462 301416 201467 301472
rect 197188 301414 201467 301416
rect 197188 301412 197194 301414
rect 200205 301411 200271 301414
rect 201401 301411 201467 301414
rect 218237 301066 218303 301069
rect 218697 301066 218763 301069
rect 263685 301066 263751 301069
rect 218237 301064 263751 301066
rect 218237 301008 218242 301064
rect 218298 301008 218702 301064
rect 218758 301008 263690 301064
rect 263746 301008 263751 301064
rect 218237 301006 263751 301008
rect 218237 301003 218303 301006
rect 218697 301003 218763 301006
rect 263685 301003 263751 301006
rect 244222 300930 244228 300932
rect 66713 300928 68908 300930
rect 66713 300872 66718 300928
rect 66774 300872 68908 300928
rect 66713 300870 68908 300872
rect 156646 300870 244228 300930
rect 66713 300867 66779 300870
rect 244222 300868 244228 300870
rect 244292 300868 244298 300932
rect 200849 300794 200915 300797
rect 202873 300794 202939 300797
rect 200849 300792 202939 300794
rect 200849 300736 200854 300792
rect 200910 300736 202878 300792
rect 202934 300736 202939 300792
rect 200849 300734 202939 300736
rect 200849 300731 200915 300734
rect 202873 300731 202939 300734
rect 219709 300794 219775 300797
rect 220169 300794 220235 300797
rect 219709 300792 220235 300794
rect 219709 300736 219714 300792
rect 219770 300736 220174 300792
rect 220230 300736 220235 300792
rect 219709 300734 220235 300736
rect 219709 300731 219775 300734
rect 220169 300731 220235 300734
rect 156646 300114 156706 300356
rect 158897 300114 158963 300117
rect 218697 300114 218763 300117
rect 156646 300112 218763 300114
rect 156646 300056 158902 300112
rect 158958 300056 218702 300112
rect 218758 300056 218763 300112
rect 156646 300054 218763 300056
rect 158897 300051 158963 300054
rect 218697 300051 218763 300054
rect 67541 299842 67607 299845
rect 67541 299840 68908 299842
rect 67541 299784 67546 299840
rect 67602 299784 68908 299840
rect 67541 299782 68908 299784
rect 67541 299779 67607 299782
rect 219709 299706 219775 299709
rect 283189 299706 283255 299709
rect 219709 299704 283255 299706
rect 219709 299648 219714 299704
rect 219770 299648 283194 299704
rect 283250 299648 283255 299704
rect 219709 299646 283255 299648
rect 219709 299643 219775 299646
rect 283189 299643 283255 299646
rect 225689 299570 225755 299573
rect 227437 299570 227503 299573
rect 302877 299570 302943 299573
rect 225689 299568 302943 299570
rect 225689 299512 225694 299568
rect 225750 299512 227442 299568
rect 227498 299512 302882 299568
rect 302938 299512 302943 299568
rect 225689 299510 302943 299512
rect 225689 299507 225755 299510
rect 227437 299507 227503 299510
rect 302877 299507 302943 299510
rect 200757 299434 200823 299437
rect 204437 299434 204503 299437
rect 204989 299434 205055 299437
rect 200757 299432 205055 299434
rect 200757 299376 200762 299432
rect 200818 299376 204442 299432
rect 204498 299376 204994 299432
rect 205050 299376 205055 299432
rect 200757 299374 205055 299376
rect 200757 299371 200823 299374
rect 204437 299371 204503 299374
rect 204989 299371 205055 299374
rect 159909 299298 159975 299301
rect 156676 299296 159975 299298
rect 156676 299240 159914 299296
rect 159970 299240 159975 299296
rect 156676 299238 159975 299240
rect 159909 299235 159975 299238
rect 66897 298754 66963 298757
rect 166349 298754 166415 298757
rect 225965 298754 226031 298757
rect 66897 298752 68908 298754
rect 66897 298696 66902 298752
rect 66958 298696 68908 298752
rect 66897 298694 68908 298696
rect 166349 298752 226031 298754
rect 166349 298696 166354 298752
rect 166410 298696 225970 298752
rect 226026 298696 226031 298752
rect 166349 298694 226031 298696
rect 66897 298691 66963 298694
rect 166349 298691 166415 298694
rect 225965 298691 226031 298694
rect 226190 298692 226196 298756
rect 226260 298754 226266 298756
rect 291193 298754 291259 298757
rect 226260 298752 291259 298754
rect 226260 298696 291198 298752
rect 291254 298696 291259 298752
rect 226260 298694 291259 298696
rect 226260 298692 226266 298694
rect 291193 298691 291259 298694
rect 582741 298754 582807 298757
rect 583520 298754 584960 298844
rect 582741 298752 584960 298754
rect 582741 298696 582746 298752
rect 582802 298696 584960 298752
rect 582741 298694 584960 298696
rect 582741 298691 582807 298694
rect 583520 298604 584960 298694
rect 159030 298210 159036 298212
rect 156676 298150 159036 298210
rect 159030 298148 159036 298150
rect 159100 298148 159106 298212
rect 209129 298210 209195 298213
rect 209405 298210 209471 298213
rect 255957 298210 256023 298213
rect 209129 298208 256023 298210
rect 209129 298152 209134 298208
rect 209190 298152 209410 298208
rect 209466 298152 255962 298208
rect 256018 298152 256023 298208
rect 209129 298150 256023 298152
rect 209129 298147 209195 298150
rect 209405 298147 209471 298150
rect 255957 298147 256023 298150
rect 66897 297666 66963 297669
rect 66897 297664 68908 297666
rect 66897 297608 66902 297664
rect 66958 297608 68908 297664
rect 66897 297606 68908 297608
rect 66897 297603 66963 297606
rect 202638 297468 202644 297532
rect 202708 297530 202714 297532
rect 209773 297530 209839 297533
rect 202708 297528 209839 297530
rect 202708 297472 209778 297528
rect 209834 297472 209839 297528
rect 202708 297470 209839 297472
rect 202708 297468 202714 297470
rect 209773 297467 209839 297470
rect 208158 297332 208164 297396
rect 208228 297394 208234 297396
rect 226333 297394 226399 297397
rect 208228 297392 226399 297394
rect 208228 297336 226338 297392
rect 226394 297336 226399 297392
rect 208228 297334 226399 297336
rect 208228 297332 208234 297334
rect 226333 297331 226399 297334
rect 158713 297122 158779 297125
rect 156676 297120 158779 297122
rect 156676 297064 158718 297120
rect 158774 297064 158779 297120
rect 156676 297062 158779 297064
rect 158713 297059 158779 297062
rect 218053 297122 218119 297125
rect 249977 297122 250043 297125
rect 218053 297120 250043 297122
rect 218053 297064 218058 297120
rect 218114 297064 249982 297120
rect 250038 297064 250043 297120
rect 218053 297062 250043 297064
rect 218053 297059 218119 297062
rect 249977 297059 250043 297062
rect 228909 296986 228975 296989
rect 275369 296986 275435 296989
rect 228909 296984 275435 296986
rect 228909 296928 228914 296984
rect 228970 296928 275374 296984
rect 275430 296928 275435 296984
rect 228909 296926 275435 296928
rect 228909 296923 228975 296926
rect 275369 296923 275435 296926
rect 160829 296850 160895 296853
rect 232589 296850 232655 296853
rect 160829 296848 232655 296850
rect 160829 296792 160834 296848
rect 160890 296792 232594 296848
rect 232650 296792 232655 296848
rect 160829 296790 232655 296792
rect 160829 296787 160895 296790
rect 232589 296787 232655 296790
rect 67173 296306 67239 296309
rect 67950 296306 67956 296308
rect 67173 296304 67956 296306
rect 67173 296248 67178 296304
rect 67234 296248 67956 296304
rect 67173 296246 67956 296248
rect 67173 296243 67239 296246
rect 67950 296244 67956 296246
rect 68020 296306 68026 296308
rect 68878 296306 68938 296548
rect 68020 296246 68938 296306
rect 68020 296244 68026 296246
rect 159909 296170 159975 296173
rect 159909 296168 161490 296170
rect 159909 296112 159914 296168
rect 159970 296112 161490 296168
rect 159909 296110 161490 296112
rect 159909 296107 159975 296110
rect 160001 296034 160067 296037
rect 156676 296032 160067 296034
rect 156676 295976 160006 296032
rect 160062 295976 160067 296032
rect 156676 295974 160067 295976
rect 161430 296034 161490 296110
rect 219198 296108 219204 296172
rect 219268 296170 219274 296172
rect 266353 296170 266419 296173
rect 219268 296168 266419 296170
rect 219268 296112 266358 296168
rect 266414 296112 266419 296168
rect 219268 296110 266419 296112
rect 219268 296108 219274 296110
rect 266353 296107 266419 296110
rect 242934 296034 242940 296036
rect 161430 295974 242940 296034
rect 160001 295971 160067 295974
rect 242934 295972 242940 295974
rect 243004 295972 243010 296036
rect 66897 295490 66963 295493
rect 66897 295488 68908 295490
rect 66897 295432 66902 295488
rect 66958 295432 68908 295488
rect 66897 295430 68908 295432
rect 66897 295427 66963 295430
rect 159950 295292 159956 295356
rect 160020 295354 160026 295356
rect 223021 295354 223087 295357
rect 160020 295352 223087 295354
rect 160020 295296 223026 295352
rect 223082 295296 223087 295352
rect 160020 295294 223087 295296
rect 160020 295292 160026 295294
rect 223021 295291 223087 295294
rect 242157 295354 242223 295357
rect 267774 295354 267780 295356
rect 242157 295352 267780 295354
rect 242157 295296 242162 295352
rect 242218 295296 267780 295352
rect 242157 295294 267780 295296
rect 242157 295291 242223 295294
rect 267774 295292 267780 295294
rect 267844 295292 267850 295356
rect 218697 295218 218763 295221
rect 228357 295218 228423 295221
rect 218697 295216 228423 295218
rect 218697 295160 218702 295216
rect 218758 295160 228362 295216
rect 228418 295160 228423 295216
rect 218697 295158 228423 295160
rect 218697 295155 218763 295158
rect 228357 295155 228423 295158
rect 178033 295082 178099 295085
rect 218053 295082 218119 295085
rect 178033 295080 218119 295082
rect 178033 295024 178038 295080
rect 178094 295024 218058 295080
rect 218114 295024 218119 295080
rect 178033 295022 218119 295024
rect 178033 295019 178099 295022
rect 218053 295019 218119 295022
rect 158713 294946 158779 294949
rect 156676 294944 158779 294946
rect 156676 294888 158718 294944
rect 158774 294888 158779 294944
rect 156676 294886 158779 294888
rect 158713 294883 158779 294886
rect 170581 294538 170647 294541
rect 177430 294538 177436 294540
rect 170581 294536 177436 294538
rect 170581 294480 170586 294536
rect 170642 294480 177436 294536
rect 170581 294478 177436 294480
rect 170581 294475 170647 294478
rect 177430 294476 177436 294478
rect 177500 294476 177506 294540
rect 201585 294538 201651 294541
rect 295333 294538 295399 294541
rect 201585 294536 295399 294538
rect 201585 294480 201590 294536
rect 201646 294480 295338 294536
rect 295394 294480 295399 294536
rect 201585 294478 295399 294480
rect 201585 294475 201651 294478
rect 295333 294475 295399 294478
rect 66253 294402 66319 294405
rect 66253 294400 68908 294402
rect 66253 294344 66258 294400
rect 66314 294344 68908 294400
rect 66253 294342 68908 294344
rect 66253 294339 66319 294342
rect 185669 293994 185735 293997
rect 241421 293994 241487 293997
rect 185669 293992 241487 293994
rect 185669 293936 185674 293992
rect 185730 293936 241426 293992
rect 241482 293936 241487 293992
rect 185669 293934 241487 293936
rect 185669 293931 185735 293934
rect 241421 293931 241487 293934
rect 242801 293994 242867 293997
rect 389173 293994 389239 293997
rect 242801 293992 389239 293994
rect 242801 293936 242806 293992
rect 242862 293936 389178 293992
rect 389234 293936 389239 293992
rect 242801 293934 389239 293936
rect 242801 293931 242867 293934
rect 389173 293931 389239 293934
rect 158805 293858 158871 293861
rect 156676 293856 158871 293858
rect 156676 293800 158810 293856
rect 158866 293800 158871 293856
rect 156676 293798 158871 293800
rect 158805 293795 158871 293798
rect 66897 293314 66963 293317
rect 199929 293314 199995 293317
rect 231117 293314 231183 293317
rect 66897 293312 68908 293314
rect -960 293178 480 293268
rect 66897 293256 66902 293312
rect 66958 293256 68908 293312
rect 66897 293254 68908 293256
rect 199929 293312 231183 293314
rect 199929 293256 199934 293312
rect 199990 293256 231122 293312
rect 231178 293256 231183 293312
rect 199929 293254 231183 293256
rect 66897 293251 66963 293254
rect 199929 293251 199995 293254
rect 231117 293251 231183 293254
rect 3509 293178 3575 293181
rect -960 293176 3575 293178
rect -960 293120 3514 293176
rect 3570 293120 3575 293176
rect -960 293118 3575 293120
rect -960 293028 480 293118
rect 3509 293115 3575 293118
rect 217542 293116 217548 293180
rect 217612 293178 217618 293180
rect 262213 293178 262279 293181
rect 217612 293176 262279 293178
rect 217612 293120 262218 293176
rect 262274 293120 262279 293176
rect 217612 293118 262279 293120
rect 217612 293116 217618 293118
rect 262213 293115 262279 293118
rect 158713 293042 158779 293045
rect 156676 293040 158779 293042
rect 156676 292984 158718 293040
rect 158774 292984 158779 293040
rect 156676 292982 158779 292984
rect 158713 292979 158779 292982
rect 191189 292634 191255 292637
rect 193857 292634 193923 292637
rect 191189 292632 193923 292634
rect 191189 292576 191194 292632
rect 191250 292576 193862 292632
rect 193918 292576 193923 292632
rect 191189 292574 193923 292576
rect 191189 292571 191255 292574
rect 193857 292571 193923 292574
rect 220721 292634 220787 292637
rect 239949 292634 240015 292637
rect 314653 292634 314719 292637
rect 315113 292634 315179 292637
rect 220721 292632 315179 292634
rect 220721 292576 220726 292632
rect 220782 292576 239954 292632
rect 240010 292576 314658 292632
rect 314714 292576 315118 292632
rect 315174 292576 315179 292632
rect 220721 292574 315179 292576
rect 220721 292571 220787 292574
rect 239949 292571 240015 292574
rect 314653 292571 314719 292574
rect 315113 292571 315179 292574
rect 66897 292226 66963 292229
rect 66897 292224 68908 292226
rect 66897 292168 66902 292224
rect 66958 292168 68908 292224
rect 66897 292166 68908 292168
rect 66897 292163 66963 292166
rect 219934 292028 219940 292092
rect 220004 292090 220010 292092
rect 230381 292090 230447 292093
rect 220004 292088 230447 292090
rect 220004 292032 230386 292088
rect 230442 292032 230447 292088
rect 220004 292030 230447 292032
rect 220004 292028 220010 292030
rect 230381 292027 230447 292030
rect 158713 291954 158779 291957
rect 156676 291952 158779 291954
rect 156676 291896 158718 291952
rect 158774 291896 158779 291952
rect 156676 291894 158779 291896
rect 158713 291891 158779 291894
rect 201677 291954 201743 291957
rect 202873 291954 202939 291957
rect 282177 291954 282243 291957
rect 201677 291952 282243 291954
rect 201677 291896 201682 291952
rect 201738 291896 202878 291952
rect 202934 291896 282182 291952
rect 282238 291896 282243 291952
rect 201677 291894 282243 291896
rect 201677 291891 201743 291894
rect 202873 291891 202939 291894
rect 282177 291891 282243 291894
rect 158069 291818 158135 291821
rect 255405 291818 255471 291821
rect 256141 291818 256207 291821
rect 158069 291816 256207 291818
rect 158069 291760 158074 291816
rect 158130 291760 255410 291816
rect 255466 291760 256146 291816
rect 256202 291760 256207 291816
rect 158069 291758 256207 291760
rect 158069 291755 158135 291758
rect 255405 291755 255471 291758
rect 256141 291755 256207 291758
rect 66897 291138 66963 291141
rect 203517 291138 203583 291141
rect 204161 291138 204227 291141
rect 66897 291136 68908 291138
rect 66897 291080 66902 291136
rect 66958 291080 68908 291136
rect 66897 291078 68908 291080
rect 203517 291136 204227 291138
rect 203517 291080 203522 291136
rect 203578 291080 204166 291136
rect 204222 291080 204227 291136
rect 203517 291078 204227 291080
rect 66897 291075 66963 291078
rect 203517 291075 203583 291078
rect 204161 291075 204227 291078
rect 303613 291138 303679 291141
rect 304257 291138 304323 291141
rect 303613 291136 304323 291138
rect 303613 291080 303618 291136
rect 303674 291080 304262 291136
rect 304318 291080 304323 291136
rect 303613 291078 304323 291080
rect 303613 291075 303679 291078
rect 304257 291075 304323 291078
rect 158713 290866 158779 290869
rect 156676 290864 158779 290866
rect 156676 290808 158718 290864
rect 158774 290808 158779 290864
rect 156676 290806 158779 290808
rect 158713 290803 158779 290806
rect 189809 290594 189875 290597
rect 220721 290594 220787 290597
rect 189809 290592 220787 290594
rect 189809 290536 189814 290592
rect 189870 290536 220726 290592
rect 220782 290536 220787 290592
rect 189809 290534 220787 290536
rect 189809 290531 189875 290534
rect 220721 290531 220787 290534
rect 211889 290458 211955 290461
rect 304257 290458 304323 290461
rect 211889 290456 304323 290458
rect 211889 290400 211894 290456
rect 211950 290400 304262 290456
rect 304318 290400 304323 290456
rect 211889 290398 304323 290400
rect 211889 290395 211955 290398
rect 304257 290395 304323 290398
rect 67357 290050 67423 290053
rect 67357 290048 68908 290050
rect 67357 289992 67362 290048
rect 67418 289992 68908 290048
rect 67357 289990 68908 289992
rect 67357 289987 67423 289990
rect 204161 289914 204227 289917
rect 211654 289914 211660 289916
rect 204161 289912 211660 289914
rect 204161 289856 204166 289912
rect 204222 289856 211660 289912
rect 204161 289854 211660 289856
rect 204161 289851 204227 289854
rect 211654 289852 211660 289854
rect 211724 289852 211730 289916
rect 221641 289914 221707 289917
rect 288525 289914 288591 289917
rect 221641 289912 288591 289914
rect 221641 289856 221646 289912
rect 221702 289856 288530 289912
rect 288586 289856 288591 289912
rect 221641 289854 288591 289856
rect 221641 289851 221707 289854
rect 288525 289851 288591 289854
rect 158805 289778 158871 289781
rect 156676 289776 158871 289778
rect 156676 289720 158810 289776
rect 158866 289720 158871 289776
rect 156676 289718 158871 289720
rect 158805 289715 158871 289718
rect 232497 289778 232563 289781
rect 236637 289778 236703 289781
rect 232497 289776 236703 289778
rect 232497 289720 232502 289776
rect 232558 289720 236642 289776
rect 236698 289720 236703 289776
rect 232497 289718 236703 289720
rect 232497 289715 232563 289718
rect 236637 289715 236703 289718
rect 240961 289778 241027 289781
rect 245745 289778 245811 289781
rect 240961 289776 245811 289778
rect 240961 289720 240966 289776
rect 241022 289720 245750 289776
rect 245806 289720 245811 289776
rect 240961 289718 245811 289720
rect 240961 289715 241027 289718
rect 245745 289715 245811 289718
rect 242801 289642 242867 289645
rect 243813 289642 243879 289645
rect 242801 289640 243879 289642
rect 242801 289584 242806 289640
rect 242862 289584 243818 289640
rect 243874 289584 243879 289640
rect 242801 289582 243879 289584
rect 242801 289579 242867 289582
rect 243813 289579 243879 289582
rect 218053 289370 218119 289373
rect 239213 289370 239279 289373
rect 218053 289368 239279 289370
rect 218053 289312 218058 289368
rect 218114 289312 239218 289368
rect 239274 289312 239279 289368
rect 218053 289310 239279 289312
rect 218053 289307 218119 289310
rect 239213 289307 239279 289310
rect 201493 289234 201559 289237
rect 242801 289234 242867 289237
rect 201493 289232 242867 289234
rect 201493 289176 201498 289232
rect 201554 289176 242806 289232
rect 242862 289176 242867 289232
rect 201493 289174 242867 289176
rect 201493 289171 201559 289174
rect 242801 289171 242867 289174
rect 235993 289098 236059 289101
rect 278773 289098 278839 289101
rect 235993 289096 278839 289098
rect 235993 289040 235998 289096
rect 236054 289040 278778 289096
rect 278834 289040 278839 289096
rect 235993 289038 278839 289040
rect 235993 289035 236059 289038
rect 278773 289035 278839 289038
rect 66621 288962 66687 288965
rect 66621 288960 68908 288962
rect 66621 288904 66626 288960
rect 66682 288904 68908 288960
rect 66621 288902 68908 288904
rect 66621 288899 66687 288902
rect 159265 288692 159331 288693
rect 159214 288690 159220 288692
rect 156676 288630 159220 288690
rect 159284 288688 159331 288692
rect 159326 288632 159331 288688
rect 159214 288628 159220 288630
rect 159284 288628 159331 288632
rect 159265 288627 159331 288628
rect 162945 288554 163011 288557
rect 222837 288554 222903 288557
rect 162945 288552 222903 288554
rect 162945 288496 162950 288552
rect 163006 288496 222842 288552
rect 222898 288496 222903 288552
rect 162945 288494 222903 288496
rect 162945 288491 163011 288494
rect 222837 288491 222903 288494
rect 245745 288554 245811 288557
rect 291285 288554 291351 288557
rect 245745 288552 291351 288554
rect 245745 288496 245750 288552
rect 245806 288496 291290 288552
rect 291346 288496 291351 288552
rect 245745 288494 291351 288496
rect 245745 288491 245811 288494
rect 291285 288491 291351 288494
rect 242893 288418 242959 288421
rect 243537 288418 243603 288421
rect 242893 288416 243603 288418
rect 242893 288360 242898 288416
rect 242954 288360 243542 288416
rect 243598 288360 243603 288416
rect 242893 288358 243603 288360
rect 242893 288355 242959 288358
rect 243537 288355 243603 288358
rect 204713 288146 204779 288149
rect 211797 288146 211863 288149
rect 204713 288144 211863 288146
rect 204713 288088 204718 288144
rect 204774 288088 211802 288144
rect 211858 288088 211863 288144
rect 204713 288086 211863 288088
rect 204713 288083 204779 288086
rect 211797 288083 211863 288086
rect 66662 287812 66668 287876
rect 66732 287874 66738 287876
rect 184381 287874 184447 287877
rect 193949 287874 194015 287877
rect 66732 287844 69460 287874
rect 184381 287872 194015 287874
rect 66732 287814 69490 287844
rect 66732 287812 66738 287814
rect 69430 287740 69490 287814
rect 184381 287816 184386 287872
rect 184442 287816 193954 287872
rect 194010 287816 194015 287872
rect 184381 287814 194015 287816
rect 184381 287811 184447 287814
rect 193949 287811 194015 287814
rect 232589 287874 232655 287877
rect 247309 287874 247375 287877
rect 232589 287872 247375 287874
rect 232589 287816 232594 287872
rect 232650 287816 247314 287872
rect 247370 287816 247375 287872
rect 232589 287814 247375 287816
rect 232589 287811 232655 287814
rect 247309 287811 247375 287814
rect 69422 287676 69428 287740
rect 69492 287676 69498 287740
rect 158069 287738 158135 287741
rect 216673 287738 216739 287741
rect 238518 287738 238524 287740
rect 158069 287736 180810 287738
rect 158069 287680 158074 287736
rect 158130 287680 180810 287736
rect 158069 287678 180810 287680
rect 158069 287675 158135 287678
rect 158713 287602 158779 287605
rect 156676 287600 158779 287602
rect 156676 287544 158718 287600
rect 158774 287544 158779 287600
rect 156676 287542 158779 287544
rect 158713 287539 158779 287542
rect 180750 287330 180810 287678
rect 216673 287736 238524 287738
rect 216673 287680 216678 287736
rect 216734 287680 238524 287736
rect 216673 287678 238524 287680
rect 216673 287675 216739 287678
rect 238518 287676 238524 287678
rect 238588 287676 238594 287740
rect 239213 287738 239279 287741
rect 278129 287738 278195 287741
rect 239213 287736 278195 287738
rect 239213 287680 239218 287736
rect 239274 287680 278134 287736
rect 278190 287680 278195 287736
rect 239213 287678 278195 287680
rect 239213 287675 239279 287678
rect 278129 287675 278195 287678
rect 194225 287466 194291 287469
rect 194225 287464 209790 287466
rect 194225 287408 194230 287464
rect 194286 287408 209790 287464
rect 194225 287406 209790 287408
rect 194225 287403 194291 287406
rect 197169 287330 197235 287333
rect 202229 287330 202295 287333
rect 180750 287328 202295 287330
rect 180750 287272 197174 287328
rect 197230 287272 202234 287328
rect 202290 287272 202295 287328
rect 180750 287270 202295 287272
rect 209730 287330 209790 287406
rect 217685 287330 217751 287333
rect 209730 287328 217751 287330
rect 209730 287272 217690 287328
rect 217746 287272 217751 287328
rect 209730 287270 217751 287272
rect 197169 287267 197235 287270
rect 202229 287267 202295 287270
rect 217685 287267 217751 287270
rect 237373 287330 237439 287333
rect 243997 287330 244063 287333
rect 237373 287328 244063 287330
rect 237373 287272 237378 287328
rect 237434 287272 244002 287328
rect 244058 287272 244063 287328
rect 237373 287270 244063 287272
rect 237373 287267 237439 287270
rect 243997 287267 244063 287270
rect 199285 287194 199351 287197
rect 204253 287194 204319 287197
rect 199285 287192 204319 287194
rect 199285 287136 199290 287192
rect 199346 287136 204258 287192
rect 204314 287136 204319 287192
rect 199285 287134 204319 287136
rect 199285 287131 199351 287134
rect 204253 287131 204319 287134
rect 229737 287194 229803 287197
rect 233182 287194 233188 287196
rect 229737 287192 233188 287194
rect 229737 287136 229742 287192
rect 229798 287136 233188 287192
rect 229737 287134 233188 287136
rect 229737 287131 229803 287134
rect 233182 287132 233188 287134
rect 233252 287132 233258 287196
rect 242893 287194 242959 287197
rect 442993 287194 443059 287197
rect 242893 287192 443059 287194
rect 242893 287136 242898 287192
rect 242954 287136 442998 287192
rect 443054 287136 443059 287192
rect 242893 287134 443059 287136
rect 242893 287131 242959 287134
rect 442993 287131 443059 287134
rect 66805 286786 66871 286789
rect 66805 286784 68908 286786
rect 66805 286728 66810 286784
rect 66866 286728 68908 286784
rect 66805 286726 68908 286728
rect 66805 286723 66871 286726
rect 158805 286514 158871 286517
rect 156676 286512 158871 286514
rect 156676 286456 158810 286512
rect 158866 286456 158871 286512
rect 156676 286454 158871 286456
rect 158805 286451 158871 286454
rect 191230 286316 191236 286380
rect 191300 286378 191306 286380
rect 200389 286378 200455 286381
rect 191300 286376 200455 286378
rect 191300 286320 200394 286376
rect 200450 286320 200455 286376
rect 191300 286318 200455 286320
rect 191300 286316 191306 286318
rect 200389 286315 200455 286318
rect 222837 286378 222903 286381
rect 234705 286378 234771 286381
rect 222837 286376 234771 286378
rect 222837 286320 222842 286376
rect 222898 286320 234710 286376
rect 234766 286320 234771 286376
rect 222837 286318 234771 286320
rect 222837 286315 222903 286318
rect 234705 286315 234771 286318
rect 273253 286378 273319 286381
rect 438894 286378 438900 286380
rect 273253 286376 438900 286378
rect 273253 286320 273258 286376
rect 273314 286320 438900 286376
rect 273253 286318 438900 286320
rect 273253 286315 273319 286318
rect 438894 286316 438900 286318
rect 438964 286316 438970 286380
rect 200246 285908 200252 285972
rect 200316 285970 200322 285972
rect 204713 285970 204779 285973
rect 200316 285968 204779 285970
rect 200316 285912 204718 285968
rect 204774 285912 204779 285968
rect 200316 285910 204779 285912
rect 200316 285908 200322 285910
rect 204713 285907 204779 285910
rect 225045 285970 225111 285973
rect 232446 285970 232452 285972
rect 225045 285968 232452 285970
rect 225045 285912 225050 285968
rect 225106 285912 232452 285968
rect 225045 285910 232452 285912
rect 225045 285907 225111 285910
rect 232446 285908 232452 285910
rect 232516 285908 232522 285972
rect 232773 285970 232839 285973
rect 259545 285970 259611 285973
rect 232773 285968 259611 285970
rect 232773 285912 232778 285968
rect 232834 285912 259550 285968
rect 259606 285912 259611 285968
rect 232773 285910 259611 285912
rect 232773 285907 232839 285910
rect 259545 285907 259611 285910
rect 173157 285834 173223 285837
rect 203701 285834 203767 285837
rect 173157 285832 203767 285834
rect 173157 285776 173162 285832
rect 173218 285776 203706 285832
rect 203762 285776 203767 285832
rect 173157 285774 203767 285776
rect 173157 285771 173223 285774
rect 203701 285771 203767 285774
rect 215937 285834 216003 285837
rect 218053 285834 218119 285837
rect 215937 285832 218119 285834
rect 215937 285776 215942 285832
rect 215998 285776 218058 285832
rect 218114 285776 218119 285832
rect 215937 285774 218119 285776
rect 215937 285771 216003 285774
rect 218053 285771 218119 285774
rect 220077 285834 220143 285837
rect 223614 285834 223620 285836
rect 220077 285832 223620 285834
rect 220077 285776 220082 285832
rect 220138 285776 223620 285832
rect 220077 285774 223620 285776
rect 220077 285771 220143 285774
rect 223614 285772 223620 285774
rect 223684 285772 223690 285836
rect 273989 285834 274055 285837
rect 229050 285832 274055 285834
rect 229050 285776 273994 285832
rect 274050 285776 274055 285832
rect 229050 285774 274055 285776
rect 66897 285698 66963 285701
rect 201125 285698 201191 285701
rect 205541 285698 205607 285701
rect 66897 285696 68908 285698
rect 66897 285640 66902 285696
rect 66958 285640 68908 285696
rect 66897 285638 68908 285640
rect 201125 285696 205607 285698
rect 201125 285640 201130 285696
rect 201186 285640 205546 285696
rect 205602 285640 205607 285696
rect 201125 285638 205607 285640
rect 66897 285635 66963 285638
rect 201125 285635 201191 285638
rect 205541 285635 205607 285638
rect 206829 285698 206895 285701
rect 207565 285698 207631 285701
rect 206829 285696 207631 285698
rect 206829 285640 206834 285696
rect 206890 285640 207570 285696
rect 207626 285640 207631 285696
rect 206829 285638 207631 285640
rect 206829 285635 206895 285638
rect 207565 285635 207631 285638
rect 211981 285698 212047 285701
rect 214005 285698 214071 285701
rect 211981 285696 214071 285698
rect 211981 285640 211986 285696
rect 212042 285640 214010 285696
rect 214066 285640 214071 285696
rect 211981 285638 214071 285640
rect 211981 285635 212047 285638
rect 214005 285635 214071 285638
rect 214741 285698 214807 285701
rect 216213 285698 216279 285701
rect 214741 285696 216279 285698
rect 214741 285640 214746 285696
rect 214802 285640 216218 285696
rect 216274 285640 216279 285696
rect 214741 285638 216279 285640
rect 214741 285635 214807 285638
rect 216213 285635 216279 285638
rect 221457 285698 221523 285701
rect 222326 285698 222332 285700
rect 221457 285696 222332 285698
rect 221457 285640 221462 285696
rect 221518 285640 222332 285696
rect 221457 285638 222332 285640
rect 221457 285635 221523 285638
rect 222326 285636 222332 285638
rect 222396 285636 222402 285700
rect 225597 285698 225663 285701
rect 226517 285698 226583 285701
rect 229050 285698 229110 285774
rect 273989 285771 274055 285774
rect 225597 285696 229110 285698
rect 225597 285640 225602 285696
rect 225658 285640 226522 285696
rect 226578 285640 229110 285696
rect 225597 285638 229110 285640
rect 236637 285698 236703 285701
rect 286174 285698 286180 285700
rect 236637 285696 286180 285698
rect 236637 285640 236642 285696
rect 236698 285640 286180 285696
rect 236637 285638 286180 285640
rect 225597 285635 225663 285638
rect 226517 285635 226583 285638
rect 236637 285635 236703 285638
rect 286174 285636 286180 285638
rect 286244 285636 286250 285700
rect 158713 285426 158779 285429
rect 156676 285424 158779 285426
rect 156676 285368 158718 285424
rect 158774 285368 158779 285424
rect 156676 285366 158779 285368
rect 158713 285363 158779 285366
rect 583520 285276 584960 285516
rect 214005 285018 214071 285021
rect 244089 285018 244155 285021
rect 214005 285016 244155 285018
rect 214005 284960 214010 285016
rect 214066 284960 244094 285016
rect 244150 284960 244155 285016
rect 214005 284958 244155 284960
rect 214005 284955 214071 284958
rect 244089 284955 244155 284958
rect 352557 285018 352623 285021
rect 425646 285018 425652 285020
rect 352557 285016 425652 285018
rect 352557 284960 352562 285016
rect 352618 284960 425652 285016
rect 352557 284958 425652 284960
rect 352557 284955 352623 284958
rect 425646 284956 425652 284958
rect 425716 284956 425722 285020
rect 191741 284882 191807 284885
rect 201493 284882 201559 284885
rect 191741 284880 201559 284882
rect 191741 284824 191746 284880
rect 191802 284824 201498 284880
rect 201554 284824 201559 284880
rect 191741 284822 201559 284824
rect 191741 284819 191807 284822
rect 201493 284819 201559 284822
rect 243997 284882 244063 284885
rect 367737 284882 367803 284885
rect 243997 284880 367803 284882
rect 243997 284824 244002 284880
rect 244058 284824 367742 284880
rect 367798 284824 367803 284880
rect 243997 284822 367803 284824
rect 243997 284819 244063 284822
rect 367737 284819 367803 284822
rect 66253 284610 66319 284613
rect 66253 284608 68908 284610
rect 66253 284552 66258 284608
rect 66314 284552 68908 284608
rect 66253 284550 68908 284552
rect 66253 284547 66319 284550
rect 199377 284474 199443 284477
rect 217317 284474 217383 284477
rect 199377 284472 217383 284474
rect 199377 284416 199382 284472
rect 199438 284416 217322 284472
rect 217378 284416 217383 284472
rect 199377 284414 217383 284416
rect 199377 284411 199443 284414
rect 217317 284411 217383 284414
rect 224309 284474 224375 284477
rect 227846 284474 227852 284476
rect 224309 284472 227852 284474
rect 224309 284416 224314 284472
rect 224370 284416 227852 284472
rect 224309 284414 227852 284416
rect 224309 284411 224375 284414
rect 227846 284412 227852 284414
rect 227916 284412 227922 284476
rect 238109 284474 238175 284477
rect 243486 284474 243492 284476
rect 238109 284472 243492 284474
rect 238109 284416 238114 284472
rect 238170 284416 243492 284472
rect 238109 284414 243492 284416
rect 238109 284411 238175 284414
rect 243486 284412 243492 284414
rect 243556 284412 243562 284476
rect 61878 284276 61884 284340
rect 61948 284338 61954 284340
rect 63401 284338 63467 284341
rect 158713 284338 158779 284341
rect 61948 284336 63467 284338
rect 61948 284280 63406 284336
rect 63462 284280 63467 284336
rect 61948 284278 63467 284280
rect 156676 284336 158779 284338
rect 156676 284280 158718 284336
rect 158774 284280 158779 284336
rect 156676 284278 158779 284280
rect 61948 284276 61954 284278
rect 63401 284275 63467 284278
rect 158713 284275 158779 284278
rect 170397 284338 170463 284341
rect 243997 284338 244063 284341
rect 170397 284336 244063 284338
rect 170397 284280 170402 284336
rect 170458 284280 244002 284336
rect 244058 284280 244063 284336
rect 170397 284278 244063 284280
rect 170397 284275 170463 284278
rect 243997 284275 244063 284278
rect 244089 284066 244155 284069
rect 271137 284066 271203 284069
rect 244089 284064 271203 284066
rect 244089 284008 244094 284064
rect 244150 284008 271142 284064
rect 271198 284008 271203 284064
rect 244089 284006 271203 284008
rect 244089 284003 244155 284006
rect 271137 284003 271203 284006
rect 214465 283932 214531 283933
rect 214414 283930 214420 283932
rect 214374 283870 214420 283930
rect 214484 283928 214531 283932
rect 214526 283872 214531 283928
rect 214414 283868 214420 283870
rect 214484 283868 214531 283872
rect 214465 283867 214531 283868
rect 216397 283932 216463 283933
rect 216397 283928 216444 283932
rect 216508 283930 216514 283932
rect 216397 283872 216402 283928
rect 216397 283868 216444 283872
rect 216508 283870 216554 283930
rect 216508 283868 216514 283870
rect 218646 283868 218652 283932
rect 218716 283930 218722 283932
rect 218789 283930 218855 283933
rect 218716 283928 218855 283930
rect 218716 283872 218794 283928
rect 218850 283872 218855 283928
rect 218716 283870 218855 283872
rect 218716 283868 218722 283870
rect 216397 283867 216463 283868
rect 218789 283867 218855 283870
rect 223757 283930 223823 283933
rect 226926 283930 226932 283932
rect 223757 283928 226932 283930
rect 223757 283872 223762 283928
rect 223818 283872 226932 283928
rect 223757 283870 226932 283872
rect 223757 283867 223823 283870
rect 226926 283868 226932 283870
rect 226996 283868 227002 283932
rect 227662 283868 227668 283932
rect 227732 283930 227738 283932
rect 227989 283930 228055 283933
rect 228214 283930 228220 283932
rect 227732 283928 228220 283930
rect 227732 283872 227994 283928
rect 228050 283872 228220 283928
rect 227732 283870 228220 283872
rect 227732 283868 227738 283870
rect 227989 283867 228055 283870
rect 228214 283868 228220 283870
rect 228284 283868 228290 283932
rect 229461 283930 229527 283933
rect 229686 283930 229692 283932
rect 229461 283928 229692 283930
rect 229461 283872 229466 283928
rect 229522 283872 229692 283928
rect 229461 283870 229692 283872
rect 229461 283867 229527 283870
rect 229686 283868 229692 283870
rect 229756 283868 229762 283932
rect 231485 283930 231551 283933
rect 231710 283930 231716 283932
rect 231485 283928 231716 283930
rect 231485 283872 231490 283928
rect 231546 283872 231716 283928
rect 231485 283870 231716 283872
rect 231485 283867 231551 283870
rect 231710 283868 231716 283870
rect 231780 283868 231786 283932
rect 236361 283930 236427 283933
rect 236494 283930 236500 283932
rect 236361 283928 236500 283930
rect 236361 283872 236366 283928
rect 236422 283872 236500 283928
rect 236361 283870 236500 283872
rect 236361 283867 236427 283870
rect 236494 283868 236500 283870
rect 236564 283930 236570 283932
rect 236729 283930 236795 283933
rect 236564 283928 236795 283930
rect 236564 283872 236734 283928
rect 236790 283872 236795 283928
rect 236564 283870 236795 283872
rect 236564 283868 236570 283870
rect 236729 283867 236795 283870
rect 246941 283794 247007 283797
rect 244076 283792 247007 283794
rect 67541 283522 67607 283525
rect 67541 283520 68908 283522
rect 67541 283464 67546 283520
rect 67602 283464 68908 283520
rect 67541 283462 68908 283464
rect 67541 283459 67607 283462
rect 159449 283250 159515 283253
rect 156676 283248 159515 283250
rect 156676 283192 159454 283248
rect 159510 283192 159515 283248
rect 156676 283190 159515 283192
rect 159449 283187 159515 283190
rect 186814 283188 186820 283252
rect 186884 283250 186890 283252
rect 200254 283250 200314 283764
rect 244076 283736 246946 283792
rect 247002 283736 247007 283792
rect 244076 283734 247007 283736
rect 246941 283731 247007 283734
rect 246849 283250 246915 283253
rect 186884 283190 200314 283250
rect 244076 283248 246915 283250
rect 244076 283192 246854 283248
rect 246910 283192 246915 283248
rect 244076 283190 246915 283192
rect 186884 283188 186890 283190
rect 246849 283187 246915 283190
rect 187601 283114 187667 283117
rect 187601 283112 200130 283114
rect 187601 283056 187606 283112
rect 187662 283056 200130 283112
rect 187601 283054 200130 283056
rect 187601 283051 187667 283054
rect 198774 282916 198780 282980
rect 198844 282978 198850 282980
rect 199285 282978 199351 282981
rect 198844 282976 199351 282978
rect 198844 282920 199290 282976
rect 199346 282920 199351 282976
rect 198844 282918 199351 282920
rect 200070 282978 200130 283054
rect 200070 282918 200284 282978
rect 198844 282916 198850 282918
rect 199285 282915 199351 282918
rect 66805 282434 66871 282437
rect 197353 282434 197419 282437
rect 244365 282434 244431 282437
rect 66805 282432 68908 282434
rect 66805 282376 66810 282432
rect 66866 282376 68908 282432
rect 66805 282374 68908 282376
rect 197353 282432 200284 282434
rect 197353 282376 197358 282432
rect 197414 282376 200284 282432
rect 197353 282374 200284 282376
rect 244076 282432 244431 282434
rect 244076 282376 244370 282432
rect 244426 282376 244431 282432
rect 244076 282374 244431 282376
rect 66805 282371 66871 282374
rect 197353 282371 197419 282374
rect 244365 282371 244431 282374
rect 158713 282162 158779 282165
rect 156676 282160 158779 282162
rect 156676 282104 158718 282160
rect 158774 282104 158779 282160
rect 156676 282102 158779 282104
rect 158713 282099 158779 282102
rect 199929 281618 199995 281621
rect 245929 281618 245995 281621
rect 199929 281616 200284 281618
rect 199929 281560 199934 281616
rect 199990 281560 200284 281616
rect 199929 281558 200284 281560
rect 244076 281616 245995 281618
rect 244076 281560 245934 281616
rect 245990 281560 245995 281616
rect 244076 281558 245995 281560
rect 199929 281555 199995 281558
rect 245929 281555 245995 281558
rect 186814 281420 186820 281484
rect 186884 281482 186890 281484
rect 187509 281482 187575 281485
rect 186884 281480 187575 281482
rect 186884 281424 187514 281480
rect 187570 281424 187575 281480
rect 186884 281422 187575 281424
rect 186884 281420 186890 281422
rect 187509 281419 187575 281422
rect 67449 281346 67515 281349
rect 67449 281344 68908 281346
rect 67449 281288 67454 281344
rect 67510 281288 68908 281344
rect 67449 281286 68908 281288
rect 67449 281283 67515 281286
rect 158713 281074 158779 281077
rect 245929 281074 245995 281077
rect 156676 281072 158779 281074
rect 156676 281016 158718 281072
rect 158774 281016 158779 281072
rect 156676 281014 158779 281016
rect 244076 281072 245995 281074
rect 244076 281016 245934 281072
rect 245990 281016 245995 281072
rect 244076 281014 245995 281016
rect 158713 281011 158779 281014
rect 245929 281011 245995 281014
rect 169201 280530 169267 280533
rect 200254 280530 200314 280772
rect 243486 280740 243492 280804
rect 243556 280802 243562 280804
rect 277393 280802 277459 280805
rect 243556 280800 277459 280802
rect 243556 280744 277398 280800
rect 277454 280744 277459 280800
rect 243556 280742 277459 280744
rect 243556 280740 243562 280742
rect 277393 280739 277459 280742
rect 169201 280528 200314 280530
rect 169201 280472 169206 280528
rect 169262 280472 200314 280528
rect 169201 280470 200314 280472
rect 169201 280467 169267 280470
rect 67173 280258 67239 280261
rect 67766 280258 67772 280260
rect 67173 280256 67772 280258
rect -960 279972 480 280212
rect 67173 280200 67178 280256
rect 67234 280200 67772 280256
rect 67173 280198 67772 280200
rect 67173 280195 67239 280198
rect 67766 280196 67772 280198
rect 67836 280258 67842 280260
rect 197353 280258 197419 280261
rect 200021 280258 200087 280261
rect 280337 280260 280403 280261
rect 244774 280258 244780 280260
rect 67836 280198 68908 280258
rect 197353 280256 200284 280258
rect 197353 280200 197358 280256
rect 197414 280200 200026 280256
rect 200082 280200 200284 280256
rect 197353 280198 200284 280200
rect 244076 280198 244780 280258
rect 67836 280196 67842 280198
rect 197353 280195 197419 280198
rect 200021 280195 200087 280198
rect 244774 280196 244780 280198
rect 244844 280196 244850 280260
rect 280286 280258 280292 280260
rect 280246 280198 280292 280258
rect 280356 280256 280403 280260
rect 280398 280200 280403 280256
rect 280286 280196 280292 280198
rect 280356 280196 280403 280200
rect 280337 280195 280403 280196
rect 158713 279986 158779 279989
rect 156676 279984 158779 279986
rect 156676 279928 158718 279984
rect 158774 279928 158779 279984
rect 156676 279926 158779 279928
rect 158713 279923 158779 279926
rect 200062 279788 200068 279852
rect 200132 279788 200138 279852
rect 173249 279714 173315 279717
rect 200070 279714 200130 279788
rect 173249 279712 200130 279714
rect 173249 279656 173254 279712
rect 173310 279656 200130 279712
rect 173249 279654 200130 279656
rect 173249 279651 173315 279654
rect 197353 279442 197419 279445
rect 248638 279442 248644 279444
rect 197353 279440 200284 279442
rect 197353 279384 197358 279440
rect 197414 279384 200284 279440
rect 197353 279382 200284 279384
rect 244076 279382 248644 279442
rect 197353 279379 197419 279382
rect 248638 279380 248644 279382
rect 248708 279442 248714 279444
rect 249701 279442 249767 279445
rect 248708 279440 249767 279442
rect 248708 279384 249706 279440
rect 249762 279384 249767 279440
rect 248708 279382 249767 279384
rect 248708 279380 248714 279382
rect 249701 279379 249767 279382
rect 66805 279170 66871 279173
rect 66805 279168 68908 279170
rect 66805 279112 66810 279168
rect 66866 279112 68908 279168
rect 66805 279110 68908 279112
rect 66805 279107 66871 279110
rect 158713 278898 158779 278901
rect 245929 278898 245995 278901
rect 156676 278896 158779 278898
rect 156676 278840 158718 278896
rect 158774 278840 158779 278896
rect 156676 278838 158779 278840
rect 244076 278896 245995 278898
rect 244076 278840 245934 278896
rect 245990 278840 245995 278896
rect 244076 278838 245995 278840
rect 158713 278835 158779 278838
rect 245929 278835 245995 278838
rect 173198 278700 173204 278764
rect 173268 278762 173274 278764
rect 178861 278762 178927 278765
rect 173268 278760 178927 278762
rect 173268 278704 178866 278760
rect 178922 278704 178927 278760
rect 173268 278702 178927 278704
rect 173268 278700 173274 278702
rect 178861 278699 178927 278702
rect 197353 278626 197419 278629
rect 197353 278624 200284 278626
rect 197353 278568 197358 278624
rect 197414 278568 200284 278624
rect 197353 278566 200284 278568
rect 197353 278563 197419 278566
rect 66897 278082 66963 278085
rect 66897 278080 68908 278082
rect 66897 278024 66902 278080
rect 66958 278024 68908 278080
rect 66897 278022 68908 278024
rect 66897 278019 66963 278022
rect 158478 278020 158484 278084
rect 158548 278082 158554 278084
rect 180006 278082 180012 278084
rect 158548 278022 180012 278082
rect 158548 278020 158554 278022
rect 180006 278020 180012 278022
rect 180076 278020 180082 278084
rect 198365 278082 198431 278085
rect 244273 278082 244339 278085
rect 246297 278082 246363 278085
rect 198365 278080 200284 278082
rect 198365 278024 198370 278080
rect 198426 278024 200284 278080
rect 198365 278022 200284 278024
rect 244076 278080 246363 278082
rect 244076 278024 244278 278080
rect 244334 278024 246302 278080
rect 246358 278024 246363 278080
rect 244076 278022 246363 278024
rect 198365 278019 198431 278022
rect 244273 278019 244339 278022
rect 246297 278019 246363 278022
rect 158478 277810 158484 277812
rect 156676 277750 158484 277810
rect 158478 277748 158484 277750
rect 158548 277748 158554 277812
rect 245929 277538 245995 277541
rect 244076 277536 245995 277538
rect 244076 277480 245934 277536
rect 245990 277480 245995 277536
rect 244076 277478 245995 277480
rect 245929 277475 245995 277478
rect 66989 277266 67055 277269
rect 67950 277266 67956 277268
rect 66989 277264 67956 277266
rect 66989 277208 66994 277264
rect 67050 277208 67956 277264
rect 66989 277206 67956 277208
rect 66989 277203 67055 277206
rect 67950 277204 67956 277206
rect 68020 277266 68026 277268
rect 68020 277206 68908 277266
rect 68020 277204 68026 277206
rect 200254 276994 200314 277236
rect 180750 276934 200314 276994
rect 158713 276722 158779 276725
rect 156676 276720 158779 276722
rect 156676 276664 158718 276720
rect 158774 276664 158779 276720
rect 156676 276662 158779 276664
rect 158713 276659 158779 276662
rect 66345 276178 66411 276181
rect 166349 276178 166415 276181
rect 180750 276178 180810 276934
rect 197353 276722 197419 276725
rect 199929 276722 199995 276725
rect 245653 276722 245719 276725
rect 197353 276720 200284 276722
rect 197353 276664 197358 276720
rect 197414 276664 199934 276720
rect 199990 276664 200284 276720
rect 197353 276662 200284 276664
rect 244076 276720 245719 276722
rect 244076 276664 245658 276720
rect 245714 276664 245719 276720
rect 244076 276662 245719 276664
rect 197353 276659 197419 276662
rect 199929 276659 199995 276662
rect 245653 276659 245719 276662
rect 66345 276176 68908 276178
rect 66345 276120 66350 276176
rect 66406 276120 68908 276176
rect 66345 276118 68908 276120
rect 166349 276176 180810 276178
rect 166349 276120 166354 276176
rect 166410 276120 180810 276176
rect 166349 276118 180810 276120
rect 66345 276115 66411 276118
rect 166349 276115 166415 276118
rect 172513 275906 172579 275909
rect 197261 275906 197327 275909
rect 245929 275906 245995 275909
rect 172513 275904 200284 275906
rect 172513 275848 172518 275904
rect 172574 275848 197266 275904
rect 197322 275848 200284 275904
rect 172513 275846 200284 275848
rect 244076 275904 245995 275906
rect 244076 275848 245934 275904
rect 245990 275848 245995 275904
rect 244076 275846 245995 275848
rect 172513 275843 172579 275846
rect 197261 275843 197327 275846
rect 245929 275843 245995 275846
rect 158713 275634 158779 275637
rect 156676 275632 158779 275634
rect 156676 275576 158718 275632
rect 158774 275576 158779 275632
rect 156676 275574 158779 275576
rect 158713 275571 158779 275574
rect 245745 275362 245811 275365
rect 244076 275360 245811 275362
rect 244076 275304 245750 275360
rect 245806 275304 245811 275360
rect 244076 275302 245811 275304
rect 245745 275299 245811 275302
rect 160870 275164 160876 275228
rect 160940 275226 160946 275228
rect 171225 275226 171291 275229
rect 160940 275224 171291 275226
rect 160940 275168 171230 275224
rect 171286 275168 171291 275224
rect 160940 275166 171291 275168
rect 160940 275164 160946 275166
rect 171225 275163 171291 275166
rect 197353 275090 197419 275093
rect 197353 275088 200284 275090
rect 68878 274682 68938 275060
rect 197353 275032 197358 275088
rect 197414 275032 200284 275088
rect 197353 275030 200284 275032
rect 197353 275027 197419 275030
rect 66118 274622 68938 274682
rect 65977 274546 66043 274549
rect 66118 274546 66178 274622
rect 158713 274546 158779 274549
rect 65977 274544 66178 274546
rect 65977 274488 65982 274544
rect 66038 274488 66178 274544
rect 65977 274486 66178 274488
rect 156676 274544 158779 274546
rect 156676 274488 158718 274544
rect 158774 274488 158779 274544
rect 156676 274486 158779 274488
rect 65977 274483 66043 274486
rect 158713 274483 158779 274486
rect 197445 274546 197511 274549
rect 245653 274546 245719 274549
rect 197445 274544 200284 274546
rect 197445 274488 197450 274544
rect 197506 274488 200284 274544
rect 197445 274486 200284 274488
rect 244076 274544 245719 274546
rect 244076 274488 245658 274544
rect 245714 274488 245719 274544
rect 244076 274486 245719 274488
rect 197445 274483 197511 274486
rect 245653 274483 245719 274486
rect 66805 274002 66871 274005
rect 66805 274000 68908 274002
rect 66805 273944 66810 274000
rect 66866 273944 68908 274000
rect 66805 273942 68908 273944
rect 66805 273939 66871 273942
rect 65977 273730 66043 273733
rect 66110 273730 66116 273732
rect 65977 273728 66116 273730
rect 65977 273672 65982 273728
rect 66038 273672 66116 273728
rect 65977 273670 66116 273672
rect 65977 273667 66043 273670
rect 66110 273668 66116 273670
rect 66180 273668 66186 273732
rect 200021 273730 200087 273733
rect 245837 273730 245903 273733
rect 200021 273728 200284 273730
rect 200021 273672 200026 273728
rect 200082 273672 200284 273728
rect 200021 273670 200284 273672
rect 244076 273728 245903 273730
rect 244076 273672 245842 273728
rect 245898 273672 245903 273728
rect 244076 273670 245903 273672
rect 200021 273667 200087 273670
rect 245837 273667 245903 273670
rect 158805 273458 158871 273461
rect 156676 273456 158871 273458
rect 156676 273400 158810 273456
rect 158866 273400 158871 273456
rect 156676 273398 158871 273400
rect 158805 273395 158871 273398
rect 173433 273322 173499 273325
rect 178677 273322 178743 273325
rect 173433 273320 178743 273322
rect 173433 273264 173438 273320
rect 173494 273264 178682 273320
rect 178738 273264 178743 273320
rect 173433 273262 178743 273264
rect 173433 273259 173499 273262
rect 178677 273259 178743 273262
rect 184749 273322 184815 273325
rect 185761 273322 185827 273325
rect 184749 273320 185827 273322
rect 184749 273264 184754 273320
rect 184810 273264 185766 273320
rect 185822 273264 185827 273320
rect 184749 273262 185827 273264
rect 184749 273259 184815 273262
rect 185761 273259 185827 273262
rect 186221 273322 186287 273325
rect 188429 273322 188495 273325
rect 186221 273320 188495 273322
rect 186221 273264 186226 273320
rect 186282 273264 188434 273320
rect 188490 273264 188495 273320
rect 186221 273262 188495 273264
rect 186221 273259 186287 273262
rect 188429 273259 188495 273262
rect 195278 273260 195284 273324
rect 195348 273322 195354 273324
rect 198774 273322 198780 273324
rect 195348 273262 198780 273322
rect 195348 273260 195354 273262
rect 198774 273260 198780 273262
rect 198844 273260 198850 273324
rect 245745 273186 245811 273189
rect 244076 273184 245811 273186
rect 244076 273128 245750 273184
rect 245806 273128 245811 273184
rect 244076 273126 245811 273128
rect 245745 273123 245811 273126
rect 66713 272914 66779 272917
rect 197353 272914 197419 272917
rect 66713 272912 68908 272914
rect 66713 272856 66718 272912
rect 66774 272856 68908 272912
rect 66713 272854 68908 272856
rect 197353 272912 200284 272914
rect 197353 272856 197358 272912
rect 197414 272856 200284 272912
rect 197353 272854 200284 272856
rect 66713 272851 66779 272854
rect 197353 272851 197419 272854
rect 176561 272506 176627 272509
rect 185342 272506 185348 272508
rect 176561 272504 185348 272506
rect 176561 272448 176566 272504
rect 176622 272448 185348 272504
rect 176561 272446 185348 272448
rect 176561 272443 176627 272446
rect 185342 272444 185348 272446
rect 185412 272444 185418 272508
rect 194501 272370 194567 272373
rect 245929 272370 245995 272373
rect 194501 272368 200284 272370
rect 156646 271962 156706 272340
rect 194501 272312 194506 272368
rect 194562 272312 200284 272368
rect 194501 272310 200284 272312
rect 244076 272368 245995 272370
rect 244076 272312 245934 272368
rect 245990 272312 245995 272368
rect 244076 272310 245995 272312
rect 194501 272307 194567 272310
rect 245929 272307 245995 272310
rect 580165 272234 580231 272237
rect 583520 272234 584960 272324
rect 580165 272232 584960 272234
rect 580165 272176 580170 272232
rect 580226 272176 584960 272232
rect 580165 272174 584960 272176
rect 580165 272171 580231 272174
rect 583520 272084 584960 272174
rect 176561 271962 176627 271965
rect 156646 271960 176627 271962
rect 156646 271904 176566 271960
rect 176622 271904 176627 271960
rect 156646 271902 176627 271904
rect 176561 271899 176627 271902
rect 66805 271826 66871 271829
rect 159633 271826 159699 271829
rect 161974 271826 161980 271828
rect 66805 271824 68908 271826
rect 66805 271768 66810 271824
rect 66866 271768 68908 271824
rect 66805 271766 68908 271768
rect 159633 271824 161980 271826
rect 159633 271768 159638 271824
rect 159694 271768 161980 271824
rect 159633 271766 161980 271768
rect 66805 271763 66871 271766
rect 159633 271763 159699 271766
rect 161974 271764 161980 271766
rect 162044 271764 162050 271828
rect 197353 271554 197419 271557
rect 245929 271554 245995 271557
rect 197353 271552 200284 271554
rect 197353 271496 197358 271552
rect 197414 271496 200284 271552
rect 197353 271494 200284 271496
rect 244076 271552 245995 271554
rect 244076 271496 245934 271552
rect 245990 271496 245995 271552
rect 244076 271494 245995 271496
rect 197353 271491 197419 271494
rect 245929 271491 245995 271494
rect 158713 271282 158779 271285
rect 156676 271280 158779 271282
rect 156676 271224 158718 271280
rect 158774 271224 158779 271280
rect 156676 271222 158779 271224
rect 158713 271219 158779 271222
rect 198406 270948 198412 271012
rect 198476 271010 198482 271012
rect 244457 271010 244523 271013
rect 198476 270950 200284 271010
rect 244076 271008 244523 271010
rect 244076 270980 244462 271008
rect 244046 270952 244462 270980
rect 244518 270952 244523 271008
rect 244046 270950 244523 270952
rect 198476 270948 198482 270950
rect 67725 270738 67791 270741
rect 67725 270736 68908 270738
rect 67725 270680 67730 270736
rect 67786 270680 68908 270736
rect 67725 270678 68908 270680
rect 67725 270675 67791 270678
rect 244046 270602 244106 270950
rect 244457 270947 244523 270950
rect 282126 270602 282132 270604
rect 244046 270542 282132 270602
rect 282126 270540 282132 270542
rect 282196 270602 282202 270604
rect 282269 270602 282335 270605
rect 282196 270600 282335 270602
rect 282196 270544 282274 270600
rect 282330 270544 282335 270600
rect 282196 270542 282335 270544
rect 282196 270540 282202 270542
rect 282269 270539 282335 270542
rect 159633 270194 159699 270197
rect 156676 270192 159699 270194
rect 156676 270136 159638 270192
rect 159694 270136 159699 270192
rect 156676 270134 159699 270136
rect 159633 270131 159699 270134
rect 199837 270194 199903 270197
rect 244273 270194 244339 270197
rect 199837 270192 200284 270194
rect 199837 270136 199842 270192
rect 199898 270136 200284 270192
rect 199837 270134 200284 270136
rect 244076 270192 244339 270194
rect 244076 270136 244278 270192
rect 244334 270136 244339 270192
rect 244076 270134 244339 270136
rect 199837 270131 199903 270134
rect 244273 270131 244339 270134
rect 168097 269786 168163 269789
rect 177481 269786 177547 269789
rect 168097 269784 177547 269786
rect 168097 269728 168102 269784
rect 168158 269728 177486 269784
rect 177542 269728 177547 269784
rect 168097 269726 177547 269728
rect 168097 269723 168163 269726
rect 177481 269723 177547 269726
rect 264329 269786 264395 269789
rect 364333 269786 364399 269789
rect 264329 269784 364399 269786
rect 264329 269728 264334 269784
rect 264390 269728 364338 269784
rect 364394 269728 364399 269784
rect 264329 269726 364399 269728
rect 264329 269723 264395 269726
rect 364333 269723 364399 269726
rect 67633 269650 67699 269653
rect 245837 269650 245903 269653
rect 67633 269648 68908 269650
rect 67633 269592 67638 269648
rect 67694 269592 68908 269648
rect 67633 269590 68908 269592
rect 244076 269648 245903 269650
rect 244076 269592 245842 269648
rect 245898 269592 245903 269648
rect 244076 269590 245903 269592
rect 67633 269587 67699 269590
rect 245837 269587 245903 269590
rect 197353 269378 197419 269381
rect 197353 269376 200284 269378
rect 197353 269320 197358 269376
rect 197414 269320 200284 269376
rect 197353 269318 200284 269320
rect 197353 269315 197419 269318
rect 253197 269242 253263 269245
rect 245702 269240 253263 269242
rect 245702 269184 253202 269240
rect 253258 269184 253263 269240
rect 245702 269182 253263 269184
rect 158713 269106 158779 269109
rect 244222 269106 244228 269108
rect 156676 269104 158779 269106
rect 156676 269048 158718 269104
rect 158774 269048 158779 269104
rect 156676 269046 158779 269048
rect 158713 269043 158779 269046
rect 244046 269046 244228 269106
rect 197445 268834 197511 268837
rect 197445 268832 200284 268834
rect 197445 268776 197450 268832
rect 197506 268776 200284 268832
rect 244046 268804 244106 269046
rect 244222 269044 244228 269046
rect 244292 269106 244298 269108
rect 245702 269106 245762 269182
rect 253197 269179 253263 269182
rect 244292 269046 245762 269106
rect 244292 269044 244298 269046
rect 197445 268774 200284 268776
rect 197445 268771 197511 268774
rect 66805 268562 66871 268565
rect 66805 268560 68908 268562
rect 66805 268504 66810 268560
rect 66866 268504 68908 268560
rect 66805 268502 68908 268504
rect 66805 268499 66871 268502
rect 157926 268364 157932 268428
rect 157996 268426 158002 268428
rect 170581 268426 170647 268429
rect 157996 268424 170647 268426
rect 157996 268368 170586 268424
rect 170642 268368 170647 268424
rect 157996 268366 170647 268368
rect 157996 268364 158002 268366
rect 170581 268363 170647 268366
rect 158253 268018 158319 268021
rect 156676 268016 158319 268018
rect 156676 267960 158258 268016
rect 158314 267960 158319 268016
rect 156676 267958 158319 267960
rect 158253 267955 158319 267958
rect 197353 268018 197419 268021
rect 197353 268016 200284 268018
rect 197353 267960 197358 268016
rect 197414 267960 200284 268016
rect 197353 267958 200284 267960
rect 244076 267958 248430 268018
rect 197353 267955 197419 267958
rect 184289 267882 184355 267885
rect 191741 267882 191807 267885
rect 184289 267880 191807 267882
rect 184289 267824 184294 267880
rect 184350 267824 191746 267880
rect 191802 267824 191807 267880
rect 184289 267822 191807 267824
rect 248370 267882 248430 267958
rect 255313 267882 255379 267885
rect 248370 267880 255379 267882
rect 248370 267824 255318 267880
rect 255374 267824 255379 267880
rect 248370 267822 255379 267824
rect 184289 267819 184355 267822
rect 191741 267819 191807 267822
rect 255313 267819 255379 267822
rect 67398 267412 67404 267476
rect 67468 267474 67474 267476
rect 67468 267414 68908 267474
rect 67468 267412 67474 267414
rect -960 267202 480 267292
rect 3509 267202 3575 267205
rect -960 267200 3575 267202
rect -960 267144 3514 267200
rect 3570 267144 3575 267200
rect -960 267142 3575 267144
rect -960 267052 480 267142
rect 3509 267139 3575 267142
rect 195973 267202 196039 267205
rect 197118 267202 197124 267204
rect 195973 267200 197124 267202
rect 195973 267144 195978 267200
rect 196034 267144 197124 267200
rect 195973 267142 197124 267144
rect 195973 267139 196039 267142
rect 197118 267140 197124 267142
rect 197188 267202 197194 267204
rect 197188 267142 200284 267202
rect 197188 267140 197194 267142
rect 244046 266930 244106 267444
rect 67173 266386 67239 266389
rect 156646 266386 156706 266900
rect 244046 266870 248430 266930
rect 197353 266658 197419 266661
rect 245745 266658 245811 266661
rect 197353 266656 200284 266658
rect 197353 266600 197358 266656
rect 197414 266600 200284 266656
rect 197353 266598 200284 266600
rect 244076 266656 245811 266658
rect 244076 266600 245750 266656
rect 245806 266600 245811 266656
rect 244076 266598 245811 266600
rect 197353 266595 197419 266598
rect 245745 266595 245811 266598
rect 166441 266386 166507 266389
rect 166901 266386 166967 266389
rect 67173 266384 68908 266386
rect 67173 266328 67178 266384
rect 67234 266328 68908 266384
rect 67173 266326 68908 266328
rect 156646 266384 166967 266386
rect 156646 266328 166446 266384
rect 166502 266328 166906 266384
rect 166962 266328 166967 266384
rect 156646 266326 166967 266328
rect 248370 266386 248430 266870
rect 262305 266386 262371 266389
rect 303613 266386 303679 266389
rect 304441 266386 304507 266389
rect 248370 266384 304507 266386
rect 248370 266328 262310 266384
rect 262366 266328 303618 266384
rect 303674 266328 304446 266384
rect 304502 266328 304507 266384
rect 248370 266326 304507 266328
rect 67173 266323 67239 266326
rect 166441 266323 166507 266326
rect 166901 266323 166967 266326
rect 262305 266323 262371 266326
rect 303613 266323 303679 266326
rect 304441 266323 304507 266326
rect 255405 266250 255471 266253
rect 262765 266250 262831 266253
rect 255405 266248 262831 266250
rect 255405 266192 255410 266248
rect 255466 266192 262770 266248
rect 262826 266192 262831 266248
rect 255405 266190 262831 266192
rect 255405 266187 255471 266190
rect 262765 266187 262831 266190
rect 378777 266250 378843 266253
rect 583017 266250 583083 266253
rect 378777 266248 583083 266250
rect 378777 266192 378782 266248
rect 378838 266192 583022 266248
rect 583078 266192 583083 266248
rect 378777 266190 583083 266192
rect 378777 266187 378843 266190
rect 583017 266187 583083 266190
rect 158713 265842 158779 265845
rect 244406 265842 244412 265844
rect 156676 265840 158779 265842
rect 156676 265784 158718 265840
rect 158774 265784 158779 265840
rect 156676 265782 158779 265784
rect 158713 265779 158779 265782
rect 195145 265570 195211 265573
rect 200254 265570 200314 265812
rect 244076 265782 244412 265842
rect 244406 265780 244412 265782
rect 244476 265842 244482 265844
rect 245653 265842 245719 265845
rect 244476 265840 245719 265842
rect 244476 265784 245658 265840
rect 245714 265784 245719 265840
rect 244476 265782 245719 265784
rect 244476 265780 244482 265782
rect 245653 265779 245719 265782
rect 255405 265570 255471 265573
rect 195145 265568 200314 265570
rect 195145 265512 195150 265568
rect 195206 265512 200314 265568
rect 195145 265510 200314 265512
rect 244046 265568 255471 265570
rect 244046 265512 255410 265568
rect 255466 265512 255471 265568
rect 244046 265510 255471 265512
rect 195145 265507 195211 265510
rect 66897 265298 66963 265301
rect 66897 265296 68908 265298
rect 66897 265240 66902 265296
rect 66958 265240 68908 265296
rect 66897 265238 68908 265240
rect 200070 265238 200284 265298
rect 244046 265268 244106 265510
rect 255405 265507 255471 265510
rect 66897 265235 66963 265238
rect 184606 265100 184612 265164
rect 184676 265162 184682 265164
rect 200070 265162 200130 265238
rect 184676 265102 200130 265162
rect 184676 265100 184682 265102
rect 177849 265026 177915 265029
rect 195145 265026 195211 265029
rect 177849 265024 195211 265026
rect 177849 264968 177854 265024
rect 177910 264968 195150 265024
rect 195206 264968 195211 265024
rect 177849 264966 195211 264968
rect 177849 264963 177915 264966
rect 195145 264963 195211 264966
rect 197118 264964 197124 265028
rect 197188 265026 197194 265028
rect 199326 265026 199332 265028
rect 197188 264966 199332 265026
rect 197188 264964 197194 264966
rect 199326 264964 199332 264966
rect 199396 264964 199402 265028
rect 190453 264890 190519 264893
rect 156646 264888 190519 264890
rect 156646 264832 190458 264888
rect 190514 264832 190519 264888
rect 156646 264830 190519 264832
rect 156646 264724 156706 264830
rect 190453 264827 190519 264830
rect 197445 264482 197511 264485
rect 246021 264482 246087 264485
rect 197445 264480 200284 264482
rect 197445 264424 197450 264480
rect 197506 264424 200284 264480
rect 197445 264422 200284 264424
rect 244076 264480 246087 264482
rect 244076 264424 246026 264480
rect 246082 264424 246087 264480
rect 244076 264422 246087 264424
rect 197445 264419 197511 264422
rect 246021 264419 246087 264422
rect 66437 264210 66503 264213
rect 66437 264208 68908 264210
rect 66437 264152 66442 264208
rect 66498 264152 68908 264208
rect 66437 264150 68908 264152
rect 66437 264147 66503 264150
rect 245837 263938 245903 263941
rect 244076 263936 245903 263938
rect 244076 263880 245842 263936
rect 245898 263880 245903 263936
rect 244076 263878 245903 263880
rect 245837 263875 245903 263878
rect 186814 263666 186820 263668
rect 156676 263606 186820 263666
rect 186814 263604 186820 263606
rect 186884 263604 186890 263668
rect 197353 263666 197419 263669
rect 197353 263664 200284 263666
rect 197353 263608 197358 263664
rect 197414 263608 200284 263664
rect 197353 263606 200284 263608
rect 197353 263603 197419 263606
rect 66897 263122 66963 263125
rect 245694 263122 245700 263124
rect 66897 263120 68908 263122
rect 66897 263064 66902 263120
rect 66958 263064 68908 263120
rect 66897 263062 68908 263064
rect 66897 263059 66963 263062
rect 174537 262986 174603 262989
rect 180190 262986 180196 262988
rect 174537 262984 180196 262986
rect 174537 262928 174542 262984
rect 174598 262928 180196 262984
rect 174537 262926 180196 262928
rect 174537 262923 174603 262926
rect 180190 262924 180196 262926
rect 180260 262924 180266 262988
rect 191649 262986 191715 262989
rect 195094 262986 195100 262988
rect 191649 262984 195100 262986
rect 191649 262928 191654 262984
rect 191710 262928 195100 262984
rect 191649 262926 195100 262928
rect 191649 262923 191715 262926
rect 195094 262924 195100 262926
rect 195164 262924 195170 262988
rect 156822 262788 156828 262852
rect 156892 262850 156898 262852
rect 198549 262850 198615 262853
rect 200254 262850 200314 263092
rect 244076 263062 245700 263122
rect 245694 263060 245700 263062
rect 245764 263060 245770 263124
rect 156892 262848 200314 262850
rect 156892 262792 198554 262848
rect 198610 262792 200314 262848
rect 156892 262790 200314 262792
rect 156892 262788 156898 262790
rect 198549 262787 198615 262790
rect 158713 262578 158779 262581
rect 156676 262576 158779 262578
rect 156676 262520 158718 262576
rect 158774 262520 158779 262576
rect 156676 262518 158779 262520
rect 158713 262515 158779 262518
rect 197997 262306 198063 262309
rect 198641 262306 198707 262309
rect 245929 262306 245995 262309
rect 197997 262304 200284 262306
rect 197997 262248 198002 262304
rect 198058 262248 198646 262304
rect 198702 262248 200284 262304
rect 197997 262246 200284 262248
rect 244076 262304 245995 262306
rect 244076 262248 245934 262304
rect 245990 262248 245995 262304
rect 244076 262246 245995 262248
rect 197997 262243 198063 262246
rect 198641 262243 198707 262246
rect 245929 262243 245995 262246
rect 163497 262170 163563 262173
rect 165061 262170 165127 262173
rect 163497 262168 165127 262170
rect 163497 262112 163502 262168
rect 163558 262112 165066 262168
rect 165122 262112 165127 262168
rect 163497 262110 165127 262112
rect 163497 262107 163563 262110
rect 165061 262107 165127 262110
rect 66529 262034 66595 262037
rect 66529 262032 68908 262034
rect 66529 261976 66534 262032
rect 66590 261976 68908 262032
rect 66529 261974 68908 261976
rect 66529 261971 66595 261974
rect 245745 261762 245811 261765
rect 244076 261760 245811 261762
rect 244076 261704 245750 261760
rect 245806 261704 245811 261760
rect 244076 261702 245811 261704
rect 245745 261699 245811 261702
rect 185342 261564 185348 261628
rect 185412 261626 185418 261628
rect 195278 261626 195284 261628
rect 185412 261566 195284 261626
rect 185412 261564 185418 261566
rect 195278 261564 195284 261566
rect 195348 261564 195354 261628
rect 158989 261490 159055 261493
rect 156676 261488 159055 261490
rect 156676 261432 158994 261488
rect 159050 261432 159055 261488
rect 156676 261430 159055 261432
rect 158989 261427 159055 261430
rect 163773 261490 163839 261493
rect 186313 261490 186379 261493
rect 163773 261488 186379 261490
rect 163773 261432 163778 261488
rect 163834 261432 186318 261488
rect 186374 261432 186379 261488
rect 163773 261430 186379 261432
rect 163773 261427 163839 261430
rect 186313 261427 186379 261430
rect 197353 261490 197419 261493
rect 246021 261490 246087 261493
rect 252737 261490 252803 261493
rect 197353 261488 200284 261490
rect 197353 261432 197358 261488
rect 197414 261432 200284 261488
rect 197353 261430 200284 261432
rect 246021 261488 252803 261490
rect 246021 261432 246026 261488
rect 246082 261432 252742 261488
rect 252798 261432 252803 261488
rect 246021 261430 252803 261432
rect 197353 261427 197419 261430
rect 246021 261427 246087 261430
rect 252737 261427 252803 261430
rect 244222 261292 244228 261356
rect 244292 261354 244298 261356
rect 299565 261354 299631 261357
rect 244292 261352 299631 261354
rect 244292 261296 299570 261352
rect 299626 261296 299631 261352
rect 244292 261294 299631 261296
rect 244292 261292 244298 261294
rect 299565 261291 299631 261294
rect 66345 260946 66411 260949
rect 195421 260946 195487 260949
rect 195830 260946 195836 260948
rect 66345 260944 68908 260946
rect 66345 260888 66350 260944
rect 66406 260888 68908 260944
rect 66345 260886 68908 260888
rect 195421 260944 195836 260946
rect 195421 260888 195426 260944
rect 195482 260888 195836 260944
rect 195421 260886 195836 260888
rect 66345 260883 66411 260886
rect 195421 260883 195487 260886
rect 195830 260884 195836 260886
rect 195900 260946 195906 260948
rect 245837 260946 245903 260949
rect 195900 260886 200284 260946
rect 244076 260944 245903 260946
rect 244076 260888 245842 260944
rect 245898 260888 245903 260944
rect 244076 260886 245903 260888
rect 195900 260884 195906 260886
rect 245837 260883 245903 260886
rect 159950 260748 159956 260812
rect 160020 260810 160026 260812
rect 160093 260810 160159 260813
rect 160020 260808 160159 260810
rect 160020 260752 160098 260808
rect 160154 260752 160159 260808
rect 160020 260750 160159 260752
rect 160020 260748 160026 260750
rect 160093 260747 160159 260750
rect 161974 260674 161980 260676
rect 156646 260614 161980 260674
rect 156646 260372 156706 260614
rect 161974 260612 161980 260614
rect 162044 260674 162050 260676
rect 162761 260674 162827 260677
rect 162044 260672 162827 260674
rect 162044 260616 162766 260672
rect 162822 260616 162827 260672
rect 162044 260614 162827 260616
rect 162044 260612 162050 260614
rect 162761 260611 162827 260614
rect 197353 260130 197419 260133
rect 247309 260130 247375 260133
rect 309041 260130 309107 260133
rect 197353 260128 200284 260130
rect 197353 260072 197358 260128
rect 197414 260072 200284 260128
rect 197353 260070 200284 260072
rect 244076 260128 309107 260130
rect 244076 260072 247314 260128
rect 247370 260072 309046 260128
rect 309102 260072 309107 260128
rect 244076 260070 309107 260072
rect 197353 260067 197419 260070
rect 247309 260067 247375 260070
rect 309041 260067 309107 260070
rect 67541 259858 67607 259861
rect 67541 259856 68908 259858
rect 67541 259800 67546 259856
rect 67602 259800 68908 259856
rect 67541 259798 68908 259800
rect 67541 259795 67607 259798
rect 243486 259796 243492 259860
rect 243556 259796 243562 259860
rect 243494 259586 243554 259796
rect 246389 259586 246455 259589
rect 243494 259584 246455 259586
rect 243494 259556 246394 259584
rect 243524 259528 246394 259556
rect 246450 259528 246455 259584
rect 243524 259526 246455 259528
rect 246389 259523 246455 259526
rect 180241 259450 180307 259453
rect 156646 259448 180307 259450
rect 156646 259392 180246 259448
rect 180302 259392 180307 259448
rect 156646 259390 180307 259392
rect 156646 259284 156706 259390
rect 180241 259387 180307 259390
rect 309041 259450 309107 259453
rect 309869 259450 309935 259453
rect 309041 259448 309935 259450
rect 309041 259392 309046 259448
rect 309102 259392 309874 259448
rect 309930 259392 309935 259448
rect 309041 259390 309935 259392
rect 309041 259387 309107 259390
rect 309869 259387 309935 259390
rect 197353 259314 197419 259317
rect 197353 259312 200284 259314
rect 197353 259256 197358 259312
rect 197414 259256 200284 259312
rect 197353 259254 200284 259256
rect 197353 259251 197419 259254
rect 583017 258906 583083 258909
rect 583520 258906 584960 258996
rect 583017 258904 584960 258906
rect 583017 258848 583022 258904
rect 583078 258848 584960 258904
rect 583017 258846 584960 258848
rect 583017 258843 583083 258846
rect 197353 258770 197419 258773
rect 245745 258770 245811 258773
rect 197353 258768 200284 258770
rect 66253 258090 66319 258093
rect 66253 258088 66362 258090
rect 66253 258032 66258 258088
rect 66314 258032 66362 258088
rect 66253 258027 66362 258032
rect 66302 257954 66362 258027
rect 68878 257954 68938 258740
rect 197353 258712 197358 258768
rect 197414 258712 200284 258768
rect 197353 258710 200284 258712
rect 244076 258768 245811 258770
rect 244076 258712 245750 258768
rect 245806 258712 245811 258768
rect 583520 258756 584960 258846
rect 244076 258710 245811 258712
rect 197353 258707 197419 258710
rect 245745 258707 245811 258710
rect 158805 258226 158871 258229
rect 244549 258226 244615 258229
rect 156676 258224 158871 258226
rect 156676 258168 158810 258224
rect 158866 258168 158871 258224
rect 156676 258166 158871 258168
rect 244076 258224 244615 258226
rect 244076 258168 244554 258224
rect 244610 258168 244615 258224
rect 244076 258166 244615 258168
rect 158805 258163 158871 258166
rect 244549 258163 244615 258166
rect 183001 258090 183067 258093
rect 182958 258088 183067 258090
rect 182958 258032 183006 258088
rect 183062 258032 183067 258088
rect 182958 258027 183067 258032
rect 66302 257894 68938 257954
rect 180241 257954 180307 257957
rect 182958 257954 183018 258027
rect 180241 257952 183018 257954
rect 180241 257896 180246 257952
rect 180302 257896 183018 257952
rect 180241 257894 183018 257896
rect 180241 257891 180307 257894
rect 66805 257682 66871 257685
rect 195329 257682 195395 257685
rect 200254 257682 200314 257924
rect 66805 257680 68908 257682
rect 66805 257624 66810 257680
rect 66866 257624 68908 257680
rect 66805 257622 68908 257624
rect 180750 257680 195395 257682
rect 180750 257624 195334 257680
rect 195390 257624 195395 257680
rect 180750 257622 195395 257624
rect 66805 257619 66871 257622
rect 174813 257274 174879 257277
rect 180750 257274 180810 257622
rect 195329 257619 195395 257622
rect 200070 257622 200314 257682
rect 200070 257546 200130 257622
rect 174813 257272 180810 257274
rect 174813 257216 174818 257272
rect 174874 257216 180810 257272
rect 174813 257214 180810 257216
rect 195286 257486 200130 257546
rect 174813 257211 174879 257214
rect 158713 257138 158779 257141
rect 156676 257136 158779 257138
rect 156676 257080 158718 257136
rect 158774 257080 158779 257136
rect 156676 257078 158779 257080
rect 158713 257075 158779 257078
rect 189073 257002 189139 257005
rect 190269 257002 190335 257005
rect 195286 257002 195346 257486
rect 197353 257410 197419 257413
rect 245745 257410 245811 257413
rect 197353 257408 200284 257410
rect 197353 257352 197358 257408
rect 197414 257352 200284 257408
rect 197353 257350 200284 257352
rect 244076 257408 245811 257410
rect 244076 257352 245750 257408
rect 245806 257352 245811 257408
rect 244076 257350 245811 257352
rect 197353 257347 197419 257350
rect 245745 257347 245811 257350
rect 189073 257000 195346 257002
rect 189073 256944 189078 257000
rect 189134 256944 190274 257000
rect 190330 256944 195346 257000
rect 189073 256942 195346 256944
rect 189073 256939 189139 256942
rect 190269 256939 190335 256942
rect 67357 256594 67423 256597
rect 197353 256594 197419 256597
rect 245653 256594 245719 256597
rect 67357 256592 68908 256594
rect 67357 256536 67362 256592
rect 67418 256536 68908 256592
rect 67357 256534 68908 256536
rect 197353 256592 200284 256594
rect 197353 256536 197358 256592
rect 197414 256536 200284 256592
rect 197353 256534 200284 256536
rect 244076 256592 245719 256594
rect 244076 256536 245658 256592
rect 245714 256536 245719 256592
rect 244076 256534 245719 256536
rect 67357 256531 67423 256534
rect 197353 256531 197419 256534
rect 245653 256531 245719 256534
rect 158713 256322 158779 256325
rect 156676 256320 158779 256322
rect 156676 256264 158718 256320
rect 158774 256264 158779 256320
rect 156676 256262 158779 256264
rect 158713 256259 158779 256262
rect 245745 256050 245811 256053
rect 244076 256048 245811 256050
rect 244076 255992 245750 256048
rect 245806 255992 245811 256048
rect 244076 255990 245811 255992
rect 245745 255987 245811 255990
rect 65977 255506 66043 255509
rect 166809 255506 166875 255509
rect 200254 255506 200314 255748
rect 65977 255504 68908 255506
rect 65977 255448 65982 255504
rect 66038 255448 68908 255504
rect 65977 255446 68908 255448
rect 166809 255504 200314 255506
rect 166809 255448 166814 255504
rect 166870 255448 200314 255504
rect 166809 255446 200314 255448
rect 65977 255443 66043 255446
rect 166809 255443 166875 255446
rect 157977 255234 158043 255237
rect 158529 255234 158595 255237
rect 156676 255232 158595 255234
rect 156676 255176 157982 255232
rect 158038 255176 158534 255232
rect 158590 255176 158595 255232
rect 156676 255174 158595 255176
rect 157977 255171 158043 255174
rect 158529 255171 158595 255174
rect 200254 254690 200314 255204
rect 244046 254693 244106 255204
rect 180750 254630 200314 254690
rect 243997 254688 244106 254693
rect 243997 254632 244002 254688
rect 244058 254632 244106 254688
rect 243997 254630 244106 254632
rect 163497 254554 163563 254557
rect 177297 254554 177363 254557
rect 163497 254552 177363 254554
rect 163497 254496 163502 254552
rect 163558 254496 177302 254552
rect 177358 254496 177363 254552
rect 163497 254494 177363 254496
rect 163497 254491 163563 254494
rect 177297 254491 177363 254494
rect 66621 254418 66687 254421
rect 66621 254416 68908 254418
rect 66621 254360 66626 254416
rect 66682 254360 68908 254416
rect 66621 254358 68908 254360
rect 66621 254355 66687 254358
rect -960 254146 480 254236
rect 2773 254146 2839 254149
rect 164141 254146 164207 254149
rect -960 254144 2839 254146
rect -960 254088 2778 254144
rect 2834 254088 2839 254144
rect -960 254086 2839 254088
rect 156676 254144 164207 254146
rect 156676 254088 164146 254144
rect 164202 254088 164207 254144
rect 156676 254086 164207 254088
rect -960 253996 480 254086
rect 2773 254083 2839 254086
rect 164141 254083 164207 254086
rect 170489 254010 170555 254013
rect 171041 254010 171107 254013
rect 180750 254010 180810 254630
rect 243997 254627 244063 254630
rect 197353 254418 197419 254421
rect 245837 254418 245903 254421
rect 197353 254416 200284 254418
rect 197353 254360 197358 254416
rect 197414 254360 200284 254416
rect 197353 254358 200284 254360
rect 244076 254416 245903 254418
rect 244076 254360 245842 254416
rect 245898 254360 245903 254416
rect 244076 254358 245903 254360
rect 197353 254355 197419 254358
rect 245837 254355 245903 254358
rect 170489 254008 180810 254010
rect 170489 253952 170494 254008
rect 170550 253952 171046 254008
rect 171102 253952 180810 254008
rect 170489 253950 180810 253952
rect 170489 253947 170555 253950
rect 171041 253947 171107 253950
rect 245929 253874 245995 253877
rect 244076 253872 245995 253874
rect 244076 253816 245934 253872
rect 245990 253816 245995 253872
rect 244076 253814 245995 253816
rect 245929 253811 245995 253814
rect 197353 253602 197419 253605
rect 197353 253600 200284 253602
rect 197353 253544 197358 253600
rect 197414 253544 200284 253600
rect 197353 253542 200284 253544
rect 197353 253539 197419 253542
rect 66805 253330 66871 253333
rect 66805 253328 68908 253330
rect 66805 253272 66810 253328
rect 66866 253272 68908 253328
rect 66805 253270 68908 253272
rect 66805 253267 66871 253270
rect 165521 253194 165587 253197
rect 194409 253194 194475 253197
rect 165521 253192 194475 253194
rect 165521 253136 165526 253192
rect 165582 253136 194414 253192
rect 194470 253136 194475 253192
rect 165521 253134 194475 253136
rect 165521 253131 165587 253134
rect 194409 253131 194475 253134
rect 158713 253058 158779 253061
rect 156676 253056 158779 253058
rect 156676 253000 158718 253056
rect 158774 253000 158779 253056
rect 156676 252998 158779 253000
rect 158713 252995 158779 252998
rect 197353 253058 197419 253061
rect 246021 253058 246087 253061
rect 197353 253056 200284 253058
rect 197353 253000 197358 253056
rect 197414 253000 200284 253056
rect 197353 252998 200284 253000
rect 244076 253056 246087 253058
rect 244076 253000 246026 253056
rect 246082 253000 246087 253056
rect 244076 252998 246087 253000
rect 197353 252995 197419 252998
rect 246021 252995 246087 252998
rect 251214 252452 251220 252516
rect 251284 252514 251290 252516
rect 251357 252514 251423 252517
rect 251284 252512 251423 252514
rect 251284 252456 251362 252512
rect 251418 252456 251423 252512
rect 251284 252454 251423 252456
rect 251284 252452 251290 252454
rect 251357 252451 251423 252454
rect 67265 252242 67331 252245
rect 245929 252242 245995 252245
rect 67265 252240 68908 252242
rect 67265 252184 67270 252240
rect 67326 252184 68908 252240
rect 244076 252240 245995 252242
rect 67265 252182 68908 252184
rect 67265 252179 67331 252182
rect 200254 251970 200314 252212
rect 244076 252184 245934 252240
rect 245990 252184 245995 252240
rect 244076 252182 245995 252184
rect 245929 252179 245995 252182
rect 156646 251290 156706 251940
rect 200070 251910 200314 251970
rect 160829 251834 160895 251837
rect 198590 251834 198596 251836
rect 160829 251832 198596 251834
rect 160829 251776 160834 251832
rect 160890 251776 198596 251832
rect 160829 251774 198596 251776
rect 160829 251771 160895 251774
rect 198590 251772 198596 251774
rect 198660 251834 198666 251836
rect 200070 251834 200130 251910
rect 198660 251774 200130 251834
rect 198660 251772 198666 251774
rect 197353 251698 197419 251701
rect 245929 251698 245995 251701
rect 197353 251696 200284 251698
rect 197353 251640 197358 251696
rect 197414 251640 200284 251696
rect 197353 251638 200284 251640
rect 244076 251696 245995 251698
rect 244076 251640 245934 251696
rect 245990 251640 245995 251696
rect 244076 251638 245995 251640
rect 197353 251635 197419 251638
rect 245929 251635 245995 251638
rect 172462 251290 172468 251292
rect 156646 251230 172468 251290
rect 172462 251228 172468 251230
rect 172532 251228 172538 251292
rect 66805 251154 66871 251157
rect 66805 251152 68908 251154
rect 66805 251096 66810 251152
rect 66866 251096 68908 251152
rect 66805 251094 68908 251096
rect 66805 251091 66871 251094
rect 158713 250882 158779 250885
rect 156676 250880 158779 250882
rect 156676 250824 158718 250880
rect 158774 250824 158779 250880
rect 156676 250822 158779 250824
rect 158713 250819 158779 250822
rect 197445 250882 197511 250885
rect 245929 250882 245995 250885
rect 197445 250880 200284 250882
rect 197445 250824 197450 250880
rect 197506 250824 200284 250880
rect 197445 250822 200284 250824
rect 244076 250880 245995 250882
rect 244076 250824 245934 250880
rect 245990 250824 245995 250880
rect 244076 250822 245995 250824
rect 197445 250819 197511 250822
rect 245929 250819 245995 250822
rect 163681 250474 163747 250477
rect 172329 250474 172395 250477
rect 163681 250472 172395 250474
rect 163681 250416 163686 250472
rect 163742 250416 172334 250472
rect 172390 250416 172395 250472
rect 163681 250414 172395 250416
rect 163681 250411 163747 250414
rect 172329 250411 172395 250414
rect 245837 250338 245903 250341
rect 244076 250336 245903 250338
rect 244076 250280 245842 250336
rect 245898 250280 245903 250336
rect 244076 250278 245903 250280
rect 245837 250275 245903 250278
rect 197353 250066 197419 250069
rect 197353 250064 200284 250066
rect 61745 249930 61811 249933
rect 68878 249930 68938 250036
rect 197353 250008 197358 250064
rect 197414 250008 200284 250064
rect 197353 250006 200284 250008
rect 197353 250003 197419 250006
rect 61745 249928 68938 249930
rect 61745 249872 61750 249928
rect 61806 249872 68938 249928
rect 61745 249870 68938 249872
rect 182449 249930 182515 249933
rect 183461 249930 183527 249933
rect 195094 249930 195100 249932
rect 182449 249928 195100 249930
rect 182449 249872 182454 249928
rect 182510 249872 183466 249928
rect 183522 249872 195100 249928
rect 182449 249870 195100 249872
rect 61745 249867 61811 249870
rect 182449 249867 182515 249870
rect 183461 249867 183527 249870
rect 195094 249868 195100 249870
rect 195164 249868 195170 249932
rect 158805 249794 158871 249797
rect 156676 249792 158871 249794
rect 156676 249736 158810 249792
rect 158866 249736 158871 249792
rect 156676 249734 158871 249736
rect 158805 249731 158871 249734
rect 251265 249794 251331 249797
rect 252369 249794 252435 249797
rect 251265 249792 252435 249794
rect 251265 249736 251270 249792
rect 251326 249736 252374 249792
rect 252430 249736 252435 249792
rect 251265 249734 252435 249736
rect 251265 249731 251331 249734
rect 252369 249731 252435 249734
rect 197353 249522 197419 249525
rect 197353 249520 200284 249522
rect 197353 249464 197358 249520
rect 197414 249464 200284 249520
rect 197353 249462 200284 249464
rect 197353 249459 197419 249462
rect 167821 249250 167887 249253
rect 174813 249250 174879 249253
rect 167821 249248 174879 249250
rect 167821 249192 167826 249248
rect 167882 249192 174818 249248
rect 174874 249192 174879 249248
rect 167821 249190 174879 249192
rect 167821 249187 167887 249190
rect 174813 249187 174879 249190
rect 159725 249114 159791 249117
rect 182449 249114 182515 249117
rect 159725 249112 182515 249114
rect 159725 249056 159730 249112
rect 159786 249056 182454 249112
rect 182510 249056 182515 249112
rect 159725 249054 182515 249056
rect 159725 249051 159791 249054
rect 182449 249051 182515 249054
rect 67766 248916 67772 248980
rect 67836 248978 67842 248980
rect 244046 248978 244106 249492
rect 251265 248978 251331 248981
rect 67836 248918 68908 248978
rect 244046 248976 251331 248978
rect 244046 248920 251270 248976
rect 251326 248920 251331 248976
rect 244046 248918 251331 248920
rect 67836 248916 67842 248918
rect 251265 248915 251331 248918
rect 158897 248706 158963 248709
rect 156676 248704 158963 248706
rect 156676 248648 158902 248704
rect 158958 248648 158963 248704
rect 156676 248646 158963 248648
rect 158897 248643 158963 248646
rect 197813 248706 197879 248709
rect 244457 248706 244523 248709
rect 197813 248704 200284 248706
rect 197813 248648 197818 248704
rect 197874 248648 200284 248704
rect 197813 248646 200284 248648
rect 244076 248704 244523 248706
rect 244076 248648 244462 248704
rect 244518 248648 244523 248704
rect 244076 248646 244523 248648
rect 197813 248643 197879 248646
rect 244457 248643 244523 248646
rect 244774 248162 244780 248164
rect 244076 248102 244780 248162
rect 244774 248100 244780 248102
rect 244844 248162 244850 248164
rect 245653 248162 245719 248165
rect 244844 248160 245719 248162
rect 244844 248104 245658 248160
rect 245714 248104 245719 248160
rect 244844 248102 245719 248104
rect 244844 248100 244850 248102
rect 245653 248099 245719 248102
rect 197353 247890 197419 247893
rect 197353 247888 200284 247890
rect 59118 247012 59124 247076
rect 59188 247074 59194 247076
rect 68878 247074 68938 247860
rect 197353 247832 197358 247888
rect 197414 247832 200284 247888
rect 197353 247830 200284 247832
rect 197353 247827 197419 247830
rect 159541 247618 159607 247621
rect 156676 247616 159607 247618
rect 156676 247560 159546 247616
rect 159602 247560 159607 247616
rect 156676 247558 159607 247560
rect 159541 247555 159607 247558
rect 245929 247346 245995 247349
rect 244076 247344 245995 247346
rect 59188 247014 68938 247074
rect 169661 247074 169727 247077
rect 171133 247074 171199 247077
rect 169661 247072 171199 247074
rect 169661 247016 169666 247072
rect 169722 247016 171138 247072
rect 171194 247016 171199 247072
rect 169661 247014 171199 247016
rect 59188 247012 59194 247014
rect 169661 247011 169727 247014
rect 171133 247011 171199 247014
rect 188286 247012 188292 247076
rect 188356 247074 188362 247076
rect 191465 247074 191531 247077
rect 200254 247074 200314 247316
rect 244076 247288 245934 247344
rect 245990 247288 245995 247344
rect 244076 247286 245995 247288
rect 245929 247283 245995 247286
rect 188356 247072 200314 247074
rect 188356 247016 191470 247072
rect 191526 247016 200314 247072
rect 188356 247014 200314 247016
rect 188356 247012 188362 247014
rect 191465 247011 191531 247014
rect 66805 246802 66871 246805
rect 66805 246800 68908 246802
rect 66805 246744 66810 246800
rect 66866 246744 68908 246800
rect 66805 246742 68908 246744
rect 66805 246739 66871 246742
rect 181437 246530 181503 246533
rect 188337 246530 188403 246533
rect 161430 246528 188403 246530
rect 156646 246258 156706 246500
rect 161430 246472 181442 246528
rect 181498 246472 188342 246528
rect 188398 246472 188403 246528
rect 161430 246470 188403 246472
rect 161430 246258 161490 246470
rect 181437 246467 181503 246470
rect 188337 246467 188403 246470
rect 197118 246468 197124 246532
rect 197188 246530 197194 246532
rect 245837 246530 245903 246533
rect 197188 246470 200284 246530
rect 244076 246528 245903 246530
rect 244076 246472 245842 246528
rect 245898 246472 245903 246528
rect 244076 246470 245903 246472
rect 197188 246468 197194 246470
rect 245837 246467 245903 246470
rect 380985 246258 381051 246261
rect 156646 246198 161490 246258
rect 364290 246256 381051 246258
rect 364290 246200 380990 246256
rect 381046 246200 381051 246256
rect 364290 246198 381051 246200
rect 245929 245986 245995 245989
rect 244076 245984 245995 245986
rect 193806 245788 193812 245852
rect 193876 245850 193882 245852
rect 197118 245850 197124 245852
rect 193876 245790 197124 245850
rect 193876 245788 193882 245790
rect 197118 245788 197124 245790
rect 197188 245788 197194 245852
rect 67633 245714 67699 245717
rect 191833 245716 191899 245717
rect 191782 245714 191788 245716
rect 67633 245712 68908 245714
rect 67633 245656 67638 245712
rect 67694 245656 68908 245712
rect 67633 245654 68908 245656
rect 191742 245654 191788 245714
rect 191852 245712 191899 245716
rect 191894 245656 191899 245712
rect 67633 245651 67699 245654
rect 191782 245652 191788 245654
rect 191852 245652 191899 245656
rect 191833 245651 191899 245652
rect 195237 245714 195303 245717
rect 195830 245714 195836 245716
rect 195237 245712 195836 245714
rect 195237 245656 195242 245712
rect 195298 245656 195836 245712
rect 195237 245654 195836 245656
rect 195237 245651 195303 245654
rect 195830 245652 195836 245654
rect 195900 245714 195906 245716
rect 200254 245714 200314 245956
rect 244076 245928 245934 245984
rect 245990 245928 245995 245984
rect 244076 245926 245995 245928
rect 245929 245923 245995 245926
rect 195900 245654 200314 245714
rect 255405 245714 255471 245717
rect 361481 245714 361547 245717
rect 364290 245714 364350 246198
rect 380985 246195 381051 246198
rect 255405 245712 364350 245714
rect 255405 245656 255410 245712
rect 255466 245656 361486 245712
rect 361542 245656 364350 245712
rect 255405 245654 364350 245656
rect 195900 245652 195906 245654
rect 255405 245651 255471 245654
rect 361481 245651 361547 245654
rect 583109 245578 583175 245581
rect 583520 245578 584960 245668
rect 583109 245576 584960 245578
rect 583109 245520 583114 245576
rect 583170 245520 584960 245576
rect 583109 245518 584960 245520
rect 583109 245515 583175 245518
rect 583520 245428 584960 245518
rect 156646 244898 156706 245412
rect 197721 245170 197787 245173
rect 198641 245170 198707 245173
rect 245653 245170 245719 245173
rect 197721 245168 200284 245170
rect 197721 245112 197726 245168
rect 197782 245112 198646 245168
rect 198702 245112 200284 245168
rect 197721 245110 200284 245112
rect 244076 245168 245719 245170
rect 244076 245112 245658 245168
rect 245714 245112 245719 245168
rect 244076 245110 245719 245112
rect 197721 245107 197787 245110
rect 198641 245107 198707 245110
rect 245653 245107 245719 245110
rect 171869 245034 171935 245037
rect 161430 245032 171935 245034
rect 161430 244976 171874 245032
rect 171930 244976 171935 245032
rect 161430 244974 171935 244976
rect 160001 244898 160067 244901
rect 161430 244898 161490 244974
rect 171869 244971 171935 244974
rect 156646 244896 161490 244898
rect 156646 244840 160006 244896
rect 160062 244840 161490 244896
rect 156646 244838 161490 244840
rect 172329 244898 172395 244901
rect 184749 244898 184815 244901
rect 172329 244896 184815 244898
rect 172329 244840 172334 244896
rect 172390 244840 184754 244896
rect 184810 244840 184815 244896
rect 172329 244838 184815 244840
rect 160001 244835 160067 244838
rect 172329 244835 172395 244838
rect 184749 244835 184815 244838
rect 66805 244626 66871 244629
rect 246297 244626 246363 244629
rect 66805 244624 68908 244626
rect 66805 244568 66810 244624
rect 66866 244568 68908 244624
rect 66805 244566 68908 244568
rect 244076 244624 246363 244626
rect 244076 244568 246302 244624
rect 246358 244568 246363 244624
rect 244076 244566 246363 244568
rect 66805 244563 66871 244566
rect 246297 244563 246363 244566
rect 158713 244354 158779 244357
rect 156676 244352 158779 244354
rect 156676 244296 158718 244352
rect 158774 244296 158779 244352
rect 156676 244294 158779 244296
rect 158713 244291 158779 244294
rect 198549 244354 198615 244357
rect 198549 244352 200284 244354
rect 198549 244296 198554 244352
rect 198610 244296 200284 244352
rect 198549 244294 200284 244296
rect 198549 244291 198615 244294
rect 197353 243810 197419 243813
rect 245837 243810 245903 243813
rect 197353 243808 200284 243810
rect 197353 243752 197358 243808
rect 197414 243752 200284 243808
rect 197353 243750 200284 243752
rect 244076 243808 245903 243810
rect 244076 243752 245842 243808
rect 245898 243752 245903 243808
rect 244076 243750 245903 243752
rect 197353 243747 197419 243750
rect 245837 243747 245903 243750
rect 66805 243538 66871 243541
rect 66805 243536 68908 243538
rect 66805 243480 66810 243536
rect 66866 243480 68908 243536
rect 66805 243478 68908 243480
rect 66805 243475 66871 243478
rect 156822 243476 156828 243540
rect 156892 243538 156898 243540
rect 172329 243538 172395 243541
rect 156892 243536 172395 243538
rect 156892 243480 172334 243536
rect 172390 243480 172395 243536
rect 156892 243478 172395 243480
rect 156892 243476 156898 243478
rect 172329 243475 172395 243478
rect 158713 243266 158779 243269
rect 156676 243264 158779 243266
rect 156676 243208 158718 243264
rect 158774 243208 158779 243264
rect 156676 243206 158779 243208
rect 158713 243203 158779 243206
rect 183093 243130 183159 243133
rect 183369 243130 183435 243133
rect 199326 243130 199332 243132
rect 183093 243128 199332 243130
rect 183093 243072 183098 243128
rect 183154 243072 183374 243128
rect 183430 243072 199332 243128
rect 183093 243070 199332 243072
rect 183093 243067 183159 243070
rect 183369 243067 183435 243070
rect 199326 243068 199332 243070
rect 199396 243068 199402 243132
rect 171685 242994 171751 242997
rect 259494 242994 259500 242996
rect 171685 242992 200284 242994
rect 171685 242936 171690 242992
rect 171746 242936 200284 242992
rect 171685 242934 200284 242936
rect 244076 242934 259500 242994
rect 171685 242931 171751 242934
rect 259494 242932 259500 242934
rect 259564 242994 259570 242996
rect 260741 242994 260807 242997
rect 259564 242992 260807 242994
rect 259564 242936 260746 242992
rect 260802 242936 260807 242992
rect 259564 242934 260807 242936
rect 259564 242932 259570 242934
rect 260741 242931 260807 242934
rect 165061 242858 165127 242861
rect 165654 242858 165660 242860
rect 165061 242856 165660 242858
rect 165061 242800 165066 242856
rect 165122 242800 165660 242856
rect 165061 242798 165660 242800
rect 165061 242795 165127 242798
rect 165654 242796 165660 242798
rect 165724 242796 165730 242860
rect 167913 242858 167979 242861
rect 168281 242858 168347 242861
rect 167913 242856 168347 242858
rect 167913 242800 167918 242856
rect 167974 242800 168286 242856
rect 168342 242800 168347 242856
rect 167913 242798 168347 242800
rect 167913 242795 167979 242798
rect 168281 242795 168347 242798
rect 246389 242450 246455 242453
rect 244076 242448 246455 242450
rect 69430 241906 69490 242420
rect 244076 242392 246394 242448
rect 246450 242392 246455 242448
rect 244076 242390 246455 242392
rect 246389 242387 246455 242390
rect 158161 242178 158227 242181
rect 156676 242176 158227 242178
rect 156676 242120 158166 242176
rect 158222 242120 158227 242176
rect 156676 242118 158227 242120
rect 158161 242115 158227 242118
rect 197353 242178 197419 242181
rect 197353 242176 200284 242178
rect 197353 242120 197358 242176
rect 197414 242120 200284 242176
rect 197353 242118 200284 242120
rect 197353 242115 197419 242118
rect 80973 242044 81039 242045
rect 154665 242044 154731 242045
rect 80973 242042 81020 242044
rect 80928 242040 81020 242042
rect 80928 241984 80978 242040
rect 80928 241982 81020 241984
rect 80973 241980 81020 241982
rect 81084 241980 81090 242044
rect 154614 241980 154620 242044
rect 154684 242042 154731 242044
rect 156689 242042 156755 242045
rect 168465 242042 168531 242045
rect 154684 242040 154776 242042
rect 154726 241984 154776 242040
rect 154684 241982 154776 241984
rect 156689 242040 168531 242042
rect 156689 241984 156694 242040
rect 156750 241984 168470 242040
rect 168526 241984 168531 242040
rect 156689 241982 168531 241984
rect 154684 241980 154731 241982
rect 80973 241979 81039 241980
rect 154665 241979 154731 241980
rect 156689 241979 156755 241982
rect 168465 241979 168531 241982
rect 69657 241906 69723 241909
rect 69430 241904 69723 241906
rect 69430 241848 69662 241904
rect 69718 241848 69723 241904
rect 69430 241846 69723 241848
rect 69657 241843 69723 241846
rect 178953 241906 179019 241909
rect 179321 241906 179387 241909
rect 199745 241906 199811 241909
rect 178953 241904 199811 241906
rect 178953 241848 178958 241904
rect 179014 241848 179326 241904
rect 179382 241848 199750 241904
rect 199806 241848 199811 241904
rect 178953 241846 199811 241848
rect 178953 241843 179019 241846
rect 179321 241843 179387 241846
rect 199745 241843 199811 241846
rect 192661 241770 192727 241773
rect 196750 241770 196756 241772
rect 192661 241768 196756 241770
rect 192661 241712 192666 241768
rect 192722 241712 196756 241768
rect 192661 241710 196756 241712
rect 192661 241707 192727 241710
rect 196750 241708 196756 241710
rect 196820 241708 196826 241772
rect 167913 241634 167979 241637
rect 192661 241634 192727 241637
rect 167913 241632 192727 241634
rect 167913 241576 167918 241632
rect 167974 241576 192666 241632
rect 192722 241576 192727 241632
rect 167913 241574 192727 241576
rect 167913 241571 167979 241574
rect 192661 241571 192727 241574
rect 198825 241634 198891 241637
rect 245745 241634 245811 241637
rect 198825 241632 200284 241634
rect 198825 241576 198830 241632
rect 198886 241576 200284 241632
rect 243524 241632 245811 241634
rect 243524 241604 245750 241632
rect 198825 241574 200284 241576
rect 243494 241576 245750 241604
rect 245806 241576 245811 241632
rect 243494 241574 245811 241576
rect 198825 241571 198891 241574
rect 67398 241436 67404 241500
rect 67468 241498 67474 241500
rect 73797 241498 73863 241501
rect 67468 241496 73863 241498
rect 67468 241440 73802 241496
rect 73858 241440 73863 241496
rect 67468 241438 73863 241440
rect 67468 241436 67474 241438
rect 73797 241435 73863 241438
rect 83958 241436 83964 241500
rect 84028 241498 84034 241500
rect 93853 241498 93919 241501
rect 94911 241498 94977 241501
rect 84028 241496 94977 241498
rect 84028 241440 93858 241496
rect 93914 241440 94916 241496
rect 94972 241440 94977 241496
rect 84028 241438 94977 241440
rect 84028 241436 84034 241438
rect 93853 241435 93919 241438
rect 94911 241435 94977 241438
rect 191557 241498 191623 241501
rect 194317 241498 194383 241501
rect 191557 241496 194383 241498
rect 191557 241440 191562 241496
rect 191618 241440 194322 241496
rect 194378 241440 194383 241496
rect 191557 241438 194383 241440
rect 191557 241435 191623 241438
rect 194317 241435 194383 241438
rect 243494 241364 243554 241574
rect 245745 241571 245811 241574
rect 243486 241300 243492 241364
rect 243556 241300 243562 241364
rect 244089 241362 244155 241365
rect 262857 241362 262923 241365
rect 244089 241360 262923 241362
rect 244089 241304 244094 241360
rect 244150 241304 262862 241360
rect 262918 241304 262923 241360
rect 244089 241302 262923 241304
rect 244089 241299 244155 241302
rect 262857 241299 262923 241302
rect 150065 241226 150131 241229
rect 151721 241226 151787 241229
rect 160686 241226 160692 241228
rect 150065 241224 160692 241226
rect -960 241090 480 241180
rect 150065 241168 150070 241224
rect 150126 241168 151726 241224
rect 151782 241168 160692 241224
rect 150065 241166 160692 241168
rect 150065 241163 150131 241166
rect 151721 241163 151787 241166
rect 160686 241164 160692 241166
rect 160756 241164 160762 241228
rect 3509 241090 3575 241093
rect -960 241088 3575 241090
rect -960 241032 3514 241088
rect 3570 241032 3575 241088
rect -960 241030 3575 241032
rect -960 240940 480 241030
rect 3509 241027 3575 241030
rect 160185 241090 160251 241093
rect 170254 241090 170260 241092
rect 160185 241088 170260 241090
rect 160185 241032 160190 241088
rect 160246 241032 170260 241088
rect 160185 241030 170260 241032
rect 160185 241027 160251 241030
rect 170254 241028 170260 241030
rect 170324 241028 170330 241092
rect 130101 240954 130167 240957
rect 161565 240954 161631 240957
rect 130101 240952 161631 240954
rect 130101 240896 130106 240952
rect 130162 240896 161570 240952
rect 161626 240896 161631 240952
rect 130101 240894 161631 240896
rect 130101 240891 130167 240894
rect 161565 240891 161631 240894
rect 170949 240954 171015 240957
rect 190453 240954 190519 240957
rect 170949 240952 190519 240954
rect 170949 240896 170954 240952
rect 171010 240896 190458 240952
rect 190514 240896 190519 240952
rect 170949 240894 190519 240896
rect 170949 240891 171015 240894
rect 190453 240891 190519 240894
rect 63217 240818 63283 240821
rect 190361 240818 190427 240821
rect 194225 240818 194291 240821
rect 246941 240818 247007 240821
rect 63217 240816 194291 240818
rect 63217 240760 63222 240816
rect 63278 240760 190366 240816
rect 190422 240760 194230 240816
rect 194286 240760 194291 240816
rect 63217 240758 194291 240760
rect 63217 240755 63283 240758
rect 190361 240755 190427 240758
rect 194225 240755 194291 240758
rect 200070 240758 200284 240818
rect 244076 240816 247007 240818
rect 244076 240760 246946 240816
rect 247002 240760 247007 240816
rect 244076 240758 247007 240760
rect 194041 240682 194107 240685
rect 199561 240682 199627 240685
rect 200070 240682 200130 240758
rect 246941 240755 247007 240758
rect 194041 240680 200130 240682
rect 194041 240624 194046 240680
rect 194102 240624 199566 240680
rect 199622 240624 200130 240680
rect 194041 240622 200130 240624
rect 194041 240619 194107 240622
rect 199561 240619 199627 240622
rect 196617 240546 196683 240549
rect 199653 240546 199719 240549
rect 196617 240544 199719 240546
rect 196617 240488 196622 240544
rect 196678 240488 199658 240544
rect 199714 240488 199719 240544
rect 196617 240486 199719 240488
rect 196617 240483 196683 240486
rect 199653 240483 199719 240486
rect 198733 240410 198799 240413
rect 198733 240408 200866 240410
rect 198733 240352 198738 240408
rect 198794 240352 200866 240408
rect 198733 240350 200866 240352
rect 198733 240347 198799 240350
rect 155542 240214 155970 240274
rect 41321 240138 41387 240141
rect 72417 240138 72483 240141
rect 72693 240138 72759 240141
rect 41321 240136 72759 240138
rect 41321 240080 41326 240136
rect 41382 240080 72422 240136
rect 72478 240080 72698 240136
rect 72754 240080 72759 240136
rect 41321 240078 72759 240080
rect 41321 240075 41387 240078
rect 72417 240075 72483 240078
rect 72693 240075 72759 240078
rect 151997 240138 152063 240141
rect 153101 240138 153167 240141
rect 155542 240138 155602 240214
rect 151997 240136 155602 240138
rect 151997 240080 152002 240136
rect 152058 240080 153106 240136
rect 153162 240080 155602 240136
rect 151997 240078 155602 240080
rect 155677 240140 155743 240141
rect 155677 240136 155724 240140
rect 155788 240138 155794 240140
rect 155910 240138 155970 240214
rect 157374 240138 157380 240140
rect 155677 240080 155682 240136
rect 151997 240075 152063 240078
rect 153101 240075 153167 240078
rect 155677 240076 155724 240080
rect 155788 240078 155834 240138
rect 155910 240078 157380 240138
rect 155788 240076 155794 240078
rect 157374 240076 157380 240078
rect 157444 240076 157450 240140
rect 199745 240138 199811 240141
rect 200205 240138 200271 240141
rect 199745 240136 200271 240138
rect 199745 240080 199750 240136
rect 199806 240080 200210 240136
rect 200266 240080 200271 240136
rect 199745 240078 200271 240080
rect 200806 240138 200866 240350
rect 256693 240274 256759 240277
rect 244076 240272 256759 240274
rect 244076 240216 256698 240272
rect 256754 240216 256759 240272
rect 244076 240214 256759 240216
rect 256693 240211 256759 240214
rect 201033 240138 201099 240141
rect 202597 240140 202663 240141
rect 202597 240138 202644 240140
rect 200806 240136 201099 240138
rect 200806 240080 201038 240136
rect 201094 240080 201099 240136
rect 200806 240078 201099 240080
rect 202552 240136 202644 240138
rect 202552 240080 202602 240136
rect 202552 240078 202644 240080
rect 155677 240075 155743 240076
rect 199745 240075 199811 240078
rect 200205 240075 200271 240078
rect 201033 240075 201099 240078
rect 202597 240076 202644 240078
rect 202708 240076 202714 240140
rect 207933 240138 207999 240141
rect 208158 240138 208164 240140
rect 207933 240136 208164 240138
rect 207933 240080 207938 240136
rect 207994 240080 208164 240136
rect 207933 240078 208164 240080
rect 202597 240075 202663 240076
rect 207933 240075 207999 240078
rect 208158 240076 208164 240078
rect 208228 240076 208234 240140
rect 208301 240138 208367 240141
rect 210693 240140 210759 240141
rect 217501 240140 217567 240141
rect 208894 240138 208900 240140
rect 208301 240136 208900 240138
rect 208301 240080 208306 240136
rect 208362 240080 208900 240136
rect 208301 240078 208900 240080
rect 208301 240075 208367 240078
rect 208894 240076 208900 240078
rect 208964 240076 208970 240140
rect 210693 240138 210740 240140
rect 210648 240136 210740 240138
rect 210648 240080 210698 240136
rect 210648 240078 210740 240080
rect 210693 240076 210740 240078
rect 210804 240076 210810 240140
rect 217501 240138 217548 240140
rect 217456 240136 217548 240138
rect 217456 240080 217506 240136
rect 217456 240078 217548 240080
rect 217501 240076 217548 240078
rect 217612 240076 217618 240140
rect 218421 240138 218487 240141
rect 219198 240138 219204 240140
rect 218421 240136 219204 240138
rect 218421 240080 218426 240136
rect 218482 240080 219204 240136
rect 218421 240078 219204 240080
rect 210693 240075 210759 240076
rect 217501 240075 217567 240076
rect 218421 240075 218487 240078
rect 219198 240076 219204 240078
rect 219268 240076 219274 240140
rect 225781 240138 225847 240141
rect 226190 240138 226196 240140
rect 225781 240136 226196 240138
rect 225781 240080 225786 240136
rect 225842 240080 226196 240136
rect 225781 240078 226196 240080
rect 225781 240075 225847 240078
rect 226190 240076 226196 240078
rect 226260 240076 226266 240140
rect 230422 240076 230428 240140
rect 230492 240138 230498 240140
rect 230565 240138 230631 240141
rect 230492 240136 230631 240138
rect 230492 240080 230570 240136
rect 230626 240080 230631 240136
rect 230492 240078 230631 240080
rect 230492 240076 230498 240078
rect 230565 240075 230631 240078
rect 231894 240076 231900 240140
rect 231964 240138 231970 240140
rect 232589 240138 232655 240141
rect 231964 240136 232655 240138
rect 231964 240080 232594 240136
rect 232650 240080 232655 240136
rect 231964 240078 232655 240080
rect 231964 240076 231970 240078
rect 232589 240075 232655 240078
rect 237414 240076 237420 240140
rect 237484 240138 237490 240140
rect 237925 240138 237991 240141
rect 237484 240136 237991 240138
rect 237484 240080 237930 240136
rect 237986 240080 237991 240136
rect 237484 240078 237991 240080
rect 237484 240076 237490 240078
rect 237925 240075 237991 240078
rect 155217 240002 155283 240005
rect 155769 240002 155835 240005
rect 155217 240000 155835 240002
rect 155217 239944 155222 240000
rect 155278 239944 155774 240000
rect 155830 239944 155835 240000
rect 155217 239942 155835 239944
rect 155217 239939 155283 239942
rect 155769 239939 155835 239942
rect 200573 240002 200639 240005
rect 201401 240002 201467 240005
rect 203006 240002 203012 240004
rect 200573 240000 203012 240002
rect 200573 239944 200578 240000
rect 200634 239944 201406 240000
rect 201462 239944 203012 240000
rect 200573 239942 203012 239944
rect 200573 239939 200639 239942
rect 201401 239939 201467 239942
rect 203006 239940 203012 239942
rect 203076 239940 203082 240004
rect 215109 240002 215175 240005
rect 220854 240002 220860 240004
rect 215109 240000 220860 240002
rect 215109 239944 215114 240000
rect 215170 239944 220860 240000
rect 215109 239942 220860 239944
rect 215109 239939 215175 239942
rect 220854 239940 220860 239942
rect 220924 239940 220930 240004
rect 236821 240002 236887 240005
rect 260097 240002 260163 240005
rect 236821 240000 260163 240002
rect 236821 239944 236826 240000
rect 236882 239944 260102 240000
rect 260158 239944 260163 240000
rect 236821 239942 260163 239944
rect 236821 239939 236887 239942
rect 260097 239939 260163 239942
rect 110689 239866 110755 239869
rect 218973 239866 219039 239869
rect 219341 239866 219407 239869
rect 110689 239864 219407 239866
rect 110689 239808 110694 239864
rect 110750 239808 218978 239864
rect 219034 239808 219346 239864
rect 219402 239808 219407 239864
rect 110689 239806 219407 239808
rect 110689 239803 110755 239806
rect 218973 239803 219039 239806
rect 219341 239803 219407 239806
rect 68369 239594 68435 239597
rect 83641 239594 83707 239597
rect 68369 239592 83707 239594
rect 68369 239536 68374 239592
rect 68430 239536 83646 239592
rect 83702 239536 83707 239592
rect 68369 239534 83707 239536
rect 68369 239531 68435 239534
rect 83641 239531 83707 239534
rect 77017 239458 77083 239461
rect 111885 239458 111951 239461
rect 77017 239456 111951 239458
rect 77017 239400 77022 239456
rect 77078 239400 111890 239456
rect 111946 239400 111951 239456
rect 77017 239398 111951 239400
rect 77017 239395 77083 239398
rect 111885 239395 111951 239398
rect 115841 239458 115907 239461
rect 179413 239458 179479 239461
rect 115841 239456 179479 239458
rect 115841 239400 115846 239456
rect 115902 239400 179418 239456
rect 179474 239400 179479 239456
rect 115841 239398 179479 239400
rect 115841 239395 115907 239398
rect 179413 239395 179479 239398
rect 226926 239396 226932 239460
rect 226996 239458 227002 239460
rect 231853 239458 231919 239461
rect 226996 239456 231919 239458
rect 226996 239400 231858 239456
rect 231914 239400 231919 239456
rect 226996 239398 231919 239400
rect 226996 239396 227002 239398
rect 231853 239395 231919 239398
rect 242157 239322 242223 239325
rect 245929 239322 245995 239325
rect 242157 239320 245995 239322
rect 242157 239264 242162 239320
rect 242218 239264 245934 239320
rect 245990 239264 245995 239320
rect 242157 239262 245995 239264
rect 242157 239259 242223 239262
rect 245929 239259 245995 239262
rect 71681 238778 71747 238781
rect 76557 238778 76623 238781
rect 71681 238776 76623 238778
rect 71681 238720 71686 238776
rect 71742 238720 76562 238776
rect 76618 238720 76623 238776
rect 71681 238718 76623 238720
rect 71681 238715 71747 238718
rect 76557 238715 76623 238718
rect 234061 238778 234127 238781
rect 305085 238778 305151 238781
rect 234061 238776 305151 238778
rect 234061 238720 234066 238776
rect 234122 238720 305090 238776
rect 305146 238720 305151 238776
rect 234061 238718 305151 238720
rect 234061 238715 234127 238718
rect 305085 238715 305151 238718
rect 153377 238642 153443 238645
rect 156638 238642 156644 238644
rect 153377 238640 156644 238642
rect 153377 238584 153382 238640
rect 153438 238584 156644 238640
rect 153377 238582 156644 238584
rect 153377 238579 153443 238582
rect 156638 238580 156644 238582
rect 156708 238580 156714 238644
rect 205817 238642 205883 238645
rect 206870 238642 206876 238644
rect 205817 238640 206876 238642
rect 205817 238584 205822 238640
rect 205878 238584 206876 238640
rect 205817 238582 206876 238584
rect 205817 238579 205883 238582
rect 206870 238580 206876 238582
rect 206940 238580 206946 238644
rect 222326 238580 222332 238644
rect 222396 238642 222402 238644
rect 223389 238642 223455 238645
rect 222396 238640 223455 238642
rect 222396 238584 223394 238640
rect 223450 238584 223455 238640
rect 222396 238582 223455 238584
rect 222396 238580 222402 238582
rect 223389 238579 223455 238582
rect 243629 238642 243695 238645
rect 244038 238642 244044 238644
rect 243629 238640 244044 238642
rect 243629 238584 243634 238640
rect 243690 238584 244044 238640
rect 243629 238582 244044 238584
rect 243629 238579 243695 238582
rect 244038 238580 244044 238582
rect 244108 238580 244114 238644
rect 67725 238506 67791 238509
rect 178953 238506 179019 238509
rect 67725 238504 179019 238506
rect 67725 238448 67730 238504
rect 67786 238448 178958 238504
rect 179014 238448 179019 238504
rect 67725 238446 179019 238448
rect 67725 238443 67791 238446
rect 178953 238443 179019 238446
rect 179413 238506 179479 238509
rect 220997 238506 221063 238509
rect 179413 238504 221063 238506
rect 179413 238448 179418 238504
rect 179474 238448 221002 238504
rect 221058 238448 221063 238504
rect 179413 238446 221063 238448
rect 179413 238443 179479 238446
rect 220997 238443 221063 238446
rect 225045 238506 225111 238509
rect 242157 238506 242223 238509
rect 225045 238504 242223 238506
rect 225045 238448 225050 238504
rect 225106 238448 242162 238504
rect 242218 238448 242223 238504
rect 225045 238446 242223 238448
rect 225045 238443 225111 238446
rect 242157 238443 242223 238446
rect 220813 238370 220879 238373
rect 226977 238370 227043 238373
rect 220813 238368 227043 238370
rect 220813 238312 220818 238368
rect 220874 238312 226982 238368
rect 227038 238312 227043 238368
rect 220813 238310 227043 238312
rect 220813 238307 220879 238310
rect 226977 238307 227043 238310
rect 232773 238370 232839 238373
rect 295241 238370 295307 238373
rect 232773 238368 295307 238370
rect 232773 238312 232778 238368
rect 232834 238312 295246 238368
rect 295302 238312 295307 238368
rect 232773 238310 295307 238312
rect 232773 238307 232839 238310
rect 295241 238307 295307 238310
rect 92565 238234 92631 238237
rect 208301 238234 208367 238237
rect 92565 238232 208367 238234
rect 92565 238176 92570 238232
rect 92626 238176 208306 238232
rect 208362 238176 208367 238232
rect 92565 238174 208367 238176
rect 92565 238171 92631 238174
rect 208301 238171 208367 238174
rect 197169 237962 197235 237965
rect 202045 237962 202111 237965
rect 197169 237960 202111 237962
rect 197169 237904 197174 237960
rect 197230 237904 202050 237960
rect 202106 237904 202111 237960
rect 197169 237902 202111 237904
rect 197169 237899 197235 237902
rect 202045 237899 202111 237902
rect 240726 237492 240732 237556
rect 240796 237554 240802 237556
rect 241697 237554 241763 237557
rect 240796 237552 241763 237554
rect 240796 237496 241702 237552
rect 241758 237496 241763 237552
rect 240796 237494 241763 237496
rect 240796 237492 240802 237494
rect 241697 237491 241763 237494
rect 152733 237418 152799 237421
rect 154062 237418 154068 237420
rect 152733 237416 154068 237418
rect 152733 237360 152738 237416
rect 152794 237360 154068 237416
rect 152733 237358 154068 237360
rect 152733 237355 152799 237358
rect 154062 237356 154068 237358
rect 154132 237356 154138 237420
rect 166717 237418 166783 237421
rect 167729 237418 167795 237421
rect 166717 237416 167795 237418
rect 166717 237360 166722 237416
rect 166778 237360 167734 237416
rect 167790 237360 167795 237416
rect 166717 237358 167795 237360
rect 166717 237355 166783 237358
rect 167729 237355 167795 237358
rect 168230 237356 168236 237420
rect 168300 237418 168306 237420
rect 168373 237418 168439 237421
rect 168300 237416 168439 237418
rect 168300 237360 168378 237416
rect 168434 237360 168439 237416
rect 168300 237358 168439 237360
rect 168300 237356 168306 237358
rect 168373 237355 168439 237358
rect 196750 237356 196756 237420
rect 196820 237418 196826 237420
rect 197169 237418 197235 237421
rect 196820 237416 197235 237418
rect 196820 237360 197174 237416
rect 197230 237360 197235 237416
rect 196820 237358 197235 237360
rect 196820 237356 196826 237358
rect 197169 237355 197235 237358
rect 200205 237418 200271 237421
rect 200205 237416 201418 237418
rect 200205 237360 200210 237416
rect 200266 237360 201418 237416
rect 200205 237358 201418 237360
rect 200205 237355 200271 237358
rect 201358 237285 201418 237358
rect 209814 237356 209820 237420
rect 209884 237418 209890 237420
rect 210693 237418 210759 237421
rect 209884 237416 210759 237418
rect 209884 237360 210698 237416
rect 210754 237360 210759 237416
rect 209884 237358 210759 237360
rect 209884 237356 209890 237358
rect 210693 237355 210759 237358
rect 216673 237418 216739 237421
rect 217501 237418 217567 237421
rect 216673 237416 217567 237418
rect 216673 237360 216678 237416
rect 216734 237360 217506 237416
rect 217562 237360 217567 237416
rect 216673 237358 217567 237360
rect 216673 237355 216739 237358
rect 217501 237355 217567 237358
rect 218145 237418 218211 237421
rect 218421 237418 218487 237421
rect 218145 237416 218487 237418
rect 218145 237360 218150 237416
rect 218206 237360 218426 237416
rect 218482 237360 218487 237416
rect 218145 237358 218487 237360
rect 218145 237355 218211 237358
rect 218421 237355 218487 237358
rect 220997 237418 221063 237421
rect 221457 237418 221523 237421
rect 220997 237416 221523 237418
rect 220997 237360 221002 237416
rect 221058 237360 221462 237416
rect 221518 237360 221523 237416
rect 220997 237358 221523 237360
rect 220997 237355 221063 237358
rect 221457 237355 221523 237358
rect 225137 237418 225203 237421
rect 225781 237418 225847 237421
rect 225137 237416 225847 237418
rect 225137 237360 225142 237416
rect 225198 237360 225786 237416
rect 225842 237360 225847 237416
rect 225137 237358 225847 237360
rect 225137 237355 225203 237358
rect 225781 237355 225847 237358
rect 227529 237418 227595 237421
rect 227662 237418 227668 237420
rect 227529 237416 227668 237418
rect 227529 237360 227534 237416
rect 227590 237360 227668 237416
rect 227529 237358 227668 237360
rect 227529 237355 227595 237358
rect 227662 237356 227668 237358
rect 227732 237356 227738 237420
rect 241646 237356 241652 237420
rect 241716 237418 241722 237420
rect 241789 237418 241855 237421
rect 241716 237416 241855 237418
rect 241716 237360 241794 237416
rect 241850 237360 241855 237416
rect 241716 237358 241855 237360
rect 241716 237356 241722 237358
rect 241789 237355 241855 237358
rect 72734 237220 72740 237284
rect 72804 237282 72810 237284
rect 101949 237282 102015 237285
rect 72804 237280 102015 237282
rect 72804 237224 101954 237280
rect 102010 237224 102015 237280
rect 72804 237222 102015 237224
rect 72804 237220 72810 237222
rect 101949 237219 102015 237222
rect 102225 237282 102291 237285
rect 188838 237282 188844 237284
rect 102225 237280 188844 237282
rect 102225 237224 102230 237280
rect 102286 237224 188844 237280
rect 102225 237222 188844 237224
rect 102225 237219 102291 237222
rect 188838 237220 188844 237222
rect 188908 237282 188914 237284
rect 188908 237222 190470 237282
rect 188908 237220 188914 237222
rect 137277 237146 137343 237149
rect 167913 237146 167979 237149
rect 137277 237144 167979 237146
rect 137277 237088 137282 237144
rect 137338 237088 167918 237144
rect 167974 237088 167979 237144
rect 137277 237086 167979 237088
rect 137277 237083 137343 237086
rect 167913 237083 167979 237086
rect 190410 236738 190470 237222
rect 195094 237220 195100 237284
rect 195164 237282 195170 237284
rect 195164 237222 200130 237282
rect 201358 237280 201467 237285
rect 201358 237224 201406 237280
rect 201462 237224 201467 237280
rect 201358 237222 201467 237224
rect 195164 237220 195170 237222
rect 200070 237146 200130 237222
rect 201401 237219 201467 237222
rect 202781 237282 202847 237285
rect 208393 237282 208459 237285
rect 202781 237280 208459 237282
rect 202781 237224 202786 237280
rect 202842 237224 208398 237280
rect 208454 237224 208459 237280
rect 202781 237222 208459 237224
rect 202781 237219 202847 237222
rect 208393 237219 208459 237222
rect 219525 237282 219591 237285
rect 260925 237282 260991 237285
rect 219525 237280 260991 237282
rect 219525 237224 219530 237280
rect 219586 237224 260930 237280
rect 260986 237224 260991 237280
rect 219525 237222 260991 237224
rect 219525 237219 219591 237222
rect 260925 237219 260991 237222
rect 207657 237146 207723 237149
rect 200070 237144 207723 237146
rect 200070 237088 207662 237144
rect 207718 237088 207723 237144
rect 200070 237086 207723 237088
rect 207657 237083 207723 237086
rect 211654 237084 211660 237148
rect 211724 237146 211730 237148
rect 219433 237146 219499 237149
rect 211724 237144 219499 237146
rect 211724 237088 219438 237144
rect 219494 237088 219499 237144
rect 211724 237086 219499 237088
rect 211724 237084 211730 237086
rect 219433 237083 219499 237086
rect 199326 236948 199332 237012
rect 199396 237010 199402 237012
rect 203517 237010 203583 237013
rect 199396 237008 203583 237010
rect 199396 236952 203522 237008
rect 203578 236952 203583 237008
rect 199396 236950 203583 236952
rect 199396 236948 199402 236950
rect 203517 236947 203583 236950
rect 196617 236738 196683 236741
rect 190410 236736 196683 236738
rect 190410 236680 196622 236736
rect 196678 236680 196683 236736
rect 190410 236678 196683 236680
rect 196617 236675 196683 236678
rect 64597 236602 64663 236605
rect 193949 236602 194015 236605
rect 64597 236600 194015 236602
rect 64597 236544 64602 236600
rect 64658 236544 193954 236600
rect 194010 236544 194015 236600
rect 64597 236542 194015 236544
rect 64597 236539 64663 236542
rect 193949 236539 194015 236542
rect 220353 236602 220419 236605
rect 229829 236602 229895 236605
rect 220353 236600 229895 236602
rect 220353 236544 220358 236600
rect 220414 236544 229834 236600
rect 229890 236544 229895 236600
rect 220353 236542 229895 236544
rect 220353 236539 220419 236542
rect 229829 236539 229895 236542
rect 101397 236058 101463 236061
rect 101949 236058 102015 236061
rect 101397 236056 102015 236058
rect 101397 236000 101402 236056
rect 101458 236000 101954 236056
rect 102010 236000 102015 236056
rect 101397 235998 102015 236000
rect 101397 235995 101463 235998
rect 101949 235995 102015 235998
rect 211889 236058 211955 236061
rect 218646 236058 218652 236060
rect 211889 236056 218652 236058
rect 211889 236000 211894 236056
rect 211950 236000 218652 236056
rect 211889 235998 218652 236000
rect 211889 235995 211955 235998
rect 218646 235996 218652 235998
rect 218716 235996 218722 236060
rect 223757 236058 223823 236061
rect 224166 236058 224172 236060
rect 223757 236056 224172 236058
rect 223757 236000 223762 236056
rect 223818 236000 224172 236056
rect 223757 235998 224172 236000
rect 223757 235995 223823 235998
rect 224166 235996 224172 235998
rect 224236 235996 224242 236060
rect 229645 236058 229711 236061
rect 336089 236058 336155 236061
rect 229645 236056 336155 236058
rect 229645 236000 229650 236056
rect 229706 236000 336094 236056
rect 336150 236000 336155 236056
rect 229645 235998 336155 236000
rect 229645 235995 229711 235998
rect 336089 235995 336155 235998
rect 142245 235922 142311 235925
rect 153377 235922 153443 235925
rect 142245 235920 153443 235922
rect 142245 235864 142250 235920
rect 142306 235864 153382 235920
rect 153438 235864 153443 235920
rect 142245 235862 153443 235864
rect 142245 235859 142311 235862
rect 153377 235859 153443 235862
rect 153561 235922 153627 235925
rect 166206 235922 166212 235924
rect 153561 235920 166212 235922
rect 153561 235864 153566 235920
rect 153622 235864 166212 235920
rect 153561 235862 166212 235864
rect 153561 235859 153627 235862
rect 166206 235860 166212 235862
rect 166276 235860 166282 235924
rect 67265 235786 67331 235789
rect 152365 235786 152431 235789
rect 67265 235784 152431 235786
rect 67265 235728 67270 235784
rect 67326 235728 152370 235784
rect 152426 235728 152431 235784
rect 67265 235726 152431 235728
rect 67265 235723 67331 235726
rect 152365 235723 152431 235726
rect 152917 235786 152983 235789
rect 156454 235786 156460 235788
rect 152917 235784 156460 235786
rect 152917 235728 152922 235784
rect 152978 235728 156460 235784
rect 152917 235726 156460 235728
rect 152917 235723 152983 235726
rect 156454 235724 156460 235726
rect 156524 235724 156530 235788
rect 180190 235724 180196 235788
rect 180260 235786 180266 235788
rect 215293 235786 215359 235789
rect 180260 235784 215359 235786
rect 180260 235728 215298 235784
rect 215354 235728 215359 235784
rect 180260 235726 215359 235728
rect 180260 235724 180266 235726
rect 215293 235723 215359 235726
rect 150617 235650 150683 235653
rect 240317 235650 240383 235653
rect 150617 235648 240383 235650
rect 150617 235592 150622 235648
rect 150678 235592 240322 235648
rect 240378 235592 240383 235648
rect 150617 235590 240383 235592
rect 150617 235587 150683 235590
rect 240317 235587 240383 235590
rect 211245 235514 211311 235517
rect 212441 235514 212507 235517
rect 213126 235514 213132 235516
rect 211245 235512 213132 235514
rect 211245 235456 211250 235512
rect 211306 235456 212446 235512
rect 212502 235456 213132 235512
rect 211245 235454 213132 235456
rect 211245 235451 211311 235454
rect 212441 235451 212507 235454
rect 213126 235452 213132 235454
rect 213196 235452 213202 235516
rect 240685 235378 240751 235381
rect 331949 235378 332015 235381
rect 240685 235376 332015 235378
rect 240685 235320 240690 235376
rect 240746 235320 331954 235376
rect 332010 235320 332015 235376
rect 240685 235318 332015 235320
rect 240685 235315 240751 235318
rect 331949 235315 332015 235318
rect 107745 235242 107811 235245
rect 140773 235242 140839 235245
rect 107745 235240 140839 235242
rect 107745 235184 107750 235240
rect 107806 235184 140778 235240
rect 140834 235184 140839 235240
rect 107745 235182 140839 235184
rect 107745 235179 107811 235182
rect 140773 235179 140839 235182
rect 155953 235242 156019 235245
rect 205633 235242 205699 235245
rect 155953 235240 205699 235242
rect 155953 235184 155958 235240
rect 156014 235184 205638 235240
rect 205694 235184 205699 235240
rect 155953 235182 205699 235184
rect 155953 235179 156019 235182
rect 205633 235179 205699 235182
rect 215293 235242 215359 235245
rect 216581 235242 216647 235245
rect 342989 235242 343055 235245
rect 215293 235240 343055 235242
rect 215293 235184 215298 235240
rect 215354 235184 216586 235240
rect 216642 235184 342994 235240
rect 343050 235184 343055 235240
rect 215293 235182 343055 235184
rect 215293 235179 215359 235182
rect 216581 235179 216647 235182
rect 342989 235179 343055 235182
rect 220077 234698 220143 234701
rect 223614 234698 223620 234700
rect 220077 234696 223620 234698
rect 220077 234640 220082 234696
rect 220138 234640 223620 234696
rect 220077 234638 223620 234640
rect 220077 234635 220143 234638
rect 223614 234636 223620 234638
rect 223684 234636 223690 234700
rect 224217 234698 224283 234701
rect 582833 234698 582899 234701
rect 224217 234696 582899 234698
rect 224217 234640 224222 234696
rect 224278 234640 582838 234696
rect 582894 234640 582899 234696
rect 224217 234638 582899 234640
rect 224217 234635 224283 234638
rect 582833 234635 582899 234638
rect 74625 234562 74691 234565
rect 155493 234562 155559 234565
rect 74625 234560 155559 234562
rect 74625 234504 74630 234560
rect 74686 234504 155498 234560
rect 155554 234504 155559 234560
rect 74625 234502 155559 234504
rect 74625 234499 74691 234502
rect 155493 234499 155559 234502
rect 155677 234562 155743 234565
rect 163681 234562 163747 234565
rect 155677 234560 163747 234562
rect 155677 234504 155682 234560
rect 155738 234504 163686 234560
rect 163742 234504 163747 234560
rect 155677 234502 163747 234504
rect 155677 234499 155743 234502
rect 163681 234499 163747 234502
rect 192661 234562 192727 234565
rect 242934 234562 242940 234564
rect 192661 234560 242940 234562
rect 192661 234504 192666 234560
rect 192722 234504 242940 234560
rect 192661 234502 242940 234504
rect 192661 234499 192727 234502
rect 242934 234500 242940 234502
rect 243004 234500 243010 234564
rect 82670 234364 82676 234428
rect 82740 234426 82746 234428
rect 103605 234426 103671 234429
rect 82740 234424 103671 234426
rect 82740 234368 103610 234424
rect 103666 234368 103671 234424
rect 82740 234366 103671 234368
rect 82740 234364 82746 234366
rect 103605 234363 103671 234366
rect 129825 234426 129891 234429
rect 177297 234426 177363 234429
rect 129825 234424 177363 234426
rect 129825 234368 129830 234424
rect 129886 234368 177302 234424
rect 177358 234368 177363 234424
rect 129825 234366 177363 234368
rect 129825 234363 129891 234366
rect 177297 234363 177363 234366
rect 182081 234426 182147 234429
rect 226149 234426 226215 234429
rect 182081 234424 226215 234426
rect 182081 234368 182086 234424
rect 182142 234368 226154 234424
rect 226210 234368 226215 234424
rect 182081 234366 226215 234368
rect 182081 234363 182147 234366
rect 226149 234363 226215 234366
rect 140773 234290 140839 234293
rect 162485 234290 162551 234293
rect 140773 234288 162551 234290
rect 140773 234232 140778 234288
rect 140834 234232 162490 234288
rect 162546 234232 162551 234288
rect 140773 234230 162551 234232
rect 140773 234227 140839 234230
rect 162485 234227 162551 234230
rect 176653 234290 176719 234293
rect 177941 234290 178007 234293
rect 201585 234290 201651 234293
rect 202413 234290 202479 234293
rect 176653 234288 202479 234290
rect 176653 234232 176658 234288
rect 176714 234232 177946 234288
rect 178002 234232 201590 234288
rect 201646 234232 202418 234288
rect 202474 234232 202479 234288
rect 176653 234230 202479 234232
rect 176653 234227 176719 234230
rect 177941 234227 178007 234230
rect 201585 234227 201651 234230
rect 202413 234227 202479 234230
rect 201493 233882 201559 233885
rect 202229 233882 202295 233885
rect 201493 233880 202295 233882
rect 201493 233824 201498 233880
rect 201554 233824 202234 233880
rect 202290 233824 202295 233880
rect 201493 233822 202295 233824
rect 201493 233819 201559 233822
rect 202229 233819 202295 233822
rect 162209 233746 162275 233749
rect 162761 233746 162827 233749
rect 162209 233744 162827 233746
rect 162209 233688 162214 233744
rect 162270 233688 162766 233744
rect 162822 233688 162827 233744
rect 162209 233686 162827 233688
rect 162209 233683 162275 233686
rect 162761 233683 162827 233686
rect 162761 233338 162827 233341
rect 182081 233338 182147 233341
rect 162761 233336 182147 233338
rect 162761 233280 162766 233336
rect 162822 233280 182086 233336
rect 182142 233280 182147 233336
rect 162761 233278 182147 233280
rect 162761 233275 162827 233278
rect 182081 233275 182147 233278
rect 227069 233338 227135 233341
rect 227621 233338 227687 233341
rect 416773 233338 416839 233341
rect 227069 233336 416839 233338
rect 227069 233280 227074 233336
rect 227130 233280 227626 233336
rect 227682 233280 416778 233336
rect 416834 233280 416839 233336
rect 227069 233278 416839 233280
rect 227069 233275 227135 233278
rect 227621 233275 227687 233278
rect 416773 233275 416839 233278
rect 60457 233202 60523 233205
rect 158713 233202 158779 233205
rect 60457 233200 158779 233202
rect 60457 233144 60462 233200
rect 60518 233144 158718 233200
rect 158774 233144 158779 233200
rect 60457 233142 158779 233144
rect 60457 233139 60523 233142
rect 158713 233139 158779 233142
rect 184289 233202 184355 233205
rect 184606 233202 184612 233204
rect 184289 233200 184612 233202
rect 184289 233144 184294 233200
rect 184350 233144 184612 233200
rect 184289 233142 184612 233144
rect 184289 233139 184355 233142
rect 184606 233140 184612 233142
rect 184676 233140 184682 233204
rect 187417 233202 187483 233205
rect 187550 233202 187556 233204
rect 187417 233200 187556 233202
rect 187417 233144 187422 233200
rect 187478 233144 187556 233200
rect 187417 233142 187556 233144
rect 187417 233139 187483 233142
rect 187550 233140 187556 233142
rect 187620 233140 187626 233204
rect 227713 233202 227779 233205
rect 355317 233202 355383 233205
rect 227713 233200 355383 233202
rect 227713 233144 227718 233200
rect 227774 233144 355322 233200
rect 355378 233144 355383 233200
rect 227713 233142 355383 233144
rect 227713 233139 227779 233142
rect 355317 233139 355383 233142
rect 91185 233066 91251 233069
rect 157333 233066 157399 233069
rect 91185 233064 157399 233066
rect 91185 233008 91190 233064
rect 91246 233008 157338 233064
rect 157394 233008 157399 233064
rect 91185 233006 157399 233008
rect 91185 233003 91251 233006
rect 157333 233003 157399 233006
rect 182817 233066 182883 233069
rect 243629 233066 243695 233069
rect 182817 233064 243695 233066
rect 182817 233008 182822 233064
rect 182878 233008 243634 233064
rect 243690 233008 243695 233064
rect 182817 233006 243695 233008
rect 182817 233003 182883 233006
rect 243629 233003 243695 233006
rect 135437 232930 135503 232933
rect 168230 232930 168236 232932
rect 135437 232928 168236 232930
rect 135437 232872 135442 232928
rect 135498 232872 168236 232928
rect 135437 232870 168236 232872
rect 135437 232867 135503 232870
rect 168230 232868 168236 232870
rect 168300 232868 168306 232932
rect 178861 232930 178927 232933
rect 228173 232930 228239 232933
rect 178861 232928 228239 232930
rect 178861 232872 178866 232928
rect 178922 232872 228178 232928
rect 228234 232872 228239 232928
rect 178861 232870 228239 232872
rect 178861 232867 178927 232870
rect 228173 232867 228239 232870
rect 238845 232930 238911 232933
rect 239397 232930 239463 232933
rect 238845 232928 239463 232930
rect 238845 232872 238850 232928
rect 238906 232872 239402 232928
rect 239458 232872 239463 232928
rect 238845 232870 239463 232872
rect 238845 232867 238911 232870
rect 239397 232867 239463 232870
rect 159173 232794 159239 232797
rect 159357 232794 159423 232797
rect 229645 232794 229711 232797
rect 159173 232792 229711 232794
rect 159173 232736 159178 232792
rect 159234 232736 159362 232792
rect 159418 232736 229650 232792
rect 229706 232736 229711 232792
rect 159173 232734 229711 232736
rect 159173 232731 159239 232734
rect 159357 232731 159423 232734
rect 229645 232731 229711 232734
rect 583293 232386 583359 232389
rect 583520 232386 584960 232476
rect 583293 232384 584960 232386
rect 583293 232328 583298 232384
rect 583354 232328 584960 232384
rect 583293 232326 584960 232328
rect 583293 232323 583359 232326
rect 583520 232236 584960 232326
rect 239397 231978 239463 231981
rect 297357 231978 297423 231981
rect 239397 231976 297423 231978
rect 239397 231920 239402 231976
rect 239458 231920 297362 231976
rect 297418 231920 297423 231976
rect 239397 231918 297423 231920
rect 239397 231915 239463 231918
rect 297357 231915 297423 231918
rect 63309 231842 63375 231845
rect 188429 231842 188495 231845
rect 188613 231842 188679 231845
rect 63309 231840 188679 231842
rect 63309 231784 63314 231840
rect 63370 231784 188434 231840
rect 188490 231784 188618 231840
rect 188674 231784 188679 231840
rect 63309 231782 188679 231784
rect 63309 231779 63375 231782
rect 188429 231779 188495 231782
rect 188613 231779 188679 231782
rect 214189 231842 214255 231845
rect 254117 231842 254183 231845
rect 214189 231840 254183 231842
rect 214189 231784 214194 231840
rect 214250 231784 254122 231840
rect 254178 231784 254183 231840
rect 214189 231782 254183 231784
rect 214189 231779 214255 231782
rect 254117 231779 254183 231782
rect 139577 231706 139643 231709
rect 155309 231706 155375 231709
rect 139577 231704 155375 231706
rect 139577 231648 139582 231704
rect 139638 231648 155314 231704
rect 155370 231648 155375 231704
rect 139577 231646 155375 231648
rect 139577 231643 139643 231646
rect 155309 231643 155375 231646
rect 155769 231706 155835 231709
rect 230565 231706 230631 231709
rect 234654 231706 234660 231708
rect 155769 231704 219450 231706
rect 155769 231648 155774 231704
rect 155830 231648 219450 231704
rect 155769 231646 219450 231648
rect 155769 231643 155835 231646
rect 147489 231570 147555 231573
rect 167637 231570 167703 231573
rect 147489 231568 167703 231570
rect 147489 231512 147494 231568
rect 147550 231512 167642 231568
rect 167698 231512 167703 231568
rect 147489 231510 167703 231512
rect 147489 231507 147555 231510
rect 167637 231507 167703 231510
rect 195237 231298 195303 231301
rect 215293 231298 215359 231301
rect 195237 231296 215359 231298
rect 195237 231240 195242 231296
rect 195298 231240 215298 231296
rect 215354 231240 215359 231296
rect 195237 231238 215359 231240
rect 219390 231298 219450 231646
rect 230565 231704 234660 231706
rect 230565 231648 230570 231704
rect 230626 231648 234660 231704
rect 230565 231646 234660 231648
rect 230565 231643 230631 231646
rect 234654 231644 234660 231646
rect 234724 231644 234730 231708
rect 238293 231298 238359 231301
rect 269849 231298 269915 231301
rect 219390 231296 269915 231298
rect 219390 231240 238298 231296
rect 238354 231240 269854 231296
rect 269910 231240 269915 231296
rect 219390 231238 269915 231240
rect 195237 231235 195303 231238
rect 215293 231235 215359 231238
rect 238293 231235 238359 231238
rect 269849 231235 269915 231238
rect 168230 231100 168236 231164
rect 168300 231162 168306 231164
rect 195646 231162 195652 231164
rect 168300 231102 195652 231162
rect 168300 231100 168306 231102
rect 195646 231100 195652 231102
rect 195716 231162 195722 231164
rect 202873 231162 202939 231165
rect 195716 231160 202939 231162
rect 195716 231104 202878 231160
rect 202934 231104 202939 231160
rect 195716 231102 202939 231104
rect 195716 231100 195722 231102
rect 202873 231099 202939 231102
rect 254117 231162 254183 231165
rect 313457 231162 313523 231165
rect 254117 231160 313523 231162
rect 254117 231104 254122 231160
rect 254178 231104 313462 231160
rect 313518 231104 313523 231160
rect 254117 231102 313523 231104
rect 254117 231099 254183 231102
rect 313457 231099 313523 231102
rect 182081 230482 182147 230485
rect 240685 230482 240751 230485
rect 182081 230480 240751 230482
rect 182081 230424 182086 230480
rect 182142 230424 240690 230480
rect 240746 230424 240751 230480
rect 182081 230422 240751 230424
rect 182081 230419 182147 230422
rect 240685 230419 240751 230422
rect 110321 230346 110387 230349
rect 163589 230346 163655 230349
rect 185342 230346 185348 230348
rect 110321 230344 163655 230346
rect 110321 230288 110326 230344
rect 110382 230288 163594 230344
rect 163650 230288 163655 230344
rect 110321 230286 163655 230288
rect 110321 230283 110387 230286
rect 163589 230283 163655 230286
rect 180750 230286 185348 230346
rect 59077 230210 59143 230213
rect 180750 230210 180810 230286
rect 185342 230284 185348 230286
rect 185412 230346 185418 230348
rect 185577 230346 185643 230349
rect 185412 230344 185643 230346
rect 185412 230288 185582 230344
rect 185638 230288 185643 230344
rect 185412 230286 185643 230288
rect 185412 230284 185418 230286
rect 185577 230283 185643 230286
rect 59077 230208 180810 230210
rect 59077 230152 59082 230208
rect 59138 230152 180810 230208
rect 59077 230150 180810 230152
rect 59077 230147 59143 230150
rect 190269 229938 190335 229941
rect 201493 229938 201559 229941
rect 190269 229936 201559 229938
rect 190269 229880 190274 229936
rect 190330 229880 201498 229936
rect 201554 229880 201559 229936
rect 190269 229878 201559 229880
rect 190269 229875 190335 229878
rect 201493 229875 201559 229878
rect 173433 229802 173499 229805
rect 194409 229802 194475 229805
rect 173433 229800 194475 229802
rect 173433 229744 173438 229800
rect 173494 229744 194414 229800
rect 194470 229744 194475 229800
rect 173433 229742 194475 229744
rect 173433 229739 173499 229742
rect 194409 229739 194475 229742
rect 195830 229740 195836 229804
rect 195900 229802 195906 229804
rect 448513 229802 448579 229805
rect 195900 229800 448579 229802
rect 195900 229744 448518 229800
rect 448574 229744 448579 229800
rect 195900 229742 448579 229744
rect 195900 229740 195906 229742
rect 448513 229739 448579 229742
rect 209681 229122 209747 229125
rect 371969 229122 372035 229125
rect 209681 229120 372035 229122
rect 209681 229064 209686 229120
rect 209742 229064 371974 229120
rect 372030 229064 372035 229120
rect 209681 229062 372035 229064
rect 209681 229059 209747 229062
rect 371969 229059 372035 229062
rect 65885 228986 65951 228989
rect 164877 228986 164943 228989
rect 65885 228984 164943 228986
rect 65885 228928 65890 228984
rect 65946 228928 164882 228984
rect 164938 228928 164943 228984
rect 65885 228926 164943 228928
rect 65885 228923 65951 228926
rect 164877 228923 164943 228926
rect 180006 228924 180012 228988
rect 180076 228986 180082 228988
rect 209037 228986 209103 228989
rect 180076 228984 209103 228986
rect 180076 228928 209042 228984
rect 209098 228928 209103 228984
rect 180076 228926 209103 228928
rect 180076 228924 180082 228926
rect 209037 228923 209103 228926
rect 231485 228986 231551 228989
rect 327073 228986 327139 228989
rect 231485 228984 327139 228986
rect 231485 228928 231490 228984
rect 231546 228928 327078 228984
rect 327134 228928 327139 228984
rect 231485 228926 327139 228928
rect 231485 228923 231551 228926
rect 327073 228923 327139 228926
rect 136541 228850 136607 228853
rect 184790 228850 184796 228852
rect 136541 228848 184796 228850
rect 136541 228792 136546 228848
rect 136602 228792 184796 228848
rect 136541 228790 184796 228792
rect 136541 228787 136607 228790
rect 184790 228788 184796 228790
rect 184860 228788 184866 228852
rect 194409 228442 194475 228445
rect 204161 228442 204227 228445
rect 194409 228440 204227 228442
rect 194409 228384 194414 228440
rect 194470 228384 204166 228440
rect 204222 228384 204227 228440
rect 194409 228382 204227 228384
rect 194409 228379 194475 228382
rect 204161 228379 204227 228382
rect 207565 228442 207631 228445
rect 232589 228442 232655 228445
rect 207565 228440 232655 228442
rect 207565 228384 207570 228440
rect 207626 228384 232594 228440
rect 232650 228384 232655 228440
rect 207565 228382 232655 228384
rect 207565 228379 207631 228382
rect 232589 228379 232655 228382
rect 61837 228306 61903 228309
rect 183461 228306 183527 228309
rect 61837 228304 183527 228306
rect 61837 228248 61842 228304
rect 61898 228248 183466 228304
rect 183522 228248 183527 228304
rect 61837 228246 183527 228248
rect 61837 228243 61903 228246
rect 183461 228243 183527 228246
rect 184790 228244 184796 228308
rect 184860 228306 184866 228308
rect 316677 228306 316743 228309
rect 184860 228304 316743 228306
rect 184860 228248 316682 228304
rect 316738 228248 316743 228304
rect 184860 228246 316743 228248
rect 184860 228244 184866 228246
rect 316677 228243 316743 228246
rect -960 227884 480 228124
rect 57789 227626 57855 227629
rect 138013 227626 138079 227629
rect 57789 227624 138079 227626
rect 57789 227568 57794 227624
rect 57850 227568 138018 227624
rect 138074 227568 138079 227624
rect 57789 227566 138079 227568
rect 57789 227563 57855 227566
rect 138013 227563 138079 227566
rect 146109 227626 146175 227629
rect 220353 227626 220419 227629
rect 146109 227624 220419 227626
rect 146109 227568 146114 227624
rect 146170 227568 220358 227624
rect 220414 227568 220419 227624
rect 146109 227566 220419 227568
rect 146109 227563 146175 227566
rect 220353 227563 220419 227566
rect 235349 227626 235415 227629
rect 271873 227626 271939 227629
rect 235349 227624 271939 227626
rect 235349 227568 235354 227624
rect 235410 227568 271878 227624
rect 271934 227568 271939 227624
rect 235349 227566 271939 227568
rect 235349 227563 235415 227566
rect 271873 227563 271939 227566
rect 91001 227490 91067 227493
rect 157926 227490 157932 227492
rect 91001 227488 157932 227490
rect 91001 227432 91006 227488
rect 91062 227432 157932 227488
rect 91001 227430 157932 227432
rect 91001 227427 91067 227430
rect 157926 227428 157932 227430
rect 157996 227428 158002 227492
rect 193857 227490 193923 227493
rect 240777 227490 240843 227493
rect 193857 227488 240843 227490
rect 193857 227432 193862 227488
rect 193918 227432 240782 227488
rect 240838 227432 240843 227488
rect 193857 227430 240843 227432
rect 193857 227427 193923 227430
rect 240777 227427 240843 227430
rect 139485 227354 139551 227357
rect 171133 227354 171199 227357
rect 172053 227354 172119 227357
rect 139485 227352 172119 227354
rect 139485 227296 139490 227352
rect 139546 227296 171138 227352
rect 171194 227296 172058 227352
rect 172114 227296 172119 227352
rect 139485 227294 172119 227296
rect 139485 227291 139551 227294
rect 171133 227291 171199 227294
rect 172053 227291 172119 227294
rect 176009 227354 176075 227357
rect 204437 227354 204503 227357
rect 176009 227352 204503 227354
rect 176009 227296 176014 227352
rect 176070 227296 204442 227352
rect 204498 227296 204503 227352
rect 176009 227294 204503 227296
rect 176009 227291 176075 227294
rect 204437 227291 204503 227294
rect 242750 226884 242756 226948
rect 242820 226946 242826 226948
rect 262305 226946 262371 226949
rect 242820 226944 262371 226946
rect 242820 226888 262310 226944
rect 262366 226888 262371 226944
rect 242820 226886 262371 226888
rect 242820 226884 242826 226886
rect 262305 226883 262371 226886
rect 271873 226946 271939 226949
rect 363689 226946 363755 226949
rect 271873 226944 363755 226946
rect 271873 226888 271878 226944
rect 271934 226888 363694 226944
rect 363750 226888 363755 226944
rect 271873 226886 363755 226888
rect 271873 226883 271939 226886
rect 363689 226883 363755 226886
rect 89805 226402 89871 226405
rect 91001 226402 91067 226405
rect 89805 226400 91067 226402
rect 89805 226344 89810 226400
rect 89866 226344 91006 226400
rect 91062 226344 91067 226400
rect 89805 226342 91067 226344
rect 89805 226339 89871 226342
rect 91001 226339 91067 226342
rect 204437 226402 204503 226405
rect 204846 226402 204852 226404
rect 204437 226400 204852 226402
rect 204437 226344 204442 226400
rect 204498 226344 204852 226400
rect 204437 226342 204852 226344
rect 204437 226339 204503 226342
rect 204846 226340 204852 226342
rect 204916 226340 204922 226404
rect 220169 226402 220235 226405
rect 227069 226402 227135 226405
rect 220169 226400 227135 226402
rect 220169 226344 220174 226400
rect 220230 226344 227074 226400
rect 227130 226344 227135 226400
rect 220169 226342 227135 226344
rect 220169 226339 220235 226342
rect 227069 226339 227135 226342
rect 101397 226266 101463 226269
rect 232773 226266 232839 226269
rect 101397 226264 232839 226266
rect 101397 226208 101402 226264
rect 101458 226208 232778 226264
rect 232834 226208 232839 226264
rect 101397 226206 232839 226208
rect 101397 226203 101463 226206
rect 232773 226203 232839 226206
rect 86861 226130 86927 226133
rect 160921 226130 160987 226133
rect 86861 226128 160987 226130
rect 86861 226072 86866 226128
rect 86922 226072 160926 226128
rect 160982 226072 160987 226128
rect 86861 226070 160987 226072
rect 86861 226067 86927 226070
rect 160921 226067 160987 226070
rect 183461 226130 183527 226133
rect 244365 226130 244431 226133
rect 183461 226128 244431 226130
rect 183461 226072 183466 226128
rect 183522 226072 244370 226128
rect 244426 226072 244431 226128
rect 183461 226070 244431 226072
rect 183461 226067 183527 226070
rect 244365 226067 244431 226070
rect 115197 225994 115263 225997
rect 180057 225994 180123 225997
rect 115197 225992 180123 225994
rect 115197 225936 115202 225992
rect 115258 225936 180062 225992
rect 180118 225936 180123 225992
rect 115197 225934 180123 225936
rect 115197 225931 115263 225934
rect 180057 225931 180123 225934
rect 204161 225994 204227 225997
rect 242801 225994 242867 225997
rect 204161 225992 242867 225994
rect 204161 225936 204166 225992
rect 204222 225936 242806 225992
rect 242862 225936 242867 225992
rect 204161 225934 242867 225936
rect 204161 225931 204227 225934
rect 242801 225931 242867 225934
rect 274081 225586 274147 225589
rect 283782 225586 283788 225588
rect 274081 225584 283788 225586
rect 274081 225528 274086 225584
rect 274142 225528 283788 225584
rect 274081 225526 283788 225528
rect 274081 225523 274147 225526
rect 283782 225524 283788 225526
rect 283852 225524 283858 225588
rect 244365 225316 244431 225317
rect 244365 225314 244412 225316
rect 244320 225312 244412 225314
rect 244320 225256 244370 225312
rect 244320 225254 244412 225256
rect 244365 225252 244412 225254
rect 244476 225252 244482 225316
rect 244365 225251 244431 225252
rect 244365 225178 244431 225181
rect 244774 225178 244780 225180
rect 244365 225176 244780 225178
rect 244365 225120 244370 225176
rect 244426 225120 244780 225176
rect 244365 225118 244780 225120
rect 244365 225115 244431 225118
rect 244774 225116 244780 225118
rect 244844 225116 244850 225180
rect 85665 225042 85731 225045
rect 86861 225042 86927 225045
rect 85665 225040 86927 225042
rect 85665 224984 85670 225040
rect 85726 224984 86866 225040
rect 86922 224984 86927 225040
rect 85665 224982 86927 224984
rect 85665 224979 85731 224982
rect 86861 224979 86927 224982
rect 196566 224980 196572 225044
rect 196636 225042 196642 225044
rect 198733 225042 198799 225045
rect 196636 225040 198799 225042
rect 196636 224984 198738 225040
rect 198794 224984 198799 225040
rect 196636 224982 198799 224984
rect 196636 224980 196642 224982
rect 198733 224979 198799 224982
rect 232497 225042 232563 225045
rect 434713 225042 434779 225045
rect 232497 225040 434779 225042
rect 232497 224984 232502 225040
rect 232558 224984 434718 225040
rect 434774 224984 434779 225040
rect 232497 224982 434779 224984
rect 232497 224979 232563 224982
rect 434713 224979 434779 224982
rect 67357 224906 67423 224909
rect 242750 224906 242756 224908
rect 67357 224904 242756 224906
rect 67357 224848 67362 224904
rect 67418 224848 242756 224904
rect 67357 224846 242756 224848
rect 67357 224843 67423 224846
rect 242750 224844 242756 224846
rect 242820 224844 242826 224908
rect 81249 224770 81315 224773
rect 157333 224770 157399 224773
rect 81249 224768 157399 224770
rect 81249 224712 81254 224768
rect 81310 224712 157338 224768
rect 157394 224712 157399 224768
rect 81249 224710 157399 224712
rect 81249 224707 81315 224710
rect 157333 224707 157399 224710
rect 135161 224362 135227 224365
rect 177941 224362 178007 224365
rect 178534 224362 178540 224364
rect 135161 224360 178540 224362
rect 135161 224304 135166 224360
rect 135222 224304 177946 224360
rect 178002 224304 178540 224360
rect 135161 224302 178540 224304
rect 135161 224299 135227 224302
rect 177941 224299 178007 224302
rect 178534 224300 178540 224302
rect 178604 224300 178610 224364
rect 160001 224226 160067 224229
rect 407205 224226 407271 224229
rect 160001 224224 407271 224226
rect 160001 224168 160006 224224
rect 160062 224168 407210 224224
rect 407266 224168 407271 224224
rect 160001 224166 407271 224168
rect 160001 224163 160067 224166
rect 407205 224163 407271 224166
rect 178033 223682 178099 223685
rect 307109 223682 307175 223685
rect 178033 223680 307175 223682
rect 178033 223624 178038 223680
rect 178094 223624 307114 223680
rect 307170 223624 307175 223680
rect 178033 223622 307175 223624
rect 178033 223619 178099 223622
rect 307109 223619 307175 223622
rect 52177 223546 52243 223549
rect 133137 223546 133203 223549
rect 52177 223544 133203 223546
rect 52177 223488 52182 223544
rect 52238 223488 133142 223544
rect 133198 223488 133203 223544
rect 52177 223486 133203 223488
rect 52177 223483 52243 223486
rect 133137 223483 133203 223486
rect 146201 223546 146267 223549
rect 238109 223546 238175 223549
rect 146201 223544 238175 223546
rect 146201 223488 146206 223544
rect 146262 223488 238114 223544
rect 238170 223488 238175 223544
rect 146201 223486 238175 223488
rect 146201 223483 146267 223486
rect 238109 223483 238175 223486
rect 76557 223410 76623 223413
rect 155217 223410 155283 223413
rect 76557 223408 155283 223410
rect 76557 223352 76562 223408
rect 76618 223352 155222 223408
rect 155278 223352 155283 223408
rect 76557 223350 155283 223352
rect 76557 223347 76623 223350
rect 155217 223347 155283 223350
rect 177389 223410 177455 223413
rect 240041 223410 240107 223413
rect 246297 223410 246363 223413
rect 177389 223408 246363 223410
rect 177389 223352 177394 223408
rect 177450 223352 240046 223408
rect 240102 223352 246302 223408
rect 246358 223352 246363 223408
rect 177389 223350 246363 223352
rect 177389 223347 177455 223350
rect 240041 223347 240107 223350
rect 246297 223347 246363 223350
rect 133689 223274 133755 223277
rect 163497 223274 163563 223277
rect 133689 223272 163563 223274
rect 133689 223216 133694 223272
rect 133750 223216 163502 223272
rect 163558 223216 163563 223272
rect 133689 223214 163563 223216
rect 133689 223211 133755 223214
rect 163497 223211 163563 223214
rect 187509 222866 187575 222869
rect 429193 222866 429259 222869
rect 187509 222864 429259 222866
rect 187509 222808 187514 222864
rect 187570 222808 429198 222864
rect 429254 222808 429259 222864
rect 187509 222806 429259 222808
rect 187509 222803 187575 222806
rect 429193 222803 429259 222806
rect 60549 222186 60615 222189
rect 259545 222186 259611 222189
rect 260741 222186 260807 222189
rect 60549 222184 260807 222186
rect 60549 222128 60554 222184
rect 60610 222128 259550 222184
rect 259606 222128 260746 222184
rect 260802 222128 260807 222184
rect 60549 222126 260807 222128
rect 60549 222123 60615 222126
rect 259545 222123 259611 222126
rect 260741 222123 260807 222126
rect 89529 222050 89595 222053
rect 248597 222052 248663 222053
rect 89529 222048 190470 222050
rect 89529 221992 89534 222048
rect 89590 221992 190470 222048
rect 89529 221990 190470 221992
rect 89529 221987 89595 221990
rect 138013 221914 138079 221917
rect 189809 221914 189875 221917
rect 138013 221912 189875 221914
rect 138013 221856 138018 221912
rect 138074 221856 189814 221912
rect 189870 221856 189875 221912
rect 138013 221854 189875 221856
rect 138013 221851 138079 221854
rect 189809 221851 189875 221854
rect 190410 221506 190470 221990
rect 248597 222048 248644 222052
rect 248708 222050 248714 222052
rect 248597 221992 248602 222048
rect 248597 221988 248644 221992
rect 248708 221990 248754 222050
rect 248708 221988 248714 221990
rect 248597 221987 248663 221988
rect 191649 221506 191715 221509
rect 323669 221506 323735 221509
rect 190410 221504 323735 221506
rect 190410 221448 191654 221504
rect 191710 221448 323674 221504
rect 323730 221448 323735 221504
rect 190410 221446 323735 221448
rect 191649 221443 191715 221446
rect 323669 221443 323735 221446
rect 75177 220826 75243 220829
rect 239397 220826 239463 220829
rect 75177 220824 239463 220826
rect 75177 220768 75182 220824
rect 75238 220768 239402 220824
rect 239458 220768 239463 220824
rect 75177 220766 239463 220768
rect 75177 220763 75243 220766
rect 239397 220763 239463 220766
rect 86217 220690 86283 220693
rect 209773 220690 209839 220693
rect 210417 220690 210483 220693
rect 86217 220688 210483 220690
rect 86217 220632 86222 220688
rect 86278 220632 209778 220688
rect 209834 220632 210422 220688
rect 210478 220632 210483 220688
rect 86217 220630 210483 220632
rect 86217 220627 86283 220630
rect 209773 220627 209839 220630
rect 210417 220627 210483 220630
rect 74533 220554 74599 220557
rect 166993 220554 167059 220557
rect 74533 220552 167059 220554
rect 74533 220496 74538 220552
rect 74594 220496 166998 220552
rect 167054 220496 167059 220552
rect 74533 220494 167059 220496
rect 74533 220491 74599 220494
rect 166993 220491 167059 220494
rect 210601 220146 210667 220149
rect 412633 220146 412699 220149
rect 210601 220144 412699 220146
rect 210601 220088 210606 220144
rect 210662 220088 412638 220144
rect 412694 220088 412699 220144
rect 210601 220086 412699 220088
rect 210601 220083 210667 220086
rect 412633 220083 412699 220086
rect 216029 219466 216095 219469
rect 276841 219466 276907 219469
rect 216029 219464 276907 219466
rect 216029 219408 216034 219464
rect 216090 219408 276846 219464
rect 276902 219408 276907 219464
rect 216029 219406 276907 219408
rect 216029 219403 216095 219406
rect 276841 219403 276907 219406
rect 64781 219330 64847 219333
rect 244365 219330 244431 219333
rect 64781 219328 244431 219330
rect 64781 219272 64786 219328
rect 64842 219272 244370 219328
rect 244426 219272 244431 219328
rect 64781 219270 244431 219272
rect 64781 219267 64847 219270
rect 244365 219267 244431 219270
rect 128353 219194 128419 219197
rect 242249 219194 242315 219197
rect 128353 219192 242315 219194
rect 128353 219136 128358 219192
rect 128414 219136 242254 219192
rect 242310 219136 242315 219192
rect 128353 219134 242315 219136
rect 128353 219131 128419 219134
rect 242249 219131 242315 219134
rect 119981 219058 120047 219061
rect 143441 219058 143507 219061
rect 119981 219056 143507 219058
rect 119981 219000 119986 219056
rect 120042 219000 143446 219056
rect 143502 219000 143507 219056
rect 119981 218998 143507 219000
rect 119981 218995 120047 218998
rect 143441 218995 143507 218998
rect 152457 219058 152523 219061
rect 208485 219058 208551 219061
rect 152457 219056 208551 219058
rect 152457 219000 152462 219056
rect 152518 219000 208490 219056
rect 208546 219000 208551 219056
rect 152457 218998 208551 219000
rect 152457 218995 152523 218998
rect 208485 218995 208551 218998
rect 583385 219058 583451 219061
rect 583520 219058 584960 219148
rect 583385 219056 584960 219058
rect 583385 219000 583390 219056
rect 583446 219000 584960 219056
rect 583385 218998 584960 219000
rect 583385 218995 583451 218998
rect 583520 218908 584960 218998
rect 39941 217970 40007 217973
rect 231117 217970 231183 217973
rect 39941 217968 231183 217970
rect 39941 217912 39946 217968
rect 40002 217912 231122 217968
rect 231178 217912 231183 217968
rect 39941 217910 231183 217912
rect 39941 217907 40007 217910
rect 231117 217907 231183 217910
rect 143349 217834 143415 217837
rect 254025 217834 254091 217837
rect 143349 217832 254091 217834
rect 143349 217776 143354 217832
rect 143410 217776 254030 217832
rect 254086 217776 254091 217832
rect 143349 217774 254091 217776
rect 143349 217771 143415 217774
rect 254025 217771 254091 217774
rect 100661 217698 100727 217701
rect 100661 217696 161490 217698
rect 100661 217640 100666 217696
rect 100722 217640 161490 217696
rect 100661 217638 161490 217640
rect 100661 217635 100727 217638
rect 161430 217290 161490 217638
rect 172421 217290 172487 217293
rect 298134 217290 298140 217292
rect 161430 217288 298140 217290
rect 161430 217232 172426 217288
rect 172482 217232 298140 217288
rect 161430 217230 298140 217232
rect 172421 217227 172487 217230
rect 298134 217228 298140 217230
rect 298204 217228 298210 217292
rect 66161 216610 66227 216613
rect 234981 216610 235047 216613
rect 66161 216608 235047 216610
rect 66161 216552 66166 216608
rect 66222 216552 234986 216608
rect 235042 216552 235047 216608
rect 66161 216550 235047 216552
rect 66161 216547 66227 216550
rect 234981 216547 235047 216550
rect 235901 216610 235967 216613
rect 270585 216610 270651 216613
rect 271781 216610 271847 216613
rect 235901 216608 271847 216610
rect 235901 216552 235906 216608
rect 235962 216552 270590 216608
rect 270646 216552 271786 216608
rect 271842 216552 271847 216608
rect 235901 216550 271847 216552
rect 235901 216547 235967 216550
rect 270585 216547 270651 216550
rect 271781 216547 271847 216550
rect 53557 216474 53623 216477
rect 218237 216474 218303 216477
rect 53557 216472 219450 216474
rect 53557 216416 53562 216472
rect 53618 216416 218242 216472
rect 218298 216416 219450 216472
rect 53557 216414 219450 216416
rect 53557 216411 53623 216414
rect 218237 216411 218303 216414
rect 219390 216066 219450 216414
rect 231945 216066 232011 216069
rect 219390 216064 232011 216066
rect 219390 216008 231950 216064
rect 232006 216008 232011 216064
rect 219390 216006 232011 216008
rect 231945 216003 232011 216006
rect 99281 215930 99347 215933
rect 251909 215930 251975 215933
rect 99281 215928 251975 215930
rect 99281 215872 99286 215928
rect 99342 215872 251914 215928
rect 251970 215872 251975 215928
rect 99281 215870 251975 215872
rect 99281 215867 99347 215870
rect 251909 215867 251975 215870
rect 271781 215930 271847 215933
rect 442022 215930 442028 215932
rect 271781 215928 442028 215930
rect 271781 215872 271786 215928
rect 271842 215872 442028 215928
rect 271781 215870 442028 215872
rect 271781 215867 271847 215870
rect 442022 215868 442028 215870
rect 442092 215868 442098 215932
rect 67950 215188 67956 215252
rect 68020 215250 68026 215252
rect 233509 215250 233575 215253
rect 68020 215248 233575 215250
rect 68020 215192 233514 215248
rect 233570 215192 233575 215248
rect 68020 215190 233575 215192
rect 68020 215188 68026 215190
rect 233509 215187 233575 215190
rect 251909 215250 251975 215253
rect 252318 215250 252324 215252
rect 251909 215248 252324 215250
rect 251909 215192 251914 215248
rect 251970 215192 252324 215248
rect 251909 215190 252324 215192
rect 251909 215187 251975 215190
rect 252318 215188 252324 215190
rect 252388 215250 252394 215252
rect 255262 215250 255268 215252
rect 252388 215190 255268 215250
rect 252388 215188 252394 215190
rect 255262 215188 255268 215190
rect 255332 215188 255338 215252
rect 111793 215114 111859 215117
rect 112989 215114 113055 215117
rect 173014 215114 173020 215116
rect 111793 215112 173020 215114
rect -960 214978 480 215068
rect 111793 215056 111798 215112
rect 111854 215056 112994 215112
rect 113050 215056 173020 215112
rect 111793 215054 173020 215056
rect 111793 215051 111859 215054
rect 112989 215051 113055 215054
rect 173014 215052 173020 215054
rect 173084 215052 173090 215116
rect 209681 215114 209747 215117
rect 209814 215114 209820 215116
rect 200070 215112 209820 215114
rect 200070 215056 209686 215112
rect 209742 215056 209820 215112
rect 200070 215054 209820 215056
rect 3325 214978 3391 214981
rect -960 214976 3391 214978
rect -960 214920 3330 214976
rect 3386 214920 3391 214976
rect -960 214918 3391 214920
rect -960 214828 480 214918
rect 3325 214915 3391 214918
rect 186129 214706 186195 214709
rect 197997 214706 198063 214709
rect 186129 214704 198063 214706
rect 186129 214648 186134 214704
rect 186190 214648 198002 214704
rect 198058 214648 198063 214704
rect 186129 214646 198063 214648
rect 186129 214643 186195 214646
rect 197997 214643 198063 214646
rect 49601 214570 49667 214573
rect 200070 214570 200130 215054
rect 209681 215051 209747 215054
rect 209814 215052 209820 215054
rect 209884 215052 209890 215116
rect 317321 215114 317387 215117
rect 219390 215112 317387 215114
rect 219390 215056 317326 215112
rect 317382 215056 317387 215112
rect 219390 215054 317387 215056
rect 208485 214978 208551 214981
rect 219390 214978 219450 215054
rect 317321 215051 317387 215054
rect 208485 214976 219450 214978
rect 208485 214920 208490 214976
rect 208546 214920 219450 214976
rect 208485 214918 219450 214920
rect 208485 214915 208551 214918
rect 235257 214706 235323 214709
rect 237414 214706 237420 214708
rect 235257 214704 237420 214706
rect 235257 214648 235262 214704
rect 235318 214648 237420 214704
rect 235257 214646 237420 214648
rect 235257 214643 235323 214646
rect 237414 214644 237420 214646
rect 237484 214644 237490 214708
rect 49601 214568 200130 214570
rect 49601 214512 49606 214568
rect 49662 214512 200130 214568
rect 49601 214510 200130 214512
rect 222101 214570 222167 214573
rect 306465 214570 306531 214573
rect 222101 214568 306531 214570
rect 222101 214512 222106 214568
rect 222162 214512 306470 214568
rect 306526 214512 306531 214568
rect 222101 214510 306531 214512
rect 49601 214507 49667 214510
rect 222101 214507 222167 214510
rect 306465 214507 306531 214510
rect 215937 214026 216003 214029
rect 215158 214024 216003 214026
rect 215158 213968 215942 214024
rect 215998 213968 216003 214024
rect 215158 213966 216003 213968
rect 56409 213890 56475 213893
rect 215158 213890 215218 213966
rect 215937 213963 216003 213966
rect 56409 213888 215218 213890
rect 56409 213832 56414 213888
rect 56470 213832 215218 213888
rect 56409 213830 215218 213832
rect 215293 213890 215359 213893
rect 292481 213890 292547 213893
rect 293217 213890 293283 213893
rect 215293 213888 293283 213890
rect 215293 213832 215298 213888
rect 215354 213832 292486 213888
rect 292542 213832 293222 213888
rect 293278 213832 293283 213888
rect 215293 213830 293283 213832
rect 56409 213827 56475 213830
rect 215293 213827 215359 213830
rect 292481 213827 292547 213830
rect 293217 213827 293283 213830
rect 117129 213754 117195 213757
rect 205633 213754 205699 213757
rect 117129 213752 205699 213754
rect 117129 213696 117134 213752
rect 117190 213696 205638 213752
rect 205694 213696 205699 213752
rect 117129 213694 205699 213696
rect 117129 213691 117195 213694
rect 205633 213691 205699 213694
rect 214557 213754 214623 213757
rect 248454 213754 248460 213756
rect 214557 213752 248460 213754
rect 214557 213696 214562 213752
rect 214618 213696 248460 213752
rect 214557 213694 248460 213696
rect 214557 213691 214623 213694
rect 248454 213692 248460 213694
rect 248524 213754 248530 213756
rect 249701 213754 249767 213757
rect 248524 213752 249767 213754
rect 248524 213696 249706 213752
rect 249762 213696 249767 213752
rect 248524 213694 249767 213696
rect 248524 213692 248530 213694
rect 249701 213691 249767 213694
rect 141417 213618 141483 213621
rect 216029 213618 216095 213621
rect 141417 213616 216095 213618
rect 141417 213560 141422 213616
rect 141478 213560 216034 213616
rect 216090 213560 216095 213616
rect 141417 213558 216095 213560
rect 141417 213555 141483 213558
rect 216029 213555 216095 213558
rect 225229 213210 225295 213213
rect 315297 213210 315363 213213
rect 225229 213208 315363 213210
rect 225229 213152 225234 213208
rect 225290 213152 315302 213208
rect 315358 213152 315363 213208
rect 225229 213150 315363 213152
rect 225229 213147 225295 213150
rect 315297 213147 315363 213150
rect 215293 212666 215359 212669
rect 216438 212666 216444 212668
rect 215293 212664 216444 212666
rect 215293 212608 215298 212664
rect 215354 212608 216444 212664
rect 215293 212606 216444 212608
rect 215293 212603 215359 212606
rect 216438 212604 216444 212606
rect 216508 212666 216514 212668
rect 221457 212666 221523 212669
rect 216508 212664 221523 212666
rect 216508 212608 221462 212664
rect 221518 212608 221523 212664
rect 216508 212606 221523 212608
rect 216508 212604 216514 212606
rect 221457 212603 221523 212606
rect 64505 212530 64571 212533
rect 193857 212532 193923 212533
rect 193806 212530 193812 212532
rect 64505 212528 193812 212530
rect 193876 212530 193923 212532
rect 213269 212530 213335 212533
rect 263593 212530 263659 212533
rect 193876 212528 193968 212530
rect 64505 212472 64510 212528
rect 64566 212472 193812 212528
rect 193918 212472 193968 212528
rect 64505 212470 193812 212472
rect 64505 212467 64571 212470
rect 193806 212468 193812 212470
rect 193876 212470 193968 212472
rect 213269 212528 263659 212530
rect 213269 212472 213274 212528
rect 213330 212472 263598 212528
rect 263654 212472 263659 212528
rect 213269 212470 263659 212472
rect 193876 212468 193923 212470
rect 193857 212467 193923 212468
rect 213269 212467 213335 212470
rect 263593 212467 263659 212470
rect 95233 212394 95299 212397
rect 96521 212394 96587 212397
rect 168414 212394 168420 212396
rect 95233 212392 168420 212394
rect 95233 212336 95238 212392
rect 95294 212336 96526 212392
rect 96582 212336 168420 212392
rect 95233 212334 168420 212336
rect 95233 212331 95299 212334
rect 96521 212331 96587 212334
rect 168414 212332 168420 212334
rect 168484 212332 168490 212396
rect 188429 211850 188495 211853
rect 253197 211850 253263 211853
rect 188429 211848 253263 211850
rect 188429 211792 188434 211848
rect 188490 211792 253202 211848
rect 253258 211792 253263 211848
rect 188429 211790 253263 211792
rect 188429 211787 188495 211790
rect 253197 211787 253263 211790
rect 196709 211170 196775 211173
rect 318241 211170 318307 211173
rect 583109 211170 583175 211173
rect 583569 211170 583635 211173
rect 196709 211168 318307 211170
rect 196709 211112 196714 211168
rect 196770 211112 318246 211168
rect 318302 211112 318307 211168
rect 196709 211110 318307 211112
rect 196709 211107 196775 211110
rect 318241 211107 318307 211110
rect 567150 211168 583635 211170
rect 567150 211112 583114 211168
rect 583170 211112 583574 211168
rect 583630 211112 583635 211168
rect 567150 211110 583635 211112
rect 131021 211034 131087 211037
rect 162117 211034 162183 211037
rect 162761 211034 162827 211037
rect 131021 211032 162827 211034
rect 131021 210976 131026 211032
rect 131082 210976 162122 211032
rect 162178 210976 162766 211032
rect 162822 210976 162827 211032
rect 131021 210974 162827 210976
rect 131021 210971 131087 210974
rect 162117 210971 162183 210974
rect 162761 210971 162827 210974
rect 240961 211034 241027 211037
rect 259361 211034 259427 211037
rect 567150 211034 567210 211110
rect 583109 211107 583175 211110
rect 583569 211107 583635 211110
rect 240961 211032 567210 211034
rect 240961 210976 240966 211032
rect 241022 210976 259366 211032
rect 259422 210976 567210 211032
rect 240961 210974 567210 210976
rect 240961 210971 241027 210974
rect 259361 210971 259427 210974
rect 102041 210898 102107 210901
rect 175181 210898 175247 210901
rect 178769 210898 178835 210901
rect 102041 210896 178835 210898
rect 102041 210840 102046 210896
rect 102102 210840 175186 210896
rect 175242 210840 178774 210896
rect 178830 210840 178835 210896
rect 102041 210838 178835 210840
rect 102041 210835 102107 210838
rect 175181 210835 175247 210838
rect 178769 210835 178835 210838
rect 162761 210762 162827 210765
rect 251265 210762 251331 210765
rect 162761 210760 251331 210762
rect 162761 210704 162766 210760
rect 162822 210704 251270 210760
rect 251326 210704 251331 210760
rect 162761 210702 251331 210704
rect 162761 210699 162827 210702
rect 251265 210699 251331 210702
rect 217317 210490 217383 210493
rect 230422 210490 230428 210492
rect 217317 210488 230428 210490
rect 217317 210432 217322 210488
rect 217378 210432 230428 210488
rect 217317 210430 230428 210432
rect 217317 210427 217383 210430
rect 230422 210428 230428 210430
rect 230492 210428 230498 210492
rect 73797 210354 73863 210357
rect 171869 210354 171935 210357
rect 73797 210352 171935 210354
rect 73797 210296 73802 210352
rect 73858 210296 171874 210352
rect 171930 210296 171935 210352
rect 73797 210294 171935 210296
rect 73797 210291 73863 210294
rect 171869 210291 171935 210294
rect 180057 210354 180123 210357
rect 201585 210354 201651 210357
rect 180057 210352 201651 210354
rect 180057 210296 180062 210352
rect 180118 210296 201590 210352
rect 201646 210296 201651 210352
rect 180057 210294 201651 210296
rect 180057 210291 180123 210294
rect 201585 210291 201651 210294
rect 203609 210354 203675 210357
rect 238753 210354 238819 210357
rect 203609 210352 238819 210354
rect 203609 210296 203614 210352
rect 203670 210296 238758 210352
rect 238814 210296 238819 210352
rect 203609 210294 238819 210296
rect 203609 210291 203675 210294
rect 238753 210291 238819 210294
rect 93945 209674 94011 209677
rect 95141 209674 95207 209677
rect 260097 209674 260163 209677
rect 93945 209672 260163 209674
rect 93945 209616 93950 209672
rect 94006 209616 95146 209672
rect 95202 209616 260102 209672
rect 260158 209616 260163 209672
rect 93945 209614 260163 209616
rect 93945 209611 94011 209614
rect 95141 209611 95207 209614
rect 260097 209611 260163 209614
rect 81341 209538 81407 209541
rect 206277 209538 206343 209541
rect 81341 209536 206343 209538
rect 81341 209480 81346 209536
rect 81402 209480 206282 209536
rect 206338 209480 206343 209536
rect 81341 209478 206343 209480
rect 81341 209475 81407 209478
rect 206277 209475 206343 209478
rect 221917 209538 221983 209541
rect 267825 209538 267891 209541
rect 221917 209536 267891 209538
rect 221917 209480 221922 209536
rect 221978 209480 267830 209536
rect 267886 209480 267891 209536
rect 221917 209478 267891 209480
rect 221917 209475 221983 209478
rect 267825 209475 267891 209478
rect 185577 208994 185643 208997
rect 374729 208994 374795 208997
rect 185577 208992 374795 208994
rect 185577 208936 185582 208992
rect 185638 208936 374734 208992
rect 374790 208936 374795 208992
rect 185577 208934 374795 208936
rect 185577 208931 185643 208934
rect 374729 208931 374795 208934
rect 233366 208388 233372 208452
rect 233436 208450 233442 208452
rect 234429 208450 234495 208453
rect 233436 208448 234495 208450
rect 233436 208392 234434 208448
rect 234490 208392 234495 208448
rect 233436 208390 234495 208392
rect 233436 208388 233442 208390
rect 234429 208387 234495 208390
rect 83457 208314 83523 208317
rect 238845 208314 238911 208317
rect 83457 208312 238911 208314
rect 83457 208256 83462 208312
rect 83518 208256 238850 208312
rect 238906 208256 238911 208312
rect 83457 208254 238911 208256
rect 83457 208251 83523 208254
rect 238845 208251 238911 208254
rect 299473 208178 299539 208181
rect 219390 208176 299539 208178
rect 219390 208120 299478 208176
rect 299534 208120 299539 208176
rect 219390 208118 299539 208120
rect 133137 208042 133203 208045
rect 216673 208042 216739 208045
rect 133137 208040 216739 208042
rect 133137 207984 133142 208040
rect 133198 207984 216678 208040
rect 216734 207984 216739 208040
rect 133137 207982 216739 207984
rect 133137 207979 133203 207982
rect 216673 207979 216739 207982
rect 212717 207906 212783 207909
rect 219390 207906 219450 208118
rect 299473 208115 299539 208118
rect 212717 207904 219450 207906
rect 212717 207848 212722 207904
rect 212778 207848 219450 207904
rect 212717 207846 219450 207848
rect 212717 207843 212783 207846
rect 238753 207770 238819 207773
rect 299749 207770 299815 207773
rect 238753 207768 299815 207770
rect 238753 207712 238758 207768
rect 238814 207712 299754 207768
rect 299810 207712 299815 207768
rect 238753 207710 299815 207712
rect 238753 207707 238819 207710
rect 299749 207707 299815 207710
rect 159214 207572 159220 207636
rect 159284 207634 159290 207636
rect 184197 207634 184263 207637
rect 159284 207632 184263 207634
rect 159284 207576 184202 207632
rect 184258 207576 184263 207632
rect 159284 207574 184263 207576
rect 159284 207572 159290 207574
rect 184197 207571 184263 207574
rect 276749 207634 276815 207637
rect 284518 207634 284524 207636
rect 276749 207632 284524 207634
rect 276749 207576 276754 207632
rect 276810 207576 284524 207632
rect 276749 207574 284524 207576
rect 276749 207571 276815 207574
rect 284518 207572 284524 207574
rect 284588 207572 284594 207636
rect 285581 207634 285647 207637
rect 290590 207634 290596 207636
rect 285581 207632 290596 207634
rect 285581 207576 285586 207632
rect 285642 207576 290596 207632
rect 285581 207574 290596 207576
rect 285581 207571 285647 207574
rect 290590 207572 290596 207574
rect 290660 207572 290666 207636
rect 299473 207634 299539 207637
rect 423990 207634 423996 207636
rect 299473 207632 423996 207634
rect 299473 207576 299478 207632
rect 299534 207576 423996 207632
rect 299473 207574 423996 207576
rect 299473 207571 299539 207574
rect 423990 207572 423996 207574
rect 424060 207572 424066 207636
rect 212717 207090 212783 207093
rect 213269 207090 213335 207093
rect 212717 207088 213335 207090
rect 212717 207032 212722 207088
rect 212778 207032 213274 207088
rect 213330 207032 213335 207088
rect 212717 207030 213335 207032
rect 212717 207027 212783 207030
rect 213269 207027 213335 207030
rect 216673 207090 216739 207093
rect 217317 207090 217383 207093
rect 216673 207088 217383 207090
rect 216673 207032 216678 207088
rect 216734 207032 217322 207088
rect 217378 207032 217383 207088
rect 216673 207030 217383 207032
rect 216673 207027 216739 207030
rect 217317 207027 217383 207030
rect 69657 206954 69723 206957
rect 204713 206954 204779 206957
rect 69657 206952 204779 206954
rect 69657 206896 69662 206952
rect 69718 206896 204718 206952
rect 204774 206896 204779 206952
rect 69657 206894 204779 206896
rect 69657 206891 69723 206894
rect 204713 206891 204779 206894
rect 82905 206818 82971 206821
rect 207105 206818 207171 206821
rect 82905 206816 207171 206818
rect 82905 206760 82910 206816
rect 82966 206760 207110 206816
rect 207166 206760 207171 206816
rect 82905 206758 207171 206760
rect 82905 206755 82971 206758
rect 207105 206755 207171 206758
rect 92473 206682 92539 206685
rect 93761 206682 93827 206685
rect 160737 206682 160803 206685
rect 92473 206680 160803 206682
rect 92473 206624 92478 206680
rect 92534 206624 93766 206680
rect 93822 206624 160742 206680
rect 160798 206624 160803 206680
rect 92473 206622 160803 206624
rect 92473 206619 92539 206622
rect 93761 206619 93827 206622
rect 160737 206619 160803 206622
rect 201585 206410 201651 206413
rect 405733 206410 405799 206413
rect 201585 206408 405799 206410
rect 201585 206352 201590 206408
rect 201646 206352 405738 206408
rect 405794 206352 405799 206408
rect 201585 206350 405799 206352
rect 201585 206347 201651 206350
rect 405733 206347 405799 206350
rect 210417 206274 210483 206277
rect 428457 206274 428523 206277
rect 210417 206272 428523 206274
rect 210417 206216 210422 206272
rect 210478 206216 428462 206272
rect 428518 206216 428523 206272
rect 210417 206214 428523 206216
rect 210417 206211 210483 206214
rect 428457 206211 428523 206214
rect 207105 205730 207171 205733
rect 207657 205730 207723 205733
rect 227713 205732 227779 205733
rect 227662 205730 227668 205732
rect 207105 205728 207723 205730
rect 207105 205672 207110 205728
rect 207166 205672 207662 205728
rect 207718 205672 207723 205728
rect 207105 205670 207723 205672
rect 227622 205670 227668 205730
rect 227732 205728 227779 205732
rect 583520 205730 584960 205820
rect 227774 205672 227779 205728
rect 207105 205667 207171 205670
rect 207657 205667 207723 205670
rect 227662 205668 227668 205670
rect 227732 205668 227779 205672
rect 227713 205667 227779 205668
rect 583342 205670 584960 205730
rect 129641 205594 129707 205597
rect 162209 205594 162275 205597
rect 214465 205596 214531 205597
rect 214414 205594 214420 205596
rect 129641 205592 162275 205594
rect 129641 205536 129646 205592
rect 129702 205536 162214 205592
rect 162270 205536 162275 205592
rect 129641 205534 162275 205536
rect 214374 205534 214420 205594
rect 214484 205592 214531 205596
rect 214526 205536 214531 205592
rect 129641 205531 129707 205534
rect 162209 205531 162275 205534
rect 214414 205532 214420 205534
rect 214484 205532 214531 205536
rect 583342 205594 583402 205670
rect 583520 205594 584960 205670
rect 583342 205580 584960 205594
rect 583342 205534 583586 205580
rect 214465 205531 214531 205532
rect 583526 205461 583586 205534
rect 583477 205456 583586 205461
rect 583477 205400 583482 205456
rect 583538 205400 583586 205456
rect 583477 205398 583586 205400
rect 583477 205395 583543 205398
rect 113081 205050 113147 205053
rect 180057 205050 180123 205053
rect 113081 205048 180123 205050
rect 113081 204992 113086 205048
rect 113142 204992 180062 205048
rect 180118 204992 180123 205048
rect 113081 204990 180123 204992
rect 113081 204987 113147 204990
rect 180057 204987 180123 204990
rect 153101 204914 153167 204917
rect 356789 204914 356855 204917
rect 153101 204912 356855 204914
rect 153101 204856 153106 204912
rect 153162 204856 356794 204912
rect 356850 204856 356855 204912
rect 153101 204854 356855 204856
rect 153101 204851 153167 204854
rect 356789 204851 356855 204854
rect 198825 204370 198891 204373
rect 436185 204370 436251 204373
rect 198825 204368 436251 204370
rect 198825 204312 198830 204368
rect 198886 204312 436190 204368
rect 436246 204312 436251 204368
rect 198825 204310 436251 204312
rect 198825 204307 198891 204310
rect 436185 204307 436251 204310
rect 148961 204234 149027 204237
rect 263593 204234 263659 204237
rect 148961 204232 263659 204234
rect 148961 204176 148966 204232
rect 149022 204176 263598 204232
rect 263654 204176 263659 204232
rect 148961 204174 263659 204176
rect 148961 204171 149027 204174
rect 263593 204171 263659 204174
rect 198825 204098 198891 204101
rect 180750 204096 198891 204098
rect 180750 204040 198830 204096
rect 198886 204040 198891 204096
rect 180750 204038 198891 204040
rect 40677 203554 40743 203557
rect 178677 203554 178743 203557
rect 180750 203554 180810 204038
rect 198825 204035 198891 204038
rect 195646 203628 195652 203692
rect 195716 203690 195722 203692
rect 300117 203690 300183 203693
rect 195716 203688 300183 203690
rect 195716 203632 300122 203688
rect 300178 203632 300183 203688
rect 195716 203630 300183 203632
rect 195716 203628 195722 203630
rect 300117 203627 300183 203630
rect 40677 203552 180810 203554
rect 40677 203496 40682 203552
rect 40738 203496 178682 203552
rect 178738 203496 180810 203552
rect 40677 203494 180810 203496
rect 263593 203554 263659 203557
rect 449893 203554 449959 203557
rect 263593 203552 449959 203554
rect 263593 203496 263598 203552
rect 263654 203496 449898 203552
rect 449954 203496 449959 203552
rect 263593 203494 449959 203496
rect 40677 203491 40743 203494
rect 178677 203491 178743 203494
rect 263593 203491 263659 203494
rect 449893 203491 449959 203494
rect 121361 202874 121427 202877
rect 160093 202874 160159 202877
rect 121361 202872 160159 202874
rect 121361 202816 121366 202872
rect 121422 202816 160098 202872
rect 160154 202816 160159 202872
rect 121361 202814 160159 202816
rect 121361 202811 121427 202814
rect 160093 202811 160159 202814
rect 180149 202466 180215 202469
rect 250437 202466 250503 202469
rect 180149 202464 250503 202466
rect 180149 202408 180154 202464
rect 180210 202408 250442 202464
rect 250498 202408 250503 202464
rect 180149 202406 250503 202408
rect 180149 202403 180215 202406
rect 250437 202403 250503 202406
rect 91001 202330 91067 202333
rect 188429 202330 188495 202333
rect 91001 202328 188495 202330
rect 91001 202272 91006 202328
rect 91062 202272 188434 202328
rect 188490 202272 188495 202328
rect 91001 202270 188495 202272
rect 91001 202267 91067 202270
rect 188429 202267 188495 202270
rect 151721 202194 151787 202197
rect 288709 202194 288775 202197
rect 151721 202192 288775 202194
rect 151721 202136 151726 202192
rect 151782 202136 288714 202192
rect 288770 202136 288775 202192
rect 151721 202134 288775 202136
rect 151721 202131 151787 202134
rect 288709 202131 288775 202134
rect -960 201922 480 202012
rect 3049 201922 3115 201925
rect -960 201920 3115 201922
rect -960 201864 3054 201920
rect 3110 201864 3115 201920
rect -960 201862 3115 201864
rect -960 201772 480 201862
rect 3049 201859 3115 201862
rect 288566 201452 288572 201516
rect 288636 201514 288642 201516
rect 288709 201514 288775 201517
rect 288636 201512 288775 201514
rect 288636 201456 288714 201512
rect 288770 201456 288775 201512
rect 288636 201454 288775 201456
rect 288636 201452 288642 201454
rect 288709 201451 288775 201454
rect 184289 201106 184355 201109
rect 210417 201106 210483 201109
rect 184289 201104 210483 201106
rect 184289 201048 184294 201104
rect 184350 201048 210422 201104
rect 210478 201048 210483 201104
rect 184289 201046 210483 201048
rect 184289 201043 184355 201046
rect 210417 201043 210483 201046
rect 171869 200970 171935 200973
rect 205081 200970 205147 200973
rect 171869 200968 205147 200970
rect 171869 200912 171874 200968
rect 171930 200912 205086 200968
rect 205142 200912 205147 200968
rect 171869 200910 205147 200912
rect 171869 200907 171935 200910
rect 205081 200907 205147 200910
rect 117221 200834 117287 200837
rect 191925 200834 191991 200837
rect 117221 200832 191991 200834
rect 117221 200776 117226 200832
rect 117282 200776 191930 200832
rect 191986 200776 191991 200832
rect 117221 200774 191991 200776
rect 117221 200771 117287 200774
rect 191925 200771 191991 200774
rect 209037 200834 209103 200837
rect 425697 200834 425763 200837
rect 209037 200832 425763 200834
rect 209037 200776 209042 200832
rect 209098 200776 425702 200832
rect 425758 200776 425763 200832
rect 209037 200774 425763 200776
rect 209037 200771 209103 200774
rect 425697 200771 425763 200774
rect 86861 200698 86927 200701
rect 173249 200698 173315 200701
rect 86861 200696 173315 200698
rect 86861 200640 86866 200696
rect 86922 200640 173254 200696
rect 173310 200640 173315 200696
rect 86861 200638 173315 200640
rect 86861 200635 86927 200638
rect 173249 200635 173315 200638
rect 204846 200636 204852 200700
rect 204916 200698 204922 200700
rect 440233 200698 440299 200701
rect 204916 200696 440299 200698
rect 204916 200640 440238 200696
rect 440294 200640 440299 200696
rect 204916 200638 440299 200640
rect 204916 200636 204922 200638
rect 440233 200635 440299 200638
rect 78673 200018 78739 200021
rect 284293 200018 284359 200021
rect 78673 200016 284359 200018
rect 78673 199960 78678 200016
rect 78734 199960 284298 200016
rect 284354 199960 284359 200016
rect 78673 199958 284359 199960
rect 78673 199955 78739 199958
rect 284293 199955 284359 199958
rect 97901 199882 97967 199885
rect 157977 199882 158043 199885
rect 97901 199880 158043 199882
rect 97901 199824 97906 199880
rect 97962 199824 157982 199880
rect 158038 199824 158043 199880
rect 97901 199822 158043 199824
rect 97901 199819 97967 199822
rect 157977 199819 158043 199822
rect 158069 199474 158135 199477
rect 167821 199474 167887 199477
rect 158069 199472 167887 199474
rect 158069 199416 158074 199472
rect 158130 199416 167826 199472
rect 167882 199416 167887 199472
rect 158069 199414 167887 199416
rect 158069 199411 158135 199414
rect 167821 199411 167887 199414
rect 193121 199474 193187 199477
rect 232497 199474 232563 199477
rect 193121 199472 232563 199474
rect 193121 199416 193126 199472
rect 193182 199416 232502 199472
rect 232558 199416 232563 199472
rect 193121 199414 232563 199416
rect 193121 199411 193187 199414
rect 232497 199411 232563 199414
rect 284293 199474 284359 199477
rect 291694 199474 291700 199476
rect 284293 199472 291700 199474
rect 284293 199416 284298 199472
rect 284354 199416 291700 199472
rect 284293 199414 291700 199416
rect 284293 199411 284359 199414
rect 291694 199412 291700 199414
rect 291764 199412 291770 199476
rect 167637 199338 167703 199341
rect 411989 199338 412055 199341
rect 167637 199336 412055 199338
rect 167637 199280 167642 199336
rect 167698 199280 411994 199336
rect 412050 199280 412055 199336
rect 167637 199278 412055 199280
rect 167637 199275 167703 199278
rect 411989 199275 412055 199278
rect 122741 198114 122807 198117
rect 171869 198114 171935 198117
rect 122741 198112 171935 198114
rect 122741 198056 122746 198112
rect 122802 198056 171874 198112
rect 171930 198056 171935 198112
rect 122741 198054 171935 198056
rect 122741 198051 122807 198054
rect 171869 198051 171935 198054
rect 172053 198114 172119 198117
rect 391197 198114 391263 198117
rect 172053 198112 391263 198114
rect 172053 198056 172058 198112
rect 172114 198056 391202 198112
rect 391258 198056 391263 198112
rect 172053 198054 391263 198056
rect 172053 198051 172119 198054
rect 391197 198051 391263 198054
rect 62757 197978 62823 197981
rect 426433 197978 426499 197981
rect 62757 197976 426499 197978
rect 62757 197920 62762 197976
rect 62818 197920 426438 197976
rect 426494 197920 426499 197976
rect 62757 197918 426499 197920
rect 62757 197915 62823 197918
rect 426433 197915 426499 197918
rect 156781 196890 156847 196893
rect 202413 196890 202479 196893
rect 156781 196888 202479 196890
rect 156781 196832 156786 196888
rect 156842 196832 202418 196888
rect 202474 196832 202479 196888
rect 156781 196830 202479 196832
rect 156781 196827 156847 196830
rect 202413 196827 202479 196830
rect 202229 196754 202295 196757
rect 296897 196754 296963 196757
rect 202229 196752 296963 196754
rect 202229 196696 202234 196752
rect 202290 196696 296902 196752
rect 296958 196696 296963 196752
rect 202229 196694 296963 196696
rect 202229 196691 202295 196694
rect 296897 196691 296963 196694
rect 72417 196618 72483 196621
rect 351177 196618 351243 196621
rect 72417 196616 351243 196618
rect 72417 196560 72422 196616
rect 72478 196560 351182 196616
rect 351238 196560 351243 196616
rect 72417 196558 351243 196560
rect 72417 196555 72483 196558
rect 351177 196555 351243 196558
rect 154481 195394 154547 195397
rect 316769 195394 316835 195397
rect 154481 195392 316835 195394
rect 154481 195336 154486 195392
rect 154542 195336 316774 195392
rect 316830 195336 316835 195392
rect 154481 195334 316835 195336
rect 154481 195331 154547 195334
rect 316769 195331 316835 195334
rect 104801 195258 104867 195261
rect 318057 195258 318123 195261
rect 104801 195256 318123 195258
rect 104801 195200 104806 195256
rect 104862 195200 318062 195256
rect 318118 195200 318123 195256
rect 104801 195198 318123 195200
rect 104801 195195 104867 195198
rect 318057 195195 318123 195198
rect 142061 194578 142127 194581
rect 380893 194578 380959 194581
rect 142061 194576 380959 194578
rect 142061 194520 142066 194576
rect 142122 194520 380898 194576
rect 380954 194520 380959 194576
rect 142061 194518 380959 194520
rect 142061 194515 142127 194518
rect 380893 194515 380959 194518
rect 107561 194442 107627 194445
rect 288433 194444 288499 194445
rect 288382 194442 288388 194444
rect 107561 194440 288388 194442
rect 288452 194440 288499 194444
rect 107561 194384 107566 194440
rect 107622 194384 288388 194440
rect 288494 194384 288499 194440
rect 107561 194382 288388 194384
rect 107561 194379 107627 194382
rect 288382 194380 288388 194382
rect 288452 194380 288499 194384
rect 288433 194379 288499 194380
rect 128997 193898 129063 193901
rect 156597 193898 156663 193901
rect 128997 193896 156663 193898
rect 128997 193840 129002 193896
rect 129058 193840 156602 193896
rect 156658 193840 156663 193896
rect 128997 193838 156663 193840
rect 128997 193835 129063 193838
rect 156597 193835 156663 193838
rect 215845 193898 215911 193901
rect 240358 193898 240364 193900
rect 215845 193896 240364 193898
rect 215845 193840 215850 193896
rect 215906 193840 240364 193896
rect 215845 193838 240364 193840
rect 215845 193835 215911 193838
rect 240358 193836 240364 193838
rect 240428 193836 240434 193900
rect 279417 193898 279483 193901
rect 287094 193898 287100 193900
rect 279417 193896 287100 193898
rect 279417 193840 279422 193896
rect 279478 193840 287100 193896
rect 279417 193838 287100 193840
rect 279417 193835 279483 193838
rect 287094 193836 287100 193838
rect 287164 193836 287170 193900
rect 15837 193218 15903 193221
rect 16481 193218 16547 193221
rect 204897 193218 204963 193221
rect 15837 193216 204963 193218
rect 15837 193160 15842 193216
rect 15898 193160 16486 193216
rect 16542 193160 204902 193216
rect 204958 193160 204963 193216
rect 15837 193158 204963 193160
rect 15837 193155 15903 193158
rect 16481 193155 16547 193158
rect 204897 193155 204963 193158
rect 169017 192674 169083 192677
rect 285029 192674 285095 192677
rect 169017 192672 285095 192674
rect 169017 192616 169022 192672
rect 169078 192616 285034 192672
rect 285090 192616 285095 192672
rect 169017 192614 285095 192616
rect 169017 192611 169083 192614
rect 285029 192611 285095 192614
rect 85573 192538 85639 192541
rect 256550 192538 256556 192540
rect 85573 192536 256556 192538
rect 85573 192480 85578 192536
rect 85634 192480 256556 192536
rect 85573 192478 256556 192480
rect 85573 192475 85639 192478
rect 256550 192476 256556 192478
rect 256620 192538 256626 192540
rect 264973 192538 265039 192541
rect 256620 192536 265039 192538
rect 256620 192480 264978 192536
rect 265034 192480 265039 192536
rect 256620 192478 265039 192480
rect 256620 192476 256626 192478
rect 264973 192475 265039 192478
rect 583109 192538 583175 192541
rect 583520 192538 584960 192628
rect 583109 192536 584960 192538
rect 583109 192480 583114 192536
rect 583170 192480 584960 192536
rect 583109 192478 584960 192480
rect 583109 192475 583175 192478
rect 583520 192388 584960 192478
rect 77150 191116 77156 191180
rect 77220 191178 77226 191180
rect 324957 191178 325023 191181
rect 77220 191176 325023 191178
rect 77220 191120 324962 191176
rect 325018 191120 325023 191176
rect 77220 191118 325023 191120
rect 77220 191116 77226 191118
rect 324957 191115 325023 191118
rect 96521 191042 96587 191045
rect 451273 191042 451339 191045
rect 96521 191040 451339 191042
rect 96521 190984 96526 191040
rect 96582 190984 451278 191040
rect 451334 190984 451339 191040
rect 96521 190982 451339 190984
rect 96521 190979 96587 190982
rect 451273 190979 451339 190982
rect 61929 190362 61995 190365
rect 220169 190362 220235 190365
rect 61929 190360 220235 190362
rect 61929 190304 61934 190360
rect 61990 190304 220174 190360
rect 220230 190304 220235 190360
rect 61929 190302 220235 190304
rect 61929 190299 61995 190302
rect 220169 190299 220235 190302
rect 223481 189954 223547 189957
rect 277894 189954 277900 189956
rect 223481 189952 277900 189954
rect 223481 189896 223486 189952
rect 223542 189896 277900 189952
rect 223481 189894 277900 189896
rect 223481 189891 223547 189894
rect 277894 189892 277900 189894
rect 277964 189892 277970 189956
rect 202413 189818 202479 189821
rect 444465 189818 444531 189821
rect 202413 189816 444531 189818
rect 202413 189760 202418 189816
rect 202474 189760 444470 189816
rect 444526 189760 444531 189816
rect 202413 189758 444531 189760
rect 202413 189755 202479 189758
rect 444465 189755 444531 189758
rect 75678 189620 75684 189684
rect 75748 189682 75754 189684
rect 448605 189682 448671 189685
rect 75748 189680 448671 189682
rect 75748 189624 448610 189680
rect 448666 189624 448671 189680
rect 75748 189622 448671 189624
rect 75748 189620 75754 189622
rect 448605 189619 448671 189622
rect -960 188866 480 188956
rect 3509 188866 3575 188869
rect -960 188864 3575 188866
rect -960 188808 3514 188864
rect 3570 188808 3575 188864
rect -960 188806 3575 188808
rect -960 188716 480 188806
rect 3509 188803 3575 188806
rect 195605 188594 195671 188597
rect 237414 188594 237420 188596
rect 195605 188592 237420 188594
rect 195605 188536 195610 188592
rect 195666 188536 237420 188592
rect 195605 188534 237420 188536
rect 195605 188531 195671 188534
rect 237414 188532 237420 188534
rect 237484 188532 237490 188596
rect 95141 188458 95207 188461
rect 299606 188458 299612 188460
rect 95141 188456 299612 188458
rect 95141 188400 95146 188456
rect 95202 188400 299612 188456
rect 95141 188398 299612 188400
rect 95141 188395 95207 188398
rect 299606 188396 299612 188398
rect 299676 188396 299682 188460
rect 69606 188260 69612 188324
rect 69676 188322 69682 188324
rect 397453 188322 397519 188325
rect 69676 188320 397519 188322
rect 69676 188264 397458 188320
rect 397514 188264 397519 188320
rect 69676 188262 397519 188264
rect 69676 188260 69682 188262
rect 397453 188259 397519 188262
rect 163497 187234 163563 187237
rect 184289 187234 184355 187237
rect 163497 187232 184355 187234
rect 163497 187176 163502 187232
rect 163558 187176 184294 187232
rect 184350 187176 184355 187232
rect 163497 187174 184355 187176
rect 163497 187171 163563 187174
rect 184289 187171 184355 187174
rect 201401 187234 201467 187237
rect 280245 187234 280311 187237
rect 201401 187232 280311 187234
rect 201401 187176 201406 187232
rect 201462 187176 280250 187232
rect 280306 187176 280311 187232
rect 201401 187174 280311 187176
rect 201401 187171 201467 187174
rect 280245 187171 280311 187174
rect 100661 187098 100727 187101
rect 303654 187098 303660 187100
rect 100661 187096 303660 187098
rect 100661 187040 100666 187096
rect 100722 187040 303660 187096
rect 100661 187038 303660 187040
rect 100661 187035 100727 187038
rect 303654 187036 303660 187038
rect 303724 187036 303730 187100
rect 90909 186962 90975 186965
rect 169017 186962 169083 186965
rect 90909 186960 169083 186962
rect 90909 186904 90914 186960
rect 90970 186904 169022 186960
rect 169078 186904 169083 186960
rect 90909 186902 169083 186904
rect 90909 186899 90975 186902
rect 169017 186899 169083 186902
rect 205081 186962 205147 186965
rect 583201 186962 583267 186965
rect 205081 186960 583267 186962
rect 205081 186904 205086 186960
rect 205142 186904 583206 186960
rect 583262 186904 583267 186960
rect 205081 186902 583267 186904
rect 205081 186899 205147 186902
rect 583201 186899 583267 186902
rect 174537 186282 174603 186285
rect 205633 186282 205699 186285
rect 174537 186280 205699 186282
rect 174537 186224 174542 186280
rect 174598 186224 205638 186280
rect 205694 186224 205699 186280
rect 174537 186222 205699 186224
rect 174537 186219 174603 186222
rect 205633 186219 205699 186222
rect 191741 185738 191807 185741
rect 320909 185738 320975 185741
rect 191741 185736 320975 185738
rect 191741 185680 191746 185736
rect 191802 185680 320914 185736
rect 320970 185680 320975 185736
rect 191741 185678 320975 185680
rect 191741 185675 191807 185678
rect 320909 185675 320975 185678
rect 93761 185602 93827 185605
rect 405825 185602 405891 185605
rect 93761 185600 405891 185602
rect 93761 185544 93766 185600
rect 93822 185544 405830 185600
rect 405886 185544 405891 185600
rect 93761 185542 405891 185544
rect 93761 185539 93827 185542
rect 405825 185539 405891 185542
rect 155718 184316 155724 184380
rect 155788 184378 155794 184380
rect 295977 184378 296043 184381
rect 155788 184376 296043 184378
rect 155788 184320 295982 184376
rect 296038 184320 296043 184376
rect 155788 184318 296043 184320
rect 155788 184316 155794 184318
rect 295977 184315 296043 184318
rect 170397 184242 170463 184245
rect 404353 184242 404419 184245
rect 170397 184240 404419 184242
rect 170397 184184 170402 184240
rect 170458 184184 404358 184240
rect 404414 184184 404419 184240
rect 170397 184182 404419 184184
rect 170397 184179 170463 184182
rect 404353 184179 404419 184182
rect 101949 183698 102015 183701
rect 166349 183698 166415 183701
rect 101949 183696 166415 183698
rect 101949 183640 101954 183696
rect 102010 183640 166354 183696
rect 166410 183640 166415 183696
rect 101949 183638 166415 183640
rect 101949 183635 102015 183638
rect 166349 183635 166415 183638
rect 225873 183698 225939 183701
rect 252645 183698 252711 183701
rect 225873 183696 252711 183698
rect 225873 183640 225878 183696
rect 225934 183640 252650 183696
rect 252706 183640 252711 183696
rect 225873 183638 252711 183640
rect 225873 183635 225939 183638
rect 252645 183635 252711 183638
rect 181529 183562 181595 183565
rect 224953 183562 225019 183565
rect 181529 183560 225019 183562
rect 181529 183504 181534 183560
rect 181590 183504 224958 183560
rect 225014 183504 225019 183560
rect 181529 183502 225019 183504
rect 181529 183499 181595 183502
rect 224953 183499 225019 183502
rect 228214 183500 228220 183564
rect 228284 183562 228290 183564
rect 228633 183562 228699 183565
rect 228284 183560 228699 183562
rect 228284 183504 228638 183560
rect 228694 183504 228699 183560
rect 228284 183502 228699 183504
rect 228284 183500 228290 183502
rect 228633 183499 228699 183502
rect 197261 183018 197327 183021
rect 228766 183018 228772 183020
rect 197261 183016 228772 183018
rect 197261 182960 197266 183016
rect 197322 182960 228772 183016
rect 197261 182958 228772 182960
rect 197261 182955 197327 182958
rect 228766 182956 228772 182958
rect 228836 182956 228842 183020
rect 271137 183018 271203 183021
rect 285622 183018 285628 183020
rect 271137 183016 285628 183018
rect 271137 182960 271142 183016
rect 271198 182960 285628 183016
rect 271137 182958 285628 182960
rect 271137 182955 271203 182958
rect 285622 182956 285628 182958
rect 285692 182956 285698 183020
rect 225597 182882 225663 182885
rect 280470 182882 280476 182884
rect 225597 182880 280476 182882
rect 225597 182824 225602 182880
rect 225658 182824 280476 182880
rect 225597 182822 280476 182824
rect 225597 182819 225663 182822
rect 280470 182820 280476 182822
rect 280540 182820 280546 182884
rect 112253 182338 112319 182341
rect 184381 182338 184447 182341
rect 112253 182336 184447 182338
rect 112253 182280 112258 182336
rect 112314 182280 184386 182336
rect 184442 182280 184447 182336
rect 112253 182278 184447 182280
rect 112253 182275 112319 182278
rect 184381 182275 184447 182278
rect 226241 182338 226307 182341
rect 242934 182338 242940 182340
rect 226241 182336 242940 182338
rect 226241 182280 226246 182336
rect 226302 182280 242940 182336
rect 226241 182278 242940 182280
rect 226241 182275 226307 182278
rect 242934 182276 242940 182278
rect 243004 182276 243010 182340
rect 103329 182202 103395 182205
rect 180333 182202 180399 182205
rect 103329 182200 180399 182202
rect 103329 182144 103334 182200
rect 103390 182144 180338 182200
rect 180394 182144 180399 182200
rect 103329 182142 180399 182144
rect 103329 182139 103395 182142
rect 180333 182139 180399 182142
rect 227713 182202 227779 182205
rect 272057 182202 272123 182205
rect 227713 182200 272123 182202
rect 227713 182144 227718 182200
rect 227774 182144 272062 182200
rect 272118 182144 272123 182200
rect 227713 182142 272123 182144
rect 227713 182139 227779 182142
rect 272057 182139 272123 182142
rect 166901 182066 166967 182069
rect 169702 182066 169708 182068
rect 166901 182064 169708 182066
rect 166901 182008 166906 182064
rect 166962 182008 169708 182064
rect 166901 182006 169708 182008
rect 166901 182003 166967 182006
rect 169702 182004 169708 182006
rect 169772 182004 169778 182068
rect 226977 181522 227043 181525
rect 278814 181522 278820 181524
rect 226977 181520 278820 181522
rect 226977 181464 226982 181520
rect 227038 181464 278820 181520
rect 226977 181462 278820 181464
rect 226977 181459 227043 181462
rect 278814 181460 278820 181462
rect 278884 181460 278890 181524
rect 194501 181386 194567 181389
rect 245837 181386 245903 181389
rect 194501 181384 245903 181386
rect 194501 181328 194506 181384
rect 194562 181328 245842 181384
rect 245898 181328 245903 181384
rect 194501 181326 245903 181328
rect 194501 181323 194567 181326
rect 245837 181323 245903 181326
rect 272057 181386 272123 181389
rect 430573 181386 430639 181389
rect 272057 181384 430639 181386
rect 272057 181328 272062 181384
rect 272118 181328 430578 181384
rect 430634 181328 430639 181384
rect 272057 181326 430639 181328
rect 272057 181323 272123 181326
rect 430573 181323 430639 181326
rect 105721 180978 105787 180981
rect 181529 180978 181595 180981
rect 105721 180976 181595 180978
rect 105721 180920 105726 180976
rect 105782 180920 181534 180976
rect 181590 180920 181595 180976
rect 105721 180918 181595 180920
rect 105721 180915 105787 180918
rect 181529 180915 181595 180918
rect 98453 180842 98519 180845
rect 169109 180842 169175 180845
rect 98453 180840 169175 180842
rect 98453 180784 98458 180840
rect 98514 180784 169114 180840
rect 169170 180784 169175 180840
rect 98453 180782 169175 180784
rect 98453 180779 98519 180782
rect 169109 180779 169175 180782
rect 169702 180780 169708 180844
rect 169772 180842 169778 180844
rect 401685 180842 401751 180845
rect 169772 180840 401751 180842
rect 169772 180784 401690 180840
rect 401746 180784 401751 180840
rect 169772 180782 401751 180784
rect 169772 180780 169778 180782
rect 401685 180779 401751 180782
rect 161974 180644 161980 180708
rect 162044 180706 162050 180708
rect 214557 180706 214623 180709
rect 162044 180704 214623 180706
rect 162044 180648 214562 180704
rect 214618 180648 214623 180704
rect 162044 180646 214623 180648
rect 162044 180644 162050 180646
rect 214557 180643 214623 180646
rect 211889 180162 211955 180165
rect 229369 180162 229435 180165
rect 211889 180160 229435 180162
rect 211889 180104 211894 180160
rect 211950 180104 229374 180160
rect 229430 180104 229435 180160
rect 211889 180102 229435 180104
rect 211889 180099 211955 180102
rect 229369 180099 229435 180102
rect 186957 180026 187023 180029
rect 244365 180026 244431 180029
rect 186957 180024 244431 180026
rect 186957 179968 186962 180024
rect 187018 179968 244370 180024
rect 244426 179968 244431 180024
rect 186957 179966 244431 179968
rect 186957 179963 187023 179966
rect 244365 179963 244431 179966
rect 264329 180026 264395 180029
rect 281574 180026 281580 180028
rect 264329 180024 281580 180026
rect 264329 179968 264334 180024
rect 264390 179968 281580 180024
rect 264329 179966 281580 179968
rect 264329 179963 264395 179966
rect 281574 179964 281580 179966
rect 281644 179964 281650 180028
rect 283557 180026 283623 180029
rect 294229 180026 294295 180029
rect 283557 180024 294295 180026
rect 283557 179968 283562 180024
rect 283618 179968 294234 180024
rect 294290 179968 294295 180024
rect 283557 179966 294295 179968
rect 283557 179963 283623 179966
rect 294229 179963 294295 179966
rect 230381 179754 230447 179757
rect 441705 179754 441771 179757
rect 230381 179752 441771 179754
rect 230381 179696 230386 179752
rect 230442 179696 441710 179752
rect 441766 179696 441771 179752
rect 230381 179694 441771 179696
rect 230381 179691 230447 179694
rect 441705 179691 441771 179694
rect 107009 179618 107075 179621
rect 173341 179618 173407 179621
rect 107009 179616 173407 179618
rect 107009 179560 107014 179616
rect 107070 179560 173346 179616
rect 173402 179560 173407 179616
rect 107009 179558 173407 179560
rect 107009 179555 107075 179558
rect 173341 179555 173407 179558
rect 221222 179556 221228 179620
rect 221292 179618 221298 179620
rect 241053 179618 241119 179621
rect 221292 179616 241119 179618
rect 221292 179560 241058 179616
rect 241114 179560 241119 179616
rect 221292 179558 241119 179560
rect 221292 179556 221298 179558
rect 241053 179555 241119 179558
rect 97441 179482 97507 179485
rect 185669 179482 185735 179485
rect 97441 179480 185735 179482
rect 97441 179424 97446 179480
rect 97502 179424 185674 179480
rect 185730 179424 185735 179480
rect 97441 179422 185735 179424
rect 97441 179419 97507 179422
rect 185669 179419 185735 179422
rect 282126 179420 282132 179484
rect 282196 179482 282202 179484
rect 282913 179482 282979 179485
rect 282196 179480 282979 179482
rect 282196 179424 282918 179480
rect 282974 179424 282979 179480
rect 282196 179422 282979 179424
rect 282196 179420 282202 179422
rect 282913 179419 282979 179422
rect 580901 179210 580967 179213
rect 583520 179210 584960 179300
rect 580901 179208 584960 179210
rect 580901 179152 580906 179208
rect 580962 179152 584960 179208
rect 580901 179150 584960 179152
rect 580901 179147 580967 179150
rect 228357 179074 228423 179077
rect 231894 179074 231900 179076
rect 228357 179072 231900 179074
rect 228357 179016 228362 179072
rect 228418 179016 231900 179072
rect 228357 179014 231900 179016
rect 228357 179011 228423 179014
rect 231894 179012 231900 179014
rect 231964 179012 231970 179076
rect 583520 179060 584960 179150
rect 192477 178938 192543 178941
rect 209037 178938 209103 178941
rect 192477 178936 209103 178938
rect 192477 178880 192482 178936
rect 192538 178880 209042 178936
rect 209098 178880 209103 178936
rect 192477 178878 209103 178880
rect 192477 178875 192543 178878
rect 209037 178875 209103 178878
rect 221457 178938 221523 178941
rect 226333 178938 226399 178941
rect 221457 178936 226399 178938
rect 221457 178880 221462 178936
rect 221518 178880 226338 178936
rect 226394 178880 226399 178936
rect 221457 178878 226399 178880
rect 221457 178875 221523 178878
rect 226333 178875 226399 178878
rect 227069 178938 227135 178941
rect 237598 178938 237604 178940
rect 227069 178936 237604 178938
rect 227069 178880 227074 178936
rect 227130 178880 237604 178936
rect 227069 178878 237604 178880
rect 227069 178875 227135 178878
rect 237598 178876 237604 178878
rect 237668 178876 237674 178940
rect 160737 178802 160803 178805
rect 197302 178802 197308 178804
rect 160737 178800 197308 178802
rect 160737 178744 160742 178800
rect 160798 178744 197308 178800
rect 160737 178742 197308 178744
rect 160737 178739 160803 178742
rect 197302 178740 197308 178742
rect 197372 178740 197378 178804
rect 209221 178802 209287 178805
rect 275369 178802 275435 178805
rect 288709 178802 288775 178805
rect 209221 178800 229110 178802
rect 209221 178744 209226 178800
rect 209282 178744 229110 178800
rect 209221 178742 229110 178744
rect 209221 178739 209287 178742
rect 35157 178666 35223 178669
rect 133137 178666 133203 178669
rect 35157 178664 133203 178666
rect 35157 178608 35162 178664
rect 35218 178608 133142 178664
rect 133198 178608 133203 178664
rect 35157 178606 133203 178608
rect 35157 178603 35223 178606
rect 133137 178603 133203 178606
rect 180241 178666 180307 178669
rect 227713 178666 227779 178669
rect 180241 178664 227779 178666
rect 180241 178608 180246 178664
rect 180302 178608 227718 178664
rect 227774 178608 227779 178664
rect 180241 178606 227779 178608
rect 229050 178666 229110 178742
rect 275369 178800 288775 178802
rect 275369 178744 275374 178800
rect 275430 178744 288714 178800
rect 288770 178744 288775 178800
rect 275369 178742 288775 178744
rect 275369 178739 275435 178742
rect 288709 178739 288775 178742
rect 230565 178666 230631 178669
rect 253933 178666 253999 178669
rect 229050 178664 253999 178666
rect 229050 178608 230570 178664
rect 230626 178608 253938 178664
rect 253994 178608 253999 178664
rect 229050 178606 253999 178608
rect 180241 178603 180307 178606
rect 227713 178603 227779 178606
rect 230565 178603 230631 178606
rect 253933 178603 253999 178606
rect 273989 178666 274055 178669
rect 291377 178666 291443 178669
rect 273989 178664 291443 178666
rect 273989 178608 273994 178664
rect 274050 178608 291382 178664
rect 291438 178608 291443 178664
rect 273989 178606 291443 178608
rect 273989 178603 274055 178606
rect 291377 178603 291443 178606
rect 167637 178258 167703 178261
rect 110646 178256 167703 178258
rect 110646 178200 167642 178256
rect 167698 178200 167703 178256
rect 110646 178198 167703 178200
rect 110646 177988 110706 178198
rect 167637 178195 167703 178198
rect 177389 178122 177455 178125
rect 118374 178120 177455 178122
rect 118374 178064 177394 178120
rect 177450 178064 177455 178120
rect 118374 178062 177455 178064
rect 118374 177988 118434 178062
rect 177389 178059 177455 178062
rect 232446 178060 232452 178124
rect 232516 178122 232522 178124
rect 233233 178122 233299 178125
rect 232516 178120 233299 178122
rect 232516 178064 233238 178120
rect 233294 178064 233299 178120
rect 232516 178062 233299 178064
rect 232516 178060 232522 178062
rect 233233 178059 233299 178062
rect 110638 177924 110644 177988
rect 110708 177924 110714 177988
rect 118366 177924 118372 177988
rect 118436 177924 118442 177988
rect 98310 177516 98316 177580
rect 98380 177578 98386 177580
rect 98453 177578 98519 177581
rect 98380 177576 98519 177578
rect 98380 177520 98458 177576
rect 98514 177520 98519 177576
rect 98380 177518 98519 177520
rect 98380 177516 98386 177518
rect 98453 177515 98519 177518
rect 100702 177516 100708 177580
rect 100772 177578 100778 177580
rect 101949 177578 102015 177581
rect 105721 177580 105787 177581
rect 105670 177578 105676 177580
rect 100772 177576 102015 177578
rect 100772 177520 101954 177576
rect 102010 177520 102015 177576
rect 100772 177518 102015 177520
rect 105630 177518 105676 177578
rect 105740 177576 105787 177580
rect 105782 177520 105787 177576
rect 100772 177516 100778 177518
rect 101949 177515 102015 177518
rect 105670 177516 105676 177518
rect 105740 177516 105787 177520
rect 108062 177516 108068 177580
rect 108132 177578 108138 177580
rect 108941 177578 109007 177581
rect 108132 177576 109007 177578
rect 108132 177520 108946 177576
rect 109002 177520 109007 177576
rect 108132 177518 109007 177520
rect 108132 177516 108138 177518
rect 105721 177515 105787 177516
rect 108941 177515 109007 177518
rect 109534 177516 109540 177580
rect 109604 177578 109610 177580
rect 110321 177578 110387 177581
rect 109604 177576 110387 177578
rect 109604 177520 110326 177576
rect 110382 177520 110387 177576
rect 109604 177518 110387 177520
rect 109604 177516 109610 177518
rect 110321 177515 110387 177518
rect 113214 177516 113220 177580
rect 113284 177578 113290 177580
rect 114461 177578 114527 177581
rect 115841 177580 115907 177581
rect 115790 177578 115796 177580
rect 113284 177576 114527 177578
rect 113284 177520 114466 177576
rect 114522 177520 114527 177576
rect 113284 177518 114527 177520
rect 115750 177518 115796 177578
rect 115860 177576 115907 177580
rect 115902 177520 115907 177576
rect 113284 177516 113290 177518
rect 114461 177515 114527 177518
rect 115790 177516 115796 177518
rect 115860 177516 115907 177520
rect 116894 177516 116900 177580
rect 116964 177578 116970 177580
rect 117221 177578 117287 177581
rect 116964 177576 117287 177578
rect 116964 177520 117226 177576
rect 117282 177520 117287 177576
rect 116964 177518 117287 177520
rect 116964 177516 116970 177518
rect 115841 177515 115907 177516
rect 117221 177515 117287 177518
rect 123150 177516 123156 177580
rect 123220 177578 123226 177580
rect 123477 177578 123543 177581
rect 123220 177576 123543 177578
rect 123220 177520 123482 177576
rect 123538 177520 123543 177576
rect 123220 177518 123543 177520
rect 123220 177516 123226 177518
rect 123477 177515 123543 177518
rect 133086 177516 133092 177580
rect 133156 177578 133162 177580
rect 133781 177578 133847 177581
rect 133156 177576 133847 177578
rect 133156 177520 133786 177576
rect 133842 177520 133847 177576
rect 133156 177518 133847 177520
rect 133156 177516 133162 177518
rect 133781 177515 133847 177518
rect 134374 177516 134380 177580
rect 134444 177578 134450 177580
rect 134793 177578 134859 177581
rect 148225 177580 148291 177581
rect 148174 177578 148180 177580
rect 134444 177576 134859 177578
rect 134444 177520 134798 177576
rect 134854 177520 134859 177576
rect 134444 177518 134859 177520
rect 148134 177518 148180 177578
rect 148244 177576 148291 177580
rect 148286 177520 148291 177576
rect 134444 177516 134450 177518
rect 134793 177515 134859 177518
rect 148174 177516 148180 177518
rect 148244 177516 148291 177520
rect 148225 177515 148291 177516
rect 112110 177380 112116 177444
rect 112180 177442 112186 177444
rect 112253 177442 112319 177445
rect 112180 177440 112319 177442
rect 112180 177384 112258 177440
rect 112314 177384 112319 177440
rect 112180 177382 112319 177384
rect 112180 177380 112186 177382
rect 112253 177379 112319 177382
rect 210417 177442 210483 177445
rect 289997 177442 290063 177445
rect 210417 177440 290063 177442
rect 210417 177384 210422 177440
rect 210478 177384 290002 177440
rect 290058 177384 290063 177440
rect 210417 177382 290063 177384
rect 210417 177379 210483 177382
rect 289997 177379 290063 177382
rect 169385 177306 169451 177309
rect 214833 177306 214899 177309
rect 169385 177304 214899 177306
rect 169385 177248 169390 177304
rect 169446 177248 214838 177304
rect 214894 177248 214899 177304
rect 169385 177246 214899 177248
rect 169385 177243 169451 177246
rect 214833 177243 214899 177246
rect 215937 177306 216003 177309
rect 440325 177306 440391 177309
rect 215937 177304 440391 177306
rect 215937 177248 215942 177304
rect 215998 177248 440330 177304
rect 440386 177248 440391 177304
rect 215937 177246 440391 177248
rect 215937 177243 216003 177246
rect 440325 177243 440391 177246
rect 104566 177108 104572 177172
rect 104636 177170 104642 177172
rect 196709 177170 196775 177173
rect 104636 177168 196775 177170
rect 104636 177112 196714 177168
rect 196770 177112 196775 177168
rect 104636 177110 196775 177112
rect 104636 177108 104642 177110
rect 196709 177107 196775 177110
rect 278773 177170 278839 177173
rect 279366 177170 279372 177172
rect 278773 177168 279372 177170
rect 278773 177112 278778 177168
rect 278834 177112 279372 177168
rect 278773 177110 279372 177112
rect 278773 177107 278839 177110
rect 279366 177108 279372 177110
rect 279436 177108 279442 177172
rect 107009 177036 107075 177037
rect 106958 177034 106964 177036
rect 106918 176974 106964 177034
rect 107028 177032 107075 177036
rect 107070 176976 107075 177032
rect 106958 176972 106964 176974
rect 107028 176972 107075 176976
rect 119470 176972 119476 177036
rect 119540 177034 119546 177036
rect 119797 177034 119863 177037
rect 119540 177032 119863 177034
rect 119540 176976 119802 177032
rect 119858 176976 119863 177032
rect 119540 176974 119863 176976
rect 119540 176972 119546 176974
rect 107009 176971 107075 176972
rect 119797 176971 119863 176974
rect 127014 176972 127020 177036
rect 127084 177034 127090 177036
rect 164969 177034 165035 177037
rect 127084 177032 165035 177034
rect 127084 176976 164974 177032
rect 165030 176976 165035 177032
rect 127084 176974 165035 176976
rect 127084 176972 127090 176974
rect 164969 176971 165035 176974
rect 97022 176836 97028 176900
rect 97092 176898 97098 176900
rect 97441 176898 97507 176901
rect 97092 176896 97507 176898
rect 97092 176840 97446 176896
rect 97502 176840 97507 176896
rect 97092 176838 97507 176840
rect 97092 176836 97098 176838
rect 97441 176835 97507 176838
rect 120758 176836 120764 176900
rect 120828 176898 120834 176900
rect 169201 176898 169267 176901
rect 120828 176896 169267 176898
rect 120828 176840 169206 176896
rect 169262 176840 169267 176896
rect 120828 176838 169267 176840
rect 120828 176836 120834 176838
rect 169201 176835 169267 176838
rect 226333 176898 226399 176901
rect 229318 176898 229324 176900
rect 226333 176896 229324 176898
rect 226333 176840 226338 176896
rect 226394 176840 229324 176896
rect 226333 176838 229324 176840
rect 226333 176835 226399 176838
rect 229318 176836 229324 176838
rect 229388 176836 229394 176900
rect 100661 176762 100727 176765
rect 102041 176764 102107 176765
rect 101990 176762 101996 176764
rect 99422 176760 100727 176762
rect 99422 176704 100666 176760
rect 100722 176704 100727 176760
rect 99422 176702 100727 176704
rect 101950 176702 101996 176762
rect 102060 176760 102107 176764
rect 103329 176762 103395 176765
rect 102102 176704 102107 176760
rect 99422 176492 99482 176702
rect 100661 176699 100727 176702
rect 101990 176700 101996 176702
rect 102060 176700 102107 176704
rect 102041 176699 102107 176700
rect 103286 176760 103395 176762
rect 103286 176704 103334 176760
rect 103390 176704 103395 176760
rect 103286 176699 103395 176704
rect 124438 176700 124444 176764
rect 124508 176762 124514 176764
rect 125041 176762 125107 176765
rect 128169 176762 128235 176765
rect 130745 176764 130811 176765
rect 132401 176764 132467 176765
rect 136081 176764 136147 176765
rect 130694 176762 130700 176764
rect 124508 176760 125107 176762
rect 124508 176704 125046 176760
rect 125102 176704 125107 176760
rect 124508 176702 125107 176704
rect 124508 176700 124514 176702
rect 125041 176699 125107 176702
rect 128126 176760 128235 176762
rect 128126 176704 128174 176760
rect 128230 176704 128235 176760
rect 128126 176699 128235 176704
rect 130654 176702 130700 176762
rect 130764 176760 130811 176764
rect 132350 176762 132356 176764
rect 130806 176704 130811 176760
rect 130694 176700 130700 176702
rect 130764 176700 130811 176704
rect 132310 176702 132356 176762
rect 132420 176760 132467 176764
rect 136030 176762 136036 176764
rect 132462 176704 132467 176760
rect 132350 176700 132356 176702
rect 132420 176700 132467 176704
rect 135990 176702 136036 176762
rect 136100 176760 136147 176764
rect 136142 176704 136147 176760
rect 136030 176700 136036 176702
rect 136100 176700 136147 176704
rect 158846 176700 158852 176764
rect 158916 176762 158922 176764
rect 158989 176762 159055 176765
rect 158916 176760 159055 176762
rect 158916 176704 158994 176760
rect 159050 176704 159055 176760
rect 158916 176702 159055 176704
rect 158916 176700 158922 176702
rect 130745 176699 130811 176700
rect 132401 176699 132467 176700
rect 136081 176699 136147 176700
rect 158989 176699 159055 176702
rect 229737 176762 229803 176765
rect 232078 176762 232084 176764
rect 229737 176760 232084 176762
rect 229737 176704 229742 176760
rect 229798 176704 232084 176760
rect 229737 176702 232084 176704
rect 229737 176699 229803 176702
rect 232078 176700 232084 176702
rect 232148 176700 232154 176764
rect 278037 176762 278103 176765
rect 284334 176762 284340 176764
rect 278037 176760 284340 176762
rect 278037 176704 278042 176760
rect 278098 176704 284340 176760
rect 278037 176702 284340 176704
rect 278037 176699 278103 176702
rect 284334 176700 284340 176702
rect 284404 176700 284410 176764
rect 103286 176492 103346 176699
rect 128126 176492 128186 176699
rect 227805 176626 227871 176629
rect 230657 176626 230723 176629
rect 227805 176624 230723 176626
rect 227805 176568 227810 176624
rect 227866 176568 230662 176624
rect 230718 176568 230723 176624
rect 227805 176566 230723 176568
rect 227805 176563 227871 176566
rect 230657 176563 230723 176566
rect 99414 176428 99420 176492
rect 99484 176428 99490 176492
rect 103278 176428 103284 176492
rect 103348 176428 103354 176492
rect 128118 176428 128124 176492
rect 128188 176428 128194 176492
rect 280061 176490 280127 176493
rect 284569 176490 284635 176493
rect 280061 176488 284635 176490
rect 280061 176432 280066 176488
rect 280122 176432 284574 176488
rect 284630 176432 284635 176488
rect 280061 176430 284635 176432
rect 280061 176427 280127 176430
rect 284569 176427 284635 176430
rect 227805 176082 227871 176085
rect 239029 176082 239095 176085
rect 227805 176080 239095 176082
rect -960 175796 480 176036
rect 227805 176024 227810 176080
rect 227866 176024 239034 176080
rect 239090 176024 239095 176080
rect 227805 176022 239095 176024
rect 227805 176019 227871 176022
rect 239029 176019 239095 176022
rect 279877 176082 279943 176085
rect 279877 176080 279986 176082
rect 279877 176024 279882 176080
rect 279938 176024 279986 176080
rect 279877 176019 279986 176024
rect 221181 175948 221247 175949
rect 224217 175948 224283 175949
rect 221181 175946 221228 175948
rect 221136 175944 221228 175946
rect 221136 175888 221186 175944
rect 221136 175886 221228 175888
rect 221181 175884 221228 175886
rect 221292 175884 221298 175948
rect 224166 175946 224172 175948
rect 224126 175886 224172 175946
rect 224236 175944 224283 175948
rect 224278 175888 224283 175944
rect 224166 175884 224172 175886
rect 224236 175884 224283 175888
rect 227662 175884 227668 175948
rect 227732 175946 227738 175948
rect 227732 175886 229202 175946
rect 227732 175884 227738 175886
rect 221181 175883 221247 175884
rect 224217 175883 224283 175884
rect 125726 175748 125732 175812
rect 125796 175810 125802 175812
rect 190361 175810 190427 175813
rect 125796 175750 132510 175810
rect 125796 175748 125802 175750
rect 129457 175676 129523 175677
rect 129406 175674 129412 175676
rect 129366 175614 129412 175674
rect 129476 175672 129523 175676
rect 129518 175616 129523 175672
rect 129406 175612 129412 175614
rect 129476 175612 129523 175616
rect 132450 175674 132510 175750
rect 190361 175808 228282 175810
rect 190361 175752 190366 175808
rect 190422 175752 228282 175808
rect 190361 175750 228282 175752
rect 190361 175747 190427 175750
rect 165153 175674 165219 175677
rect 132450 175672 165219 175674
rect 132450 175616 165158 175672
rect 165214 175616 165219 175672
rect 132450 175614 165219 175616
rect 129457 175611 129523 175612
rect 165153 175611 165219 175614
rect 213913 175674 213979 175677
rect 213913 175672 217028 175674
rect 213913 175616 213918 175672
rect 213974 175616 217028 175672
rect 228222 175644 228282 175750
rect 213913 175614 217028 175616
rect 213913 175611 213979 175614
rect 121862 175476 121868 175540
rect 121932 175538 121938 175540
rect 167913 175538 167979 175541
rect 121932 175536 167979 175538
rect 121932 175480 167918 175536
rect 167974 175480 167979 175536
rect 121932 175478 167979 175480
rect 121932 175476 121938 175478
rect 167913 175475 167979 175478
rect 114318 175340 114324 175404
rect 114388 175402 114394 175404
rect 166533 175402 166599 175405
rect 114388 175400 166599 175402
rect 114388 175344 166538 175400
rect 166594 175344 166599 175400
rect 114388 175342 166599 175344
rect 114388 175340 114394 175342
rect 166533 175339 166599 175342
rect 164877 175266 164943 175269
rect 214557 175266 214623 175269
rect 229142 175266 229202 175886
rect 277894 175748 277900 175812
rect 277964 175810 277970 175812
rect 279601 175810 279667 175813
rect 277964 175808 279667 175810
rect 277964 175752 279606 175808
rect 279662 175752 279667 175808
rect 277964 175750 279667 175752
rect 277964 175748 277970 175750
rect 279601 175747 279667 175750
rect 264973 175674 265039 175677
rect 264973 175672 268180 175674
rect 264973 175616 264978 175672
rect 265034 175616 268180 175672
rect 264973 175614 268180 175616
rect 264973 175611 265039 175614
rect 279926 175538 279986 176019
rect 281809 175538 281875 175541
rect 279926 175536 281875 175538
rect 279926 175508 281814 175536
rect 279956 175480 281814 175508
rect 281870 175480 281875 175536
rect 279956 175478 281875 175480
rect 281809 175475 281875 175478
rect 164877 175264 214623 175266
rect 164877 175208 164882 175264
rect 164938 175208 214562 175264
rect 214618 175208 214623 175264
rect 164877 175206 214623 175208
rect 228988 175206 229202 175266
rect 265065 175266 265131 175269
rect 265065 175264 268180 175266
rect 265065 175208 265070 175264
rect 265126 175208 268180 175264
rect 265065 175206 268180 175208
rect 164877 175203 164943 175206
rect 214557 175203 214623 175206
rect 265065 175203 265131 175206
rect 203609 175130 203675 175133
rect 214557 175130 214623 175133
rect 203609 175128 214623 175130
rect 203609 175072 203614 175128
rect 203670 175072 214562 175128
rect 214618 175072 214623 175128
rect 203609 175070 214623 175072
rect 203609 175067 203675 175070
rect 214557 175067 214623 175070
rect 213913 174994 213979 174997
rect 213913 174992 217028 174994
rect 213913 174936 213918 174992
rect 213974 174936 217028 174992
rect 213913 174934 217028 174936
rect 213913 174931 213979 174934
rect 265709 174858 265775 174861
rect 265709 174856 268180 174858
rect 265709 174800 265714 174856
rect 265770 174800 268180 174856
rect 265709 174798 268180 174800
rect 265709 174795 265775 174798
rect 230565 174722 230631 174725
rect 282821 174722 282887 174725
rect 228988 174720 230631 174722
rect 228988 174664 230570 174720
rect 230626 174664 230631 174720
rect 228988 174662 230631 174664
rect 279956 174720 282887 174722
rect 279956 174664 282826 174720
rect 282882 174664 282887 174720
rect 279956 174662 282887 174664
rect 230565 174659 230631 174662
rect 282821 174659 282887 174662
rect 238017 174586 238083 174589
rect 245929 174586 245995 174589
rect 238017 174584 245995 174586
rect 238017 174528 238022 174584
rect 238078 174528 245934 174584
rect 245990 174528 245995 174584
rect 238017 174526 245995 174528
rect 238017 174523 238083 174526
rect 245929 174523 245995 174526
rect 229134 174388 229140 174452
rect 229204 174450 229210 174452
rect 230565 174450 230631 174453
rect 229204 174448 230631 174450
rect 229204 174392 230570 174448
rect 230626 174392 230631 174448
rect 229204 174390 230631 174392
rect 229204 174388 229210 174390
rect 230565 174387 230631 174390
rect 258030 174390 268180 174450
rect 214005 174314 214071 174317
rect 241697 174314 241763 174317
rect 214005 174312 217028 174314
rect 214005 174256 214010 174312
rect 214066 174256 217028 174312
rect 214005 174254 217028 174256
rect 228988 174312 241763 174314
rect 228988 174256 241702 174312
rect 241758 174256 241763 174312
rect 228988 174254 241763 174256
rect 214005 174251 214071 174254
rect 241697 174251 241763 174254
rect 249241 174314 249307 174317
rect 258030 174314 258090 174390
rect 249241 174312 258090 174314
rect 249241 174256 249246 174312
rect 249302 174256 258090 174312
rect 249241 174254 258090 174256
rect 279601 174314 279667 174317
rect 282729 174314 282795 174317
rect 279601 174312 282795 174314
rect 279601 174256 279606 174312
rect 279662 174256 282734 174312
rect 282790 174256 282795 174312
rect 279601 174254 282795 174256
rect 249241 174251 249307 174254
rect 279601 174251 279667 174254
rect 282729 174251 282795 174254
rect 229185 174042 229251 174045
rect 232037 174042 232103 174045
rect 229185 174040 232103 174042
rect 229185 173984 229190 174040
rect 229246 173984 232042 174040
rect 232098 173984 232103 174040
rect 229185 173982 232103 173984
rect 229185 173979 229251 173982
rect 232037 173979 232103 173982
rect 264973 174042 265039 174045
rect 282821 174042 282887 174045
rect 264973 174040 268180 174042
rect 264973 173984 264978 174040
rect 265034 173984 268180 174040
rect 264973 173982 268180 173984
rect 279956 174040 282887 174042
rect 279956 173984 282826 174040
rect 282882 173984 282887 174040
rect 279956 173982 282887 173984
rect 264973 173979 265039 173982
rect 282821 173979 282887 173982
rect 171777 173906 171843 173909
rect 215385 173906 215451 173909
rect 171777 173904 215451 173906
rect 171777 173848 171782 173904
rect 171838 173848 215390 173904
rect 215446 173848 215451 173904
rect 171777 173846 215451 173848
rect 171777 173843 171843 173846
rect 215385 173843 215451 173846
rect 229093 173770 229159 173773
rect 228988 173768 229159 173770
rect 228988 173712 229098 173768
rect 229154 173712 229159 173768
rect 228988 173710 229159 173712
rect 229093 173707 229159 173710
rect 279325 173770 279391 173773
rect 279325 173768 279434 173770
rect 279325 173712 279330 173768
rect 279386 173712 279434 173768
rect 279325 173707 279434 173712
rect 213913 173634 213979 173637
rect 265065 173634 265131 173637
rect 213913 173632 217028 173634
rect 213913 173576 213918 173632
rect 213974 173576 217028 173632
rect 213913 173574 217028 173576
rect 265065 173632 268180 173634
rect 265065 173576 265070 173632
rect 265126 173576 268180 173632
rect 265065 173574 268180 173576
rect 213913 173571 213979 173574
rect 265065 173571 265131 173574
rect 230749 173362 230815 173365
rect 228988 173360 230815 173362
rect 228988 173304 230754 173360
rect 230810 173304 230815 173360
rect 228988 173302 230815 173304
rect 230749 173299 230815 173302
rect 279374 173196 279434 173707
rect 258030 173030 268180 173090
rect 214005 172954 214071 172957
rect 242249 172954 242315 172957
rect 258030 172954 258090 173030
rect 281441 172954 281507 172957
rect 214005 172952 217028 172954
rect 214005 172896 214010 172952
rect 214066 172896 217028 172952
rect 214005 172894 217028 172896
rect 242249 172952 258090 172954
rect 242249 172896 242254 172952
rect 242310 172896 258090 172952
rect 242249 172894 258090 172896
rect 279926 172952 281507 172954
rect 279926 172896 281446 172952
rect 281502 172896 281507 172952
rect 279926 172894 281507 172896
rect 214005 172891 214071 172894
rect 242249 172891 242315 172894
rect 244273 172818 244339 172821
rect 228988 172816 244339 172818
rect 228988 172760 244278 172816
rect 244334 172760 244339 172816
rect 228988 172758 244339 172760
rect 244273 172755 244339 172758
rect 264973 172682 265039 172685
rect 264973 172680 268180 172682
rect 264973 172624 264978 172680
rect 265034 172624 268180 172680
rect 264973 172622 268180 172624
rect 264973 172619 265039 172622
rect 279926 172516 279986 172894
rect 281441 172891 281507 172894
rect 252737 172410 252803 172413
rect 228988 172408 252803 172410
rect 228988 172352 252742 172408
rect 252798 172352 252803 172408
rect 228988 172350 252803 172352
rect 252737 172347 252803 172350
rect 213913 172274 213979 172277
rect 265065 172274 265131 172277
rect 279325 172274 279391 172277
rect 213913 172272 217028 172274
rect 213913 172216 213918 172272
rect 213974 172216 217028 172272
rect 213913 172214 217028 172216
rect 265065 172272 268180 172274
rect 265065 172216 265070 172272
rect 265126 172216 268180 172272
rect 265065 172214 268180 172216
rect 279325 172272 279434 172274
rect 279325 172216 279330 172272
rect 279386 172216 279434 172272
rect 213913 172211 213979 172214
rect 265065 172211 265131 172214
rect 279325 172211 279434 172216
rect 231761 171866 231827 171869
rect 228988 171864 231827 171866
rect 228988 171808 231766 171864
rect 231822 171808 231827 171864
rect 228988 171806 231827 171808
rect 231761 171803 231827 171806
rect 164724 171594 165354 171600
rect 167821 171594 167887 171597
rect 164724 171592 167887 171594
rect 164724 171540 167826 171592
rect 165294 171536 167826 171540
rect 167882 171536 167887 171592
rect 165294 171534 167887 171536
rect 167821 171531 167887 171534
rect 214097 171594 214163 171597
rect 253473 171594 253539 171597
rect 268150 171594 268210 171836
rect 279374 171700 279434 172211
rect 214097 171592 217028 171594
rect 214097 171536 214102 171592
rect 214158 171536 217028 171592
rect 214097 171534 217028 171536
rect 253473 171592 268210 171594
rect 253473 171536 253478 171592
rect 253534 171536 268210 171592
rect 253473 171534 268210 171536
rect 214097 171531 214163 171534
rect 253473 171531 253539 171534
rect 231577 171458 231643 171461
rect 228988 171456 231643 171458
rect 228988 171400 231582 171456
rect 231638 171400 231643 171456
rect 228988 171398 231643 171400
rect 231577 171395 231643 171398
rect 264973 171458 265039 171461
rect 264973 171456 268180 171458
rect 264973 171400 264978 171456
rect 265034 171400 268180 171456
rect 264973 171398 268180 171400
rect 264973 171395 265039 171398
rect 213913 171050 213979 171053
rect 264973 171050 265039 171053
rect 213913 171048 217028 171050
rect 213913 170992 213918 171048
rect 213974 170992 217028 171048
rect 213913 170990 217028 170992
rect 264973 171048 268180 171050
rect 264973 170992 264978 171048
rect 265034 170992 268180 171048
rect 264973 170990 268180 170992
rect 213913 170987 213979 170990
rect 264973 170987 265039 170990
rect 229277 170914 229343 170917
rect 281809 170914 281875 170917
rect 228988 170912 229343 170914
rect 228988 170856 229282 170912
rect 229338 170856 229343 170912
rect 228988 170854 229343 170856
rect 279956 170912 281875 170914
rect 279956 170856 281814 170912
rect 281870 170856 281875 170912
rect 279956 170854 281875 170856
rect 229277 170851 229343 170854
rect 281809 170851 281875 170854
rect 279366 170580 279372 170644
rect 279436 170580 279442 170644
rect 230749 170506 230815 170509
rect 228988 170504 230815 170506
rect 228988 170448 230754 170504
rect 230810 170448 230815 170504
rect 228988 170446 230815 170448
rect 230749 170443 230815 170446
rect 214005 170370 214071 170373
rect 229737 170370 229803 170373
rect 238937 170370 239003 170373
rect 214005 170368 217028 170370
rect 214005 170312 214010 170368
rect 214066 170312 217028 170368
rect 214005 170310 217028 170312
rect 229737 170368 239003 170370
rect 229737 170312 229742 170368
rect 229798 170312 238942 170368
rect 238998 170312 239003 170368
rect 229737 170310 239003 170312
rect 214005 170307 214071 170310
rect 229737 170307 229803 170310
rect 238937 170307 239003 170310
rect 260097 170234 260163 170237
rect 268150 170234 268210 170476
rect 260097 170232 268210 170234
rect 260097 170176 260102 170232
rect 260158 170176 268210 170232
rect 279374 170204 279434 170580
rect 260097 170174 268210 170176
rect 260097 170171 260163 170174
rect 264237 170098 264303 170101
rect 264237 170096 268180 170098
rect 264237 170040 264242 170096
rect 264298 170040 268180 170096
rect 264237 170038 268180 170040
rect 264237 170035 264303 170038
rect 231761 169962 231827 169965
rect 228988 169960 231827 169962
rect 228988 169904 231766 169960
rect 231822 169904 231827 169960
rect 228988 169902 231827 169904
rect 231761 169899 231827 169902
rect 213913 169690 213979 169693
rect 264973 169690 265039 169693
rect 213913 169688 217028 169690
rect 213913 169632 213918 169688
rect 213974 169632 217028 169688
rect 213913 169630 217028 169632
rect 264973 169688 268180 169690
rect 264973 169632 264978 169688
rect 265034 169632 268180 169688
rect 264973 169630 268180 169632
rect 213913 169627 213979 169630
rect 264973 169627 265039 169630
rect 234705 169554 234771 169557
rect 228988 169552 234771 169554
rect 228988 169496 234710 169552
rect 234766 169496 234771 169552
rect 228988 169494 234771 169496
rect 234705 169491 234771 169494
rect 282821 169418 282887 169421
rect 279956 169416 282887 169418
rect 279956 169360 282826 169416
rect 282882 169360 282887 169416
rect 279956 169358 282887 169360
rect 282821 169355 282887 169358
rect 214005 169010 214071 169013
rect 231209 169010 231275 169013
rect 268150 169010 268210 169252
rect 279417 169146 279483 169149
rect 214005 169008 217028 169010
rect 214005 168952 214010 169008
rect 214066 168952 217028 169008
rect 214005 168950 217028 168952
rect 228988 169008 231275 169010
rect 228988 168952 231214 169008
rect 231270 168952 231275 169008
rect 228988 168950 231275 168952
rect 214005 168947 214071 168950
rect 231209 168947 231275 168950
rect 258030 168950 268210 169010
rect 279374 169144 279483 169146
rect 279374 169088 279422 169144
rect 279478 169088 279483 169144
rect 279374 169083 279483 169088
rect 231761 168602 231827 168605
rect 228988 168600 231827 168602
rect 228988 168544 231766 168600
rect 231822 168544 231827 168600
rect 228988 168542 231827 168544
rect 231761 168539 231827 168542
rect 234613 168602 234679 168605
rect 236494 168602 236500 168604
rect 234613 168600 236500 168602
rect 234613 168544 234618 168600
rect 234674 168544 236500 168600
rect 234613 168542 236500 168544
rect 234613 168539 234679 168542
rect 236494 168540 236500 168542
rect 236564 168540 236570 168604
rect 251817 168602 251883 168605
rect 258030 168602 258090 168950
rect 265065 168874 265131 168877
rect 265065 168872 268180 168874
rect 265065 168816 265070 168872
rect 265126 168816 268180 168872
rect 265065 168814 268180 168816
rect 265065 168811 265131 168814
rect 279374 168708 279434 169083
rect 251817 168600 258090 168602
rect 251817 168544 251822 168600
rect 251878 168544 258090 168600
rect 251817 168542 258090 168544
rect 251817 168539 251883 168542
rect 236085 168466 236151 168469
rect 236678 168466 236684 168468
rect 236085 168464 236684 168466
rect 236085 168408 236090 168464
rect 236146 168408 236684 168464
rect 236085 168406 236684 168408
rect 236085 168403 236151 168406
rect 236678 168404 236684 168406
rect 236748 168404 236754 168468
rect 236821 168466 236887 168469
rect 236821 168464 268180 168466
rect 236821 168408 236826 168464
rect 236882 168408 268180 168464
rect 236821 168406 268180 168408
rect 236821 168403 236887 168406
rect 213913 168330 213979 168333
rect 213913 168328 217028 168330
rect 213913 168272 213918 168328
rect 213974 168272 217028 168328
rect 213913 168270 217028 168272
rect 213913 168267 213979 168270
rect 231393 168058 231459 168061
rect 228988 168056 231459 168058
rect 228988 168000 231398 168056
rect 231454 168000 231459 168056
rect 228988 167998 231459 168000
rect 231393 167995 231459 167998
rect 264973 167922 265039 167925
rect 282821 167922 282887 167925
rect 264973 167920 268180 167922
rect 264973 167864 264978 167920
rect 265034 167864 268180 167920
rect 264973 167862 268180 167864
rect 279956 167920 282887 167922
rect 279956 167864 282826 167920
rect 282882 167864 282887 167920
rect 279956 167862 282887 167864
rect 264973 167859 265039 167862
rect 282821 167859 282887 167862
rect 214005 167650 214071 167653
rect 231761 167650 231827 167653
rect 214005 167648 217028 167650
rect 214005 167592 214010 167648
rect 214066 167592 217028 167648
rect 214005 167590 217028 167592
rect 228988 167648 231827 167650
rect 228988 167592 231766 167648
rect 231822 167592 231827 167648
rect 228988 167590 231827 167592
rect 214005 167587 214071 167590
rect 231761 167587 231827 167590
rect 238385 167650 238451 167653
rect 244406 167650 244412 167652
rect 238385 167648 244412 167650
rect 238385 167592 238390 167648
rect 238446 167592 244412 167648
rect 238385 167590 244412 167592
rect 238385 167587 238451 167590
rect 244406 167588 244412 167590
rect 244476 167588 244482 167652
rect 265065 167514 265131 167517
rect 265065 167512 268180 167514
rect 265065 167456 265070 167512
rect 265126 167456 268180 167512
rect 265065 167454 268180 167456
rect 265065 167451 265131 167454
rect 247033 167106 247099 167109
rect 282729 167106 282795 167109
rect 228988 167104 247099 167106
rect 228988 167048 247038 167104
rect 247094 167048 247099 167104
rect 228988 167046 247099 167048
rect 247033 167043 247099 167046
rect 264976 167046 268180 167106
rect 279956 167104 282795 167106
rect 279956 167048 282734 167104
rect 282790 167048 282795 167104
rect 279956 167046 282795 167048
rect 213913 166970 213979 166973
rect 262857 166970 262923 166973
rect 264976 166970 265036 167046
rect 282729 167043 282795 167046
rect 213913 166968 217028 166970
rect 213913 166912 213918 166968
rect 213974 166912 217028 166968
rect 213913 166910 217028 166912
rect 262857 166968 265036 166970
rect 262857 166912 262862 166968
rect 262918 166912 265036 166968
rect 262857 166910 265036 166912
rect 213913 166907 213979 166910
rect 262857 166907 262923 166910
rect 279509 166834 279575 166837
rect 279509 166832 279618 166834
rect 279509 166776 279514 166832
rect 279570 166776 279618 166832
rect 279509 166771 279618 166776
rect 231761 166698 231827 166701
rect 228988 166696 231827 166698
rect 228988 166640 231766 166696
rect 231822 166640 231827 166696
rect 228988 166638 231827 166640
rect 231761 166635 231827 166638
rect 214005 166426 214071 166429
rect 268150 166426 268210 166668
rect 214005 166424 217028 166426
rect 214005 166368 214010 166424
rect 214066 166368 217028 166424
rect 214005 166366 217028 166368
rect 258030 166366 268210 166426
rect 279558 166396 279618 166771
rect 214005 166363 214071 166366
rect 235533 166290 235599 166293
rect 237373 166290 237439 166293
rect 235533 166288 237439 166290
rect 235533 166232 235538 166288
rect 235594 166232 237378 166288
rect 237434 166232 237439 166288
rect 235533 166230 237439 166232
rect 235533 166227 235599 166230
rect 237373 166227 237439 166230
rect 231117 166154 231183 166157
rect 228988 166152 231183 166154
rect 228988 166096 231122 166152
rect 231178 166096 231183 166152
rect 228988 166094 231183 166096
rect 231117 166091 231183 166094
rect 250437 166018 250503 166021
rect 258030 166018 258090 166366
rect 264973 166290 265039 166293
rect 264973 166288 268180 166290
rect 264973 166232 264978 166288
rect 265034 166232 268180 166288
rect 264973 166230 268180 166232
rect 264973 166227 265039 166230
rect 250437 166016 258090 166018
rect 250437 165960 250442 166016
rect 250498 165960 258090 166016
rect 250437 165958 258090 165960
rect 250437 165955 250503 165958
rect 265617 165882 265683 165885
rect 582465 165882 582531 165885
rect 583520 165882 584960 165972
rect 265617 165880 268180 165882
rect 265617 165824 265622 165880
rect 265678 165824 268180 165880
rect 265617 165822 268180 165824
rect 582465 165880 584960 165882
rect 582465 165824 582470 165880
rect 582526 165824 584960 165880
rect 582465 165822 584960 165824
rect 265617 165819 265683 165822
rect 582465 165819 582531 165822
rect 214833 165746 214899 165749
rect 237598 165746 237604 165748
rect 214833 165744 217028 165746
rect 214833 165688 214838 165744
rect 214894 165688 217028 165744
rect 214833 165686 217028 165688
rect 228988 165686 237604 165746
rect 214833 165683 214899 165686
rect 237598 165684 237604 165686
rect 237668 165684 237674 165748
rect 583520 165732 584960 165822
rect 282821 165610 282887 165613
rect 279956 165608 282887 165610
rect 279956 165552 282826 165608
rect 282882 165552 282887 165608
rect 279956 165550 282887 165552
rect 282821 165547 282887 165550
rect 265065 165338 265131 165341
rect 265065 165336 268180 165338
rect 265065 165280 265070 165336
rect 265126 165280 268180 165336
rect 265065 165278 268180 165280
rect 265065 165275 265131 165278
rect 234613 165202 234679 165205
rect 228988 165200 234679 165202
rect 228988 165144 234618 165200
rect 234674 165144 234679 165200
rect 228988 165142 234679 165144
rect 234613 165139 234679 165142
rect 213913 165066 213979 165069
rect 213913 165064 217028 165066
rect 213913 165008 213918 165064
rect 213974 165008 217028 165064
rect 213913 165006 217028 165008
rect 213913 165003 213979 165006
rect 264973 164930 265039 164933
rect 280245 164930 280311 164933
rect 264973 164928 268180 164930
rect 264973 164872 264978 164928
rect 265034 164872 268180 164928
rect 264973 164870 268180 164872
rect 279956 164928 280311 164930
rect 279956 164872 280250 164928
rect 280306 164872 280311 164928
rect 279956 164870 280311 164872
rect 264973 164867 265039 164870
rect 280245 164867 280311 164870
rect 231485 164794 231551 164797
rect 228988 164792 231551 164794
rect 228988 164736 231490 164792
rect 231546 164736 231551 164792
rect 228988 164734 231551 164736
rect 231485 164731 231551 164734
rect 238017 164522 238083 164525
rect 238017 164520 268180 164522
rect 238017 164464 238022 164520
rect 238078 164464 268180 164520
rect 238017 164462 268180 164464
rect 238017 164459 238083 164462
rect 214005 164386 214071 164389
rect 229185 164386 229251 164389
rect 214005 164384 217028 164386
rect 214005 164328 214010 164384
rect 214066 164328 217028 164384
rect 214005 164326 217028 164328
rect 228988 164384 229251 164386
rect 228988 164328 229190 164384
rect 229246 164328 229251 164384
rect 228988 164326 229251 164328
rect 214005 164323 214071 164326
rect 229185 164323 229251 164326
rect 265249 164114 265315 164117
rect 281809 164114 281875 164117
rect 265249 164112 268180 164114
rect 265249 164056 265254 164112
rect 265310 164056 268180 164112
rect 265249 164054 268180 164056
rect 279956 164112 281875 164114
rect 279956 164056 281814 164112
rect 281870 164056 281875 164112
rect 279956 164054 281875 164056
rect 265249 164051 265315 164054
rect 281809 164051 281875 164054
rect 231761 163842 231827 163845
rect 228988 163840 231827 163842
rect 228988 163784 231766 163840
rect 231822 163784 231827 163840
rect 228988 163782 231827 163784
rect 231761 163779 231827 163782
rect 214465 163706 214531 163709
rect 265065 163706 265131 163709
rect 214465 163704 217028 163706
rect 214465 163648 214470 163704
rect 214526 163648 217028 163704
rect 214465 163646 217028 163648
rect 265065 163704 268180 163706
rect 265065 163648 265070 163704
rect 265126 163648 268180 163704
rect 265065 163646 268180 163648
rect 214465 163643 214531 163646
rect 265065 163643 265131 163646
rect 239029 163434 239095 163437
rect 228988 163432 239095 163434
rect 228988 163376 239034 163432
rect 239090 163376 239095 163432
rect 228988 163374 239095 163376
rect 239029 163371 239095 163374
rect 282177 163298 282243 163301
rect 258030 163238 268180 163298
rect 279956 163296 282243 163298
rect 279956 163240 282182 163296
rect 282238 163240 282243 163296
rect 279956 163238 282243 163240
rect 257429 163162 257495 163165
rect 258030 163162 258090 163238
rect 282177 163235 282243 163238
rect 257429 163160 258090 163162
rect 257429 163104 257434 163160
rect 257490 163104 258090 163160
rect 257429 163102 258090 163104
rect 257429 163099 257495 163102
rect 213913 163026 213979 163029
rect 213913 163024 217028 163026
rect -960 162890 480 162980
rect 213913 162968 213918 163024
rect 213974 162968 217028 163024
rect 213913 162966 217028 162968
rect 213913 162963 213979 162966
rect 3509 162890 3575 162893
rect 231669 162890 231735 162893
rect -960 162888 3575 162890
rect -960 162832 3514 162888
rect 3570 162832 3575 162888
rect -960 162830 3575 162832
rect 228988 162888 231735 162890
rect 228988 162832 231674 162888
rect 231730 162832 231735 162888
rect 228988 162830 231735 162832
rect -960 162740 480 162830
rect 3509 162827 3575 162830
rect 231669 162827 231735 162830
rect 264973 162890 265039 162893
rect 264973 162888 268180 162890
rect 264973 162832 264978 162888
rect 265034 162832 268180 162888
rect 264973 162830 268180 162832
rect 264973 162827 265039 162830
rect 282821 162618 282887 162621
rect 279956 162616 282887 162618
rect 279956 162560 282826 162616
rect 282882 162560 282887 162616
rect 279956 162558 282887 162560
rect 282821 162555 282887 162558
rect 249885 162482 249951 162485
rect 228988 162480 249951 162482
rect 228988 162424 249890 162480
rect 249946 162424 249951 162480
rect 228988 162422 249951 162424
rect 249885 162419 249951 162422
rect 213913 162346 213979 162349
rect 265065 162346 265131 162349
rect 213913 162344 217028 162346
rect 213913 162288 213918 162344
rect 213974 162288 217028 162344
rect 213913 162286 217028 162288
rect 265065 162344 268180 162346
rect 265065 162288 265070 162344
rect 265126 162288 268180 162344
rect 265065 162286 268180 162288
rect 213913 162283 213979 162286
rect 265065 162283 265131 162286
rect 229829 162074 229895 162077
rect 242934 162074 242940 162076
rect 229829 162072 242940 162074
rect 229829 162016 229834 162072
rect 229890 162016 242940 162072
rect 229829 162014 242940 162016
rect 229829 162011 229895 162014
rect 242934 162012 242940 162014
rect 243004 162012 243010 162076
rect 230933 161938 230999 161941
rect 228988 161936 230999 161938
rect 228988 161880 230938 161936
rect 230994 161880 230999 161936
rect 228988 161878 230999 161880
rect 230933 161875 230999 161878
rect 258901 161938 258967 161941
rect 258901 161936 268180 161938
rect 258901 161880 258906 161936
rect 258962 161880 268180 161936
rect 258901 161878 268180 161880
rect 258901 161875 258967 161878
rect 214005 161802 214071 161805
rect 282269 161802 282335 161805
rect 214005 161800 217028 161802
rect 214005 161744 214010 161800
rect 214066 161744 217028 161800
rect 214005 161742 217028 161744
rect 279956 161800 282335 161802
rect 279956 161744 282274 161800
rect 282330 161744 282335 161800
rect 279956 161742 282335 161744
rect 214005 161739 214071 161742
rect 282269 161739 282335 161742
rect 240358 161530 240364 161532
rect 228988 161470 240364 161530
rect 240358 161468 240364 161470
rect 240428 161468 240434 161532
rect 264973 161530 265039 161533
rect 264973 161528 268180 161530
rect 264973 161472 264978 161528
rect 265034 161472 268180 161528
rect 264973 161470 268180 161472
rect 264973 161467 265039 161470
rect 213913 161122 213979 161125
rect 265065 161122 265131 161125
rect 280337 161122 280403 161125
rect 213913 161120 217028 161122
rect 213913 161064 213918 161120
rect 213974 161064 217028 161120
rect 213913 161062 217028 161064
rect 265065 161120 268180 161122
rect 265065 161064 265070 161120
rect 265126 161064 268180 161120
rect 265065 161062 268180 161064
rect 279956 161120 280403 161122
rect 279956 161064 280342 161120
rect 280398 161064 280403 161120
rect 279956 161062 280403 161064
rect 213913 161059 213979 161062
rect 265065 161059 265131 161062
rect 280337 161059 280403 161062
rect 230657 160986 230723 160989
rect 228988 160984 230723 160986
rect 228988 160928 230662 160984
rect 230718 160928 230723 160984
rect 228988 160926 230723 160928
rect 230657 160923 230723 160926
rect 264973 160714 265039 160717
rect 264973 160712 268180 160714
rect 264973 160656 264978 160712
rect 265034 160656 268180 160712
rect 264973 160654 268180 160656
rect 264973 160651 265039 160654
rect 286174 160652 286180 160716
rect 286244 160714 286250 160716
rect 441613 160714 441679 160717
rect 286244 160712 441679 160714
rect 286244 160656 441618 160712
rect 441674 160656 441679 160712
rect 286244 160654 441679 160656
rect 286244 160652 286250 160654
rect 441613 160651 441679 160654
rect 233366 160578 233372 160580
rect 228988 160518 233372 160578
rect 233366 160516 233372 160518
rect 233436 160516 233442 160580
rect 214005 160442 214071 160445
rect 214005 160440 217028 160442
rect 214005 160384 214010 160440
rect 214066 160384 217028 160440
rect 214005 160382 217028 160384
rect 214005 160379 214071 160382
rect 282637 160306 282703 160309
rect 258030 160246 268180 160306
rect 279956 160304 282703 160306
rect 279956 160248 282642 160304
rect 282698 160248 282703 160304
rect 279956 160246 282703 160248
rect 233734 160108 233740 160172
rect 233804 160170 233810 160172
rect 236678 160170 236684 160172
rect 233804 160110 236684 160170
rect 233804 160108 233810 160110
rect 236678 160108 236684 160110
rect 236748 160108 236754 160172
rect 240726 160108 240732 160172
rect 240796 160170 240802 160172
rect 258030 160170 258090 160246
rect 282637 160243 282703 160246
rect 240796 160110 258090 160170
rect 240796 160108 240802 160110
rect 251173 160034 251239 160037
rect 228988 160032 251239 160034
rect 228988 159976 251178 160032
rect 251234 159976 251239 160032
rect 228988 159974 251239 159976
rect 251173 159971 251239 159974
rect 213913 159762 213979 159765
rect 265065 159762 265131 159765
rect 213913 159760 217028 159762
rect 213913 159704 213918 159760
rect 213974 159704 217028 159760
rect 213913 159702 217028 159704
rect 265065 159760 268180 159762
rect 265065 159704 265070 159760
rect 265126 159704 268180 159760
rect 265065 159702 268180 159704
rect 213913 159699 213979 159702
rect 265065 159699 265131 159702
rect 231761 159626 231827 159629
rect 228988 159624 231827 159626
rect 228988 159568 231766 159624
rect 231822 159568 231827 159624
rect 228988 159566 231827 159568
rect 231761 159563 231827 159566
rect 282821 159490 282887 159493
rect 279956 159488 282887 159490
rect 279956 159432 282826 159488
rect 282882 159432 282887 159488
rect 279956 159430 282887 159432
rect 282821 159427 282887 159430
rect 214005 159082 214071 159085
rect 231117 159082 231183 159085
rect 214005 159080 217028 159082
rect 214005 159024 214010 159080
rect 214066 159024 217028 159080
rect 214005 159022 217028 159024
rect 228988 159080 231183 159082
rect 228988 159024 231122 159080
rect 231178 159024 231183 159080
rect 228988 159022 231183 159024
rect 214005 159019 214071 159022
rect 231117 159019 231183 159022
rect 249057 159082 249123 159085
rect 268150 159082 268210 159324
rect 249057 159080 268210 159082
rect 249057 159024 249062 159080
rect 249118 159024 268210 159080
rect 249057 159022 268210 159024
rect 249057 159019 249123 159022
rect 264973 158946 265039 158949
rect 264973 158944 268180 158946
rect 264973 158888 264978 158944
rect 265034 158888 268180 158944
rect 264973 158886 268180 158888
rect 264973 158883 265039 158886
rect 282729 158810 282795 158813
rect 279956 158808 282795 158810
rect 279956 158752 282734 158808
rect 282790 158752 282795 158808
rect 279956 158750 282795 158752
rect 282729 158747 282795 158750
rect 230749 158674 230815 158677
rect 228988 158672 230815 158674
rect 228988 158616 230754 158672
rect 230810 158616 230815 158672
rect 228988 158614 230815 158616
rect 230749 158611 230815 158614
rect 265065 158538 265131 158541
rect 265065 158536 268180 158538
rect 265065 158480 265070 158536
rect 265126 158480 268180 158536
rect 265065 158478 268180 158480
rect 265065 158475 265131 158478
rect 213913 158402 213979 158405
rect 213913 158400 217028 158402
rect 213913 158344 213918 158400
rect 213974 158344 217028 158400
rect 213913 158342 217028 158344
rect 213913 158339 213979 158342
rect 230565 158130 230631 158133
rect 228988 158128 230631 158130
rect 228988 158072 230570 158128
rect 230626 158072 230631 158128
rect 228988 158070 230631 158072
rect 230565 158067 230631 158070
rect 231669 157994 231735 157997
rect 235533 157994 235599 157997
rect 231669 157992 235599 157994
rect 231669 157936 231674 157992
rect 231730 157936 235538 157992
rect 235594 157936 235599 157992
rect 231669 157934 235599 157936
rect 231669 157931 231735 157934
rect 235533 157931 235599 157934
rect 232681 157858 232747 157861
rect 268150 157858 268210 158100
rect 282085 157994 282151 157997
rect 279956 157992 282151 157994
rect 279956 157936 282090 157992
rect 282146 157936 282151 157992
rect 279956 157934 282151 157936
rect 282085 157931 282151 157934
rect 232681 157856 268210 157858
rect 232681 157800 232686 157856
rect 232742 157800 268210 157856
rect 232681 157798 268210 157800
rect 232681 157795 232747 157798
rect 214833 157722 214899 157725
rect 230841 157722 230907 157725
rect 214833 157720 217028 157722
rect 214833 157664 214838 157720
rect 214894 157664 217028 157720
rect 214833 157662 217028 157664
rect 228988 157720 230907 157722
rect 228988 157664 230846 157720
rect 230902 157664 230907 157720
rect 228988 157662 230907 157664
rect 214833 157659 214899 157662
rect 230841 157659 230907 157662
rect 264973 157722 265039 157725
rect 264973 157720 268180 157722
rect 264973 157664 264978 157720
rect 265034 157664 268180 157720
rect 264973 157662 268180 157664
rect 264973 157659 265039 157662
rect 283782 157314 283788 157316
rect 279956 157254 283788 157314
rect 283782 157252 283788 157254
rect 283852 157252 283858 157316
rect 213913 157178 213979 157181
rect 233182 157178 233188 157180
rect 213913 157176 217028 157178
rect 213913 157120 213918 157176
rect 213974 157120 217028 157176
rect 213913 157118 217028 157120
rect 228988 157118 233188 157178
rect 213913 157115 213979 157118
rect 233182 157116 233188 157118
rect 233252 157116 233258 157180
rect 265801 157178 265867 157181
rect 265801 157176 268180 157178
rect 265801 157120 265806 157176
rect 265862 157120 268180 157176
rect 265801 157118 268180 157120
rect 265801 157115 265867 157118
rect 248505 156770 248571 156773
rect 228988 156768 248571 156770
rect 228988 156712 248510 156768
rect 248566 156712 248571 156768
rect 228988 156710 248571 156712
rect 248505 156707 248571 156710
rect 265065 156770 265131 156773
rect 265065 156768 268180 156770
rect 265065 156712 265070 156768
rect 265126 156712 268180 156768
rect 265065 156710 268180 156712
rect 265065 156707 265131 156710
rect 214005 156498 214071 156501
rect 214005 156496 217028 156498
rect 214005 156440 214010 156496
rect 214066 156440 217028 156496
rect 214005 156438 217028 156440
rect 214005 156435 214071 156438
rect 264973 156362 265039 156365
rect 264973 156360 268180 156362
rect 264973 156304 264978 156360
rect 265034 156304 268180 156360
rect 264973 156302 268180 156304
rect 264973 156299 265039 156302
rect 230422 156226 230428 156228
rect 228988 156166 230428 156226
rect 230422 156164 230428 156166
rect 230492 156164 230498 156228
rect 279926 156090 279986 156468
rect 304993 156090 305059 156093
rect 279926 156088 305059 156090
rect 279926 156032 304998 156088
rect 305054 156032 305059 156088
rect 279926 156030 305059 156032
rect 304993 156027 305059 156030
rect 265157 155954 265223 155957
rect 265157 155952 268180 155954
rect 265157 155896 265162 155952
rect 265218 155896 268180 155952
rect 265157 155894 268180 155896
rect 265157 155891 265223 155894
rect 213913 155818 213979 155821
rect 229369 155818 229435 155821
rect 213913 155816 217028 155818
rect 213913 155760 213918 155816
rect 213974 155760 217028 155816
rect 213913 155758 217028 155760
rect 228988 155816 229435 155818
rect 228988 155760 229374 155816
rect 229430 155760 229435 155816
rect 228988 155758 229435 155760
rect 213913 155755 213979 155758
rect 229369 155755 229435 155758
rect 282545 155682 282611 155685
rect 279956 155680 282611 155682
rect 279956 155624 282550 155680
rect 282606 155624 282611 155680
rect 279956 155622 282611 155624
rect 282545 155619 282611 155622
rect 231301 155274 231367 155277
rect 228988 155272 231367 155274
rect 228988 155216 231306 155272
rect 231362 155216 231367 155272
rect 228988 155214 231367 155216
rect 231301 155211 231367 155214
rect 233877 155274 233943 155277
rect 268150 155274 268210 155516
rect 233877 155272 268210 155274
rect 233877 155216 233882 155272
rect 233938 155216 268210 155272
rect 233877 155214 268210 155216
rect 233877 155211 233943 155214
rect 214005 155138 214071 155141
rect 214005 155136 217028 155138
rect 214005 155080 214010 155136
rect 214066 155080 217028 155136
rect 214005 155078 217028 155080
rect 214005 155075 214071 155078
rect 238109 154866 238175 154869
rect 228988 154864 238175 154866
rect 228988 154808 238114 154864
rect 238170 154808 238175 154864
rect 228988 154806 238175 154808
rect 238109 154803 238175 154806
rect 251909 154866 251975 154869
rect 268150 154866 268210 155108
rect 281574 155002 281580 155004
rect 279956 154942 281580 155002
rect 281574 154940 281580 154942
rect 281644 154940 281650 155004
rect 251909 154864 268210 154866
rect 251909 154808 251914 154864
rect 251970 154808 268210 154864
rect 251909 154806 268210 154808
rect 251909 154803 251975 154806
rect 264973 154594 265039 154597
rect 264973 154592 268180 154594
rect 264973 154536 264978 154592
rect 265034 154536 268180 154592
rect 264973 154534 268180 154536
rect 264973 154531 265039 154534
rect 214005 154458 214071 154461
rect 214005 154456 217028 154458
rect 214005 154400 214010 154456
rect 214066 154400 217028 154456
rect 214005 154398 217028 154400
rect 214005 154395 214071 154398
rect 231669 154322 231735 154325
rect 228988 154320 231735 154322
rect 228988 154264 231674 154320
rect 231730 154264 231735 154320
rect 228988 154262 231735 154264
rect 231669 154259 231735 154262
rect 265985 154186 266051 154189
rect 282821 154186 282887 154189
rect 265985 154184 268180 154186
rect 265985 154128 265990 154184
rect 266046 154128 268180 154184
rect 265985 154126 268180 154128
rect 279956 154184 282887 154186
rect 279956 154128 282826 154184
rect 282882 154128 282887 154184
rect 279956 154126 282887 154128
rect 265985 154123 266051 154126
rect 282821 154123 282887 154126
rect 231761 153914 231827 153917
rect 228988 153912 231827 153914
rect 228988 153856 231766 153912
rect 231822 153856 231827 153912
rect 228988 153854 231827 153856
rect 231761 153851 231827 153854
rect 213913 153778 213979 153781
rect 230565 153778 230631 153781
rect 244222 153778 244228 153780
rect 213913 153776 217028 153778
rect 213913 153720 213918 153776
rect 213974 153720 217028 153776
rect 213913 153718 217028 153720
rect 230565 153776 244228 153778
rect 230565 153720 230570 153776
rect 230626 153720 244228 153776
rect 230565 153718 244228 153720
rect 213913 153715 213979 153718
rect 230565 153715 230631 153718
rect 244222 153716 244228 153718
rect 244292 153716 244298 153780
rect 264973 153778 265039 153781
rect 264973 153776 268180 153778
rect 264973 153720 264978 153776
rect 265034 153720 268180 153776
rect 264973 153718 268180 153720
rect 264973 153715 265039 153718
rect 282126 153716 282132 153780
rect 282196 153778 282202 153780
rect 291285 153778 291351 153781
rect 282196 153776 291351 153778
rect 282196 153720 291290 153776
rect 291346 153720 291351 153776
rect 282196 153718 291351 153720
rect 282196 153716 282202 153718
rect 291285 153715 291351 153718
rect 282361 153506 282427 153509
rect 279956 153504 282427 153506
rect 279956 153448 282366 153504
rect 282422 153448 282427 153504
rect 279956 153446 282427 153448
rect 282361 153443 282427 153446
rect 231577 153370 231643 153373
rect 228988 153368 231643 153370
rect 228988 153312 231582 153368
rect 231638 153312 231643 153368
rect 228988 153310 231643 153312
rect 231577 153307 231643 153310
rect 258030 153310 268180 153370
rect 243905 153234 243971 153237
rect 258030 153234 258090 153310
rect 243905 153232 258090 153234
rect 243905 153176 243910 153232
rect 243966 153176 258090 153232
rect 243905 153174 258090 153176
rect 243905 153171 243971 153174
rect 213913 153098 213979 153101
rect 213913 153096 217028 153098
rect 213913 153040 213918 153096
rect 213974 153040 217028 153096
rect 213913 153038 217028 153040
rect 213913 153035 213979 153038
rect 254577 152962 254643 152965
rect 228988 152960 254643 152962
rect 228988 152904 254582 152960
rect 254638 152904 254643 152960
rect 228988 152902 254643 152904
rect 254577 152899 254643 152902
rect 264973 152962 265039 152965
rect 264973 152960 268180 152962
rect 264973 152904 264978 152960
rect 265034 152904 268180 152960
rect 264973 152902 268180 152904
rect 264973 152899 265039 152902
rect 282821 152690 282887 152693
rect 279956 152688 282887 152690
rect 279956 152632 282826 152688
rect 282882 152632 282887 152688
rect 279956 152630 282887 152632
rect 282821 152627 282887 152630
rect 582741 152690 582807 152693
rect 583520 152690 584960 152780
rect 582741 152688 584960 152690
rect 582741 152632 582746 152688
rect 582802 152632 584960 152688
rect 582741 152630 584960 152632
rect 582741 152627 582807 152630
rect 214465 152554 214531 152557
rect 229829 152554 229895 152557
rect 214465 152552 217028 152554
rect 214465 152496 214470 152552
rect 214526 152496 217028 152552
rect 214465 152494 217028 152496
rect 228988 152552 229895 152554
rect 228988 152496 229834 152552
rect 229890 152496 229895 152552
rect 228988 152494 229895 152496
rect 214465 152491 214531 152494
rect 229829 152491 229895 152494
rect 264329 152554 264395 152557
rect 264329 152552 268180 152554
rect 264329 152496 264334 152552
rect 264390 152496 268180 152552
rect 583520 152540 584960 152630
rect 264329 152494 268180 152496
rect 264329 152491 264395 152494
rect 230565 152010 230631 152013
rect 228988 152008 230631 152010
rect 228988 151952 230570 152008
rect 230626 151952 230631 152008
rect 228988 151950 230631 151952
rect 230565 151947 230631 151950
rect 258030 151950 268180 152010
rect 213361 151874 213427 151877
rect 254761 151874 254827 151877
rect 258030 151874 258090 151950
rect 281717 151874 281783 151877
rect 213361 151872 217028 151874
rect 213361 151816 213366 151872
rect 213422 151816 217028 151872
rect 213361 151814 217028 151816
rect 254761 151872 258090 151874
rect 254761 151816 254766 151872
rect 254822 151816 258090 151872
rect 254761 151814 258090 151816
rect 279956 151872 281783 151874
rect 279956 151816 281722 151872
rect 281778 151816 281783 151872
rect 279956 151814 281783 151816
rect 213361 151811 213427 151814
rect 254761 151811 254827 151814
rect 281717 151811 281783 151814
rect 231894 151602 231900 151604
rect 228988 151542 231900 151602
rect 231894 151540 231900 151542
rect 231964 151540 231970 151604
rect 268150 151330 268210 151572
rect 258030 151270 268210 151330
rect 214649 151194 214715 151197
rect 214649 151192 217028 151194
rect 214649 151136 214654 151192
rect 214710 151136 217028 151192
rect 214649 151134 217028 151136
rect 214649 151131 214715 151134
rect 170254 150996 170260 151060
rect 170324 151058 170330 151060
rect 215886 151058 215892 151060
rect 170324 150998 215892 151058
rect 170324 150996 170330 150998
rect 215886 150996 215892 150998
rect 215956 150996 215962 151060
rect 230657 151058 230723 151061
rect 228988 151056 230723 151058
rect 228988 151000 230662 151056
rect 230718 151000 230723 151056
rect 228988 150998 230723 151000
rect 230657 150995 230723 150998
rect 233182 150996 233188 151060
rect 233252 151058 233258 151060
rect 241646 151058 241652 151060
rect 233252 150998 241652 151058
rect 233252 150996 233258 150998
rect 241646 150996 241652 150998
rect 241716 150996 241722 151060
rect 250529 150922 250595 150925
rect 258030 150922 258090 151270
rect 264973 151194 265039 151197
rect 282729 151194 282795 151197
rect 264973 151192 268180 151194
rect 264973 151136 264978 151192
rect 265034 151136 268180 151192
rect 264973 151134 268180 151136
rect 279956 151192 282795 151194
rect 279956 151136 282734 151192
rect 282790 151136 282795 151192
rect 279956 151134 282795 151136
rect 264973 151131 265039 151134
rect 282729 151131 282795 151134
rect 250529 150920 258090 150922
rect 250529 150864 250534 150920
rect 250590 150864 258090 150920
rect 250529 150862 258090 150864
rect 250529 150859 250595 150862
rect 265065 150786 265131 150789
rect 265065 150784 268180 150786
rect 265065 150728 265070 150784
rect 265126 150728 268180 150784
rect 265065 150726 268180 150728
rect 265065 150723 265131 150726
rect 232078 150650 232084 150652
rect 228988 150590 232084 150650
rect 232078 150588 232084 150590
rect 232148 150588 232154 150652
rect 213913 150514 213979 150517
rect 213913 150512 217028 150514
rect 213913 150456 213918 150512
rect 213974 150456 217028 150512
rect 213913 150454 217028 150456
rect 213913 150451 213979 150454
rect 282821 150378 282887 150381
rect 279956 150376 282887 150378
rect 229134 150106 229140 150108
rect 228988 150046 229140 150106
rect 229134 150044 229140 150046
rect 229204 150044 229210 150108
rect 242433 150106 242499 150109
rect 268150 150106 268210 150348
rect 279956 150320 282826 150376
rect 282882 150320 282887 150376
rect 279956 150318 282887 150320
rect 282821 150315 282887 150318
rect 242433 150104 268210 150106
rect 242433 150048 242438 150104
rect 242494 150048 268210 150104
rect 242433 150046 268210 150048
rect 242433 150043 242499 150046
rect 264973 149970 265039 149973
rect 264973 149968 268180 149970
rect -960 149834 480 149924
rect 264973 149912 264978 149968
rect 265034 149912 268180 149968
rect 264973 149910 268180 149912
rect 264973 149907 265039 149910
rect 2773 149834 2839 149837
rect -960 149832 2839 149834
rect -960 149776 2778 149832
rect 2834 149776 2839 149832
rect -960 149774 2839 149776
rect -960 149684 480 149774
rect 2773 149771 2839 149774
rect 214005 149834 214071 149837
rect 214005 149832 217028 149834
rect 214005 149776 214010 149832
rect 214066 149776 217028 149832
rect 214005 149774 217028 149776
rect 214005 149771 214071 149774
rect 231117 149698 231183 149701
rect 228988 149696 231183 149698
rect 228988 149640 231122 149696
rect 231178 149640 231183 149696
rect 228988 149638 231183 149640
rect 231117 149635 231183 149638
rect 257521 149698 257587 149701
rect 265065 149698 265131 149701
rect 281901 149698 281967 149701
rect 257521 149696 265131 149698
rect 257521 149640 257526 149696
rect 257582 149640 265070 149696
rect 265126 149640 265131 149696
rect 257521 149638 265131 149640
rect 279956 149696 281967 149698
rect 279956 149640 281906 149696
rect 281962 149640 281967 149696
rect 279956 149638 281967 149640
rect 257521 149635 257587 149638
rect 265065 149635 265131 149638
rect 281901 149635 281967 149638
rect 265157 149562 265223 149565
rect 265157 149560 268180 149562
rect 265157 149504 265162 149560
rect 265218 149504 268180 149560
rect 265157 149502 268180 149504
rect 265157 149499 265223 149502
rect 213913 149154 213979 149157
rect 230565 149154 230631 149157
rect 213913 149152 217028 149154
rect 213913 149096 213918 149152
rect 213974 149096 217028 149152
rect 213913 149094 217028 149096
rect 228988 149152 230631 149154
rect 228988 149096 230570 149152
rect 230626 149096 230631 149152
rect 228988 149094 230631 149096
rect 213913 149091 213979 149094
rect 230565 149091 230631 149094
rect 231301 149154 231367 149157
rect 233734 149154 233740 149156
rect 231301 149152 233740 149154
rect 231301 149096 231306 149152
rect 231362 149096 233740 149152
rect 231301 149094 233740 149096
rect 231301 149091 231367 149094
rect 233734 149092 233740 149094
rect 233804 149092 233810 149156
rect 265065 149018 265131 149021
rect 265065 149016 268180 149018
rect 265065 148960 265070 149016
rect 265126 148960 268180 149016
rect 265065 148958 268180 148960
rect 265065 148955 265131 148958
rect 282729 148882 282795 148885
rect 279956 148880 282795 148882
rect 279956 148824 282734 148880
rect 282790 148824 282795 148880
rect 279956 148822 282795 148824
rect 282729 148819 282795 148822
rect 242985 148746 243051 148749
rect 228988 148744 243051 148746
rect 228988 148688 242990 148744
rect 243046 148688 243051 148744
rect 228988 148686 243051 148688
rect 242985 148683 243051 148686
rect 265709 148610 265775 148613
rect 265709 148608 268180 148610
rect 265709 148552 265714 148608
rect 265770 148552 268180 148608
rect 265709 148550 268180 148552
rect 265709 148547 265775 148550
rect 214557 148474 214623 148477
rect 214557 148472 217028 148474
rect 214557 148416 214562 148472
rect 214618 148416 217028 148472
rect 214557 148414 217028 148416
rect 214557 148411 214623 148414
rect 230749 148202 230815 148205
rect 228988 148200 230815 148202
rect 228988 148144 230754 148200
rect 230810 148144 230815 148200
rect 228988 148142 230815 148144
rect 230749 148139 230815 148142
rect 258030 148142 268180 148202
rect 234102 148004 234108 148068
rect 234172 148066 234178 148068
rect 258030 148066 258090 148142
rect 282821 148066 282887 148069
rect 234172 148006 258090 148066
rect 279956 148064 282887 148066
rect 279956 148008 282826 148064
rect 282882 148008 282887 148064
rect 279956 148006 282887 148008
rect 234172 148004 234178 148006
rect 282821 148003 282887 148006
rect 213913 147930 213979 147933
rect 213913 147928 217028 147930
rect 213913 147872 213918 147928
rect 213974 147872 217028 147928
rect 213913 147870 217028 147872
rect 213913 147867 213979 147870
rect 230565 147794 230631 147797
rect 228988 147792 230631 147794
rect 228988 147736 230570 147792
rect 230626 147736 230631 147792
rect 228988 147734 230631 147736
rect 230565 147731 230631 147734
rect 264973 147794 265039 147797
rect 264973 147792 268180 147794
rect 264973 147736 264978 147792
rect 265034 147736 268180 147792
rect 264973 147734 268180 147736
rect 264973 147731 265039 147734
rect 298134 147732 298140 147796
rect 298204 147794 298210 147796
rect 299381 147794 299447 147797
rect 298204 147792 299447 147794
rect 298204 147736 299386 147792
rect 299442 147736 299447 147792
rect 298204 147734 299447 147736
rect 298204 147732 298210 147734
rect 299381 147731 299447 147734
rect 265065 147386 265131 147389
rect 282821 147386 282887 147389
rect 265065 147384 268180 147386
rect 265065 147328 265070 147384
rect 265126 147328 268180 147384
rect 265065 147326 268180 147328
rect 279956 147384 282887 147386
rect 279956 147328 282826 147384
rect 282882 147328 282887 147384
rect 279956 147326 282887 147328
rect 265065 147323 265131 147326
rect 282821 147323 282887 147326
rect 213269 147250 213335 147253
rect 230749 147250 230815 147253
rect 213269 147248 217028 147250
rect 213269 147192 213274 147248
rect 213330 147192 217028 147248
rect 213269 147190 217028 147192
rect 228988 147248 230815 147250
rect 228988 147192 230754 147248
rect 230810 147192 230815 147248
rect 228988 147190 230815 147192
rect 213269 147187 213335 147190
rect 230749 147187 230815 147190
rect 231158 146916 231164 146980
rect 231228 146978 231234 146980
rect 240869 146978 240935 146981
rect 231228 146976 240935 146978
rect 231228 146920 240874 146976
rect 240930 146920 240935 146976
rect 231228 146918 240935 146920
rect 231228 146916 231234 146918
rect 240869 146915 240935 146918
rect 231761 146842 231827 146845
rect 228988 146840 231827 146842
rect 228988 146784 231766 146840
rect 231822 146784 231827 146840
rect 228988 146782 231827 146784
rect 231761 146779 231827 146782
rect 242341 146706 242407 146709
rect 268150 146706 268210 146948
rect 242341 146704 268210 146706
rect 242341 146648 242346 146704
rect 242402 146648 268210 146704
rect 242341 146646 268210 146648
rect 242341 146643 242407 146646
rect 213913 146570 213979 146573
rect 282729 146570 282795 146573
rect 213913 146568 217028 146570
rect 213913 146512 213918 146568
rect 213974 146512 217028 146568
rect 213913 146510 217028 146512
rect 279956 146568 282795 146570
rect 279956 146512 282734 146568
rect 282790 146512 282795 146568
rect 279956 146510 282795 146512
rect 213913 146507 213979 146510
rect 282729 146507 282795 146510
rect 264973 146434 265039 146437
rect 264973 146432 268180 146434
rect 264973 146376 264978 146432
rect 265034 146376 268180 146432
rect 264973 146374 268180 146376
rect 264973 146371 265039 146374
rect 229737 146298 229803 146301
rect 228988 146296 229803 146298
rect 228988 146240 229742 146296
rect 229798 146240 229803 146296
rect 228988 146238 229803 146240
rect 229737 146235 229803 146238
rect 265065 146026 265131 146029
rect 265065 146024 268180 146026
rect 265065 145968 265070 146024
rect 265126 145968 268180 146024
rect 265065 145966 268180 145968
rect 265065 145963 265131 145966
rect 214005 145890 214071 145893
rect 233785 145890 233851 145893
rect 282821 145890 282887 145893
rect 214005 145888 217028 145890
rect 214005 145832 214010 145888
rect 214066 145832 217028 145888
rect 214005 145830 217028 145832
rect 228988 145888 233851 145890
rect 228988 145832 233790 145888
rect 233846 145832 233851 145888
rect 228988 145830 233851 145832
rect 279956 145888 282887 145890
rect 279956 145832 282826 145888
rect 282882 145832 282887 145888
rect 279956 145830 282887 145832
rect 214005 145827 214071 145830
rect 233785 145827 233851 145830
rect 282821 145827 282887 145830
rect 231669 145754 231735 145757
rect 248413 145754 248479 145757
rect 265157 145754 265223 145757
rect 231669 145752 248479 145754
rect 231669 145696 231674 145752
rect 231730 145696 248418 145752
rect 248474 145696 248479 145752
rect 231669 145694 248479 145696
rect 231669 145691 231735 145694
rect 248413 145691 248479 145694
rect 258030 145752 265223 145754
rect 258030 145696 265162 145752
rect 265218 145696 265223 145752
rect 258030 145694 265223 145696
rect 245193 145618 245259 145621
rect 258030 145618 258090 145694
rect 265157 145691 265223 145694
rect 245193 145616 258090 145618
rect 245193 145560 245198 145616
rect 245254 145560 258090 145616
rect 245193 145558 258090 145560
rect 263133 145618 263199 145621
rect 395981 145618 396047 145621
rect 405917 145618 405983 145621
rect 263133 145616 268180 145618
rect 263133 145560 263138 145616
rect 263194 145560 268180 145616
rect 263133 145558 268180 145560
rect 395981 145616 405983 145618
rect 395981 145560 395986 145616
rect 396042 145560 405922 145616
rect 405978 145560 405983 145616
rect 395981 145558 405983 145560
rect 245193 145555 245259 145558
rect 263133 145555 263199 145558
rect 395981 145555 396047 145558
rect 405917 145555 405983 145558
rect 411437 145618 411503 145621
rect 582649 145618 582715 145621
rect 411437 145616 582715 145618
rect 411437 145560 411442 145616
rect 411498 145560 582654 145616
rect 582710 145560 582715 145616
rect 411437 145558 582715 145560
rect 411437 145555 411503 145558
rect 582649 145555 582715 145558
rect 231301 145346 231367 145349
rect 228988 145344 231367 145346
rect 228988 145288 231306 145344
rect 231362 145288 231367 145344
rect 228988 145286 231367 145288
rect 231301 145283 231367 145286
rect 213913 145210 213979 145213
rect 264973 145210 265039 145213
rect 213913 145208 217028 145210
rect 213913 145152 213918 145208
rect 213974 145152 217028 145208
rect 213913 145150 217028 145152
rect 264973 145208 268180 145210
rect 264973 145152 264978 145208
rect 265034 145152 268180 145208
rect 264973 145150 268180 145152
rect 213913 145147 213979 145150
rect 264973 145147 265039 145150
rect 282545 145074 282611 145077
rect 279956 145072 282611 145074
rect 279956 145016 282550 145072
rect 282606 145016 282611 145072
rect 279956 145014 282611 145016
rect 282545 145011 282611 145014
rect 230657 144938 230723 144941
rect 228988 144936 230723 144938
rect 228988 144880 230662 144936
rect 230718 144880 230723 144936
rect 228988 144878 230723 144880
rect 230657 144875 230723 144878
rect 265065 144802 265131 144805
rect 279325 144802 279391 144805
rect 265065 144800 268180 144802
rect 265065 144744 265070 144800
rect 265126 144744 268180 144800
rect 265065 144742 268180 144744
rect 279325 144800 279434 144802
rect 279325 144744 279330 144800
rect 279386 144744 279434 144800
rect 265065 144739 265131 144742
rect 279325 144739 279434 144744
rect 215937 144530 216003 144533
rect 215937 144528 217028 144530
rect 215937 144472 215942 144528
rect 215998 144472 217028 144528
rect 215937 144470 217028 144472
rect 215937 144467 216003 144470
rect 231669 144394 231735 144397
rect 228988 144392 231735 144394
rect 228988 144336 231674 144392
rect 231730 144336 231735 144392
rect 228988 144334 231735 144336
rect 231669 144331 231735 144334
rect 264973 144394 265039 144397
rect 264973 144392 268180 144394
rect 264973 144336 264978 144392
rect 265034 144336 268180 144392
rect 264973 144334 268180 144336
rect 264973 144331 265039 144334
rect 279374 144228 279434 144739
rect 229645 144122 229711 144125
rect 245929 144122 245995 144125
rect 229645 144120 245995 144122
rect 229645 144064 229650 144120
rect 229706 144064 245934 144120
rect 245990 144064 245995 144120
rect 229645 144062 245995 144064
rect 229645 144059 229711 144062
rect 245929 144059 245995 144062
rect 231761 143986 231827 143989
rect 228988 143984 231827 143986
rect 228988 143928 231766 143984
rect 231822 143928 231827 143984
rect 228988 143926 231827 143928
rect 231761 143923 231827 143926
rect 213913 143850 213979 143853
rect 265157 143850 265223 143853
rect 213913 143848 217028 143850
rect 213913 143792 213918 143848
rect 213974 143792 217028 143848
rect 213913 143790 217028 143792
rect 265157 143848 268180 143850
rect 265157 143792 265162 143848
rect 265218 143792 268180 143848
rect 265157 143790 268180 143792
rect 213913 143787 213979 143790
rect 265157 143787 265223 143790
rect 282453 143578 282519 143581
rect 279956 143576 282519 143578
rect 279956 143520 282458 143576
rect 282514 143520 282519 143576
rect 279956 143518 282519 143520
rect 282453 143515 282519 143518
rect 231761 143442 231827 143445
rect 228988 143440 231827 143442
rect 228988 143384 231766 143440
rect 231822 143384 231827 143440
rect 228988 143382 231827 143384
rect 231761 143379 231827 143382
rect 265801 143442 265867 143445
rect 409873 143444 409939 143445
rect 409822 143442 409828 143444
rect 265801 143440 268180 143442
rect 265801 143384 265806 143440
rect 265862 143384 268180 143440
rect 265801 143382 268180 143384
rect 409746 143382 409828 143442
rect 409892 143442 409939 143444
rect 410885 143442 410951 143445
rect 409892 143440 410951 143442
rect 409934 143384 410890 143440
rect 410946 143384 410951 143440
rect 265801 143379 265867 143382
rect 409822 143380 409828 143382
rect 409892 143382 410951 143384
rect 409892 143380 409939 143382
rect 409873 143379 409939 143380
rect 410885 143379 410951 143382
rect 417366 143380 417372 143444
rect 417436 143442 417442 143444
rect 420913 143442 420979 143445
rect 422109 143442 422175 143445
rect 417436 143440 422175 143442
rect 417436 143384 420918 143440
rect 420974 143384 422114 143440
rect 422170 143384 422175 143440
rect 417436 143382 422175 143384
rect 417436 143380 417442 143382
rect 420913 143379 420979 143382
rect 422109 143379 422175 143382
rect 214005 143306 214071 143309
rect 214005 143304 217028 143306
rect 214005 143248 214010 143304
rect 214066 143248 217028 143304
rect 214005 143246 217028 143248
rect 214005 143243 214071 143246
rect 230381 143034 230447 143037
rect 228988 143032 230447 143034
rect 228988 142976 230386 143032
rect 230442 142976 230447 143032
rect 228988 142974 230447 142976
rect 230381 142971 230447 142974
rect 230974 142700 230980 142764
rect 231044 142762 231050 142764
rect 255957 142762 256023 142765
rect 231044 142760 256023 142762
rect 231044 142704 255962 142760
rect 256018 142704 256023 142760
rect 231044 142702 256023 142704
rect 231044 142700 231050 142702
rect 255957 142699 256023 142702
rect 256141 142762 256207 142765
rect 268150 142762 268210 143004
rect 282821 142762 282887 142765
rect 256141 142760 268210 142762
rect 256141 142704 256146 142760
rect 256202 142704 268210 142760
rect 256141 142702 268210 142704
rect 279956 142760 282887 142762
rect 279956 142704 282826 142760
rect 282882 142704 282887 142760
rect 279956 142702 282887 142704
rect 256141 142699 256207 142702
rect 282821 142699 282887 142702
rect 213913 142626 213979 142629
rect 264605 142626 264671 142629
rect 213913 142624 217028 142626
rect 213913 142568 213918 142624
rect 213974 142568 217028 142624
rect 213913 142566 217028 142568
rect 264605 142624 268180 142626
rect 264605 142568 264610 142624
rect 264666 142568 268180 142624
rect 264605 142566 268180 142568
rect 213913 142563 213979 142566
rect 264605 142563 264671 142566
rect 233182 142490 233188 142492
rect 228988 142430 233188 142490
rect 233182 142428 233188 142430
rect 233252 142428 233258 142492
rect 356697 142490 356763 142493
rect 406285 142490 406351 142493
rect 356697 142488 406351 142490
rect 356697 142432 356702 142488
rect 356758 142432 406290 142488
rect 406346 142432 406351 142488
rect 356697 142430 406351 142432
rect 356697 142427 356763 142430
rect 406285 142427 406351 142430
rect 396717 142354 396783 142357
rect 427813 142354 427879 142357
rect 396717 142352 427879 142354
rect 396717 142296 396722 142352
rect 396778 142296 427818 142352
rect 427874 142296 427879 142352
rect 396717 142294 427879 142296
rect 396717 142291 396783 142294
rect 427813 142291 427879 142294
rect 264973 142218 265039 142221
rect 395521 142218 395587 142221
rect 400765 142218 400831 142221
rect 431953 142220 432019 142221
rect 431902 142218 431908 142220
rect 264973 142216 268180 142218
rect 264973 142160 264978 142216
rect 265034 142160 268180 142216
rect 264973 142158 268180 142160
rect 395521 142216 400831 142218
rect 395521 142160 395526 142216
rect 395582 142160 400770 142216
rect 400826 142160 400831 142216
rect 395521 142158 400831 142160
rect 431826 142158 431908 142218
rect 431972 142218 432019 142220
rect 432965 142218 433031 142221
rect 431972 142216 433031 142218
rect 432014 142160 432970 142216
rect 433026 142160 433031 142216
rect 264973 142155 265039 142158
rect 395521 142155 395587 142158
rect 400765 142155 400831 142158
rect 431902 142156 431908 142158
rect 431972 142158 433031 142160
rect 431972 142156 432019 142158
rect 431953 142155 432019 142156
rect 432965 142155 433031 142158
rect 238702 142082 238708 142084
rect 228988 142022 238708 142082
rect 238702 142020 238708 142022
rect 238772 142020 238778 142084
rect 282821 142082 282887 142085
rect 279956 142080 282887 142082
rect 279956 142024 282826 142080
rect 282882 142024 282887 142080
rect 279956 142022 282887 142024
rect 282821 142019 282887 142022
rect 213913 141946 213979 141949
rect 213913 141944 217028 141946
rect 213913 141888 213918 141944
rect 213974 141888 217028 141944
rect 213913 141886 217028 141888
rect 213913 141883 213979 141886
rect 265893 141810 265959 141813
rect 265893 141808 268180 141810
rect 265893 141752 265898 141808
rect 265954 141752 268180 141808
rect 265893 141750 268180 141752
rect 265893 141747 265959 141750
rect 229645 141674 229711 141677
rect 228988 141672 229711 141674
rect 228988 141616 229650 141672
rect 229706 141616 229711 141672
rect 228988 141614 229711 141616
rect 229645 141611 229711 141614
rect 247861 141402 247927 141405
rect 265157 141402 265223 141405
rect 247861 141400 265223 141402
rect 247861 141344 247866 141400
rect 247922 141344 265162 141400
rect 265218 141344 265223 141400
rect 247861 141342 265223 141344
rect 247861 141339 247927 141342
rect 265157 141339 265223 141342
rect 214557 141266 214623 141269
rect 266077 141266 266143 141269
rect 282729 141266 282795 141269
rect 214557 141264 217028 141266
rect 214557 141208 214562 141264
rect 214618 141208 217028 141264
rect 214557 141206 217028 141208
rect 266077 141264 268180 141266
rect 266077 141208 266082 141264
rect 266138 141208 268180 141264
rect 266077 141206 268180 141208
rect 279956 141264 282795 141266
rect 279956 141208 282734 141264
rect 282790 141208 282795 141264
rect 279956 141206 282795 141208
rect 214557 141203 214623 141206
rect 266077 141203 266143 141206
rect 282729 141203 282795 141206
rect 248638 141130 248644 141132
rect 228988 141070 248644 141130
rect 248638 141068 248644 141070
rect 248708 141068 248714 141132
rect 264973 140858 265039 140861
rect 303613 140860 303679 140861
rect 264973 140856 268180 140858
rect 264973 140800 264978 140856
rect 265034 140800 268180 140856
rect 264973 140798 268180 140800
rect 303613 140856 303660 140860
rect 303724 140858 303730 140860
rect 329097 140858 329163 140861
rect 426525 140858 426591 140861
rect 303613 140800 303618 140856
rect 264973 140795 265039 140798
rect 303613 140796 303660 140800
rect 303724 140798 303770 140858
rect 329097 140856 426591 140858
rect 329097 140800 329102 140856
rect 329158 140800 426530 140856
rect 426586 140800 426591 140856
rect 329097 140798 426591 140800
rect 303724 140796 303730 140798
rect 303613 140795 303679 140796
rect 329097 140795 329163 140798
rect 426525 140795 426591 140798
rect 435357 140858 435423 140861
rect 440509 140858 440575 140861
rect 441705 140860 441771 140861
rect 435357 140856 440575 140858
rect 435357 140800 435362 140856
rect 435418 140800 440514 140856
rect 440570 140800 440575 140856
rect 435357 140798 440575 140800
rect 435357 140795 435423 140798
rect 440509 140795 440575 140798
rect 441654 140796 441660 140860
rect 441724 140858 441771 140860
rect 441724 140856 441816 140858
rect 441766 140800 441816 140856
rect 441724 140798 441816 140800
rect 441724 140796 441771 140798
rect 441705 140795 441771 140796
rect 229093 140722 229159 140725
rect 228988 140720 229159 140722
rect 228988 140664 229098 140720
rect 229154 140664 229159 140720
rect 228988 140662 229159 140664
rect 229093 140659 229159 140662
rect 213913 140586 213979 140589
rect 213913 140584 217028 140586
rect 213913 140528 213918 140584
rect 213974 140528 217028 140584
rect 213913 140526 217028 140528
rect 213913 140523 213979 140526
rect 266854 140388 266860 140452
rect 266924 140450 266930 140452
rect 282821 140450 282887 140453
rect 266924 140390 268180 140450
rect 279956 140448 282887 140450
rect 279956 140392 282826 140448
rect 282882 140392 282887 140448
rect 279956 140390 282887 140392
rect 266924 140388 266930 140390
rect 282821 140387 282887 140390
rect 245745 140178 245811 140181
rect 228988 140176 245811 140178
rect 228988 140120 245750 140176
rect 245806 140120 245811 140176
rect 228988 140118 245811 140120
rect 245745 140115 245811 140118
rect 264973 140042 265039 140045
rect 433977 140042 434043 140045
rect 440417 140042 440483 140045
rect 264973 140040 268180 140042
rect 264973 139984 264978 140040
rect 265034 139984 268180 140040
rect 264973 139982 268180 139984
rect 433977 140040 440483 140042
rect 433977 139984 433982 140040
rect 434038 139984 440422 140040
rect 440478 139984 440483 140040
rect 433977 139982 440483 139984
rect 264973 139979 265039 139982
rect 433977 139979 434043 139982
rect 440417 139979 440483 139982
rect 213177 139906 213243 139909
rect 213177 139904 217028 139906
rect 213177 139848 213182 139904
rect 213238 139848 217028 139904
rect 213177 139846 217028 139848
rect 213177 139843 213243 139846
rect 231894 139770 231900 139772
rect 228988 139710 231900 139770
rect 231894 139708 231900 139710
rect 231964 139708 231970 139772
rect 280102 139770 280108 139772
rect 279956 139710 280108 139770
rect 280102 139708 280108 139710
rect 280172 139708 280178 139772
rect 419022 139708 419028 139772
rect 419092 139770 419098 139772
rect 420545 139770 420611 139773
rect 419092 139768 420611 139770
rect 419092 139712 420550 139768
rect 420606 139712 420611 139768
rect 419092 139710 420611 139712
rect 419092 139708 419098 139710
rect 420545 139707 420611 139710
rect 419901 139634 419967 139637
rect 420678 139634 420684 139636
rect 258030 139574 268180 139634
rect 419901 139632 420684 139634
rect 419901 139576 419906 139632
rect 419962 139576 420684 139632
rect 419901 139574 420684 139576
rect 239397 139498 239463 139501
rect 258030 139498 258090 139574
rect 419901 139571 419967 139574
rect 420678 139572 420684 139574
rect 420748 139572 420754 139636
rect 239397 139496 258090 139498
rect 239397 139440 239402 139496
rect 239458 139440 258090 139496
rect 239397 139438 258090 139440
rect 322197 139498 322263 139501
rect 418705 139498 418771 139501
rect 322197 139496 418771 139498
rect 322197 139440 322202 139496
rect 322258 139440 418710 139496
rect 418766 139440 418771 139496
rect 322197 139438 418771 139440
rect 239397 139435 239463 139438
rect 322197 139435 322263 139438
rect 418705 139435 418771 139438
rect 420545 139498 420611 139501
rect 421046 139498 421052 139500
rect 420545 139496 421052 139498
rect 420545 139440 420550 139496
rect 420606 139440 421052 139496
rect 420545 139438 421052 139440
rect 420545 139435 420611 139438
rect 421046 139436 421052 139438
rect 421116 139436 421122 139500
rect 426382 139436 426388 139500
rect 426452 139498 426458 139500
rect 426893 139498 426959 139501
rect 426452 139496 426959 139498
rect 426452 139440 426898 139496
rect 426954 139440 426959 139496
rect 426452 139438 426959 139440
rect 426452 139436 426458 139438
rect 426893 139435 426959 139438
rect 427854 139436 427860 139500
rect 427924 139498 427930 139500
rect 428733 139498 428799 139501
rect 427924 139496 428799 139498
rect 427924 139440 428738 139496
rect 428794 139440 428799 139496
rect 427924 139438 428799 139440
rect 427924 139436 427930 139438
rect 428733 139435 428799 139438
rect 429142 139436 429148 139500
rect 429212 139498 429218 139500
rect 429469 139498 429535 139501
rect 429212 139496 429535 139498
rect 429212 139440 429474 139496
rect 429530 139440 429535 139496
rect 429212 139438 429535 139440
rect 429212 139436 429218 139438
rect 429469 139435 429535 139438
rect 434989 139500 435055 139501
rect 439037 139500 439103 139501
rect 434989 139496 435036 139500
rect 435100 139498 435106 139500
rect 434989 139440 434994 139496
rect 434989 139436 435036 139440
rect 435100 139438 435146 139498
rect 439037 139496 439084 139500
rect 439148 139498 439154 139500
rect 439037 139440 439042 139496
rect 435100 139436 435106 139438
rect 439037 139436 439084 139440
rect 439148 139438 439194 139498
rect 439148 139436 439154 139438
rect 434989 139435 435055 139436
rect 439037 139435 439103 139436
rect 380893 139362 380959 139365
rect 397545 139362 397611 139365
rect 580165 139362 580231 139365
rect 583520 139362 584960 139452
rect 380893 139360 393330 139362
rect 380893 139304 380898 139360
rect 380954 139304 393330 139360
rect 380893 139302 393330 139304
rect 380893 139299 380959 139302
rect 214005 139226 214071 139229
rect 234654 139226 234660 139228
rect 214005 139224 217028 139226
rect 214005 139168 214010 139224
rect 214066 139168 217028 139224
rect 214005 139166 217028 139168
rect 228988 139166 234660 139226
rect 214005 139163 214071 139166
rect 234654 139164 234660 139166
rect 234724 139164 234730 139228
rect 264329 139226 264395 139229
rect 264329 139224 268180 139226
rect 264329 139168 264334 139224
rect 264390 139168 268180 139224
rect 264329 139166 268180 139168
rect 264329 139163 264395 139166
rect 281717 138954 281783 138957
rect 279956 138952 281783 138954
rect 279956 138896 281722 138952
rect 281778 138896 281783 138952
rect 279956 138894 281783 138896
rect 393270 138954 393330 139302
rect 397545 139360 400108 139362
rect 397545 139304 397550 139360
rect 397606 139304 400108 139360
rect 397545 139302 400108 139304
rect 580165 139360 584960 139362
rect 580165 139304 580170 139360
rect 580226 139304 584960 139360
rect 580165 139302 584960 139304
rect 397545 139299 397611 139302
rect 580165 139299 580231 139302
rect 583520 139212 584960 139302
rect 393270 138894 400138 138954
rect 281717 138891 281783 138894
rect 237414 138818 237420 138820
rect 228988 138758 237420 138818
rect 237414 138756 237420 138758
rect 237484 138756 237490 138820
rect 213913 138682 213979 138685
rect 264973 138682 265039 138685
rect 352649 138682 352715 138685
rect 380893 138682 380959 138685
rect 213913 138680 217028 138682
rect 213913 138624 213918 138680
rect 213974 138624 217028 138680
rect 213913 138622 217028 138624
rect 264973 138680 268180 138682
rect 264973 138624 264978 138680
rect 265034 138624 268180 138680
rect 264973 138622 268180 138624
rect 352649 138680 380959 138682
rect 352649 138624 352654 138680
rect 352710 138624 380898 138680
rect 380954 138624 380959 138680
rect 352649 138622 380959 138624
rect 213913 138619 213979 138622
rect 264973 138619 265039 138622
rect 352649 138619 352715 138622
rect 380893 138619 380959 138622
rect 231761 138274 231827 138277
rect 282637 138274 282703 138277
rect 228988 138272 231827 138274
rect 228988 138216 231766 138272
rect 231822 138216 231827 138272
rect 228988 138214 231827 138216
rect 231761 138211 231827 138214
rect 258030 138214 268180 138274
rect 279956 138272 282703 138274
rect 279956 138216 282642 138272
rect 282698 138216 282703 138272
rect 400078 138244 400138 138894
rect 439822 138682 439882 138924
rect 441654 138682 441660 138684
rect 439822 138622 441660 138682
rect 441654 138620 441660 138622
rect 441724 138682 441730 138684
rect 447317 138682 447383 138685
rect 441724 138680 447383 138682
rect 441724 138624 447322 138680
rect 447378 138624 447383 138680
rect 441724 138622 447383 138624
rect 441724 138620 441730 138622
rect 447317 138619 447383 138622
rect 442165 138274 442231 138277
rect 439852 138272 442231 138274
rect 279956 138214 282703 138216
rect 439852 138216 442170 138272
rect 442226 138216 442231 138272
rect 439852 138214 442231 138216
rect 243537 138138 243603 138141
rect 258030 138138 258090 138214
rect 282637 138211 282703 138214
rect 442165 138211 442231 138214
rect 243537 138136 258090 138138
rect 243537 138080 243542 138136
rect 243598 138080 258090 138136
rect 243537 138078 258090 138080
rect 243537 138075 243603 138078
rect 214097 138002 214163 138005
rect 214097 138000 217028 138002
rect 214097 137944 214102 138000
rect 214158 137944 217028 138000
rect 214097 137942 217028 137944
rect 214097 137939 214163 137942
rect 231761 137866 231827 137869
rect 228988 137864 231827 137866
rect 228988 137808 231766 137864
rect 231822 137808 231827 137864
rect 228988 137806 231827 137808
rect 231761 137803 231827 137806
rect 262765 137594 262831 137597
rect 268150 137594 268210 137836
rect 335353 137730 335419 137733
rect 399845 137730 399911 137733
rect 335353 137728 399911 137730
rect 335353 137672 335358 137728
rect 335414 137672 399850 137728
rect 399906 137672 399911 137728
rect 335353 137670 399911 137672
rect 335353 137667 335419 137670
rect 399845 137667 399911 137670
rect 262765 137592 268210 137594
rect 262765 137536 262770 137592
rect 262826 137536 268210 137592
rect 262765 137534 268210 137536
rect 262765 137531 262831 137534
rect 282821 137458 282887 137461
rect 258030 137398 268180 137458
rect 279956 137456 282887 137458
rect 279956 137400 282826 137456
rect 282882 137400 282887 137456
rect 279956 137398 282887 137400
rect 213913 137322 213979 137325
rect 229686 137322 229692 137324
rect 213913 137320 217028 137322
rect 213913 137264 213918 137320
rect 213974 137264 217028 137320
rect 213913 137262 217028 137264
rect 228988 137262 229692 137322
rect 213913 137259 213979 137262
rect 229686 137260 229692 137262
rect 229756 137260 229762 137324
rect 236494 137260 236500 137324
rect 236564 137322 236570 137324
rect 258030 137322 258090 137398
rect 282821 137395 282887 137398
rect 236564 137262 258090 137322
rect 397913 137322 397979 137325
rect 397913 137320 400108 137322
rect 397913 137264 397918 137320
rect 397974 137264 400108 137320
rect 397913 137262 400108 137264
rect 236564 137260 236570 137262
rect 397913 137259 397979 137262
rect 229870 137124 229876 137188
rect 229940 137186 229946 137188
rect 262765 137186 262831 137189
rect 442901 137186 442967 137189
rect 229940 137184 262831 137186
rect 229940 137128 262770 137184
rect 262826 137128 262831 137184
rect 229940 137126 262831 137128
rect 439852 137184 442967 137186
rect 439852 137128 442906 137184
rect 442962 137128 442967 137184
rect 439852 137126 442967 137128
rect 229940 137124 229946 137126
rect 262765 137123 262831 137126
rect 442901 137123 442967 137126
rect 264973 137050 265039 137053
rect 264973 137048 268180 137050
rect 264973 136992 264978 137048
rect 265034 136992 268180 137048
rect 264973 136990 268180 136992
rect 264973 136987 265039 136990
rect 229737 136914 229803 136917
rect 228988 136912 229803 136914
rect -960 136778 480 136868
rect 228988 136856 229742 136912
rect 229798 136856 229803 136912
rect 228988 136854 229803 136856
rect 229737 136851 229803 136854
rect 3509 136778 3575 136781
rect -960 136776 3575 136778
rect -960 136720 3514 136776
rect 3570 136720 3575 136776
rect -960 136718 3575 136720
rect -960 136628 480 136718
rect 3509 136715 3575 136718
rect 211981 136642 212047 136645
rect 282177 136642 282243 136645
rect 211981 136640 217028 136642
rect 211981 136584 211986 136640
rect 212042 136584 217028 136640
rect 279956 136640 282243 136642
rect 211981 136582 217028 136584
rect 211981 136579 212047 136582
rect 230565 136370 230631 136373
rect 228988 136368 230631 136370
rect 228988 136312 230570 136368
rect 230626 136312 230631 136368
rect 228988 136310 230631 136312
rect 230565 136307 230631 136310
rect 262673 136370 262739 136373
rect 268150 136370 268210 136612
rect 279956 136584 282182 136640
rect 282238 136584 282243 136640
rect 279956 136582 282243 136584
rect 282177 136579 282243 136582
rect 262673 136368 268210 136370
rect 262673 136312 262678 136368
rect 262734 136312 268210 136368
rect 262673 136310 268210 136312
rect 262673 136307 262739 136310
rect 264973 136234 265039 136237
rect 397637 136234 397703 136237
rect 442901 136234 442967 136237
rect 264973 136232 268180 136234
rect 264973 136176 264978 136232
rect 265034 136176 268180 136232
rect 264973 136174 268180 136176
rect 397637 136232 400108 136234
rect 397637 136176 397642 136232
rect 397698 136176 400108 136232
rect 397637 136174 400108 136176
rect 439852 136232 442967 136234
rect 439852 136176 442906 136232
rect 442962 136176 442967 136232
rect 439852 136174 442967 136176
rect 264973 136171 265039 136174
rect 397637 136171 397703 136174
rect 442901 136171 442967 136174
rect 231209 135962 231275 135965
rect 228988 135960 231275 135962
rect 206369 135554 206435 135557
rect 216998 135554 217058 135932
rect 228988 135904 231214 135960
rect 231270 135904 231275 135960
rect 228988 135902 231275 135904
rect 231209 135899 231275 135902
rect 245285 135962 245351 135965
rect 282821 135962 282887 135965
rect 245285 135960 262874 135962
rect 245285 135904 245290 135960
rect 245346 135904 262874 135960
rect 245285 135902 262874 135904
rect 279956 135960 282887 135962
rect 279956 135904 282826 135960
rect 282882 135904 282887 135960
rect 279956 135902 282887 135904
rect 245285 135899 245351 135902
rect 235257 135826 235323 135829
rect 262673 135826 262739 135829
rect 235257 135824 262739 135826
rect 235257 135768 235262 135824
rect 235318 135768 262678 135824
rect 262734 135768 262739 135824
rect 235257 135766 262739 135768
rect 235257 135763 235323 135766
rect 262673 135763 262739 135766
rect 206369 135552 217058 135554
rect 206369 135496 206374 135552
rect 206430 135496 217058 135552
rect 206369 135494 217058 135496
rect 262814 135554 262874 135902
rect 282821 135899 282887 135902
rect 265065 135690 265131 135693
rect 265065 135688 268180 135690
rect 265065 135632 265070 135688
rect 265126 135632 268180 135688
rect 265065 135630 268180 135632
rect 265065 135627 265131 135630
rect 262814 135494 267750 135554
rect 206369 135491 206435 135494
rect 231301 135418 231367 135421
rect 228988 135416 231367 135418
rect 228988 135360 231306 135416
rect 231362 135360 231367 135416
rect 228988 135358 231367 135360
rect 267690 135418 267750 135494
rect 397545 135418 397611 135421
rect 267690 135358 268210 135418
rect 231301 135355 231367 135358
rect 214833 135282 214899 135285
rect 214833 135280 217028 135282
rect 214833 135224 214838 135280
rect 214894 135224 217028 135280
rect 268150 135252 268210 135358
rect 397545 135416 400108 135418
rect 397545 135360 397550 135416
rect 397606 135360 400108 135416
rect 397545 135358 400108 135360
rect 397545 135355 397611 135358
rect 214833 135222 217028 135224
rect 214833 135219 214899 135222
rect 282821 135146 282887 135149
rect 279956 135144 282887 135146
rect 279956 135088 282826 135144
rect 282882 135088 282887 135144
rect 279956 135086 282887 135088
rect 282821 135083 282887 135086
rect 400254 135084 400260 135148
rect 400324 135084 400330 135148
rect 442901 135146 442967 135149
rect 439852 135144 442967 135146
rect 439852 135088 442906 135144
rect 442962 135088 442967 135144
rect 439852 135086 442967 135088
rect 231761 135010 231827 135013
rect 228988 135008 231827 135010
rect 228988 134952 231766 135008
rect 231822 134952 231827 135008
rect 228988 134950 231827 134952
rect 231761 134947 231827 134950
rect 262806 134812 262812 134876
rect 262876 134874 262882 134876
rect 262876 134814 268180 134874
rect 262876 134812 262882 134814
rect 397637 134738 397703 134741
rect 400262 134738 400322 135084
rect 442901 135083 442967 135086
rect 397637 134736 400322 134738
rect 397637 134680 397642 134736
rect 397698 134708 400322 134736
rect 397698 134680 400292 134708
rect 397637 134678 400292 134680
rect 397637 134675 397703 134678
rect 213913 134602 213979 134605
rect 213913 134600 217028 134602
rect 213913 134544 213918 134600
rect 213974 134544 217028 134600
rect 213913 134542 217028 134544
rect 213913 134539 213979 134542
rect 231158 134466 231164 134468
rect 228988 134406 231164 134466
rect 231158 134404 231164 134406
rect 231228 134404 231234 134468
rect 266997 134466 267063 134469
rect 282453 134466 282519 134469
rect 266997 134464 268180 134466
rect 266997 134408 267002 134464
rect 267058 134408 268180 134464
rect 266997 134406 268180 134408
rect 279956 134464 282519 134466
rect 279956 134408 282458 134464
rect 282514 134408 282519 134464
rect 279956 134406 282519 134408
rect 266997 134403 267063 134406
rect 282453 134403 282519 134406
rect 376753 134466 376819 134469
rect 395429 134466 395495 134469
rect 443177 134466 443243 134469
rect 376753 134464 395495 134466
rect 376753 134408 376758 134464
rect 376814 134408 395434 134464
rect 395490 134408 395495 134464
rect 376753 134406 395495 134408
rect 439852 134464 443243 134466
rect 439852 134408 443182 134464
rect 443238 134408 443243 134464
rect 439852 134406 443243 134408
rect 376753 134403 376819 134406
rect 395429 134403 395495 134406
rect 443177 134403 443243 134406
rect 231485 134058 231551 134061
rect 228988 134056 231551 134058
rect 228988 134000 231490 134056
rect 231546 134000 231551 134056
rect 228988 133998 231551 134000
rect 231485 133995 231551 133998
rect 258030 133998 268180 134058
rect 189717 133922 189783 133925
rect 189717 133920 217028 133922
rect 189717 133864 189722 133920
rect 189778 133864 217028 133920
rect 189717 133862 217028 133864
rect 189717 133859 189783 133862
rect 249006 133860 249012 133924
rect 249076 133922 249082 133924
rect 258030 133922 258090 133998
rect 249076 133862 258090 133922
rect 249076 133860 249082 133862
rect 229737 133650 229803 133653
rect 230422 133650 230428 133652
rect 229737 133648 230428 133650
rect 229737 133592 229742 133648
rect 229798 133592 230428 133648
rect 229737 133590 230428 133592
rect 229737 133587 229803 133590
rect 230422 133588 230428 133590
rect 230492 133588 230498 133652
rect 284518 133650 284524 133652
rect 242249 133514 242315 133517
rect 228988 133512 242315 133514
rect 228988 133456 242254 133512
rect 242310 133456 242315 133512
rect 228988 133454 242315 133456
rect 242249 133451 242315 133454
rect 214005 133378 214071 133381
rect 214005 133376 217028 133378
rect 214005 133320 214010 133376
rect 214066 133320 217028 133376
rect 214005 133318 217028 133320
rect 214005 133315 214071 133318
rect 262765 133242 262831 133245
rect 268150 133242 268210 133620
rect 279956 133590 284524 133650
rect 284518 133588 284524 133590
rect 284588 133588 284594 133652
rect 397545 133514 397611 133517
rect 397545 133512 400108 133514
rect 397545 133456 397550 133512
rect 397606 133456 400108 133512
rect 397545 133454 400108 133456
rect 397545 133451 397611 133454
rect 279325 133378 279391 133381
rect 279325 133376 279434 133378
rect 279325 133320 279330 133376
rect 279386 133320 279434 133376
rect 279325 133315 279434 133320
rect 262765 133240 268210 133242
rect 262765 133184 262770 133240
rect 262826 133184 268210 133240
rect 262765 133182 268210 133184
rect 262765 133179 262831 133182
rect 231485 133106 231551 133109
rect 228988 133104 231551 133106
rect 228988 133048 231490 133104
rect 231546 133048 231551 133104
rect 228988 133046 231551 133048
rect 231485 133043 231551 133046
rect 258030 133046 268180 133106
rect 253197 132970 253263 132973
rect 258030 132970 258090 133046
rect 253197 132968 258090 132970
rect 253197 132912 253202 132968
rect 253258 132912 258090 132968
rect 253197 132910 258090 132912
rect 253197 132907 253263 132910
rect 246665 132834 246731 132837
rect 262765 132834 262831 132837
rect 246665 132832 262831 132834
rect 246665 132776 246670 132832
rect 246726 132776 262770 132832
rect 262826 132776 262831 132832
rect 279374 132804 279434 133315
rect 442901 133242 442967 133245
rect 439852 133240 442967 133242
rect 439852 133184 442906 133240
rect 442962 133184 442967 133240
rect 439852 133182 442967 133184
rect 442901 133179 442967 133182
rect 246665 132774 262831 132776
rect 246665 132771 246731 132774
rect 262765 132771 262831 132774
rect 213913 132698 213979 132701
rect 264973 132698 265039 132701
rect 395429 132698 395495 132701
rect 213913 132696 217028 132698
rect 213913 132640 213918 132696
rect 213974 132640 217028 132696
rect 213913 132638 217028 132640
rect 264973 132696 268180 132698
rect 264973 132640 264978 132696
rect 265034 132640 268180 132696
rect 264973 132638 268180 132640
rect 395429 132696 400108 132698
rect 395429 132640 395434 132696
rect 395490 132640 400108 132696
rect 395429 132638 400108 132640
rect 213913 132635 213979 132638
rect 264973 132635 265039 132638
rect 395429 132635 395495 132638
rect 231393 132562 231459 132565
rect 228988 132560 231459 132562
rect 228988 132504 231398 132560
rect 231454 132504 231459 132560
rect 228988 132502 231459 132504
rect 231393 132499 231459 132502
rect 253473 132426 253539 132429
rect 442901 132426 442967 132429
rect 238710 132424 253539 132426
rect 238710 132368 253478 132424
rect 253534 132368 253539 132424
rect 238710 132366 253539 132368
rect 439852 132424 442967 132426
rect 439852 132368 442906 132424
rect 442962 132368 442967 132424
rect 439852 132366 442967 132368
rect 238710 132154 238770 132366
rect 253473 132363 253539 132366
rect 442901 132363 442967 132366
rect 228988 132094 238770 132154
rect 213913 132018 213979 132021
rect 268150 132018 268210 132260
rect 282126 132154 282132 132156
rect 279956 132094 282132 132154
rect 282126 132092 282132 132094
rect 282196 132092 282202 132156
rect 439957 132018 440023 132021
rect 213913 132016 217028 132018
rect 213913 131960 213918 132016
rect 213974 131960 217028 132016
rect 213913 131958 217028 131960
rect 258030 131958 268210 132018
rect 439822 132016 440023 132018
rect 439822 131960 439962 132016
rect 440018 131960 440023 132016
rect 439822 131958 440023 131960
rect 213913 131955 213979 131958
rect 169017 131746 169083 131749
rect 191189 131746 191255 131749
rect 169017 131744 191255 131746
rect 169017 131688 169022 131744
rect 169078 131688 191194 131744
rect 191250 131688 191255 131744
rect 169017 131686 191255 131688
rect 169017 131683 169083 131686
rect 191189 131683 191255 131686
rect 231761 131610 231827 131613
rect 258030 131610 258090 131958
rect 265065 131882 265131 131885
rect 265065 131880 268180 131882
rect 265065 131824 265070 131880
rect 265126 131824 268180 131880
rect 265065 131822 268180 131824
rect 265065 131819 265131 131822
rect 398465 131746 398531 131749
rect 398465 131744 400108 131746
rect 398465 131688 398470 131744
rect 398526 131688 400108 131744
rect 439822 131716 439882 131958
rect 439957 131955 440023 131958
rect 398465 131686 400108 131688
rect 398465 131683 398531 131686
rect 228988 131608 231827 131610
rect 228988 131552 231766 131608
rect 231822 131552 231827 131608
rect 228988 131550 231827 131552
rect 231761 131547 231827 131550
rect 238710 131550 258090 131610
rect 229921 131474 229987 131477
rect 238710 131474 238770 131550
rect 229921 131472 238770 131474
rect 229921 131416 229926 131472
rect 229982 131416 238770 131472
rect 229921 131414 238770 131416
rect 264973 131474 265039 131477
rect 264973 131472 268180 131474
rect 264973 131416 264978 131472
rect 265034 131416 268180 131472
rect 264973 131414 268180 131416
rect 229921 131411 229987 131414
rect 264973 131411 265039 131414
rect 214649 131338 214715 131341
rect 282821 131338 282887 131341
rect 214649 131336 217028 131338
rect 214649 131280 214654 131336
rect 214710 131280 217028 131336
rect 214649 131278 217028 131280
rect 279956 131336 282887 131338
rect 279956 131280 282826 131336
rect 282882 131280 282887 131336
rect 279956 131278 282887 131280
rect 214649 131275 214715 131278
rect 282821 131275 282887 131278
rect 231393 131202 231459 131205
rect 228988 131200 231459 131202
rect 228988 131144 231398 131200
rect 231454 131144 231459 131200
rect 228988 131142 231459 131144
rect 231393 131139 231459 131142
rect 213913 130658 213979 130661
rect 231117 130658 231183 130661
rect 213913 130656 217028 130658
rect 213913 130600 213918 130656
rect 213974 130600 217028 130656
rect 213913 130598 217028 130600
rect 228988 130656 231183 130658
rect 228988 130600 231122 130656
rect 231178 130600 231183 130656
rect 228988 130598 231183 130600
rect 213913 130595 213979 130598
rect 231117 130595 231183 130598
rect 258574 130596 258580 130660
rect 258644 130658 258650 130660
rect 268150 130658 268210 131036
rect 398833 130930 398899 130933
rect 398833 130928 400108 130930
rect 398833 130872 398838 130928
rect 398894 130872 400108 130928
rect 398833 130870 400108 130872
rect 398833 130867 398899 130870
rect 282269 130658 282335 130661
rect 441981 130658 442047 130661
rect 258644 130598 268210 130658
rect 279956 130656 282335 130658
rect 279956 130600 282274 130656
rect 282330 130600 282335 130656
rect 279956 130598 282335 130600
rect 439852 130656 442047 130658
rect 439852 130600 441986 130656
rect 442042 130600 442047 130656
rect 439852 130598 442047 130600
rect 258644 130596 258650 130598
rect 282269 130595 282335 130598
rect 441981 130595 442047 130598
rect 231761 130250 231827 130253
rect 228988 130248 231827 130250
rect 228988 130192 231766 130248
rect 231822 130192 231827 130248
rect 228988 130190 231827 130192
rect 231761 130187 231827 130190
rect 242750 130188 242756 130252
rect 242820 130250 242826 130252
rect 268150 130250 268210 130492
rect 242820 130190 268210 130250
rect 242820 130188 242826 130190
rect 264094 130052 264100 130116
rect 264164 130114 264170 130116
rect 264164 130054 268180 130114
rect 264164 130052 264170 130054
rect 214005 129978 214071 129981
rect 214005 129976 217028 129978
rect 214005 129920 214010 129976
rect 214066 129920 217028 129976
rect 214005 129918 217028 129920
rect 214005 129915 214071 129918
rect 231025 129842 231091 129845
rect 282637 129842 282703 129845
rect 228988 129840 231091 129842
rect 228988 129784 231030 129840
rect 231086 129784 231091 129840
rect 228988 129782 231091 129784
rect 279956 129840 282703 129842
rect 279956 129784 282642 129840
rect 282698 129784 282703 129840
rect 279956 129782 282703 129784
rect 231025 129779 231091 129782
rect 282637 129779 282703 129782
rect 264973 129706 265039 129709
rect 398649 129706 398715 129709
rect 442901 129706 442967 129709
rect 264973 129704 268180 129706
rect 264973 129648 264978 129704
rect 265034 129648 268180 129704
rect 264973 129646 268180 129648
rect 398649 129704 400108 129706
rect 398649 129648 398654 129704
rect 398710 129648 400108 129704
rect 398649 129646 400108 129648
rect 439852 129704 442967 129706
rect 439852 129648 442906 129704
rect 442962 129648 442967 129704
rect 439852 129646 442967 129648
rect 264973 129643 265039 129646
rect 398649 129643 398715 129646
rect 442901 129643 442967 129646
rect 66069 129298 66135 129301
rect 68142 129298 68816 129304
rect 66069 129296 68816 129298
rect 66069 129240 66074 129296
rect 66130 129244 68816 129296
rect 214005 129298 214071 129301
rect 231301 129298 231367 129301
rect 214005 129296 217028 129298
rect 66130 129240 68202 129244
rect 66069 129238 68202 129240
rect 214005 129240 214010 129296
rect 214066 129240 217028 129296
rect 214005 129238 217028 129240
rect 228988 129296 231367 129298
rect 228988 129240 231306 129296
rect 231362 129240 231367 129296
rect 228988 129238 231367 129240
rect 66069 129235 66135 129238
rect 214005 129235 214071 129238
rect 231301 129235 231367 129238
rect 232446 128964 232452 129028
rect 232516 129026 232522 129028
rect 268150 129026 268210 129268
rect 281625 129026 281691 129029
rect 232516 128966 268210 129026
rect 279956 129024 281691 129026
rect 279956 128968 281630 129024
rect 281686 128968 281691 129024
rect 279956 128966 281691 128968
rect 232516 128964 232522 128966
rect 281625 128963 281691 128966
rect 397545 129026 397611 129029
rect 397545 129024 400108 129026
rect 397545 128968 397550 129024
rect 397606 128968 400108 129024
rect 397545 128966 400108 128968
rect 397545 128963 397611 128966
rect 230749 128890 230815 128893
rect 228988 128888 230815 128890
rect 228988 128832 230754 128888
rect 230810 128832 230815 128888
rect 228988 128830 230815 128832
rect 230749 128827 230815 128830
rect 258030 128830 268180 128890
rect 213913 128754 213979 128757
rect 240869 128754 240935 128757
rect 258030 128754 258090 128830
rect 440417 128754 440483 128757
rect 213913 128752 217028 128754
rect 213913 128696 213918 128752
rect 213974 128696 217028 128752
rect 213913 128694 217028 128696
rect 240869 128752 258090 128754
rect 240869 128696 240874 128752
rect 240930 128696 258090 128752
rect 240869 128694 258090 128696
rect 439852 128752 440483 128754
rect 439852 128696 440422 128752
rect 440478 128696 440483 128752
rect 439852 128694 440483 128696
rect 213913 128691 213979 128694
rect 240869 128691 240935 128694
rect 440417 128691 440483 128694
rect 265617 128482 265683 128485
rect 265617 128480 268180 128482
rect 265617 128424 265622 128480
rect 265678 128424 268180 128480
rect 265617 128422 268180 128424
rect 265617 128419 265683 128422
rect 231669 128346 231735 128349
rect 282821 128346 282887 128349
rect 228988 128344 231735 128346
rect 228988 128288 231674 128344
rect 231730 128288 231735 128344
rect 228988 128286 231735 128288
rect 279956 128344 282887 128346
rect 279956 128288 282826 128344
rect 282882 128288 282887 128344
rect 279956 128286 282887 128288
rect 231669 128283 231735 128286
rect 282821 128283 282887 128286
rect 397545 128210 397611 128213
rect 397545 128208 400108 128210
rect 397545 128152 397550 128208
rect 397606 128152 400108 128208
rect 397545 128150 400108 128152
rect 397545 128147 397611 128150
rect 65517 128074 65583 128077
rect 68142 128074 68816 128080
rect 65517 128072 68816 128074
rect 65517 128016 65522 128072
rect 65578 128020 68816 128072
rect 213913 128074 213979 128077
rect 231669 128074 231735 128077
rect 238017 128074 238083 128077
rect 213913 128072 217028 128074
rect 65578 128016 68202 128020
rect 65517 128014 68202 128016
rect 213913 128016 213918 128072
rect 213974 128016 217028 128072
rect 213913 128014 217028 128016
rect 231669 128072 238083 128074
rect 231669 128016 231674 128072
rect 231730 128016 238022 128072
rect 238078 128016 238083 128072
rect 231669 128014 238083 128016
rect 65517 128011 65583 128014
rect 213913 128011 213979 128014
rect 231669 128011 231735 128014
rect 238017 128011 238083 128014
rect 230657 127938 230723 127941
rect 228988 127936 230723 127938
rect 228988 127880 230662 127936
rect 230718 127880 230723 127936
rect 228988 127878 230723 127880
rect 230657 127875 230723 127878
rect 264973 127938 265039 127941
rect 264973 127936 268180 127938
rect 264973 127880 264978 127936
rect 265034 127880 268180 127936
rect 264973 127878 268180 127880
rect 264973 127875 265039 127878
rect 442901 127802 442967 127805
rect 439852 127800 442967 127802
rect 439852 127744 442906 127800
rect 442962 127744 442967 127800
rect 439852 127742 442967 127744
rect 442901 127739 442967 127742
rect 282821 127530 282887 127533
rect 258030 127470 268180 127530
rect 279956 127528 282887 127530
rect 279956 127472 282826 127528
rect 282882 127472 282887 127528
rect 279956 127470 282887 127472
rect 231761 127394 231827 127397
rect 228988 127392 231827 127394
rect 199469 127258 199535 127261
rect 216998 127258 217058 127364
rect 228988 127336 231766 127392
rect 231822 127336 231827 127392
rect 228988 127334 231827 127336
rect 231761 127331 231827 127334
rect 244038 127332 244044 127396
rect 244108 127394 244114 127396
rect 258030 127394 258090 127470
rect 282821 127467 282887 127470
rect 244108 127334 258090 127394
rect 244108 127332 244114 127334
rect 199469 127256 217058 127258
rect 199469 127200 199474 127256
rect 199530 127200 217058 127256
rect 199469 127198 217058 127200
rect 199469 127195 199535 127198
rect 265065 127122 265131 127125
rect 397545 127122 397611 127125
rect 265065 127120 268180 127122
rect 265065 127064 265070 127120
rect 265126 127064 268180 127120
rect 265065 127062 268180 127064
rect 397545 127120 400108 127122
rect 397545 127064 397550 127120
rect 397606 127064 400108 127120
rect 397545 127062 400108 127064
rect 265065 127059 265131 127062
rect 397545 127059 397611 127062
rect 262857 126986 262923 126989
rect 228988 126984 262923 126986
rect 228988 126928 262862 126984
rect 262918 126928 262923 126984
rect 228988 126926 262923 126928
rect 262857 126923 262923 126926
rect 231209 126850 231275 126853
rect 235441 126850 235507 126853
rect 281533 126850 281599 126853
rect 231209 126848 235507 126850
rect 231209 126792 231214 126848
rect 231270 126792 235446 126848
rect 235502 126792 235507 126848
rect 231209 126790 235507 126792
rect 279956 126848 281599 126850
rect 279956 126792 281538 126848
rect 281594 126792 281599 126848
rect 279956 126790 281599 126792
rect 231209 126787 231275 126790
rect 235441 126787 235507 126790
rect 281533 126787 281599 126790
rect 213913 126714 213979 126717
rect 442901 126714 442967 126717
rect 213913 126712 217028 126714
rect 213913 126656 213918 126712
rect 213974 126656 217028 126712
rect 439852 126712 442967 126714
rect 213913 126654 217028 126656
rect 213913 126651 213979 126654
rect 231301 126442 231367 126445
rect 228988 126440 231367 126442
rect 228988 126384 231306 126440
rect 231362 126384 231367 126440
rect 228988 126382 231367 126384
rect 231301 126379 231367 126382
rect 260046 126380 260052 126444
rect 260116 126442 260122 126444
rect 268150 126442 268210 126684
rect 439852 126656 442906 126712
rect 442962 126656 442967 126712
rect 439852 126654 442967 126656
rect 442901 126651 442967 126654
rect 260116 126382 268210 126442
rect 260116 126380 260122 126382
rect 64965 126306 65031 126309
rect 68142 126306 68816 126312
rect 64965 126304 68816 126306
rect 64965 126248 64970 126304
rect 65026 126252 68816 126304
rect 264973 126306 265039 126309
rect 397545 126306 397611 126309
rect 264973 126304 268180 126306
rect 65026 126248 68202 126252
rect 64965 126246 68202 126248
rect 264973 126248 264978 126304
rect 265034 126248 268180 126304
rect 264973 126246 268180 126248
rect 397545 126304 400108 126306
rect 397545 126248 397550 126304
rect 397606 126248 400108 126304
rect 397545 126246 400108 126248
rect 64965 126243 65031 126246
rect 264973 126243 265039 126246
rect 397545 126243 397611 126246
rect 216029 126034 216095 126037
rect 230565 126034 230631 126037
rect 282821 126034 282887 126037
rect 216029 126032 217028 126034
rect 216029 125976 216034 126032
rect 216090 125976 217028 126032
rect 216029 125974 217028 125976
rect 228988 126032 230631 126034
rect 228988 125976 230570 126032
rect 230626 125976 230631 126032
rect 228988 125974 230631 125976
rect 279956 126032 282887 126034
rect 279956 125976 282826 126032
rect 282882 125976 282887 126032
rect 279956 125974 282887 125976
rect 216029 125971 216095 125974
rect 230565 125971 230631 125974
rect 282821 125971 282887 125974
rect 580165 126034 580231 126037
rect 583520 126034 584960 126124
rect 580165 126032 584960 126034
rect 580165 125976 580170 126032
rect 580226 125976 584960 126032
rect 580165 125974 584960 125976
rect 580165 125971 580231 125974
rect 265709 125898 265775 125901
rect 440417 125898 440483 125901
rect 265709 125896 268180 125898
rect 265709 125840 265714 125896
rect 265770 125840 268180 125896
rect 265709 125838 268180 125840
rect 439852 125896 440483 125898
rect 439852 125840 440422 125896
rect 440478 125840 440483 125896
rect 583520 125884 584960 125974
rect 439852 125838 440483 125840
rect 265709 125835 265775 125838
rect 440417 125835 440483 125838
rect 64781 125626 64847 125629
rect 64965 125626 65031 125629
rect 64781 125624 65031 125626
rect 64781 125568 64786 125624
rect 64842 125568 64970 125624
rect 65026 125568 65031 125624
rect 64781 125566 65031 125568
rect 64781 125563 64847 125566
rect 64965 125563 65031 125566
rect 237005 125490 237071 125493
rect 228988 125488 237071 125490
rect 228988 125432 237010 125488
rect 237066 125432 237071 125488
rect 228988 125430 237071 125432
rect 237005 125427 237071 125430
rect 214005 125354 214071 125357
rect 265065 125354 265131 125357
rect 214005 125352 217028 125354
rect 214005 125296 214010 125352
rect 214066 125296 217028 125352
rect 214005 125294 217028 125296
rect 265065 125352 268180 125354
rect 265065 125296 265070 125352
rect 265126 125296 268180 125352
rect 265065 125294 268180 125296
rect 214005 125291 214071 125294
rect 265065 125291 265131 125294
rect 66161 125218 66227 125221
rect 68142 125218 68816 125224
rect 282177 125218 282243 125221
rect 66161 125216 68816 125218
rect 66161 125160 66166 125216
rect 66222 125164 68816 125216
rect 279956 125216 282243 125218
rect 66222 125160 68202 125164
rect 66161 125158 68202 125160
rect 279956 125160 282182 125216
rect 282238 125160 282243 125216
rect 279956 125158 282243 125160
rect 66161 125155 66227 125158
rect 282177 125155 282243 125158
rect 397545 125218 397611 125221
rect 397545 125216 400108 125218
rect 397545 125160 397550 125216
rect 397606 125160 400108 125216
rect 397545 125158 400108 125160
rect 397545 125155 397611 125158
rect 231485 125082 231551 125085
rect 442206 125082 442212 125084
rect 228988 125080 231551 125082
rect 228988 125024 231490 125080
rect 231546 125024 231551 125080
rect 228988 125022 231551 125024
rect 439852 125022 442212 125082
rect 231485 125019 231551 125022
rect 442206 125020 442212 125022
rect 442276 125020 442282 125084
rect 199377 124810 199443 124813
rect 209221 124810 209287 124813
rect 199377 124808 209287 124810
rect 199377 124752 199382 124808
rect 199438 124752 209226 124808
rect 209282 124752 209287 124808
rect 199377 124750 209287 124752
rect 199377 124747 199443 124750
rect 209221 124747 209287 124750
rect 231301 124810 231367 124813
rect 243905 124810 243971 124813
rect 231301 124808 243971 124810
rect 231301 124752 231306 124808
rect 231362 124752 243910 124808
rect 243966 124752 243971 124808
rect 231301 124750 243971 124752
rect 231301 124747 231367 124750
rect 243905 124747 243971 124750
rect 213913 124674 213979 124677
rect 213913 124672 217028 124674
rect 213913 124616 213918 124672
rect 213974 124616 217028 124672
rect 213913 124614 217028 124616
rect 213913 124611 213979 124614
rect 244774 124612 244780 124676
rect 244844 124674 244850 124676
rect 268150 124674 268210 124916
rect 244844 124614 268210 124674
rect 244844 124612 244850 124614
rect 230749 124538 230815 124541
rect 228988 124536 230815 124538
rect 228988 124480 230754 124536
rect 230810 124480 230815 124536
rect 228988 124478 230815 124480
rect 230749 124475 230815 124478
rect 264973 124538 265039 124541
rect 281625 124538 281691 124541
rect 264973 124536 268180 124538
rect 264973 124480 264978 124536
rect 265034 124480 268180 124536
rect 264973 124478 268180 124480
rect 279956 124536 281691 124538
rect 279956 124480 281630 124536
rect 281686 124480 281691 124536
rect 279956 124478 281691 124480
rect 264973 124475 265039 124478
rect 281625 124475 281691 124478
rect 397637 124402 397703 124405
rect 397637 124400 400108 124402
rect 397637 124344 397642 124400
rect 397698 124344 400108 124400
rect 397637 124342 400108 124344
rect 397637 124339 397703 124342
rect 213913 124130 213979 124133
rect 231669 124130 231735 124133
rect 213913 124128 217028 124130
rect 213913 124072 213918 124128
rect 213974 124072 217028 124128
rect 213913 124070 217028 124072
rect 228988 124128 231735 124130
rect 228988 124072 231674 124128
rect 231730 124072 231735 124128
rect 228988 124070 231735 124072
rect 213913 124067 213979 124070
rect 231669 124067 231735 124070
rect 264973 124130 265039 124133
rect 442901 124130 442967 124133
rect 264973 124128 268180 124130
rect 264973 124072 264978 124128
rect 265034 124072 268180 124128
rect 264973 124070 268180 124072
rect 439852 124128 442967 124130
rect 439852 124072 442906 124128
rect 442962 124072 442967 124128
rect 439852 124070 442967 124072
rect 264973 124067 265039 124070
rect 442901 124067 442967 124070
rect -960 123572 480 123812
rect 265065 123722 265131 123725
rect 282085 123722 282151 123725
rect 265065 123720 268180 123722
rect 265065 123664 265070 123720
rect 265126 123664 268180 123720
rect 265065 123662 268180 123664
rect 279956 123720 282151 123722
rect 279956 123664 282090 123720
rect 282146 123664 282151 123720
rect 279956 123662 282151 123664
rect 265065 123659 265131 123662
rect 282085 123659 282151 123662
rect 67633 123586 67699 123589
rect 68142 123586 68816 123592
rect 230013 123586 230079 123589
rect 67633 123584 68816 123586
rect 67633 123528 67638 123584
rect 67694 123532 68816 123584
rect 228988 123584 230079 123586
rect 67694 123528 68202 123532
rect 67633 123526 68202 123528
rect 228988 123528 230018 123584
rect 230074 123528 230079 123584
rect 228988 123526 230079 123528
rect 67633 123523 67699 123526
rect 230013 123523 230079 123526
rect 184289 123450 184355 123453
rect 213453 123450 213519 123453
rect 234153 123450 234219 123453
rect 265893 123450 265959 123453
rect 184289 123448 200130 123450
rect 184289 123392 184294 123448
rect 184350 123392 200130 123448
rect 184289 123390 200130 123392
rect 184289 123387 184355 123390
rect 200070 123314 200130 123390
rect 213453 123448 217028 123450
rect 213453 123392 213458 123448
rect 213514 123392 217028 123448
rect 213453 123390 217028 123392
rect 234153 123448 265959 123450
rect 234153 123392 234158 123448
rect 234214 123392 265898 123448
rect 265954 123392 265959 123448
rect 234153 123390 265959 123392
rect 213453 123387 213519 123390
rect 234153 123387 234219 123390
rect 265893 123387 265959 123390
rect 214414 123314 214420 123316
rect 200070 123254 214420 123314
rect 214414 123252 214420 123254
rect 214484 123252 214490 123316
rect 229737 123314 229803 123317
rect 397545 123314 397611 123317
rect 442809 123314 442875 123317
rect 229737 123312 268180 123314
rect 229737 123256 229742 123312
rect 229798 123256 268180 123312
rect 229737 123254 268180 123256
rect 397545 123312 400108 123314
rect 397545 123256 397550 123312
rect 397606 123256 400108 123312
rect 397545 123254 400108 123256
rect 439852 123312 442875 123314
rect 439852 123256 442814 123312
rect 442870 123256 442875 123312
rect 439852 123254 442875 123256
rect 229737 123251 229803 123254
rect 397545 123251 397611 123254
rect 442809 123251 442875 123254
rect 230974 123178 230980 123180
rect 228988 123118 230980 123178
rect 230974 123116 230980 123118
rect 231044 123116 231050 123180
rect 282637 123042 282703 123045
rect 279956 123040 282703 123042
rect 279956 122984 282642 123040
rect 282698 122984 282703 123040
rect 279956 122982 282703 122984
rect 282637 122979 282703 122982
rect 267089 122906 267155 122909
rect 267089 122904 268180 122906
rect 267089 122848 267094 122904
rect 267150 122848 268180 122904
rect 267089 122846 268180 122848
rect 267089 122843 267155 122846
rect 214005 122770 214071 122773
rect 214005 122768 217028 122770
rect 214005 122712 214010 122768
rect 214066 122712 217028 122768
rect 214005 122710 217028 122712
rect 214005 122707 214071 122710
rect 65977 122634 66043 122637
rect 68142 122634 68816 122640
rect 231761 122634 231827 122637
rect 65977 122632 68816 122634
rect 65977 122576 65982 122632
rect 66038 122580 68816 122632
rect 228988 122632 231827 122634
rect 66038 122576 68202 122580
rect 65977 122574 68202 122576
rect 228988 122576 231766 122632
rect 231822 122576 231827 122632
rect 228988 122574 231827 122576
rect 65977 122571 66043 122574
rect 231761 122571 231827 122574
rect 397545 122362 397611 122365
rect 397545 122360 400108 122362
rect 231025 122226 231091 122229
rect 228988 122224 231091 122226
rect 228988 122168 231030 122224
rect 231086 122168 231091 122224
rect 228988 122166 231091 122168
rect 231025 122163 231091 122166
rect 213913 122090 213979 122093
rect 234061 122090 234127 122093
rect 268150 122090 268210 122332
rect 397545 122304 397550 122360
rect 397606 122304 400108 122360
rect 397545 122302 400108 122304
rect 397545 122299 397611 122302
rect 282821 122226 282887 122229
rect 279956 122224 282887 122226
rect 279956 122168 282826 122224
rect 282882 122168 282887 122224
rect 279956 122166 282887 122168
rect 282821 122163 282887 122166
rect 442993 122090 443059 122093
rect 213913 122088 217028 122090
rect 213913 122032 213918 122088
rect 213974 122032 217028 122088
rect 213913 122030 217028 122032
rect 234061 122088 268210 122090
rect 234061 122032 234066 122088
rect 234122 122032 268210 122088
rect 234061 122030 268210 122032
rect 439852 122088 443059 122090
rect 439852 122032 442998 122088
rect 443054 122032 443059 122088
rect 439852 122030 443059 122032
rect 213913 122027 213979 122030
rect 234061 122027 234127 122030
rect 442993 122027 443059 122030
rect 264973 121954 265039 121957
rect 264973 121952 268180 121954
rect 264973 121896 264978 121952
rect 265034 121896 268180 121952
rect 264973 121894 268180 121896
rect 264973 121891 265039 121894
rect 231209 121682 231275 121685
rect 228988 121680 231275 121682
rect 228988 121624 231214 121680
rect 231270 121624 231275 121680
rect 228988 121622 231275 121624
rect 231209 121619 231275 121622
rect 246297 121682 246363 121685
rect 246297 121680 268210 121682
rect 246297 121624 246302 121680
rect 246358 121624 268210 121680
rect 246297 121622 268210 121624
rect 246297 121619 246363 121622
rect 268150 121516 268210 121622
rect 214005 121410 214071 121413
rect 258901 121410 258967 121413
rect 280153 121410 280219 121413
rect 214005 121408 217028 121410
rect 214005 121352 214010 121408
rect 214066 121352 217028 121408
rect 214005 121350 217028 121352
rect 238710 121408 258967 121410
rect 238710 121352 258906 121408
rect 258962 121352 258967 121408
rect 238710 121350 258967 121352
rect 279956 121408 280219 121410
rect 279956 121352 280158 121408
rect 280214 121352 280219 121408
rect 279956 121350 280219 121352
rect 214005 121347 214071 121350
rect 238710 121274 238770 121350
rect 258901 121347 258967 121350
rect 280153 121347 280219 121350
rect 398189 121410 398255 121413
rect 442901 121410 442967 121413
rect 398189 121408 400108 121410
rect 398189 121352 398194 121408
rect 398250 121352 400108 121408
rect 398189 121350 400108 121352
rect 439852 121408 442967 121410
rect 439852 121352 442906 121408
rect 442962 121352 442967 121408
rect 439852 121350 442967 121352
rect 398189 121347 398255 121350
rect 442901 121347 442967 121350
rect 228988 121214 238770 121274
rect 265065 121138 265131 121141
rect 265065 121136 268180 121138
rect 265065 121080 265070 121136
rect 265126 121080 268180 121136
rect 265065 121078 268180 121080
rect 265065 121075 265131 121078
rect 67449 120866 67515 120869
rect 68142 120866 68816 120872
rect 263133 120866 263199 120869
rect 67449 120864 68816 120866
rect 67449 120808 67454 120864
rect 67510 120812 68816 120864
rect 258030 120864 263199 120866
rect 67510 120808 68202 120812
rect 67449 120806 68202 120808
rect 258030 120808 263138 120864
rect 263194 120808 263199 120864
rect 258030 120806 263199 120808
rect 67449 120803 67515 120806
rect 213913 120730 213979 120733
rect 231761 120730 231827 120733
rect 258030 120730 258090 120806
rect 263133 120803 263199 120806
rect 213913 120728 217028 120730
rect 213913 120672 213918 120728
rect 213974 120672 217028 120728
rect 213913 120670 217028 120672
rect 228988 120728 231827 120730
rect 228988 120672 231766 120728
rect 231822 120672 231827 120728
rect 228988 120670 231827 120672
rect 213913 120667 213979 120670
rect 231761 120667 231827 120670
rect 238710 120670 258090 120730
rect 262857 120730 262923 120733
rect 262857 120728 268180 120730
rect 262857 120672 262862 120728
rect 262918 120672 268180 120728
rect 262857 120670 268180 120672
rect 231209 120594 231275 120597
rect 238710 120594 238770 120670
rect 262857 120667 262923 120670
rect 231209 120592 238770 120594
rect 231209 120536 231214 120592
rect 231270 120536 238770 120592
rect 231209 120534 238770 120536
rect 231209 120531 231275 120534
rect 231485 120322 231551 120325
rect 228988 120320 231551 120322
rect 228988 120264 231490 120320
rect 231546 120264 231551 120320
rect 228988 120262 231551 120264
rect 231485 120259 231551 120262
rect 262949 120322 263015 120325
rect 262949 120320 268180 120322
rect 262949 120264 262954 120320
rect 263010 120264 268180 120320
rect 262949 120262 268180 120264
rect 262949 120259 263015 120262
rect 279374 120189 279434 120700
rect 398741 120594 398807 120597
rect 398741 120592 400108 120594
rect 398741 120536 398746 120592
rect 398802 120536 400108 120592
rect 398741 120534 400108 120536
rect 398741 120531 398807 120534
rect 439262 120532 439268 120596
rect 439332 120594 439338 120596
rect 439630 120594 439636 120596
rect 439332 120534 439636 120594
rect 439332 120532 439338 120534
rect 439630 120532 439636 120534
rect 439700 120532 439706 120596
rect 442625 120322 442691 120325
rect 439852 120320 442691 120322
rect 439852 120264 442630 120320
rect 442686 120264 442691 120320
rect 439852 120262 442691 120264
rect 442625 120259 442691 120262
rect 279325 120184 279434 120189
rect 279325 120128 279330 120184
rect 279386 120128 279434 120184
rect 279325 120126 279434 120128
rect 279325 120123 279391 120126
rect 214005 120050 214071 120053
rect 231669 120050 231735 120053
rect 240726 120050 240732 120052
rect 214005 120048 217028 120050
rect 214005 119992 214010 120048
rect 214066 119992 217028 120048
rect 214005 119990 217028 119992
rect 231669 120048 240732 120050
rect 231669 119992 231674 120048
rect 231730 119992 240732 120048
rect 231669 119990 240732 119992
rect 214005 119987 214071 119990
rect 231669 119987 231735 119990
rect 240726 119988 240732 119990
rect 240796 119988 240802 120052
rect 282821 119914 282887 119917
rect 279956 119912 282887 119914
rect 279956 119856 282826 119912
rect 282882 119856 282887 119912
rect 279956 119854 282887 119856
rect 282821 119851 282887 119854
rect 231761 119778 231827 119781
rect 228988 119776 231827 119778
rect 228988 119720 231766 119776
rect 231822 119720 231827 119776
rect 228988 119718 231827 119720
rect 231761 119715 231827 119718
rect 264973 119778 265039 119781
rect 397545 119778 397611 119781
rect 264973 119776 268180 119778
rect 264973 119720 264978 119776
rect 265034 119720 268180 119776
rect 264973 119718 268180 119720
rect 397545 119776 400108 119778
rect 397545 119720 397550 119776
rect 397606 119720 400108 119776
rect 397545 119718 400108 119720
rect 264973 119715 265039 119718
rect 397545 119715 397611 119718
rect 213913 119506 213979 119509
rect 442901 119506 442967 119509
rect 213913 119504 217028 119506
rect 213913 119448 213918 119504
rect 213974 119448 217028 119504
rect 213913 119446 217028 119448
rect 439852 119504 442967 119506
rect 439852 119448 442906 119504
rect 442962 119448 442967 119504
rect 439852 119446 442967 119448
rect 213913 119443 213979 119446
rect 442901 119443 442967 119446
rect 174537 119370 174603 119373
rect 211981 119370 212047 119373
rect 231669 119370 231735 119373
rect 174537 119368 212047 119370
rect 174537 119312 174542 119368
rect 174598 119312 211986 119368
rect 212042 119312 212047 119368
rect 174537 119310 212047 119312
rect 228988 119368 231735 119370
rect 228988 119312 231674 119368
rect 231730 119312 231735 119368
rect 228988 119310 231735 119312
rect 174537 119307 174603 119310
rect 211981 119307 212047 119310
rect 231669 119307 231735 119310
rect 261477 119370 261543 119373
rect 261477 119368 268180 119370
rect 261477 119312 261482 119368
rect 261538 119312 268180 119368
rect 261477 119310 268180 119312
rect 261477 119307 261543 119310
rect 280429 119234 280495 119237
rect 279956 119232 280495 119234
rect 279956 119176 280434 119232
rect 280490 119176 280495 119232
rect 279956 119174 280495 119176
rect 280429 119171 280495 119174
rect 230657 118962 230723 118965
rect 228988 118960 230723 118962
rect 228988 118904 230662 118960
rect 230718 118904 230723 118960
rect 228988 118902 230723 118904
rect 230657 118899 230723 118902
rect 258030 118902 268180 118962
rect 213269 118826 213335 118829
rect 239489 118826 239555 118829
rect 258030 118826 258090 118902
rect 213269 118824 217028 118826
rect 213269 118768 213274 118824
rect 213330 118768 217028 118824
rect 213269 118766 217028 118768
rect 239489 118824 258090 118826
rect 239489 118768 239494 118824
rect 239550 118768 258090 118824
rect 239489 118766 258090 118768
rect 213269 118763 213335 118766
rect 239489 118763 239555 118766
rect 249057 118690 249123 118693
rect 441705 118690 441771 118693
rect 238710 118688 249123 118690
rect 238710 118632 249062 118688
rect 249118 118632 249123 118688
rect 238710 118630 249123 118632
rect 439852 118688 441771 118690
rect 439852 118632 441710 118688
rect 441766 118632 441771 118688
rect 439852 118630 441771 118632
rect 238710 118418 238770 118630
rect 249057 118627 249123 118630
rect 441705 118627 441771 118630
rect 264973 118554 265039 118557
rect 397545 118554 397611 118557
rect 264973 118552 268180 118554
rect 264973 118496 264978 118552
rect 265034 118496 268180 118552
rect 264973 118494 268180 118496
rect 397545 118552 400108 118554
rect 397545 118496 397550 118552
rect 397606 118496 400108 118552
rect 397545 118494 400108 118496
rect 264973 118491 265039 118494
rect 397545 118491 397611 118494
rect 282821 118418 282887 118421
rect 228988 118358 238770 118418
rect 279956 118416 282887 118418
rect 279956 118360 282826 118416
rect 282882 118360 282887 118416
rect 279956 118358 282887 118360
rect 282821 118355 282887 118358
rect 214005 118146 214071 118149
rect 214005 118144 217028 118146
rect 214005 118088 214010 118144
rect 214066 118088 217028 118144
rect 214005 118086 217028 118088
rect 214005 118083 214071 118086
rect 193857 118010 193923 118013
rect 209313 118010 209379 118013
rect 238201 118010 238267 118013
rect 193857 118008 209379 118010
rect 193857 117952 193862 118008
rect 193918 117952 209318 118008
rect 209374 117952 209379 118008
rect 193857 117950 209379 117952
rect 228988 118008 238267 118010
rect 228988 117952 238206 118008
rect 238262 117952 238267 118008
rect 228988 117950 238267 117952
rect 193857 117947 193923 117950
rect 209313 117947 209379 117950
rect 238201 117947 238267 117950
rect 260097 117874 260163 117877
rect 268150 117874 268210 118116
rect 260097 117872 268210 117874
rect 260097 117816 260102 117872
rect 260158 117816 268210 117872
rect 260097 117814 268210 117816
rect 397637 117874 397703 117877
rect 397637 117872 400108 117874
rect 397637 117816 397642 117872
rect 397698 117816 400108 117872
rect 397637 117814 400108 117816
rect 260097 117811 260163 117814
rect 397637 117811 397703 117814
rect 258030 117678 268180 117738
rect 242157 117602 242223 117605
rect 258030 117602 258090 117678
rect 282821 117602 282887 117605
rect 440509 117602 440575 117605
rect 242157 117600 258090 117602
rect 242157 117544 242162 117600
rect 242218 117544 258090 117600
rect 242157 117542 258090 117544
rect 279956 117600 282887 117602
rect 279956 117544 282826 117600
rect 282882 117544 282887 117600
rect 279956 117542 282887 117544
rect 439852 117600 440575 117602
rect 439852 117544 440514 117600
rect 440570 117544 440575 117600
rect 439852 117542 440575 117544
rect 242157 117539 242223 117542
rect 282821 117539 282887 117542
rect 440509 117539 440575 117542
rect 213913 117466 213979 117469
rect 230565 117466 230631 117469
rect 213913 117464 217028 117466
rect 213913 117408 213918 117464
rect 213974 117408 217028 117464
rect 213913 117406 217028 117408
rect 228988 117464 230631 117466
rect 228988 117408 230570 117464
rect 230626 117408 230631 117464
rect 228988 117406 230631 117408
rect 213913 117403 213979 117406
rect 230565 117403 230631 117406
rect 265065 117194 265131 117197
rect 291101 117194 291167 117197
rect 361614 117194 361620 117196
rect 265065 117192 268180 117194
rect 265065 117136 265070 117192
rect 265126 117136 268180 117192
rect 265065 117134 268180 117136
rect 291101 117192 361620 117194
rect 291101 117136 291106 117192
rect 291162 117136 361620 117192
rect 291101 117134 361620 117136
rect 265065 117131 265131 117134
rect 291101 117131 291167 117134
rect 361614 117132 361620 117134
rect 361684 117132 361690 117196
rect 230841 117058 230907 117061
rect 228988 117056 230907 117058
rect 228988 117000 230846 117056
rect 230902 117000 230907 117056
rect 228988 116998 230907 117000
rect 230841 116995 230907 116998
rect 282821 116922 282887 116925
rect 279956 116920 282887 116922
rect 279956 116864 282826 116920
rect 282882 116864 282887 116920
rect 279956 116862 282887 116864
rect 282821 116859 282887 116862
rect 214005 116786 214071 116789
rect 397545 116786 397611 116789
rect 214005 116784 217028 116786
rect 214005 116728 214010 116784
rect 214066 116728 217028 116784
rect 214005 116726 217028 116728
rect 258030 116726 268180 116786
rect 397545 116784 400108 116786
rect 397545 116728 397550 116784
rect 397606 116728 400108 116784
rect 397545 116726 400108 116728
rect 214005 116723 214071 116726
rect 232773 116650 232839 116653
rect 258030 116650 258090 116726
rect 397545 116723 397611 116726
rect 441705 116650 441771 116653
rect 232773 116648 258090 116650
rect 232773 116592 232778 116648
rect 232834 116592 258090 116648
rect 232773 116590 258090 116592
rect 439852 116648 441771 116650
rect 439852 116592 441710 116648
rect 441766 116592 441771 116648
rect 439852 116590 441771 116592
rect 232773 116587 232839 116590
rect 441705 116587 441771 116590
rect 231761 116514 231827 116517
rect 256233 116514 256299 116517
rect 228988 116512 231827 116514
rect 228988 116456 231766 116512
rect 231822 116456 231827 116512
rect 228988 116454 231827 116456
rect 231761 116451 231827 116454
rect 238710 116512 256299 116514
rect 238710 116456 256238 116512
rect 256294 116456 256299 116512
rect 238710 116454 256299 116456
rect 231393 116378 231459 116381
rect 238710 116378 238770 116454
rect 256233 116451 256299 116454
rect 231393 116376 238770 116378
rect 231393 116320 231398 116376
rect 231454 116320 238770 116376
rect 231393 116318 238770 116320
rect 264973 116378 265039 116381
rect 264973 116376 268180 116378
rect 264973 116320 264978 116376
rect 265034 116320 268180 116376
rect 264973 116318 268180 116320
rect 231393 116315 231459 116318
rect 264973 116315 265039 116318
rect 213913 116106 213979 116109
rect 231669 116106 231735 116109
rect 282269 116106 282335 116109
rect 213913 116104 217028 116106
rect 213913 116048 213918 116104
rect 213974 116048 217028 116104
rect 213913 116046 217028 116048
rect 228988 116104 231735 116106
rect 228988 116048 231674 116104
rect 231730 116048 231735 116104
rect 228988 116046 231735 116048
rect 279956 116104 282335 116106
rect 279956 116048 282274 116104
rect 282330 116048 282335 116104
rect 279956 116046 282335 116048
rect 213913 116043 213979 116046
rect 231669 116043 231735 116046
rect 282269 116043 282335 116046
rect 267641 115970 267707 115973
rect 267641 115968 268180 115970
rect 267641 115912 267646 115968
rect 267702 115912 268180 115968
rect 267641 115910 268180 115912
rect 267641 115907 267707 115910
rect 397361 115834 397427 115837
rect 397361 115832 400108 115834
rect 397361 115776 397366 115832
rect 397422 115776 400108 115832
rect 397361 115774 400108 115776
rect 397361 115771 397427 115774
rect 239857 115562 239923 115565
rect 228988 115560 239923 115562
rect 228988 115504 239862 115560
rect 239918 115504 239923 115560
rect 228988 115502 239923 115504
rect 239857 115499 239923 115502
rect 265065 115562 265131 115565
rect 442901 115562 442967 115565
rect 265065 115560 268180 115562
rect 265065 115504 265070 115560
rect 265126 115504 268180 115560
rect 265065 115502 268180 115504
rect 439852 115560 442967 115562
rect 439852 115504 442906 115560
rect 442962 115504 442967 115560
rect 439852 115502 442967 115504
rect 265065 115499 265131 115502
rect 442901 115499 442967 115502
rect 214005 115426 214071 115429
rect 281717 115426 281783 115429
rect 214005 115424 217028 115426
rect 214005 115368 214010 115424
rect 214066 115368 217028 115424
rect 214005 115366 217028 115368
rect 279956 115424 281783 115426
rect 279956 115368 281722 115424
rect 281778 115368 281783 115424
rect 279956 115366 281783 115368
rect 214005 115363 214071 115366
rect 281717 115363 281783 115366
rect 231485 115154 231551 115157
rect 228988 115152 231551 115154
rect 228988 115096 231490 115152
rect 231546 115096 231551 115152
rect 228988 115094 231551 115096
rect 231485 115091 231551 115094
rect 239673 115154 239739 115157
rect 259269 115154 259335 115157
rect 239673 115152 259335 115154
rect 239673 115096 239678 115152
rect 239734 115096 259274 115152
rect 259330 115096 259335 115152
rect 239673 115094 259335 115096
rect 239673 115091 239739 115094
rect 259269 115091 259335 115094
rect 264973 115154 265039 115157
rect 264973 115152 268180 115154
rect 264973 115096 264978 115152
rect 265034 115096 268180 115152
rect 264973 115094 268180 115096
rect 264973 115091 265039 115094
rect 213913 114882 213979 114885
rect 397545 114882 397611 114885
rect 213913 114880 217028 114882
rect 213913 114824 213918 114880
rect 213974 114824 217028 114880
rect 213913 114822 217028 114824
rect 397545 114880 400108 114882
rect 397545 114824 397550 114880
rect 397606 114824 400108 114880
rect 397545 114822 400108 114824
rect 213913 114819 213979 114822
rect 397545 114819 397611 114822
rect 440509 114746 440575 114749
rect 439852 114744 440575 114746
rect 439852 114688 440514 114744
rect 440570 114688 440575 114744
rect 439852 114686 440575 114688
rect 440509 114683 440575 114686
rect 231117 114610 231183 114613
rect 228988 114608 231183 114610
rect 228988 114552 231122 114608
rect 231178 114552 231183 114608
rect 228988 114550 231183 114552
rect 231117 114547 231183 114550
rect 254669 114610 254735 114613
rect 282453 114610 282519 114613
rect 254669 114608 268180 114610
rect 254669 114552 254674 114608
rect 254730 114552 268180 114608
rect 254669 114550 268180 114552
rect 279956 114608 282519 114610
rect 279956 114552 282458 114608
rect 282514 114552 282519 114608
rect 279956 114550 282519 114552
rect 254669 114547 254735 114550
rect 282453 114547 282519 114550
rect 214005 114202 214071 114205
rect 231485 114202 231551 114205
rect 214005 114200 217028 114202
rect 214005 114144 214010 114200
rect 214066 114144 217028 114200
rect 214005 114142 217028 114144
rect 228988 114200 231551 114202
rect 228988 114144 231490 114200
rect 231546 114144 231551 114200
rect 228988 114142 231551 114144
rect 214005 114139 214071 114142
rect 231485 114139 231551 114142
rect 268150 113930 268210 114172
rect 397545 114066 397611 114069
rect 397545 114064 400108 114066
rect 397545 114008 397550 114064
rect 397606 114008 400108 114064
rect 397545 114006 400108 114008
rect 397545 114003 397611 114006
rect 258030 113870 268210 113930
rect 230657 113658 230723 113661
rect 228988 113656 230723 113658
rect 228988 113600 230662 113656
rect 230718 113600 230723 113656
rect 228988 113598 230723 113600
rect 230657 113595 230723 113598
rect 213913 113522 213979 113525
rect 213913 113520 217028 113522
rect 213913 113464 213918 113520
rect 213974 113464 217028 113520
rect 213913 113462 217028 113464
rect 213913 113459 213979 113462
rect 233734 113460 233740 113524
rect 233804 113522 233810 113524
rect 258030 113522 258090 113870
rect 264973 113794 265039 113797
rect 282269 113794 282335 113797
rect 442349 113794 442415 113797
rect 264973 113792 268180 113794
rect 264973 113736 264978 113792
rect 265034 113736 268180 113792
rect 264973 113734 268180 113736
rect 279956 113792 282335 113794
rect 279956 113736 282274 113792
rect 282330 113736 282335 113792
rect 279956 113734 282335 113736
rect 439852 113792 442415 113794
rect 439852 113736 442354 113792
rect 442410 113736 442415 113792
rect 439852 113734 442415 113736
rect 264973 113731 265039 113734
rect 282269 113731 282335 113734
rect 442349 113731 442415 113734
rect 233804 113462 258090 113522
rect 233804 113460 233810 113462
rect 244917 113386 244983 113389
rect 244917 113384 268180 113386
rect 244917 113328 244922 113384
rect 244978 113328 268180 113384
rect 244917 113326 268180 113328
rect 244917 113323 244983 113326
rect 231669 113250 231735 113253
rect 228988 113248 231735 113250
rect 228988 113192 231674 113248
rect 231730 113192 231735 113248
rect 228988 113190 231735 113192
rect 231669 113187 231735 113190
rect 282821 113114 282887 113117
rect 279956 113112 282887 113114
rect 279956 113056 282826 113112
rect 282882 113056 282887 113112
rect 279956 113054 282887 113056
rect 282821 113051 282887 113054
rect 397637 113114 397703 113117
rect 397637 113112 400108 113114
rect 397637 113056 397642 113112
rect 397698 113056 400108 113112
rect 397637 113054 400108 113056
rect 397637 113051 397703 113054
rect 439262 113052 439268 113116
rect 439332 113052 439338 113116
rect 439270 112948 439330 113052
rect 214005 112842 214071 112845
rect 214005 112840 217028 112842
rect 214005 112784 214010 112840
rect 214066 112784 217028 112840
rect 214005 112782 217028 112784
rect 214005 112779 214071 112782
rect 231025 112706 231091 112709
rect 268150 112706 268210 112948
rect 583017 112842 583083 112845
rect 583520 112842 584960 112932
rect 583017 112840 584960 112842
rect 583017 112784 583022 112840
rect 583078 112784 584960 112840
rect 583017 112782 584960 112784
rect 583017 112779 583083 112782
rect 228988 112704 231091 112706
rect 228988 112648 231030 112704
rect 231086 112648 231091 112704
rect 228988 112646 231091 112648
rect 231025 112643 231091 112646
rect 258030 112646 268210 112706
rect 583520 112692 584960 112782
rect 231761 112298 231827 112301
rect 228988 112296 231827 112298
rect 228988 112240 231766 112296
rect 231822 112240 231827 112296
rect 228988 112238 231827 112240
rect 231761 112235 231827 112238
rect 213913 112162 213979 112165
rect 231117 112162 231183 112165
rect 258030 112162 258090 112646
rect 265249 112570 265315 112573
rect 265249 112568 268180 112570
rect 265249 112512 265254 112568
rect 265310 112512 268180 112568
rect 265249 112510 268180 112512
rect 265249 112507 265315 112510
rect 282821 112298 282887 112301
rect 279956 112296 282887 112298
rect 279956 112240 282826 112296
rect 282882 112240 282887 112296
rect 279956 112238 282887 112240
rect 282821 112235 282887 112238
rect 213913 112160 217028 112162
rect 213913 112104 213918 112160
rect 213974 112104 217028 112160
rect 213913 112102 217028 112104
rect 231117 112160 258090 112162
rect 231117 112104 231122 112160
rect 231178 112104 258090 112160
rect 231117 112102 258090 112104
rect 213913 112099 213979 112102
rect 231117 112099 231183 112102
rect 264973 112026 265039 112029
rect 397729 112026 397795 112029
rect 264973 112024 268180 112026
rect 264973 111968 264978 112024
rect 265034 111968 268180 112024
rect 264973 111966 268180 111968
rect 397729 112024 400108 112026
rect 397729 111968 397734 112024
rect 397790 111968 400108 112024
rect 397729 111966 400108 111968
rect 264973 111963 265039 111966
rect 397729 111963 397795 111966
rect 164724 111754 165354 111760
rect 167821 111754 167887 111757
rect 231301 111754 231367 111757
rect 442165 111754 442231 111757
rect 164724 111752 167887 111754
rect 164724 111700 167826 111752
rect 165294 111696 167826 111700
rect 167882 111696 167887 111752
rect 165294 111694 167887 111696
rect 228988 111752 231367 111754
rect 228988 111696 231306 111752
rect 231362 111696 231367 111752
rect 228988 111694 231367 111696
rect 439852 111752 442231 111754
rect 439852 111696 442170 111752
rect 442226 111696 442231 111752
rect 439852 111694 442231 111696
rect 167821 111691 167887 111694
rect 231301 111691 231367 111694
rect 442165 111691 442231 111694
rect 265065 111618 265131 111621
rect 285622 111618 285628 111620
rect 265065 111616 268180 111618
rect 265065 111560 265070 111616
rect 265126 111560 268180 111616
rect 265065 111558 268180 111560
rect 279956 111558 285628 111618
rect 265065 111555 265131 111558
rect 285622 111556 285628 111558
rect 285692 111556 285698 111620
rect 214005 111482 214071 111485
rect 214005 111480 217028 111482
rect 214005 111424 214010 111480
rect 214066 111424 217028 111480
rect 214005 111422 217028 111424
rect 214005 111419 214071 111422
rect 230565 111346 230631 111349
rect 228988 111344 230631 111346
rect 228988 111288 230570 111344
rect 230626 111288 230631 111344
rect 228988 111286 230631 111288
rect 230565 111283 230631 111286
rect 397453 111346 397519 111349
rect 397453 111344 400108 111346
rect 397453 111288 397458 111344
rect 397514 111288 400108 111344
rect 397453 111286 400108 111288
rect 397453 111283 397519 111286
rect 264973 111210 265039 111213
rect 264973 111208 268180 111210
rect 264973 111152 264978 111208
rect 265034 111152 268180 111208
rect 264973 111150 268180 111152
rect 264973 111147 265039 111150
rect 231669 111074 231735 111077
rect 250529 111074 250595 111077
rect 442349 111074 442415 111077
rect 231669 111072 250595 111074
rect 231669 111016 231674 111072
rect 231730 111016 250534 111072
rect 250590 111016 250595 111072
rect 231669 111014 250595 111016
rect 439852 111072 442415 111074
rect 439852 111016 442354 111072
rect 442410 111016 442415 111072
rect 439852 111014 442415 111016
rect 231669 111011 231735 111014
rect 250529 111011 250595 111014
rect 442349 111011 442415 111014
rect 213913 110802 213979 110805
rect 231761 110802 231827 110805
rect 213913 110800 217028 110802
rect -960 110666 480 110756
rect 213913 110744 213918 110800
rect 213974 110744 217028 110800
rect 213913 110742 217028 110744
rect 228988 110800 231827 110802
rect 228988 110744 231766 110800
rect 231822 110744 231827 110800
rect 228988 110742 231827 110744
rect 213913 110739 213979 110742
rect 231761 110739 231827 110742
rect 242249 110802 242315 110805
rect 282269 110802 282335 110805
rect 242249 110800 268180 110802
rect 242249 110744 242254 110800
rect 242310 110744 268180 110800
rect 242249 110742 268180 110744
rect 279956 110800 282335 110802
rect 279956 110744 282274 110800
rect 282330 110744 282335 110800
rect 279956 110742 282335 110744
rect 242249 110739 242315 110742
rect 282269 110739 282335 110742
rect 3141 110666 3207 110669
rect -960 110664 3207 110666
rect -960 110608 3146 110664
rect 3202 110608 3207 110664
rect -960 110606 3207 110608
rect -960 110516 480 110606
rect 3141 110603 3207 110606
rect 254761 110394 254827 110397
rect 228988 110392 254827 110394
rect 228988 110336 254766 110392
rect 254822 110336 254827 110392
rect 228988 110334 254827 110336
rect 254761 110331 254827 110334
rect 267733 110394 267799 110397
rect 267733 110392 268180 110394
rect 267733 110336 267738 110392
rect 267794 110336 268180 110392
rect 267733 110334 268180 110336
rect 267733 110331 267799 110334
rect 214005 110258 214071 110261
rect 397545 110258 397611 110261
rect 214005 110256 217028 110258
rect 214005 110200 214010 110256
rect 214066 110200 217028 110256
rect 214005 110198 217028 110200
rect 397545 110256 400108 110258
rect 397545 110200 397550 110256
rect 397606 110200 400108 110256
rect 397545 110198 400108 110200
rect 214005 110195 214071 110198
rect 397545 110195 397611 110198
rect 164724 110122 165354 110128
rect 167821 110122 167887 110125
rect 441797 110122 441863 110125
rect 164724 110120 167887 110122
rect 164724 110068 167826 110120
rect 165294 110064 167826 110068
rect 167882 110064 167887 110120
rect 165294 110062 167887 110064
rect 439852 110120 441863 110122
rect 439852 110064 441802 110120
rect 441858 110064 441863 110120
rect 439852 110062 441863 110064
rect 167821 110059 167887 110062
rect 441797 110059 441863 110062
rect 265065 109986 265131 109989
rect 265065 109984 268180 109986
rect 265065 109928 265070 109984
rect 265126 109928 268180 109984
rect 265065 109926 268180 109928
rect 265065 109923 265131 109926
rect 231669 109850 231735 109853
rect 228988 109848 231735 109850
rect 228988 109792 231674 109848
rect 231730 109792 231735 109848
rect 228988 109790 231735 109792
rect 231669 109787 231735 109790
rect 168230 109652 168236 109716
rect 168300 109714 168306 109716
rect 192661 109714 192727 109717
rect 168300 109712 192727 109714
rect 168300 109656 192666 109712
rect 192722 109656 192727 109712
rect 168300 109654 192727 109656
rect 168300 109652 168306 109654
rect 192661 109651 192727 109654
rect 213913 109578 213979 109581
rect 264973 109578 265039 109581
rect 213913 109576 217028 109578
rect 213913 109520 213918 109576
rect 213974 109520 217028 109576
rect 213913 109518 217028 109520
rect 264973 109576 268180 109578
rect 264973 109520 264978 109576
rect 265034 109520 268180 109576
rect 264973 109518 268180 109520
rect 213913 109515 213979 109518
rect 264973 109515 265039 109518
rect 231761 109442 231827 109445
rect 228988 109440 231827 109442
rect 228988 109384 231766 109440
rect 231822 109384 231827 109440
rect 228988 109382 231827 109384
rect 279926 109442 279986 109956
rect 287094 109442 287100 109444
rect 279926 109382 287100 109442
rect 231761 109379 231827 109382
rect 287094 109380 287100 109382
rect 287164 109380 287170 109444
rect 282821 109306 282887 109309
rect 279956 109304 282887 109306
rect 279956 109248 282826 109304
rect 282882 109248 282887 109304
rect 279956 109246 282887 109248
rect 282821 109243 282887 109246
rect 397453 109306 397519 109309
rect 397453 109304 400108 109306
rect 397453 109248 397458 109304
rect 397514 109248 400108 109304
rect 397453 109246 400108 109248
rect 397453 109243 397519 109246
rect 440325 109170 440391 109173
rect 439852 109168 440391 109170
rect 439852 109112 440330 109168
rect 440386 109112 440391 109168
rect 439852 109110 440391 109112
rect 440325 109107 440391 109110
rect 257521 109034 257587 109037
rect 238710 109032 257587 109034
rect 238710 108976 257526 109032
rect 257582 108976 257587 109032
rect 238710 108974 257587 108976
rect 214005 108898 214071 108901
rect 238710 108898 238770 108974
rect 257521 108971 257587 108974
rect 266261 109034 266327 109037
rect 266261 109032 267842 109034
rect 266261 108976 266266 109032
rect 266322 108976 267842 109032
rect 266261 108974 267842 108976
rect 266261 108971 266327 108974
rect 267782 108900 267842 108974
rect 214005 108896 217028 108898
rect 214005 108840 214010 108896
rect 214066 108840 217028 108896
rect 214005 108838 217028 108840
rect 228988 108838 238770 108898
rect 214005 108835 214071 108838
rect 267774 108836 267780 108900
rect 267844 108836 267850 108900
rect 164724 108762 165354 108768
rect 167729 108762 167795 108765
rect 164724 108760 167795 108762
rect 164724 108708 167734 108760
rect 165294 108704 167734 108708
rect 167790 108704 167795 108760
rect 165294 108702 167795 108704
rect 167729 108699 167795 108702
rect 264237 108762 264303 108765
rect 268150 108762 268210 109004
rect 264237 108760 268210 108762
rect 264237 108704 264242 108760
rect 264298 108704 268210 108760
rect 264237 108702 268210 108704
rect 264237 108699 264303 108702
rect 264421 108626 264487 108629
rect 264421 108624 268180 108626
rect 264421 108568 264426 108624
rect 264482 108568 268180 108624
rect 264421 108566 268180 108568
rect 264421 108563 264487 108566
rect 231761 108490 231827 108493
rect 282177 108490 282243 108493
rect 228988 108488 231827 108490
rect 228988 108432 231766 108488
rect 231822 108432 231827 108488
rect 228988 108430 231827 108432
rect 279956 108488 282243 108490
rect 279956 108432 282182 108488
rect 282238 108432 282243 108488
rect 279956 108430 282243 108432
rect 231761 108427 231827 108430
rect 282177 108427 282243 108430
rect 213913 108218 213979 108221
rect 397453 108218 397519 108221
rect 442901 108218 442967 108221
rect 213913 108216 217028 108218
rect 213913 108160 213918 108216
rect 213974 108160 217028 108216
rect 213913 108158 217028 108160
rect 258030 108158 268180 108218
rect 397453 108216 400108 108218
rect 397453 108160 397458 108216
rect 397514 108160 400108 108216
rect 397453 108158 400108 108160
rect 439852 108216 442967 108218
rect 439852 108160 442906 108216
rect 442962 108160 442967 108216
rect 439852 108158 442967 108160
rect 213913 108155 213979 108158
rect 246573 108082 246639 108085
rect 258030 108082 258090 108158
rect 397453 108155 397519 108158
rect 442901 108155 442967 108158
rect 246573 108080 258090 108082
rect 246573 108024 246578 108080
rect 246634 108024 258090 108080
rect 246573 108022 258090 108024
rect 246573 108019 246639 108022
rect 231485 107946 231551 107949
rect 228988 107944 231551 107946
rect 228988 107888 231490 107944
rect 231546 107888 231551 107944
rect 228988 107886 231551 107888
rect 231485 107883 231551 107886
rect 253289 107810 253355 107813
rect 282361 107810 282427 107813
rect 253289 107808 268180 107810
rect 253289 107752 253294 107808
rect 253350 107752 268180 107808
rect 253289 107750 268180 107752
rect 279956 107808 282427 107810
rect 279956 107752 282366 107808
rect 282422 107752 282427 107808
rect 279956 107750 282427 107752
rect 253289 107747 253355 107750
rect 282361 107747 282427 107750
rect 214005 107538 214071 107541
rect 245193 107538 245259 107541
rect 214005 107536 217028 107538
rect 214005 107480 214010 107536
rect 214066 107480 217028 107536
rect 214005 107478 217028 107480
rect 228988 107536 245259 107538
rect 228988 107480 245198 107536
rect 245254 107480 245259 107536
rect 228988 107478 245259 107480
rect 214005 107475 214071 107478
rect 245193 107475 245259 107478
rect 397545 107538 397611 107541
rect 397545 107536 400108 107538
rect 397545 107480 397550 107536
rect 397606 107480 400108 107536
rect 397545 107478 400108 107480
rect 397545 107475 397611 107478
rect 230933 107130 230999 107133
rect 228988 107128 230999 107130
rect 228988 107072 230938 107128
rect 230994 107072 230999 107128
rect 228988 107070 230999 107072
rect 230933 107067 230999 107070
rect 267958 107068 267964 107132
rect 268028 107130 268034 107132
rect 268150 107130 268210 107372
rect 442533 107266 442599 107269
rect 439852 107264 442599 107266
rect 439852 107208 442538 107264
rect 442594 107208 442599 107264
rect 439852 107206 442599 107208
rect 442533 107203 442599 107206
rect 268028 107070 268210 107130
rect 268028 107068 268034 107070
rect 264973 106994 265039 106997
rect 281625 106994 281691 106997
rect 264973 106992 268180 106994
rect 264973 106936 264978 106992
rect 265034 106936 268180 106992
rect 264973 106934 268180 106936
rect 279956 106992 281691 106994
rect 279956 106936 281630 106992
rect 281686 106936 281691 106992
rect 279956 106934 281691 106936
rect 264973 106931 265039 106934
rect 281625 106931 281691 106934
rect 166257 106858 166323 106861
rect 213913 106858 213979 106861
rect 166257 106856 200130 106858
rect 166257 106800 166262 106856
rect 166318 106800 200130 106856
rect 166257 106798 200130 106800
rect 166257 106795 166323 106798
rect 200070 106722 200130 106798
rect 213913 106856 217028 106858
rect 213913 106800 213918 106856
rect 213974 106800 217028 106856
rect 213913 106798 217028 106800
rect 213913 106795 213979 106798
rect 216121 106722 216187 106725
rect 200070 106720 216187 106722
rect 200070 106664 216126 106720
rect 216182 106664 216187 106720
rect 200070 106662 216187 106664
rect 216121 106659 216187 106662
rect 397453 106722 397519 106725
rect 397453 106720 400108 106722
rect 397453 106664 397458 106720
rect 397514 106664 400108 106720
rect 397453 106662 400108 106664
rect 397453 106659 397519 106662
rect 231577 106586 231643 106589
rect 228988 106584 231643 106586
rect 228988 106528 231582 106584
rect 231638 106528 231643 106584
rect 228988 106526 231643 106528
rect 231577 106523 231643 106526
rect 262949 106450 263015 106453
rect 440233 106450 440299 106453
rect 262949 106448 268180 106450
rect 262949 106392 262954 106448
rect 263010 106392 268180 106448
rect 262949 106390 268180 106392
rect 439852 106448 440299 106450
rect 439852 106392 440238 106448
rect 440294 106392 440299 106448
rect 439852 106390 440299 106392
rect 262949 106387 263015 106390
rect 440233 106387 440299 106390
rect 213361 106178 213427 106181
rect 234102 106178 234108 106180
rect 213361 106176 217028 106178
rect 213361 106120 213366 106176
rect 213422 106120 217028 106176
rect 213361 106118 217028 106120
rect 228988 106118 234108 106178
rect 213361 106115 213427 106118
rect 234102 106116 234108 106118
rect 234172 106116 234178 106180
rect 281809 106178 281875 106181
rect 279956 106176 281875 106178
rect 279956 106120 281814 106176
rect 281870 106120 281875 106176
rect 279956 106118 281875 106120
rect 281809 106115 281875 106118
rect 264973 106042 265039 106045
rect 264973 106040 268180 106042
rect 264973 105984 264978 106040
rect 265034 105984 268180 106040
rect 264973 105982 268180 105984
rect 264973 105979 265039 105982
rect 231393 105634 231459 105637
rect 228988 105632 231459 105634
rect 170581 105226 170647 105229
rect 216998 105226 217058 105604
rect 228988 105576 231398 105632
rect 231454 105576 231459 105632
rect 228988 105574 231459 105576
rect 231393 105571 231459 105574
rect 233877 105634 233943 105637
rect 246665 105634 246731 105637
rect 233877 105632 246731 105634
rect 233877 105576 233882 105632
rect 233938 105576 246670 105632
rect 246726 105576 246731 105632
rect 233877 105574 246731 105576
rect 233877 105571 233943 105574
rect 246665 105571 246731 105574
rect 250713 105634 250779 105637
rect 264094 105634 264100 105636
rect 250713 105632 264100 105634
rect 250713 105576 250718 105632
rect 250774 105576 264100 105632
rect 250713 105574 264100 105576
rect 250713 105571 250779 105574
rect 264094 105572 264100 105574
rect 264164 105572 264170 105636
rect 265065 105634 265131 105637
rect 397453 105634 397519 105637
rect 265065 105632 268180 105634
rect 265065 105576 265070 105632
rect 265126 105576 268180 105632
rect 265065 105574 268180 105576
rect 397453 105632 400108 105634
rect 397453 105576 397458 105632
rect 397514 105576 400108 105632
rect 397453 105574 400108 105576
rect 265065 105571 265131 105574
rect 397453 105571 397519 105574
rect 232589 105498 232655 105501
rect 258993 105498 259059 105501
rect 280286 105498 280292 105500
rect 232589 105496 259059 105498
rect 232589 105440 232594 105496
rect 232650 105440 258998 105496
rect 259054 105440 259059 105496
rect 232589 105438 259059 105440
rect 279956 105438 280292 105498
rect 232589 105435 232655 105438
rect 258993 105435 259059 105438
rect 280286 105436 280292 105438
rect 280356 105436 280362 105500
rect 442022 105362 442028 105364
rect 439852 105302 442028 105362
rect 442022 105300 442028 105302
rect 442092 105300 442098 105364
rect 231577 105226 231643 105229
rect 170581 105224 217058 105226
rect 170581 105168 170586 105224
rect 170642 105168 217058 105224
rect 170581 105166 217058 105168
rect 228988 105224 231643 105226
rect 228988 105168 231582 105224
rect 231638 105168 231643 105224
rect 228988 105166 231643 105168
rect 170581 105163 170647 105166
rect 231577 105163 231643 105166
rect 264329 105226 264395 105229
rect 264329 105224 268180 105226
rect 264329 105168 264334 105224
rect 264390 105168 268180 105224
rect 264329 105166 268180 105168
rect 264329 105163 264395 105166
rect 213913 104954 213979 104957
rect 213913 104952 217028 104954
rect 213913 104896 213918 104952
rect 213974 104896 217028 104952
rect 213913 104894 217028 104896
rect 213913 104891 213979 104894
rect 197302 104756 197308 104820
rect 197372 104818 197378 104820
rect 198641 104818 198707 104821
rect 242341 104818 242407 104821
rect 197372 104816 198707 104818
rect 197372 104760 198646 104816
rect 198702 104760 198707 104816
rect 197372 104758 198707 104760
rect 197372 104756 197378 104758
rect 198641 104755 198707 104758
rect 230614 104816 242407 104818
rect 230614 104760 242346 104816
rect 242402 104760 242407 104816
rect 397453 104818 397519 104821
rect 397453 104816 400108 104818
rect 230614 104758 242407 104760
rect 230614 104682 230674 104758
rect 242341 104755 242407 104758
rect 228988 104622 230674 104682
rect 230749 104682 230815 104685
rect 235349 104682 235415 104685
rect 230749 104680 235415 104682
rect 230749 104624 230754 104680
rect 230810 104624 235354 104680
rect 235410 104624 235415 104680
rect 230749 104622 235415 104624
rect 230749 104619 230815 104622
rect 235349 104619 235415 104622
rect 268150 104546 268210 104788
rect 397453 104760 397458 104816
rect 397514 104760 400108 104816
rect 397453 104758 400108 104760
rect 397453 104755 397519 104758
rect 258030 104486 268210 104546
rect 231761 104274 231827 104277
rect 228988 104272 231827 104274
rect 192569 103866 192635 103869
rect 216998 103866 217058 104244
rect 228988 104216 231766 104272
rect 231822 104216 231827 104272
rect 228988 104214 231827 104216
rect 231761 104211 231827 104214
rect 242525 104138 242591 104141
rect 258030 104138 258090 104486
rect 242525 104136 258090 104138
rect 242525 104080 242530 104136
rect 242586 104080 258090 104136
rect 242525 104078 258090 104080
rect 242525 104075 242591 104078
rect 238109 104002 238175 104005
rect 268150 104002 268210 104380
rect 279374 104277 279434 104652
rect 441981 104410 442047 104413
rect 439852 104408 442047 104410
rect 439852 104352 441986 104408
rect 442042 104352 442047 104408
rect 439852 104350 442047 104352
rect 441981 104347 442047 104350
rect 279325 104272 279434 104277
rect 279325 104216 279330 104272
rect 279386 104216 279434 104272
rect 279325 104214 279434 104216
rect 279325 104211 279391 104214
rect 382917 104138 382983 104141
rect 397637 104138 397703 104141
rect 382917 104136 400138 104138
rect 382917 104080 382922 104136
rect 382978 104080 397642 104136
rect 397698 104080 400138 104136
rect 382917 104078 400138 104080
rect 382917 104075 382983 104078
rect 397637 104075 397703 104078
rect 281901 104002 281967 104005
rect 238109 104000 268210 104002
rect 238109 103944 238114 104000
rect 238170 103944 268210 104000
rect 238109 103942 268210 103944
rect 279956 104000 281967 104002
rect 279956 103944 281906 104000
rect 281962 103944 281967 104000
rect 279956 103942 281967 103944
rect 238109 103939 238175 103942
rect 281901 103939 281967 103942
rect 192569 103864 217058 103866
rect 192569 103808 192574 103864
rect 192630 103808 217058 103864
rect 192569 103806 217058 103808
rect 264973 103866 265039 103869
rect 264973 103864 268180 103866
rect 264973 103808 264978 103864
rect 265034 103808 268180 103864
rect 264973 103806 268180 103808
rect 192569 103803 192635 103806
rect 264973 103803 265039 103806
rect 231485 103730 231551 103733
rect 228988 103728 231551 103730
rect 228988 103672 231490 103728
rect 231546 103672 231551 103728
rect 400078 103700 400138 104078
rect 228988 103670 231551 103672
rect 231485 103667 231551 103670
rect 213913 103594 213979 103597
rect 442901 103594 442967 103597
rect 213913 103592 217028 103594
rect 213913 103536 213918 103592
rect 213974 103536 217028 103592
rect 213913 103534 217028 103536
rect 439852 103592 442967 103594
rect 439852 103536 442906 103592
rect 442962 103536 442967 103592
rect 439852 103534 442967 103536
rect 213913 103531 213979 103534
rect 442901 103531 442967 103534
rect 264973 103458 265039 103461
rect 264973 103456 268180 103458
rect 264973 103400 264978 103456
rect 265034 103400 268180 103456
rect 264973 103398 268180 103400
rect 264973 103395 265039 103398
rect 231209 103322 231275 103325
rect 228988 103320 231275 103322
rect 228988 103264 231214 103320
rect 231270 103264 231275 103320
rect 228988 103262 231275 103264
rect 231209 103259 231275 103262
rect 281717 103186 281783 103189
rect 279956 103184 281783 103186
rect 279956 103128 281722 103184
rect 281778 103128 281783 103184
rect 279956 103126 281783 103128
rect 281717 103123 281783 103126
rect 258030 102990 268180 103050
rect 214005 102914 214071 102917
rect 214005 102912 217028 102914
rect 214005 102856 214010 102912
rect 214066 102856 217028 102912
rect 214005 102854 217028 102856
rect 214005 102851 214071 102854
rect 237966 102852 237972 102916
rect 238036 102914 238042 102916
rect 258030 102914 258090 102990
rect 238036 102854 258090 102914
rect 397453 102914 397519 102917
rect 397453 102912 400108 102914
rect 397453 102856 397458 102912
rect 397514 102856 400108 102912
rect 397453 102854 400108 102856
rect 238036 102852 238042 102854
rect 397453 102851 397519 102854
rect 231393 102778 231459 102781
rect 228988 102776 231459 102778
rect 228988 102720 231398 102776
rect 231454 102720 231459 102776
rect 228988 102718 231459 102720
rect 231393 102715 231459 102718
rect 231669 102778 231735 102781
rect 264513 102778 264579 102781
rect 231669 102776 264579 102778
rect 231669 102720 231674 102776
rect 231730 102720 264518 102776
rect 264574 102720 264579 102776
rect 231669 102718 264579 102720
rect 231669 102715 231735 102718
rect 264513 102715 264579 102718
rect 377397 102778 377463 102781
rect 398782 102778 398788 102780
rect 377397 102776 398788 102778
rect 377397 102720 377402 102776
rect 377458 102720 398788 102776
rect 377397 102718 398788 102720
rect 377397 102715 377463 102718
rect 398782 102716 398788 102718
rect 398852 102716 398858 102780
rect 264881 102642 264947 102645
rect 442717 102642 442783 102645
rect 264881 102640 268180 102642
rect 264881 102584 264886 102640
rect 264942 102584 268180 102640
rect 264881 102582 268180 102584
rect 439852 102640 442783 102642
rect 439852 102584 442722 102640
rect 442778 102584 442783 102640
rect 439852 102582 442783 102584
rect 264881 102579 264947 102582
rect 442717 102579 442783 102582
rect 67541 102370 67607 102373
rect 68142 102370 68816 102376
rect 231761 102370 231827 102373
rect 282821 102370 282887 102373
rect 67541 102368 68816 102370
rect 67541 102312 67546 102368
rect 67602 102316 68816 102368
rect 228988 102368 231827 102370
rect 67602 102312 68202 102316
rect 67541 102310 68202 102312
rect 228988 102312 231766 102368
rect 231822 102312 231827 102368
rect 228988 102310 231827 102312
rect 279956 102368 282887 102370
rect 279956 102312 282826 102368
rect 282882 102312 282887 102368
rect 279956 102310 282887 102312
rect 67541 102307 67607 102310
rect 231761 102307 231827 102310
rect 282821 102307 282887 102310
rect 213913 102234 213979 102237
rect 213913 102232 217028 102234
rect 213913 102176 213918 102232
rect 213974 102176 217028 102232
rect 213913 102174 217028 102176
rect 213913 102171 213979 102174
rect 262990 102172 262996 102236
rect 263060 102234 263066 102236
rect 263060 102174 268180 102234
rect 263060 102172 263066 102174
rect 231485 101826 231551 101829
rect 228988 101824 231551 101826
rect 228988 101768 231490 101824
rect 231546 101768 231551 101824
rect 228988 101766 231551 101768
rect 231485 101763 231551 101766
rect 264973 101826 265039 101829
rect 264973 101824 268180 101826
rect 264973 101768 264978 101824
rect 265034 101768 268180 101824
rect 264973 101766 268180 101768
rect 264973 101763 265039 101766
rect 284334 101690 284340 101692
rect 279956 101630 284340 101690
rect 284334 101628 284340 101630
rect 284404 101628 284410 101692
rect 397453 101690 397519 101693
rect 441613 101690 441679 101693
rect 397453 101688 400108 101690
rect 397453 101632 397458 101688
rect 397514 101632 400108 101688
rect 397453 101630 400108 101632
rect 439852 101688 441679 101690
rect 439852 101632 441618 101688
rect 441674 101632 441679 101688
rect 439852 101630 441679 101632
rect 397453 101627 397519 101630
rect 441613 101627 441679 101630
rect 213913 101554 213979 101557
rect 213913 101552 217028 101554
rect 213913 101496 213918 101552
rect 213974 101496 217028 101552
rect 213913 101494 217028 101496
rect 213913 101491 213979 101494
rect 164969 101418 165035 101421
rect 187141 101418 187207 101421
rect 231761 101418 231827 101421
rect 257613 101418 257679 101421
rect 164969 101416 187207 101418
rect 164969 101360 164974 101416
rect 165030 101360 187146 101416
rect 187202 101360 187207 101416
rect 164969 101358 187207 101360
rect 228988 101416 231827 101418
rect 228988 101360 231766 101416
rect 231822 101360 231827 101416
rect 228988 101358 231827 101360
rect 164969 101355 165035 101358
rect 187141 101355 187207 101358
rect 231761 101355 231827 101358
rect 238710 101416 257679 101418
rect 238710 101360 257618 101416
rect 257674 101360 257679 101416
rect 238710 101358 257679 101360
rect 231209 101282 231275 101285
rect 238710 101282 238770 101358
rect 257613 101355 257679 101358
rect 298737 101418 298803 101421
rect 298737 101416 412650 101418
rect 298737 101360 298742 101416
rect 298798 101360 412650 101416
rect 298737 101358 412650 101360
rect 298737 101355 298803 101358
rect 231209 101280 238770 101282
rect 231209 101224 231214 101280
rect 231270 101224 238770 101280
rect 231209 101222 238770 101224
rect 265065 101282 265131 101285
rect 367737 101282 367803 101285
rect 265065 101280 268180 101282
rect 265065 101224 265070 101280
rect 265126 101224 268180 101280
rect 265065 101222 268180 101224
rect 367737 101280 401426 101282
rect 367737 101224 367742 101280
rect 367798 101224 401426 101280
rect 367737 101222 401426 101224
rect 231209 101219 231275 101222
rect 265065 101219 265131 101222
rect 367737 101219 367803 101222
rect 214557 101010 214623 101013
rect 214557 101008 217028 101010
rect 214557 100952 214562 101008
rect 214618 100952 217028 101008
rect 214557 100950 217028 100952
rect 214557 100947 214623 100950
rect 230473 100874 230539 100877
rect 228988 100872 230539 100874
rect 228988 100816 230478 100872
rect 230534 100816 230539 100872
rect 228988 100814 230539 100816
rect 230473 100811 230539 100814
rect 247769 100874 247835 100877
rect 281717 100874 281783 100877
rect 247769 100872 268180 100874
rect 247769 100816 247774 100872
rect 247830 100816 268180 100872
rect 247769 100814 268180 100816
rect 279956 100872 281783 100874
rect 279956 100816 281722 100872
rect 281778 100816 281783 100872
rect 279956 100814 281783 100816
rect 247769 100811 247835 100814
rect 281717 100811 281783 100814
rect 397545 100874 397611 100877
rect 397545 100872 400108 100874
rect 397545 100816 397550 100872
rect 397606 100816 400108 100872
rect 397545 100814 400108 100816
rect 397545 100811 397611 100814
rect 67357 100738 67423 100741
rect 68142 100738 68816 100744
rect 67357 100736 68816 100738
rect 67357 100680 67362 100736
rect 67418 100684 68816 100736
rect 401366 100741 401426 101222
rect 412590 100874 412650 101358
rect 412590 100814 424978 100874
rect 401366 100736 401475 100741
rect 67418 100680 68202 100684
rect 67357 100678 68202 100680
rect 401366 100680 401414 100736
rect 401470 100680 401475 100736
rect 401366 100678 401475 100680
rect 67357 100675 67423 100678
rect 401409 100675 401475 100678
rect 421649 100738 421715 100741
rect 423990 100738 423996 100740
rect 421649 100736 423996 100738
rect 421649 100680 421654 100736
rect 421710 100680 423996 100736
rect 421649 100678 423996 100680
rect 421649 100675 421715 100678
rect 423990 100676 423996 100678
rect 424060 100676 424066 100740
rect 424918 100738 424978 100814
rect 425053 100738 425119 100741
rect 424918 100736 425119 100738
rect 424918 100680 425058 100736
rect 425114 100680 425119 100736
rect 424918 100678 425119 100680
rect 425053 100675 425119 100678
rect 425646 100676 425652 100740
rect 425716 100738 425722 100740
rect 428641 100738 428707 100741
rect 425716 100736 428707 100738
rect 425716 100680 428646 100736
rect 428702 100680 428707 100736
rect 425716 100678 428707 100680
rect 425716 100676 425722 100678
rect 428641 100675 428707 100678
rect 279366 100540 279372 100604
rect 279436 100540 279442 100604
rect 231761 100466 231827 100469
rect 228988 100464 231827 100466
rect 228988 100408 231766 100464
rect 231822 100408 231827 100464
rect 228988 100406 231827 100408
rect 231761 100403 231827 100406
rect 267181 100466 267247 100469
rect 267181 100464 268180 100466
rect 267181 100408 267186 100464
rect 267242 100408 268180 100464
rect 267181 100406 268180 100408
rect 267181 100403 267247 100406
rect 213913 100330 213979 100333
rect 213913 100328 217028 100330
rect 213913 100272 213918 100328
rect 213974 100272 217028 100328
rect 213913 100270 217028 100272
rect 213913 100267 213979 100270
rect 279374 100164 279434 100540
rect 173433 100058 173499 100061
rect 215293 100058 215359 100061
rect 173433 100056 215359 100058
rect 173433 100000 173438 100056
rect 173494 100000 215298 100056
rect 215354 100000 215359 100056
rect 173433 99998 215359 100000
rect 173433 99995 173499 99998
rect 215293 99995 215359 99998
rect 242341 100058 242407 100061
rect 262990 100058 262996 100060
rect 242341 100056 262996 100058
rect 242341 100000 242346 100056
rect 242402 100000 262996 100056
rect 242341 99998 262996 100000
rect 242341 99995 242407 99998
rect 262990 99996 262996 99998
rect 263060 99996 263066 100060
rect 265065 100058 265131 100061
rect 265065 100056 268180 100058
rect 265065 100000 265070 100056
rect 265126 100000 268180 100056
rect 265065 99998 268180 100000
rect 265065 99995 265131 99998
rect 231669 99922 231735 99925
rect 228988 99920 231735 99922
rect 228988 99864 231674 99920
rect 231730 99864 231735 99920
rect 228988 99862 231735 99864
rect 231669 99859 231735 99862
rect 392577 99786 392643 99789
rect 404445 99786 404511 99789
rect 392577 99784 404511 99786
rect 392577 99728 392582 99784
rect 392638 99728 404450 99784
rect 404506 99728 404511 99784
rect 392577 99726 404511 99728
rect 392577 99723 392643 99726
rect 404445 99723 404511 99726
rect 214465 99650 214531 99653
rect 264973 99650 265039 99653
rect 385677 99650 385743 99653
rect 404537 99650 404603 99653
rect 405549 99650 405615 99653
rect 214465 99648 217028 99650
rect 214465 99592 214470 99648
rect 214526 99592 217028 99648
rect 214465 99590 217028 99592
rect 264973 99648 268180 99650
rect 264973 99592 264978 99648
rect 265034 99592 268180 99648
rect 264973 99590 268180 99592
rect 385677 99648 405615 99650
rect 385677 99592 385682 99648
rect 385738 99592 404542 99648
rect 404598 99592 405554 99648
rect 405610 99592 405615 99648
rect 385677 99590 405615 99592
rect 214465 99587 214531 99590
rect 264973 99587 265039 99590
rect 385677 99587 385743 99590
rect 404537 99587 404603 99590
rect 405549 99587 405615 99590
rect 230565 99514 230631 99517
rect 228988 99512 230631 99514
rect 228988 99456 230570 99512
rect 230626 99456 230631 99512
rect 228988 99454 230631 99456
rect 230565 99451 230631 99454
rect 387057 99514 387123 99517
rect 422109 99514 422175 99517
rect 387057 99512 422175 99514
rect 387057 99456 387062 99512
rect 387118 99456 422114 99512
rect 422170 99456 422175 99512
rect 387057 99454 422175 99456
rect 387057 99451 387123 99454
rect 422109 99451 422175 99454
rect 425881 99514 425947 99517
rect 439270 99514 439330 100572
rect 425881 99512 439330 99514
rect 425881 99456 425886 99512
rect 425942 99456 439330 99512
rect 425881 99454 439330 99456
rect 580165 99514 580231 99517
rect 583520 99514 584960 99604
rect 580165 99512 584960 99514
rect 580165 99456 580170 99512
rect 580226 99456 584960 99512
rect 580165 99454 584960 99456
rect 425881 99451 425947 99454
rect 580165 99451 580231 99454
rect 282821 99378 282887 99381
rect 279956 99376 282887 99378
rect 279956 99320 282826 99376
rect 282882 99320 282887 99376
rect 279956 99318 282887 99320
rect 282821 99315 282887 99318
rect 292665 99378 292731 99381
rect 293217 99378 293283 99381
rect 397453 99378 397519 99381
rect 292665 99376 397519 99378
rect 292665 99320 292670 99376
rect 292726 99320 293222 99376
rect 293278 99320 397458 99376
rect 397514 99320 397519 99376
rect 292665 99318 397519 99320
rect 292665 99315 292731 99318
rect 293217 99315 293283 99318
rect 397453 99315 397519 99318
rect 398782 99316 398788 99380
rect 398852 99378 398858 99380
rect 407573 99378 407639 99381
rect 398852 99376 407639 99378
rect 398852 99320 407578 99376
rect 407634 99320 407639 99376
rect 583520 99364 584960 99454
rect 398852 99318 407639 99320
rect 398852 99316 398858 99318
rect 407573 99315 407639 99318
rect 267774 99180 267780 99244
rect 267844 99242 267850 99244
rect 388437 99242 388503 99245
rect 429653 99242 429719 99245
rect 267844 99182 268180 99242
rect 388437 99240 429719 99242
rect 388437 99184 388442 99240
rect 388498 99184 429658 99240
rect 429714 99184 429719 99240
rect 388437 99182 429719 99184
rect 267844 99180 267850 99182
rect 388437 99179 388503 99182
rect 429653 99179 429719 99182
rect 214005 98970 214071 98973
rect 230749 98970 230815 98973
rect 214005 98968 217028 98970
rect 214005 98912 214010 98968
rect 214066 98912 217028 98968
rect 214005 98910 217028 98912
rect 228988 98968 230815 98970
rect 228988 98912 230754 98968
rect 230810 98912 230815 98968
rect 228988 98910 230815 98912
rect 214005 98907 214071 98910
rect 230749 98907 230815 98910
rect 210601 98698 210667 98701
rect 215937 98698 216003 98701
rect 210601 98696 216003 98698
rect 210601 98640 210606 98696
rect 210662 98640 215942 98696
rect 215998 98640 216003 98696
rect 210601 98638 216003 98640
rect 210601 98635 210667 98638
rect 215937 98635 216003 98638
rect 231393 98698 231459 98701
rect 261661 98698 261727 98701
rect 231393 98696 261727 98698
rect 231393 98640 231398 98696
rect 231454 98640 261666 98696
rect 261722 98640 261727 98696
rect 231393 98638 261727 98640
rect 231393 98635 231459 98638
rect 261661 98635 261727 98638
rect 264973 98698 265039 98701
rect 264973 98696 268180 98698
rect 264973 98640 264978 98696
rect 265034 98640 268180 98696
rect 264973 98638 268180 98640
rect 264973 98635 265039 98638
rect 230749 98562 230815 98565
rect 281993 98562 282059 98565
rect 228988 98560 230815 98562
rect 228988 98504 230754 98560
rect 230810 98504 230815 98560
rect 228988 98502 230815 98504
rect 279956 98560 282059 98562
rect 279956 98504 281998 98560
rect 282054 98504 282059 98560
rect 279956 98502 282059 98504
rect 230749 98499 230815 98502
rect 281993 98499 282059 98502
rect 213913 98290 213979 98293
rect 265801 98290 265867 98293
rect 213913 98288 217028 98290
rect 213913 98232 213918 98288
rect 213974 98232 217028 98288
rect 213913 98230 217028 98232
rect 265801 98288 268180 98290
rect 265801 98232 265806 98288
rect 265862 98232 268180 98288
rect 265801 98230 268180 98232
rect 213913 98227 213979 98230
rect 265801 98227 265867 98230
rect 231025 98018 231091 98021
rect 228988 98016 231091 98018
rect 228988 97960 231030 98016
rect 231086 97960 231091 98016
rect 228988 97958 231091 97960
rect 231025 97955 231091 97958
rect 265065 97882 265131 97885
rect 282821 97882 282887 97885
rect 265065 97880 268180 97882
rect 265065 97824 265070 97880
rect 265126 97824 268180 97880
rect 265065 97822 268180 97824
rect 279956 97880 282887 97882
rect 279956 97824 282826 97880
rect 282882 97824 282887 97880
rect 279956 97822 282887 97824
rect 265065 97819 265131 97822
rect 282821 97819 282887 97822
rect 394049 97746 394115 97749
rect 427813 97746 427879 97749
rect 394049 97744 427879 97746
rect -960 97610 480 97700
rect 394049 97688 394054 97744
rect 394110 97688 427818 97744
rect 427874 97688 427879 97744
rect 394049 97686 427879 97688
rect 394049 97683 394115 97686
rect 427813 97683 427879 97686
rect 3509 97610 3575 97613
rect -960 97608 3575 97610
rect -960 97552 3514 97608
rect 3570 97552 3575 97608
rect -960 97550 3575 97552
rect -960 97460 480 97550
rect 3509 97547 3575 97550
rect 213913 97610 213979 97613
rect 231393 97610 231459 97613
rect 213913 97608 217028 97610
rect 213913 97552 213918 97608
rect 213974 97552 217028 97608
rect 213913 97550 217028 97552
rect 228988 97608 231459 97610
rect 228988 97552 231398 97608
rect 231454 97552 231459 97608
rect 228988 97550 231459 97552
rect 213913 97547 213979 97550
rect 231393 97547 231459 97550
rect 264094 97412 264100 97476
rect 264164 97474 264170 97476
rect 264164 97414 268180 97474
rect 264164 97412 264170 97414
rect 238710 97142 258090 97202
rect 229134 97066 229140 97068
rect 228988 97006 229140 97066
rect 229134 97004 229140 97006
rect 229204 97004 229210 97068
rect 214741 96930 214807 96933
rect 214741 96928 217028 96930
rect 214741 96872 214746 96928
rect 214802 96872 217028 96928
rect 214741 96870 217028 96872
rect 214741 96867 214807 96870
rect 229093 96794 229159 96797
rect 238710 96794 238770 97142
rect 229093 96792 238770 96794
rect 229093 96736 229098 96792
rect 229154 96736 238770 96792
rect 229093 96734 238770 96736
rect 258030 96794 258090 97142
rect 264973 97066 265039 97069
rect 282729 97066 282795 97069
rect 264973 97064 268180 97066
rect 264973 97008 264978 97064
rect 265034 97008 268180 97064
rect 264973 97006 268180 97008
rect 279956 97064 282795 97066
rect 279956 97008 282734 97064
rect 282790 97008 282795 97064
rect 279956 97006 282795 97008
rect 264973 97003 265039 97006
rect 282729 97003 282795 97006
rect 432597 96930 432663 96933
rect 438485 96930 438551 96933
rect 432597 96928 438551 96930
rect 432597 96872 432602 96928
rect 432658 96872 438490 96928
rect 438546 96872 438551 96928
rect 432597 96870 438551 96872
rect 432597 96867 432663 96870
rect 438485 96867 438551 96870
rect 258030 96734 268210 96794
rect 229093 96731 229159 96734
rect 231301 96658 231367 96661
rect 228988 96656 231367 96658
rect 228988 96600 231306 96656
rect 231362 96600 231367 96656
rect 268150 96628 268210 96734
rect 228988 96598 231367 96600
rect 231301 96595 231367 96598
rect 361481 96522 361547 96525
rect 416405 96522 416471 96525
rect 361481 96520 416471 96522
rect 361481 96464 361486 96520
rect 361542 96464 416410 96520
rect 416466 96464 416471 96520
rect 361481 96462 416471 96464
rect 361481 96459 361547 96462
rect 416405 96459 416471 96462
rect 214833 96386 214899 96389
rect 282821 96386 282887 96389
rect 214833 96384 217028 96386
rect 214833 96328 214838 96384
rect 214894 96328 217028 96384
rect 214833 96326 217028 96328
rect 279956 96384 282887 96386
rect 279956 96328 282826 96384
rect 282882 96328 282887 96384
rect 279956 96326 282887 96328
rect 214833 96323 214899 96326
rect 282821 96323 282887 96326
rect 230473 96250 230539 96253
rect 228988 96248 230539 96250
rect 228988 96192 230478 96248
rect 230534 96192 230539 96248
rect 228988 96190 230539 96192
rect 230473 96187 230539 96190
rect 225045 95980 225111 95981
rect 226425 95980 226491 95981
rect 225045 95976 225092 95980
rect 225156 95978 225162 95980
rect 226374 95978 226380 95980
rect 225045 95920 225050 95976
rect 225045 95916 225092 95920
rect 225156 95918 225202 95978
rect 226334 95918 226380 95978
rect 226444 95976 226491 95980
rect 226486 95920 226491 95976
rect 225156 95916 225162 95918
rect 226374 95916 226380 95918
rect 226444 95916 226491 95920
rect 226926 95916 226932 95980
rect 226996 95978 227002 95980
rect 229001 95978 229067 95981
rect 226996 95976 229067 95978
rect 226996 95920 229006 95976
rect 229062 95920 229067 95976
rect 226996 95918 229067 95920
rect 226996 95916 227002 95918
rect 225045 95915 225111 95916
rect 226425 95915 226491 95916
rect 229001 95915 229067 95918
rect 241513 95706 241579 95709
rect 242750 95706 242756 95708
rect 241513 95704 242756 95706
rect 241513 95648 241518 95704
rect 241574 95648 242756 95704
rect 241513 95646 242756 95648
rect 241513 95643 241579 95646
rect 242750 95644 242756 95646
rect 242820 95644 242826 95708
rect 229001 95570 229067 95573
rect 267825 95570 267891 95573
rect 229001 95568 267891 95570
rect 229001 95512 229006 95568
rect 229062 95512 267830 95568
rect 267886 95512 267891 95568
rect 229001 95510 267891 95512
rect 229001 95507 229067 95510
rect 267825 95507 267891 95510
rect 228541 95298 228607 95301
rect 268150 95298 268210 96220
rect 429837 95842 429903 95845
rect 442206 95842 442212 95844
rect 429837 95840 442212 95842
rect 429837 95784 429842 95840
rect 429898 95784 442212 95840
rect 429837 95782 442212 95784
rect 429837 95779 429903 95782
rect 442206 95780 442212 95782
rect 442276 95780 442282 95844
rect 228541 95296 268210 95298
rect 228541 95240 228546 95296
rect 228602 95240 268210 95296
rect 228541 95238 268210 95240
rect 410057 95298 410123 95301
rect 582465 95298 582531 95301
rect 410057 95296 582531 95298
rect 410057 95240 410062 95296
rect 410118 95240 582470 95296
rect 582526 95240 582531 95296
rect 410057 95238 582531 95240
rect 228541 95235 228607 95238
rect 410057 95235 410123 95238
rect 582465 95235 582531 95238
rect 393957 95162 394023 95165
rect 437197 95162 437263 95165
rect 393957 95160 437263 95162
rect 393957 95104 393962 95160
rect 394018 95104 437202 95160
rect 437258 95104 437263 95160
rect 393957 95102 437263 95104
rect 393957 95099 394023 95102
rect 437197 95099 437263 95102
rect 67541 95026 67607 95029
rect 165521 95026 165587 95029
rect 67541 95024 165587 95026
rect 67541 94968 67546 95024
rect 67602 94968 165526 95024
rect 165582 94968 165587 95024
rect 67541 94966 165587 94968
rect 67541 94963 67607 94966
rect 165521 94963 165587 94966
rect 113173 94756 113239 94757
rect 130745 94756 130811 94757
rect 113136 94692 113142 94756
rect 113206 94754 113239 94756
rect 113206 94752 113298 94754
rect 113234 94696 113298 94752
rect 113206 94694 113298 94696
rect 113206 94692 113239 94694
rect 130680 94692 130686 94756
rect 130750 94754 130811 94756
rect 130750 94752 130842 94754
rect 130806 94696 130842 94752
rect 130750 94694 130842 94696
rect 130750 94692 130811 94694
rect 151486 94692 151492 94756
rect 151556 94754 151562 94756
rect 151760 94754 151766 94756
rect 151556 94694 151766 94754
rect 151556 94692 151562 94694
rect 151760 94692 151766 94694
rect 151830 94692 151836 94756
rect 220813 94754 220879 94757
rect 230422 94754 230428 94756
rect 220813 94752 230428 94754
rect 220813 94696 220818 94752
rect 220874 94696 230428 94752
rect 220813 94694 230428 94696
rect 113173 94691 113239 94692
rect 130745 94691 130811 94692
rect 220813 94691 220879 94694
rect 230422 94692 230428 94694
rect 230492 94692 230498 94756
rect 186957 94618 187023 94621
rect 224217 94618 224283 94621
rect 186957 94616 224283 94618
rect 186957 94560 186962 94616
rect 187018 94560 224222 94616
rect 224278 94560 224283 94616
rect 186957 94558 224283 94560
rect 186957 94555 187023 94558
rect 224217 94555 224283 94558
rect 225597 94618 225663 94621
rect 264881 94618 264947 94621
rect 225597 94616 264947 94618
rect 225597 94560 225602 94616
rect 225658 94560 264886 94616
rect 264942 94560 264947 94616
rect 225597 94558 264947 94560
rect 225597 94555 225663 94558
rect 264881 94555 264947 94558
rect 267590 94556 267596 94620
rect 267660 94618 267666 94620
rect 270493 94618 270559 94621
rect 267660 94616 270559 94618
rect 267660 94560 270498 94616
rect 270554 94560 270559 94616
rect 267660 94558 270559 94560
rect 267660 94556 267666 94558
rect 270493 94555 270559 94558
rect 162853 94482 162919 94485
rect 206369 94482 206435 94485
rect 162853 94480 206435 94482
rect 162853 94424 162858 94480
rect 162914 94424 206374 94480
rect 206430 94424 206435 94480
rect 162853 94422 206435 94424
rect 162853 94419 162919 94422
rect 206369 94419 206435 94422
rect 214414 94420 214420 94484
rect 214484 94482 214490 94484
rect 271873 94482 271939 94485
rect 214484 94480 271939 94482
rect 214484 94424 271878 94480
rect 271934 94424 271939 94480
rect 214484 94422 271939 94424
rect 214484 94420 214490 94422
rect 271873 94419 271939 94422
rect 349797 94482 349863 94485
rect 393313 94482 393379 94485
rect 349797 94480 393379 94482
rect 349797 94424 349802 94480
rect 349858 94424 393318 94480
rect 393374 94424 393379 94480
rect 349797 94422 393379 94424
rect 349797 94419 349863 94422
rect 393313 94419 393379 94422
rect 100886 93876 100892 93940
rect 100956 93938 100962 93940
rect 202413 93938 202479 93941
rect 100956 93936 202479 93938
rect 100956 93880 202418 93936
rect 202474 93880 202479 93936
rect 100956 93878 202479 93880
rect 100956 93876 100962 93878
rect 202413 93875 202479 93878
rect 99230 93740 99236 93804
rect 99300 93802 99306 93804
rect 205173 93802 205239 93805
rect 99300 93800 205239 93802
rect 99300 93744 205178 93800
rect 205234 93744 205239 93800
rect 99300 93742 205239 93744
rect 99300 93740 99306 93742
rect 205173 93739 205239 93742
rect 206461 93802 206527 93805
rect 408585 93802 408651 93805
rect 206461 93800 408651 93802
rect 206461 93744 206466 93800
rect 206522 93744 408590 93800
rect 408646 93744 408651 93800
rect 206461 93742 408651 93744
rect 206461 93739 206527 93742
rect 408585 93739 408651 93742
rect 118182 93604 118188 93668
rect 118252 93666 118258 93668
rect 196801 93666 196867 93669
rect 118252 93664 196867 93666
rect 118252 93608 196806 93664
rect 196862 93608 196867 93664
rect 118252 93606 196867 93608
rect 118252 93604 118258 93606
rect 196801 93603 196867 93606
rect 228766 93604 228772 93668
rect 228836 93666 228842 93668
rect 260741 93666 260807 93669
rect 228836 93664 260807 93666
rect 228836 93608 260746 93664
rect 260802 93608 260807 93664
rect 228836 93606 260807 93608
rect 228836 93604 228842 93606
rect 260741 93603 260807 93606
rect 110086 93468 110092 93532
rect 110156 93530 110162 93532
rect 169293 93530 169359 93533
rect 110156 93528 169359 93530
rect 110156 93472 169298 93528
rect 169354 93472 169359 93528
rect 110156 93470 169359 93472
rect 110156 93468 110162 93470
rect 169293 93467 169359 93470
rect 119705 93396 119771 93397
rect 123017 93396 123083 93397
rect 119654 93394 119660 93396
rect 119614 93334 119660 93394
rect 119724 93392 119771 93396
rect 122966 93394 122972 93396
rect 119766 93336 119771 93392
rect 119654 93332 119660 93334
rect 119724 93332 119771 93336
rect 122926 93334 122972 93394
rect 123036 93392 123083 93396
rect 123078 93336 123083 93392
rect 122966 93332 122972 93334
rect 123036 93332 123083 93336
rect 119705 93331 119771 93332
rect 123017 93331 123083 93332
rect 103278 93196 103284 93260
rect 103348 93258 103354 93260
rect 103421 93258 103487 93261
rect 103348 93256 103487 93258
rect 103348 93200 103426 93256
rect 103482 93200 103487 93256
rect 103348 93198 103487 93200
rect 103348 93196 103354 93198
rect 103421 93195 103487 93198
rect 218789 93122 218855 93125
rect 229921 93122 229987 93125
rect 218789 93120 229987 93122
rect 218789 93064 218794 93120
rect 218850 93064 229926 93120
rect 229982 93064 229987 93120
rect 218789 93062 229987 93064
rect 218789 93059 218855 93062
rect 229921 93059 229987 93062
rect 74809 92444 74875 92445
rect 74758 92442 74764 92444
rect 74718 92382 74764 92442
rect 74828 92440 74875 92444
rect 74870 92384 74875 92440
rect 74758 92380 74764 92382
rect 74828 92380 74875 92384
rect 97206 92380 97212 92444
rect 97276 92442 97282 92444
rect 97349 92442 97415 92445
rect 97276 92440 97415 92442
rect 97276 92384 97354 92440
rect 97410 92384 97415 92440
rect 97276 92382 97415 92384
rect 97276 92380 97282 92382
rect 74809 92379 74875 92380
rect 97349 92379 97415 92382
rect 99966 92380 99972 92444
rect 100036 92442 100042 92444
rect 100109 92442 100175 92445
rect 100036 92440 100175 92442
rect 100036 92384 100114 92440
rect 100170 92384 100175 92440
rect 100036 92382 100175 92384
rect 100036 92380 100042 92382
rect 100109 92379 100175 92382
rect 102726 92380 102732 92444
rect 102796 92442 102802 92444
rect 103145 92442 103211 92445
rect 102796 92440 103211 92442
rect 102796 92384 103150 92440
rect 103206 92384 103211 92440
rect 102796 92382 103211 92384
rect 102796 92380 102802 92382
rect 103145 92379 103211 92382
rect 108062 92380 108068 92444
rect 108132 92442 108138 92444
rect 108573 92442 108639 92445
rect 116761 92444 116827 92445
rect 124121 92444 124187 92445
rect 134425 92444 134491 92445
rect 151353 92444 151419 92445
rect 116710 92442 116716 92444
rect 108132 92440 108639 92442
rect 108132 92384 108578 92440
rect 108634 92384 108639 92440
rect 108132 92382 108639 92384
rect 116670 92382 116716 92442
rect 116780 92440 116827 92444
rect 124070 92442 124076 92444
rect 116822 92384 116827 92440
rect 108132 92380 108138 92382
rect 108573 92379 108639 92382
rect 116710 92380 116716 92382
rect 116780 92380 116827 92384
rect 124030 92382 124076 92442
rect 124140 92440 124187 92444
rect 134374 92442 134380 92444
rect 124182 92384 124187 92440
rect 124070 92380 124076 92382
rect 124140 92380 124187 92384
rect 134334 92382 134380 92442
rect 134444 92440 134491 92444
rect 151302 92442 151308 92444
rect 134486 92384 134491 92440
rect 134374 92380 134380 92382
rect 134444 92380 134491 92384
rect 151262 92382 151308 92442
rect 151372 92440 151419 92444
rect 151414 92384 151419 92440
rect 151302 92380 151308 92382
rect 151372 92380 151419 92384
rect 116761 92379 116827 92380
rect 124121 92379 124187 92380
rect 134425 92379 134491 92380
rect 151353 92379 151419 92380
rect 209313 92442 209379 92445
rect 425421 92442 425487 92445
rect 209313 92440 425487 92442
rect 209313 92384 209318 92440
rect 209374 92384 425426 92440
rect 425482 92384 425487 92440
rect 209313 92382 425487 92384
rect 209313 92379 209379 92382
rect 425421 92379 425487 92382
rect 106774 92244 106780 92308
rect 106844 92306 106850 92308
rect 209129 92306 209195 92309
rect 106844 92304 209195 92306
rect 106844 92248 209134 92304
rect 209190 92248 209195 92304
rect 106844 92246 209195 92248
rect 106844 92244 106850 92246
rect 209129 92243 209195 92246
rect 253054 92244 253060 92308
rect 253124 92306 253130 92308
rect 275921 92306 275987 92309
rect 253124 92304 275987 92306
rect 253124 92248 275926 92304
rect 275982 92248 275987 92304
rect 253124 92246 275987 92248
rect 253124 92244 253130 92246
rect 275921 92243 275987 92246
rect 88057 92172 88123 92173
rect 88006 92170 88012 92172
rect 87966 92110 88012 92170
rect 88076 92168 88123 92172
rect 88118 92112 88123 92168
rect 88006 92108 88012 92110
rect 88076 92108 88123 92112
rect 133086 92108 133092 92172
rect 133156 92170 133162 92172
rect 178677 92170 178743 92173
rect 133156 92168 178743 92170
rect 133156 92112 178682 92168
rect 178738 92112 178743 92168
rect 133156 92110 178743 92112
rect 133156 92108 133162 92110
rect 88057 92107 88123 92108
rect 178677 92107 178743 92110
rect 91318 91972 91324 92036
rect 91388 92034 91394 92036
rect 91645 92034 91711 92037
rect 91388 92032 91711 92034
rect 91388 91976 91650 92032
rect 91706 91976 91711 92032
rect 91388 91974 91711 91976
rect 91388 91972 91394 91974
rect 91645 91971 91711 91974
rect 109166 91700 109172 91764
rect 109236 91762 109242 91764
rect 110137 91762 110203 91765
rect 109236 91760 110203 91762
rect 109236 91704 110142 91760
rect 110198 91704 110203 91760
rect 109236 91702 110203 91704
rect 109236 91700 109242 91702
rect 110137 91699 110203 91702
rect 120574 91700 120580 91764
rect 120644 91762 120650 91764
rect 121177 91762 121243 91765
rect 120644 91760 121243 91762
rect 120644 91704 121182 91760
rect 121238 91704 121243 91760
rect 120644 91702 121243 91704
rect 120644 91700 120650 91702
rect 121177 91699 121243 91702
rect 136030 91700 136036 91764
rect 136100 91762 136106 91764
rect 136449 91762 136515 91765
rect 136100 91760 136515 91762
rect 136100 91704 136454 91760
rect 136510 91704 136515 91760
rect 136100 91702 136515 91704
rect 136100 91700 136106 91702
rect 136449 91699 136515 91702
rect 221457 91762 221523 91765
rect 254761 91762 254827 91765
rect 221457 91760 254827 91762
rect 221457 91704 221462 91760
rect 221518 91704 254766 91760
rect 254822 91704 254827 91760
rect 221457 91702 254827 91704
rect 221457 91699 221523 91702
rect 254761 91699 254827 91702
rect 101990 91564 101996 91628
rect 102060 91626 102066 91628
rect 210509 91626 210575 91629
rect 102060 91624 210575 91626
rect 102060 91568 210514 91624
rect 210570 91568 210575 91624
rect 102060 91566 210575 91568
rect 102060 91564 102066 91566
rect 210509 91563 210575 91566
rect 126697 91492 126763 91493
rect 126646 91490 126652 91492
rect 126606 91430 126652 91490
rect 126716 91488 126763 91492
rect 126758 91432 126763 91488
rect 126646 91428 126652 91430
rect 126716 91428 126763 91432
rect 126697 91427 126763 91428
rect 85798 91292 85804 91356
rect 85868 91354 85874 91356
rect 86861 91354 86927 91357
rect 95049 91356 95115 91357
rect 94998 91354 95004 91356
rect 85868 91352 86927 91354
rect 85868 91296 86866 91352
rect 86922 91296 86927 91352
rect 85868 91294 86927 91296
rect 94958 91294 95004 91354
rect 95068 91352 95115 91356
rect 95110 91296 95115 91352
rect 85868 91292 85874 91294
rect 86861 91291 86927 91294
rect 94998 91292 95004 91294
rect 95068 91292 95115 91296
rect 98494 91292 98500 91356
rect 98564 91354 98570 91356
rect 98729 91354 98795 91357
rect 98564 91352 98795 91354
rect 98564 91296 98734 91352
rect 98790 91296 98795 91352
rect 98564 91294 98795 91296
rect 98564 91292 98570 91294
rect 95049 91291 95115 91292
rect 98729 91291 98795 91294
rect 110638 91292 110644 91356
rect 110708 91354 110714 91356
rect 111701 91354 111767 91357
rect 110708 91352 111767 91354
rect 110708 91296 111706 91352
rect 111762 91296 111767 91352
rect 110708 91294 111767 91296
rect 110708 91292 110714 91294
rect 111701 91291 111767 91294
rect 113214 91292 113220 91356
rect 113284 91354 113290 91356
rect 114369 91354 114435 91357
rect 115473 91356 115539 91357
rect 115422 91354 115428 91356
rect 113284 91352 114435 91354
rect 113284 91296 114374 91352
rect 114430 91296 114435 91352
rect 113284 91294 114435 91296
rect 115382 91294 115428 91354
rect 115492 91352 115539 91356
rect 115534 91296 115539 91352
rect 113284 91292 113290 91294
rect 114369 91291 114435 91294
rect 115422 91292 115428 91294
rect 115492 91292 115539 91296
rect 115473 91291 115539 91292
rect 115749 91356 115815 91357
rect 115749 91352 115796 91356
rect 115860 91354 115866 91356
rect 115749 91296 115754 91352
rect 115749 91292 115796 91296
rect 115860 91294 115906 91354
rect 115860 91292 115866 91294
rect 124438 91292 124444 91356
rect 124508 91354 124514 91356
rect 125501 91354 125567 91357
rect 124508 91352 125567 91354
rect 124508 91296 125506 91352
rect 125562 91296 125567 91352
rect 124508 91294 125567 91296
rect 124508 91292 124514 91294
rect 115749 91291 115815 91292
rect 125501 91291 125567 91294
rect 125726 91292 125732 91356
rect 125796 91354 125802 91356
rect 126697 91354 126763 91357
rect 151537 91356 151603 91357
rect 151486 91354 151492 91356
rect 125796 91352 126763 91354
rect 125796 91296 126702 91352
rect 126758 91296 126763 91352
rect 125796 91294 126763 91296
rect 151446 91294 151492 91354
rect 151556 91352 151603 91356
rect 151598 91296 151603 91352
rect 125796 91292 125802 91294
rect 126697 91291 126763 91294
rect 151486 91292 151492 91294
rect 151556 91292 151603 91296
rect 151537 91291 151603 91292
rect 84326 91156 84332 91220
rect 84396 91218 84402 91220
rect 85481 91218 85547 91221
rect 86769 91220 86835 91221
rect 86718 91218 86724 91220
rect 84396 91216 85547 91218
rect 84396 91160 85486 91216
rect 85542 91160 85547 91216
rect 84396 91158 85547 91160
rect 86678 91158 86724 91218
rect 86788 91216 86835 91220
rect 86830 91160 86835 91216
rect 84396 91156 84402 91158
rect 85481 91155 85547 91158
rect 86718 91156 86724 91158
rect 86788 91156 86835 91160
rect 88926 91156 88932 91220
rect 88996 91218 89002 91220
rect 89069 91218 89135 91221
rect 88996 91216 89135 91218
rect 88996 91160 89074 91216
rect 89130 91160 89135 91216
rect 88996 91158 89135 91160
rect 88996 91156 89002 91158
rect 86769 91155 86835 91156
rect 89069 91155 89135 91158
rect 90214 91156 90220 91220
rect 90284 91218 90290 91220
rect 91001 91218 91067 91221
rect 90284 91216 91067 91218
rect 90284 91160 91006 91216
rect 91062 91160 91067 91216
rect 90284 91158 91067 91160
rect 90284 91156 90290 91158
rect 91001 91155 91067 91158
rect 92606 91156 92612 91220
rect 92676 91218 92682 91220
rect 93669 91218 93735 91221
rect 92676 91216 93735 91218
rect 92676 91160 93674 91216
rect 93730 91160 93735 91216
rect 92676 91158 93735 91160
rect 92676 91156 92682 91158
rect 93669 91155 93735 91158
rect 93894 91156 93900 91220
rect 93964 91218 93970 91220
rect 95141 91218 95207 91221
rect 93964 91216 95207 91218
rect 93964 91160 95146 91216
rect 95202 91160 95207 91216
rect 93964 91158 95207 91160
rect 93964 91156 93970 91158
rect 95141 91155 95207 91158
rect 96286 91156 96292 91220
rect 96356 91218 96362 91220
rect 96521 91218 96587 91221
rect 96356 91216 96587 91218
rect 96356 91160 96526 91216
rect 96582 91160 96587 91216
rect 96356 91158 96587 91160
rect 96356 91156 96362 91158
rect 96521 91155 96587 91158
rect 96654 91156 96660 91220
rect 96724 91218 96730 91220
rect 97809 91218 97875 91221
rect 96724 91216 97875 91218
rect 96724 91160 97814 91216
rect 97870 91160 97875 91216
rect 96724 91158 97875 91160
rect 96724 91156 96730 91158
rect 97809 91155 97875 91158
rect 98126 91156 98132 91220
rect 98196 91218 98202 91220
rect 99281 91218 99347 91221
rect 100569 91220 100635 91221
rect 100518 91218 100524 91220
rect 98196 91216 99347 91218
rect 98196 91160 99286 91216
rect 99342 91160 99347 91216
rect 98196 91158 99347 91160
rect 100478 91158 100524 91218
rect 100588 91216 100635 91220
rect 100630 91160 100635 91216
rect 98196 91156 98202 91158
rect 99281 91155 99347 91158
rect 100518 91156 100524 91158
rect 100588 91156 100635 91160
rect 101806 91156 101812 91220
rect 101876 91218 101882 91220
rect 102041 91218 102107 91221
rect 104249 91220 104315 91221
rect 104198 91218 104204 91220
rect 101876 91216 102107 91218
rect 101876 91160 102046 91216
rect 102102 91160 102107 91216
rect 101876 91158 102107 91160
rect 104158 91158 104204 91218
rect 104268 91216 104315 91220
rect 104310 91160 104315 91216
rect 101876 91156 101882 91158
rect 100569 91155 100635 91156
rect 102041 91155 102107 91158
rect 104198 91156 104204 91158
rect 104268 91156 104315 91160
rect 104566 91156 104572 91220
rect 104636 91218 104642 91220
rect 104801 91218 104867 91221
rect 105537 91220 105603 91221
rect 105486 91218 105492 91220
rect 104636 91216 104867 91218
rect 104636 91160 104806 91216
rect 104862 91160 104867 91216
rect 104636 91158 104867 91160
rect 105446 91158 105492 91218
rect 105556 91216 105603 91220
rect 105598 91160 105603 91216
rect 104636 91156 104642 91158
rect 104249 91155 104315 91156
rect 104801 91155 104867 91158
rect 105486 91156 105492 91158
rect 105556 91156 105603 91160
rect 105670 91156 105676 91220
rect 105740 91218 105746 91220
rect 106181 91218 106247 91221
rect 105740 91216 106247 91218
rect 105740 91160 106186 91216
rect 106242 91160 106247 91216
rect 105740 91158 106247 91160
rect 105740 91156 105746 91158
rect 105537 91155 105603 91156
rect 106181 91155 106247 91158
rect 106406 91156 106412 91220
rect 106476 91218 106482 91220
rect 107469 91218 107535 91221
rect 106476 91216 107535 91218
rect 106476 91160 107474 91216
rect 107530 91160 107535 91216
rect 106476 91158 107535 91160
rect 106476 91156 106482 91158
rect 107469 91155 107535 91158
rect 107694 91156 107700 91220
rect 107764 91218 107770 91220
rect 108481 91218 108547 91221
rect 107764 91216 108547 91218
rect 107764 91160 108486 91216
rect 108542 91160 108547 91216
rect 107764 91158 108547 91160
rect 107764 91156 107770 91158
rect 108481 91155 108547 91158
rect 109534 91156 109540 91220
rect 109604 91218 109610 91220
rect 110321 91218 110387 91221
rect 109604 91216 110387 91218
rect 109604 91160 110326 91216
rect 110382 91160 110387 91216
rect 109604 91158 110387 91160
rect 109604 91156 109610 91158
rect 110321 91155 110387 91158
rect 111190 91156 111196 91220
rect 111260 91218 111266 91220
rect 111609 91218 111675 91221
rect 111260 91216 111675 91218
rect 111260 91160 111614 91216
rect 111670 91160 111675 91216
rect 111260 91158 111675 91160
rect 111260 91156 111266 91158
rect 111609 91155 111675 91158
rect 111926 91156 111932 91220
rect 111996 91156 112002 91220
rect 112294 91156 112300 91220
rect 112364 91218 112370 91220
rect 112989 91218 113055 91221
rect 112364 91216 113055 91218
rect 112364 91160 112994 91216
rect 113050 91160 113055 91216
rect 112364 91158 113055 91160
rect 112364 91156 112370 91158
rect 111934 91082 111994 91156
rect 112989 91155 113055 91158
rect 114318 91156 114324 91220
rect 114388 91218 114394 91220
rect 114461 91218 114527 91221
rect 114388 91216 114527 91218
rect 114388 91160 114466 91216
rect 114522 91160 114527 91216
rect 114388 91158 114527 91160
rect 114388 91156 114394 91158
rect 114461 91155 114527 91158
rect 114870 91156 114876 91220
rect 114940 91218 114946 91220
rect 115841 91218 115907 91221
rect 117129 91220 117195 91221
rect 117078 91218 117084 91220
rect 114940 91216 115907 91218
rect 114940 91160 115846 91216
rect 115902 91160 115907 91216
rect 114940 91158 115907 91160
rect 117038 91158 117084 91218
rect 117148 91216 117195 91220
rect 117190 91160 117195 91216
rect 114940 91156 114946 91158
rect 115841 91155 115907 91158
rect 117078 91156 117084 91158
rect 117148 91156 117195 91160
rect 117998 91156 118004 91220
rect 118068 91218 118074 91220
rect 118601 91218 118667 91221
rect 118068 91216 118667 91218
rect 118068 91160 118606 91216
rect 118662 91160 118667 91216
rect 118068 91158 118667 91160
rect 118068 91156 118074 91158
rect 117129 91155 117195 91156
rect 118601 91155 118667 91158
rect 119286 91156 119292 91220
rect 119356 91218 119362 91220
rect 119981 91218 120047 91221
rect 119356 91216 120047 91218
rect 119356 91160 119986 91216
rect 120042 91160 120047 91216
rect 119356 91158 120047 91160
rect 119356 91156 119362 91158
rect 119981 91155 120047 91158
rect 120206 91156 120212 91220
rect 120276 91218 120282 91220
rect 121361 91218 121427 91221
rect 120276 91216 121427 91218
rect 120276 91160 121366 91216
rect 121422 91160 121427 91216
rect 120276 91158 121427 91160
rect 120276 91156 120282 91158
rect 121361 91155 121427 91158
rect 121678 91156 121684 91220
rect 121748 91218 121754 91220
rect 121821 91218 121887 91221
rect 121748 91216 121887 91218
rect 121748 91160 121826 91216
rect 121882 91160 121887 91216
rect 121748 91158 121887 91160
rect 121748 91156 121754 91158
rect 121821 91155 121887 91158
rect 122046 91156 122052 91220
rect 122116 91218 122122 91220
rect 122741 91218 122807 91221
rect 122116 91216 122807 91218
rect 122116 91160 122746 91216
rect 122802 91160 122807 91216
rect 122116 91158 122807 91160
rect 122116 91156 122122 91158
rect 122741 91155 122807 91158
rect 123150 91156 123156 91220
rect 123220 91218 123226 91220
rect 124029 91218 124095 91221
rect 125409 91220 125475 91221
rect 125358 91218 125364 91220
rect 123220 91216 124095 91218
rect 123220 91160 124034 91216
rect 124090 91160 124095 91216
rect 123220 91158 124095 91160
rect 125318 91158 125364 91218
rect 125428 91216 125475 91220
rect 125470 91160 125475 91216
rect 123220 91156 123226 91158
rect 124029 91155 124095 91158
rect 125358 91156 125364 91158
rect 125428 91156 125475 91160
rect 126462 91156 126468 91220
rect 126532 91218 126538 91220
rect 126789 91218 126855 91221
rect 126532 91216 126855 91218
rect 126532 91160 126794 91216
rect 126850 91160 126855 91216
rect 126532 91158 126855 91160
rect 126532 91156 126538 91158
rect 125409 91155 125475 91156
rect 126789 91155 126855 91158
rect 127566 91156 127572 91220
rect 127636 91218 127642 91220
rect 128261 91218 128327 91221
rect 127636 91216 128327 91218
rect 127636 91160 128266 91216
rect 128322 91160 128327 91216
rect 127636 91158 128327 91160
rect 127636 91156 127642 91158
rect 128261 91155 128327 91158
rect 129406 91156 129412 91220
rect 129476 91218 129482 91220
rect 129641 91218 129707 91221
rect 132401 91220 132467 91221
rect 151721 91220 151787 91221
rect 132350 91218 132356 91220
rect 129476 91216 129707 91218
rect 129476 91160 129646 91216
rect 129702 91160 129707 91216
rect 129476 91158 129707 91160
rect 132310 91158 132356 91218
rect 132420 91216 132467 91220
rect 151670 91218 151676 91220
rect 132462 91160 132467 91216
rect 129476 91156 129482 91158
rect 129641 91155 129707 91158
rect 132350 91156 132356 91158
rect 132420 91156 132467 91160
rect 151630 91158 151676 91218
rect 151740 91216 151787 91220
rect 151782 91160 151787 91216
rect 151670 91156 151676 91158
rect 151740 91156 151787 91160
rect 152038 91156 152044 91220
rect 152108 91218 152114 91220
rect 152457 91218 152523 91221
rect 152108 91216 152523 91218
rect 152108 91160 152462 91216
rect 152518 91160 152523 91216
rect 152108 91158 152523 91160
rect 152108 91156 152114 91158
rect 132401 91155 132467 91156
rect 151721 91155 151787 91156
rect 152457 91155 152523 91158
rect 182909 91082 182975 91085
rect 111934 91080 182975 91082
rect 111934 91024 182914 91080
rect 182970 91024 182975 91080
rect 111934 91022 182975 91024
rect 182909 91019 182975 91022
rect 224718 91020 224724 91084
rect 224788 91082 224794 91084
rect 281625 91082 281691 91085
rect 224788 91080 281691 91082
rect 224788 91024 281630 91080
rect 281686 91024 281691 91080
rect 224788 91022 281691 91024
rect 224788 91020 224794 91022
rect 281625 91019 281691 91022
rect 153193 90946 153259 90949
rect 162853 90946 162919 90949
rect 153193 90944 162919 90946
rect 153193 90888 153198 90944
rect 153254 90888 162858 90944
rect 162914 90888 162919 90944
rect 153193 90886 162919 90888
rect 153193 90883 153259 90886
rect 162853 90883 162919 90886
rect 177389 90538 177455 90541
rect 211889 90538 211955 90541
rect 177389 90536 211955 90538
rect 177389 90480 177394 90536
rect 177450 90480 211894 90536
rect 211950 90480 211955 90536
rect 177389 90478 211955 90480
rect 177389 90475 177455 90478
rect 211889 90475 211955 90478
rect 88057 90402 88123 90405
rect 161933 90402 161999 90405
rect 88057 90400 161999 90402
rect 88057 90344 88062 90400
rect 88118 90344 161938 90400
rect 161994 90344 161999 90400
rect 88057 90342 161999 90344
rect 88057 90339 88123 90342
rect 161933 90339 161999 90342
rect 202229 90402 202295 90405
rect 281625 90402 281691 90405
rect 420678 90402 420684 90404
rect 202229 90400 420684 90402
rect 202229 90344 202234 90400
rect 202290 90344 281630 90400
rect 281686 90344 420684 90400
rect 202229 90342 420684 90344
rect 202229 90339 202295 90342
rect 281625 90339 281691 90342
rect 420678 90340 420684 90342
rect 420748 90340 420754 90404
rect 110137 89722 110203 89725
rect 200941 89722 201007 89725
rect 110137 89720 201007 89722
rect 110137 89664 110142 89720
rect 110198 89664 200946 89720
rect 201002 89664 201007 89720
rect 110137 89662 201007 89664
rect 110137 89659 110203 89662
rect 200941 89659 201007 89662
rect 91645 89586 91711 89589
rect 167821 89586 167887 89589
rect 91645 89584 167887 89586
rect 91645 89528 91650 89584
rect 91706 89528 167826 89584
rect 167882 89528 167887 89584
rect 91645 89526 167887 89528
rect 91645 89523 91711 89526
rect 167821 89523 167887 89526
rect 136449 89450 136515 89453
rect 162117 89450 162183 89453
rect 136449 89448 162183 89450
rect 136449 89392 136454 89448
rect 136510 89392 162122 89448
rect 162178 89392 162183 89448
rect 136449 89390 162183 89392
rect 136449 89387 136515 89390
rect 162117 89387 162183 89390
rect 169293 89178 169359 89181
rect 214557 89178 214623 89181
rect 169293 89176 214623 89178
rect 169293 89120 169298 89176
rect 169354 89120 214562 89176
rect 214618 89120 214623 89176
rect 169293 89118 214623 89120
rect 169293 89115 169359 89118
rect 214557 89115 214623 89118
rect 217317 89178 217383 89181
rect 245694 89178 245700 89180
rect 217317 89176 245700 89178
rect 217317 89120 217322 89176
rect 217378 89120 245700 89176
rect 217317 89118 245700 89120
rect 217317 89115 217383 89118
rect 245694 89116 245700 89118
rect 245764 89116 245770 89180
rect 186957 89042 187023 89045
rect 261845 89042 261911 89045
rect 186957 89040 261911 89042
rect 186957 88984 186962 89040
rect 187018 88984 261850 89040
rect 261906 88984 261911 89040
rect 186957 88982 261911 88984
rect 186957 88979 187023 88982
rect 261845 88979 261911 88982
rect 104249 88226 104315 88229
rect 181621 88226 181687 88229
rect 104249 88224 181687 88226
rect 104249 88168 104254 88224
rect 104310 88168 181626 88224
rect 181682 88168 181687 88224
rect 104249 88166 181687 88168
rect 104249 88163 104315 88166
rect 181621 88163 181687 88166
rect 393313 88226 393379 88229
rect 430665 88226 430731 88229
rect 393313 88224 430731 88226
rect 393313 88168 393318 88224
rect 393374 88168 430670 88224
rect 430726 88168 430731 88224
rect 393313 88166 430731 88168
rect 393313 88163 393379 88166
rect 430665 88163 430731 88166
rect 161933 88090 161999 88093
rect 211981 88090 212047 88093
rect 161933 88088 212047 88090
rect 161933 88032 161938 88088
rect 161994 88032 211986 88088
rect 212042 88032 212047 88088
rect 161933 88030 212047 88032
rect 161933 88027 161999 88030
rect 211981 88027 212047 88030
rect 115473 87954 115539 87957
rect 164969 87954 165035 87957
rect 115473 87952 165035 87954
rect 115473 87896 115478 87952
rect 115534 87896 164974 87952
rect 165030 87896 165035 87952
rect 115473 87894 165035 87896
rect 115473 87891 115539 87894
rect 164969 87891 165035 87894
rect 211797 87682 211863 87685
rect 250713 87682 250779 87685
rect 211797 87680 250779 87682
rect 211797 87624 211802 87680
rect 211858 87624 250718 87680
rect 250774 87624 250779 87680
rect 211797 87622 250779 87624
rect 211797 87619 211863 87622
rect 250713 87619 250779 87622
rect 177297 87546 177363 87549
rect 226425 87546 226491 87549
rect 177297 87544 226491 87546
rect 177297 87488 177302 87544
rect 177358 87488 226430 87544
rect 226486 87488 226491 87544
rect 177297 87486 226491 87488
rect 177297 87483 177363 87486
rect 226425 87483 226491 87486
rect 291694 86940 291700 87004
rect 291764 87002 291770 87004
rect 298093 87002 298159 87005
rect 291764 87000 298159 87002
rect 291764 86944 298098 87000
rect 298154 86944 298159 87000
rect 291764 86942 298159 86944
rect 291764 86940 291770 86942
rect 298093 86939 298159 86942
rect 89713 86866 89779 86869
rect 214833 86866 214899 86869
rect 89713 86864 214899 86866
rect 89713 86808 89718 86864
rect 89774 86808 214838 86864
rect 214894 86808 214899 86864
rect 89713 86806 214899 86808
rect 89713 86803 89779 86806
rect 214833 86803 214899 86806
rect 98729 86730 98795 86733
rect 166533 86730 166599 86733
rect 98729 86728 166599 86730
rect 98729 86672 98734 86728
rect 98790 86672 166538 86728
rect 166594 86672 166599 86728
rect 98729 86670 166599 86672
rect 98729 86667 98795 86670
rect 166533 86667 166599 86670
rect 133781 86594 133847 86597
rect 169201 86594 169267 86597
rect 133781 86592 169267 86594
rect 133781 86536 133786 86592
rect 133842 86536 169206 86592
rect 169262 86536 169267 86592
rect 133781 86534 169267 86536
rect 133781 86531 133847 86534
rect 169201 86531 169267 86534
rect 215886 86124 215892 86188
rect 215956 86186 215962 86188
rect 278037 86186 278103 86189
rect 215956 86184 278103 86186
rect 215956 86128 278042 86184
rect 278098 86128 278103 86184
rect 215956 86126 278103 86128
rect 215956 86124 215962 86126
rect 278037 86123 278103 86126
rect 582373 86186 582439 86189
rect 583520 86186 584960 86276
rect 582373 86184 584960 86186
rect 582373 86128 582378 86184
rect 582434 86128 584960 86184
rect 582373 86126 584960 86128
rect 582373 86123 582439 86126
rect 583520 86036 584960 86126
rect 89069 85506 89135 85509
rect 181713 85506 181779 85509
rect 89069 85504 181779 85506
rect 89069 85448 89074 85504
rect 89130 85448 181718 85504
rect 181774 85448 181779 85504
rect 89069 85446 181779 85448
rect 89069 85443 89135 85446
rect 181713 85443 181779 85446
rect 105537 85370 105603 85373
rect 198089 85370 198155 85373
rect 105537 85368 198155 85370
rect 105537 85312 105542 85368
rect 105598 85312 198094 85368
rect 198150 85312 198155 85368
rect 105537 85310 198155 85312
rect 105537 85307 105603 85310
rect 198089 85307 198155 85310
rect 100569 85234 100635 85237
rect 162025 85234 162091 85237
rect 100569 85232 162091 85234
rect 100569 85176 100574 85232
rect 100630 85176 162030 85232
rect 162086 85176 162091 85232
rect 100569 85174 162091 85176
rect 100569 85171 100635 85174
rect 162025 85171 162091 85174
rect 222929 84962 222995 84965
rect 236729 84962 236795 84965
rect 222929 84960 236795 84962
rect 222929 84904 222934 84960
rect 222990 84904 236734 84960
rect 236790 84904 236795 84960
rect 222929 84902 236795 84904
rect 222929 84899 222995 84902
rect 236729 84899 236795 84902
rect -960 84690 480 84780
rect 191046 84764 191052 84828
rect 191116 84826 191122 84828
rect 314009 84826 314075 84829
rect 191116 84824 314075 84826
rect 191116 84768 314014 84824
rect 314070 84768 314075 84824
rect 191116 84766 314075 84768
rect 191116 84764 191122 84766
rect 314009 84763 314075 84766
rect 3509 84690 3575 84693
rect -960 84688 3575 84690
rect -960 84632 3514 84688
rect 3570 84632 3575 84688
rect -960 84630 3575 84632
rect -960 84540 480 84630
rect 3509 84627 3575 84630
rect 86769 84146 86835 84149
rect 173433 84146 173499 84149
rect 86769 84144 173499 84146
rect 86769 84088 86774 84144
rect 86830 84088 173438 84144
rect 173494 84088 173499 84144
rect 86769 84086 173499 84088
rect 86769 84083 86835 84086
rect 173433 84083 173499 84086
rect 96521 84010 96587 84013
rect 180333 84010 180399 84013
rect 96521 84008 180399 84010
rect 96521 83952 96526 84008
rect 96582 83952 180338 84008
rect 180394 83952 180399 84008
rect 96521 83950 180399 83952
rect 96521 83947 96587 83950
rect 180333 83947 180399 83950
rect 220169 83466 220235 83469
rect 241145 83466 241211 83469
rect 220169 83464 241211 83466
rect 220169 83408 220174 83464
rect 220230 83408 241150 83464
rect 241206 83408 241211 83464
rect 220169 83406 241211 83408
rect 220169 83403 220235 83406
rect 241145 83403 241211 83406
rect 66161 82786 66227 82789
rect 177389 82786 177455 82789
rect 66161 82784 177455 82786
rect 66161 82728 66166 82784
rect 66222 82728 177394 82784
rect 177450 82728 177455 82784
rect 66161 82726 177455 82728
rect 66161 82723 66227 82726
rect 177389 82723 177455 82726
rect 231301 82786 231367 82789
rect 313917 82786 313983 82789
rect 231301 82784 313983 82786
rect 231301 82728 231306 82784
rect 231362 82728 313922 82784
rect 313978 82728 313983 82784
rect 231301 82726 313983 82728
rect 231301 82723 231367 82726
rect 313917 82723 313983 82726
rect 106181 82650 106247 82653
rect 185669 82650 185735 82653
rect 106181 82648 185735 82650
rect 106181 82592 106186 82648
rect 106242 82592 185674 82648
rect 185730 82592 185735 82648
rect 106181 82590 185735 82592
rect 106181 82587 106247 82590
rect 185669 82587 185735 82590
rect 106181 82106 106247 82109
rect 235441 82106 235507 82109
rect 106181 82104 235507 82106
rect 106181 82048 106186 82104
rect 106242 82048 235446 82104
rect 235502 82048 235507 82104
rect 106181 82046 235507 82048
rect 106181 82043 106247 82046
rect 235441 82043 235507 82046
rect 64781 81426 64847 81429
rect 192569 81426 192635 81429
rect 64781 81424 192635 81426
rect 64781 81368 64786 81424
rect 64842 81368 192574 81424
rect 192630 81368 192635 81424
rect 64781 81366 192635 81368
rect 64781 81363 64847 81366
rect 192569 81363 192635 81366
rect 113081 80882 113147 80885
rect 244774 80882 244780 80884
rect 113081 80880 244780 80882
rect 113081 80824 113086 80880
rect 113142 80824 244780 80880
rect 113081 80822 244780 80824
rect 113081 80819 113147 80822
rect 244774 80820 244780 80822
rect 244844 80820 244850 80884
rect 12341 80746 12407 80749
rect 264094 80746 264100 80748
rect 12341 80744 264100 80746
rect 12341 80688 12346 80744
rect 12402 80688 264100 80744
rect 12341 80686 264100 80688
rect 12341 80683 12407 80686
rect 264094 80684 264100 80686
rect 264164 80684 264170 80748
rect 97809 80066 97875 80069
rect 199469 80066 199535 80069
rect 97809 80064 199535 80066
rect 97809 80008 97814 80064
rect 97870 80008 199474 80064
rect 199530 80008 199535 80064
rect 97809 80006 199535 80008
rect 97809 80003 97875 80006
rect 199469 80003 199535 80006
rect 228357 79658 228423 79661
rect 237966 79658 237972 79660
rect 228357 79656 237972 79658
rect 228357 79600 228362 79656
rect 228418 79600 237972 79656
rect 228357 79598 237972 79600
rect 228357 79595 228423 79598
rect 237966 79596 237972 79598
rect 238036 79596 238042 79660
rect 5441 79522 5507 79525
rect 228541 79522 228607 79525
rect 5441 79520 228607 79522
rect 5441 79464 5446 79520
rect 5502 79464 228546 79520
rect 228602 79464 228607 79520
rect 5441 79462 228607 79464
rect 5441 79459 5507 79462
rect 228541 79459 228607 79462
rect 36537 79386 36603 79389
rect 265801 79386 265867 79389
rect 36537 79384 265867 79386
rect 36537 79328 36542 79384
rect 36598 79328 265806 79384
rect 265862 79328 265867 79384
rect 36537 79326 265867 79328
rect 36537 79323 36603 79326
rect 265801 79323 265867 79326
rect 107561 78026 107627 78029
rect 229870 78026 229876 78028
rect 107561 78024 229876 78026
rect 107561 77968 107566 78024
rect 107622 77968 229876 78024
rect 107561 77966 229876 77968
rect 107561 77963 107627 77966
rect 229870 77964 229876 77966
rect 229940 77964 229946 78028
rect 17861 77890 17927 77893
rect 257521 77890 257587 77893
rect 17861 77888 257587 77890
rect 17861 77832 17866 77888
rect 17922 77832 257526 77888
rect 257582 77832 257587 77888
rect 17861 77830 257587 77832
rect 17861 77827 17927 77830
rect 257521 77827 257587 77830
rect 62021 77210 62087 77213
rect 198181 77210 198247 77213
rect 62021 77208 198247 77210
rect 62021 77152 62026 77208
rect 62082 77152 198186 77208
rect 198242 77152 198247 77208
rect 62021 77150 198247 77152
rect 62021 77147 62087 77150
rect 198181 77147 198247 77150
rect 117221 76666 117287 76669
rect 236637 76666 236703 76669
rect 117221 76664 236703 76666
rect 117221 76608 117226 76664
rect 117282 76608 236642 76664
rect 236698 76608 236703 76664
rect 117221 76606 236703 76608
rect 117221 76603 117287 76606
rect 236637 76603 236703 76606
rect 86861 76530 86927 76533
rect 246573 76530 246639 76533
rect 86861 76528 246639 76530
rect 86861 76472 86866 76528
rect 86922 76472 246578 76528
rect 246634 76472 246639 76528
rect 86861 76470 246639 76472
rect 86861 76467 86927 76470
rect 246573 76467 246639 76470
rect 87597 75306 87663 75309
rect 242341 75306 242407 75309
rect 87597 75304 242407 75306
rect 87597 75248 87602 75304
rect 87658 75248 242346 75304
rect 242402 75248 242407 75304
rect 87597 75246 242407 75248
rect 87597 75243 87663 75246
rect 242341 75243 242407 75246
rect 19149 75170 19215 75173
rect 253473 75170 253539 75173
rect 19149 75168 253539 75170
rect 19149 75112 19154 75168
rect 19210 75112 253478 75168
rect 253534 75112 253539 75168
rect 19149 75110 253539 75112
rect 19149 75107 19215 75110
rect 253473 75107 253539 75110
rect 115289 74490 115355 74493
rect 169017 74490 169083 74493
rect 115289 74488 169083 74490
rect 115289 74432 115294 74488
rect 115350 74432 169022 74488
rect 169078 74432 169083 74488
rect 115289 74430 169083 74432
rect 115289 74427 115355 74430
rect 169017 74427 169083 74430
rect 35801 73810 35867 73813
rect 258901 73810 258967 73813
rect 35801 73808 258967 73810
rect 35801 73752 35806 73808
rect 35862 73752 258906 73808
rect 258962 73752 258967 73808
rect 35801 73750 258967 73752
rect 35801 73747 35867 73750
rect 258901 73747 258967 73750
rect 319437 73810 319503 73813
rect 421046 73810 421052 73812
rect 319437 73808 421052 73810
rect 319437 73752 319442 73808
rect 319498 73752 421052 73808
rect 319437 73750 421052 73752
rect 319437 73747 319503 73750
rect 421046 73748 421052 73750
rect 421116 73748 421122 73812
rect 582373 72994 582439 72997
rect 583520 72994 584960 73084
rect 582373 72992 584960 72994
rect 582373 72936 582378 72992
rect 582434 72936 584960 72992
rect 582373 72934 584960 72936
rect 582373 72931 582439 72934
rect 583520 72844 584960 72934
rect 22001 72586 22067 72589
rect 267181 72586 267247 72589
rect 22001 72584 267247 72586
rect 22001 72528 22006 72584
rect 22062 72528 267186 72584
rect 267242 72528 267247 72584
rect 22001 72526 267247 72528
rect 22001 72523 22067 72526
rect 267181 72523 267247 72526
rect 50981 72450 51047 72453
rect 297357 72450 297423 72453
rect 50981 72448 297423 72450
rect 50981 72392 50986 72448
rect 51042 72392 297362 72448
rect 297418 72392 297423 72448
rect 50981 72390 297423 72392
rect 50981 72387 51047 72390
rect 297357 72387 297423 72390
rect 32397 71770 32463 71773
rect 443085 71770 443151 71773
rect 6870 71768 443151 71770
rect -960 71634 480 71724
rect 6870 71712 32402 71768
rect 32458 71712 443090 71768
rect 443146 71712 443151 71768
rect 6870 71710 443151 71712
rect 6870 71634 6930 71710
rect 32397 71707 32463 71710
rect 443085 71707 443151 71710
rect -960 71574 6930 71634
rect -960 71484 480 71574
rect 50981 71090 51047 71093
rect 258574 71090 258580 71092
rect 50981 71088 258580 71090
rect 50981 71032 50986 71088
rect 51042 71032 258580 71088
rect 50981 71030 258580 71032
rect 50981 71027 51047 71030
rect 258574 71028 258580 71030
rect 258644 71028 258650 71092
rect 93761 69730 93827 69733
rect 260189 69730 260255 69733
rect 93761 69728 260255 69730
rect 93761 69672 93766 69728
rect 93822 69672 260194 69728
rect 260250 69672 260255 69728
rect 93761 69670 260255 69672
rect 93761 69667 93827 69670
rect 260189 69667 260255 69670
rect 15101 69594 15167 69597
rect 261569 69594 261635 69597
rect 15101 69592 261635 69594
rect 15101 69536 15106 69592
rect 15162 69536 261574 69592
rect 261630 69536 261635 69592
rect 15101 69534 261635 69536
rect 15101 69531 15167 69534
rect 261569 69531 261635 69534
rect 125501 68370 125567 68373
rect 254577 68370 254643 68373
rect 125501 68368 254643 68370
rect 125501 68312 125506 68368
rect 125562 68312 254582 68368
rect 254638 68312 254643 68368
rect 125501 68310 254643 68312
rect 125501 68307 125567 68310
rect 254577 68307 254643 68310
rect 95141 68234 95207 68237
rect 267089 68234 267155 68237
rect 95141 68232 267155 68234
rect 95141 68176 95146 68232
rect 95202 68176 267094 68232
rect 267150 68176 267155 68232
rect 95141 68174 267155 68176
rect 95141 68171 95207 68174
rect 267089 68171 267155 68174
rect 116577 67554 116643 67557
rect 168230 67554 168236 67556
rect 116577 67552 168236 67554
rect 116577 67496 116582 67552
rect 116638 67496 168236 67552
rect 116577 67494 168236 67496
rect 116577 67491 116643 67494
rect 168230 67492 168236 67494
rect 168300 67492 168306 67556
rect 122097 66874 122163 66877
rect 265709 66874 265775 66877
rect 122097 66872 265775 66874
rect 122097 66816 122102 66872
rect 122158 66816 265714 66872
rect 265770 66816 265775 66872
rect 122097 66814 265775 66816
rect 122097 66811 122163 66814
rect 265709 66811 265775 66814
rect 64781 65650 64847 65653
rect 255957 65650 256023 65653
rect 64781 65648 256023 65650
rect 64781 65592 64786 65648
rect 64842 65592 255962 65648
rect 256018 65592 256023 65648
rect 64781 65590 256023 65592
rect 64781 65587 64847 65590
rect 255957 65587 256023 65590
rect 48221 65514 48287 65517
rect 249149 65514 249215 65517
rect 48221 65512 249215 65514
rect 48221 65456 48226 65512
rect 48282 65456 249154 65512
rect 249210 65456 249215 65512
rect 48221 65454 249215 65456
rect 48221 65451 48287 65454
rect 249149 65451 249215 65454
rect 352557 65514 352623 65517
rect 431718 65514 431724 65516
rect 352557 65512 431724 65514
rect 352557 65456 352562 65512
rect 352618 65456 431724 65512
rect 352557 65454 431724 65456
rect 352557 65451 352623 65454
rect 431718 65452 431724 65454
rect 431788 65452 431794 65516
rect 77201 64290 77267 64293
rect 246481 64290 246547 64293
rect 77201 64288 246547 64290
rect 77201 64232 77206 64288
rect 77262 64232 246486 64288
rect 246542 64232 246547 64288
rect 77201 64230 246547 64232
rect 77201 64227 77267 64230
rect 246481 64227 246547 64230
rect 42701 64154 42767 64157
rect 257429 64154 257495 64157
rect 42701 64152 257495 64154
rect 42701 64096 42706 64152
rect 42762 64096 257434 64152
rect 257490 64096 257495 64152
rect 42701 64094 257495 64096
rect 42701 64091 42767 64094
rect 257429 64091 257495 64094
rect 287646 64092 287652 64156
rect 287716 64154 287722 64156
rect 302877 64154 302943 64157
rect 287716 64152 302943 64154
rect 287716 64096 302882 64152
rect 302938 64096 302943 64152
rect 287716 64094 302943 64096
rect 287716 64092 287722 64094
rect 302877 64091 302943 64094
rect 79961 62794 80027 62797
rect 267958 62794 267964 62796
rect 79961 62792 267964 62794
rect 79961 62736 79966 62792
rect 80022 62736 267964 62792
rect 79961 62734 267964 62736
rect 79961 62731 80027 62734
rect 267958 62732 267964 62734
rect 268028 62732 268034 62796
rect 273989 62794 274055 62797
rect 288566 62794 288572 62796
rect 273989 62792 288572 62794
rect 273989 62736 273994 62792
rect 274050 62736 288572 62792
rect 273989 62734 288572 62736
rect 273989 62731 274055 62734
rect 288566 62732 288572 62734
rect 288636 62732 288642 62796
rect 75821 61434 75887 61437
rect 249006 61434 249012 61436
rect 75821 61432 249012 61434
rect 75821 61376 75826 61432
rect 75882 61376 249012 61432
rect 75821 61374 249012 61376
rect 75821 61371 75887 61374
rect 249006 61372 249012 61374
rect 249076 61372 249082 61436
rect 288341 60484 288407 60485
rect 288341 60480 288388 60484
rect 288452 60482 288458 60484
rect 288341 60424 288346 60480
rect 288341 60420 288388 60424
rect 288452 60422 288498 60482
rect 288452 60420 288458 60422
rect 288341 60419 288407 60420
rect 82721 59938 82787 59941
rect 262806 59938 262812 59940
rect 82721 59936 262812 59938
rect 82721 59880 82726 59936
rect 82782 59880 262812 59936
rect 82721 59878 262812 59880
rect 82721 59875 82787 59878
rect 262806 59876 262812 59878
rect 262876 59876 262882 59940
rect 582649 59666 582715 59669
rect 583520 59666 584960 59756
rect 582649 59664 584960 59666
rect 582649 59608 582654 59664
rect 582710 59608 584960 59664
rect 582649 59606 584960 59608
rect 582649 59603 582715 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 3049 58578 3115 58581
rect -960 58576 3115 58578
rect -960 58520 3054 58576
rect 3110 58520 3115 58576
rect -960 58518 3115 58520
rect -960 58428 480 58518
rect 3049 58515 3115 58518
rect 78581 58578 78647 58581
rect 266997 58578 267063 58581
rect 78581 58576 267063 58578
rect 78581 58520 78586 58576
rect 78642 58520 267002 58576
rect 267058 58520 267063 58576
rect 78581 58518 267063 58520
rect 78581 58515 78647 58518
rect 266997 58515 267063 58518
rect 57881 57218 57947 57221
rect 247677 57218 247743 57221
rect 57881 57216 247743 57218
rect 57881 57160 57886 57216
rect 57942 57160 247682 57216
rect 247738 57160 247743 57216
rect 57881 57158 247743 57160
rect 57881 57155 57947 57158
rect 247677 57155 247743 57158
rect 262949 57218 263015 57221
rect 409822 57218 409828 57220
rect 262949 57216 409828 57218
rect 262949 57160 262954 57216
rect 263010 57160 409828 57216
rect 262949 57158 409828 57160
rect 262949 57155 263015 57158
rect 409822 57156 409828 57158
rect 409892 57156 409898 57220
rect 10961 55858 11027 55861
rect 260046 55858 260052 55860
rect 10961 55856 260052 55858
rect 10961 55800 10966 55856
rect 11022 55800 260052 55856
rect 10961 55798 260052 55800
rect 10961 55795 11027 55798
rect 260046 55796 260052 55798
rect 260116 55796 260122 55860
rect 206277 55178 206343 55181
rect 260373 55178 260439 55181
rect 206277 55176 260439 55178
rect 206277 55120 206282 55176
rect 206338 55120 260378 55176
rect 260434 55120 260439 55176
rect 206277 55118 260439 55120
rect 206277 55115 206343 55118
rect 260373 55115 260439 55118
rect 23381 54498 23447 54501
rect 233734 54498 233740 54500
rect 23381 54496 233740 54498
rect 23381 54440 23386 54496
rect 23442 54440 233740 54496
rect 23381 54438 233740 54440
rect 23381 54435 23447 54438
rect 233734 54436 233740 54438
rect 233804 54436 233810 54500
rect 259453 53954 259519 53957
rect 260373 53954 260439 53957
rect 259453 53952 260439 53954
rect 259453 53896 259458 53952
rect 259514 53896 260378 53952
rect 260434 53896 260439 53952
rect 259453 53894 260439 53896
rect 259453 53891 259519 53894
rect 260373 53891 260439 53894
rect 58617 53138 58683 53141
rect 221457 53138 221523 53141
rect 58617 53136 221523 53138
rect 58617 53080 58622 53136
rect 58678 53080 221462 53136
rect 221518 53080 221523 53136
rect 58617 53078 221523 53080
rect 58617 53075 58683 53078
rect 221457 53075 221523 53078
rect 252502 53076 252508 53140
rect 252572 53138 252578 53140
rect 429142 53138 429148 53140
rect 252572 53078 429148 53138
rect 252572 53076 252578 53078
rect 429142 53076 429148 53078
rect 429212 53076 429218 53140
rect 53741 51778 53807 51781
rect 251817 51778 251883 51781
rect 53741 51776 251883 51778
rect 53741 51720 53746 51776
rect 53802 51720 251822 51776
rect 251878 51720 251883 51776
rect 53741 51718 251883 51720
rect 53741 51715 53807 51718
rect 251817 51715 251883 51718
rect 249793 50964 249859 50965
rect 249742 50962 249748 50964
rect 249702 50902 249748 50962
rect 249812 50960 249859 50964
rect 249854 50904 249859 50960
rect 249742 50900 249748 50902
rect 249812 50900 249859 50904
rect 249793 50899 249859 50900
rect 28901 50282 28967 50285
rect 254669 50282 254735 50285
rect 28901 50280 254735 50282
rect 28901 50224 28906 50280
rect 28962 50224 254674 50280
rect 254730 50224 254735 50280
rect 28901 50222 254735 50224
rect 28901 50219 28967 50222
rect 254669 50219 254735 50222
rect 27521 48922 27587 48925
rect 247769 48922 247835 48925
rect 27521 48920 247835 48922
rect 27521 48864 27526 48920
rect 27582 48864 247774 48920
rect 247830 48864 247835 48920
rect 27521 48862 247835 48864
rect 27521 48859 27587 48862
rect 247769 48859 247835 48862
rect 582925 46338 582991 46341
rect 583520 46338 584960 46428
rect 582925 46336 584960 46338
rect 582925 46280 582930 46336
rect 582986 46280 584960 46336
rect 582925 46278 584960 46280
rect 582925 46275 582991 46278
rect 53649 46202 53715 46205
rect 249149 46202 249215 46205
rect 53649 46200 249215 46202
rect 53649 46144 53654 46200
rect 53710 46144 249154 46200
rect 249210 46144 249215 46200
rect 583520 46188 584960 46278
rect 53649 46142 249215 46144
rect 53649 46139 53715 46142
rect 249149 46139 249215 46142
rect -960 45522 480 45612
rect -960 45462 674 45522
rect -960 45372 480 45462
rect 614 45250 674 45462
rect 430 45190 674 45250
rect 430 44842 490 45190
rect 141417 44842 141483 44845
rect 180149 44842 180215 44845
rect 430 44782 6930 44842
rect 6870 44298 6930 44782
rect 141417 44840 180215 44842
rect 141417 44784 141422 44840
rect 141478 44784 180154 44840
rect 180210 44784 180215 44840
rect 141417 44782 180215 44784
rect 141417 44779 141483 44782
rect 180149 44779 180215 44782
rect 188429 44842 188495 44845
rect 296069 44842 296135 44845
rect 188429 44840 296135 44842
rect 188429 44784 188434 44840
rect 188490 44784 296074 44840
rect 296130 44784 296135 44840
rect 188429 44782 296135 44784
rect 188429 44779 188495 44782
rect 296069 44779 296135 44782
rect 47577 44298 47643 44301
rect 6870 44296 47643 44298
rect 6870 44240 47582 44296
rect 47638 44240 47643 44296
rect 6870 44238 47643 44240
rect 47577 44235 47643 44238
rect 37181 42122 37247 42125
rect 232446 42122 232452 42124
rect 37181 42120 232452 42122
rect 37181 42064 37186 42120
rect 37242 42064 232452 42120
rect 37181 42062 232452 42064
rect 37181 42059 37247 42062
rect 232446 42060 232452 42062
rect 232516 42060 232522 42124
rect 144821 39266 144887 39269
rect 399477 39266 399543 39269
rect 144821 39264 399543 39266
rect 144821 39208 144826 39264
rect 144882 39208 399482 39264
rect 399538 39208 399543 39264
rect 144821 39206 399543 39208
rect 144821 39203 144887 39206
rect 399477 39203 399543 39206
rect 6821 38042 6887 38045
rect 226374 38042 226380 38044
rect 6821 38040 226380 38042
rect 6821 37984 6826 38040
rect 6882 37984 226380 38040
rect 6821 37982 226380 37984
rect 6821 37979 6887 37982
rect 226374 37980 226380 37982
rect 226444 37980 226450 38044
rect 66110 37844 66116 37908
rect 66180 37906 66186 37908
rect 325049 37906 325115 37909
rect 66180 37904 325115 37906
rect 66180 37848 325054 37904
rect 325110 37848 325115 37904
rect 66180 37846 325115 37848
rect 66180 37844 66186 37846
rect 325049 37843 325115 37846
rect 54477 36546 54543 36549
rect 267774 36546 267780 36548
rect 54477 36544 267780 36546
rect 54477 36488 54482 36544
rect 54538 36488 267780 36544
rect 54477 36486 267780 36488
rect 54477 36483 54543 36486
rect 267774 36484 267780 36486
rect 267844 36484 267850 36548
rect 46841 35186 46907 35189
rect 177297 35186 177363 35189
rect 46841 35184 177363 35186
rect 46841 35128 46846 35184
rect 46902 35128 177302 35184
rect 177358 35128 177363 35184
rect 46841 35126 177363 35128
rect 46841 35123 46907 35126
rect 177297 35123 177363 35126
rect 186814 35124 186820 35188
rect 186884 35186 186890 35188
rect 302969 35186 303035 35189
rect 186884 35184 303035 35186
rect 186884 35128 302974 35184
rect 303030 35128 303035 35184
rect 186884 35126 303035 35128
rect 186884 35124 186890 35126
rect 302969 35123 303035 35126
rect 302969 34642 303035 34645
rect 304257 34642 304323 34645
rect 302969 34640 304323 34642
rect 302969 34584 302974 34640
rect 303030 34584 304262 34640
rect 304318 34584 304323 34640
rect 302969 34582 304323 34584
rect 302969 34579 303035 34582
rect 304257 34579 304323 34582
rect 61878 33764 61884 33828
rect 61948 33826 61954 33828
rect 251817 33826 251883 33829
rect 61948 33824 251883 33826
rect 61948 33768 251822 33824
rect 251878 33768 251883 33824
rect 61948 33766 251883 33768
rect 61948 33764 61954 33766
rect 251817 33763 251883 33766
rect 300117 33826 300183 33829
rect 417366 33826 417372 33828
rect 300117 33824 417372 33826
rect 300117 33768 300122 33824
rect 300178 33768 417372 33824
rect 300117 33766 417372 33768
rect 300117 33763 300183 33766
rect 417366 33764 417372 33766
rect 417436 33764 417442 33828
rect 295333 33146 295399 33149
rect 296069 33146 296135 33149
rect 426382 33146 426388 33148
rect 295333 33144 426388 33146
rect 295333 33088 295338 33144
rect 295394 33088 296074 33144
rect 296130 33088 426388 33144
rect 295333 33086 426388 33088
rect 295333 33083 295399 33086
rect 296069 33083 296135 33086
rect 426382 33084 426388 33086
rect 426452 33084 426458 33148
rect 582741 33146 582807 33149
rect 583520 33146 584960 33236
rect 582741 33144 584960 33146
rect 582741 33088 582746 33144
rect 582802 33088 584960 33144
rect 582741 33086 584960 33088
rect 582741 33083 582807 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 2865 32466 2931 32469
rect -960 32464 2931 32466
rect -960 32408 2870 32464
rect 2926 32408 2931 32464
rect -960 32406 2931 32408
rect -960 32316 480 32406
rect 2865 32403 2931 32406
rect 176561 30290 176627 30293
rect 273253 30290 273319 30293
rect 273897 30290 273963 30293
rect 176561 30288 273963 30290
rect 176561 30232 176566 30288
rect 176622 30232 273258 30288
rect 273314 30232 273902 30288
rect 273958 30232 273963 30288
rect 176561 30230 273963 30232
rect 176561 30227 176627 30230
rect 273253 30227 273319 30230
rect 273897 30227 273963 30230
rect 169518 26828 169524 26892
rect 169588 26890 169594 26892
rect 242893 26890 242959 26893
rect 169588 26888 242959 26890
rect 169588 26832 242898 26888
rect 242954 26832 242959 26888
rect 169588 26830 242959 26832
rect 169588 26828 169594 26830
rect 242893 26827 242959 26830
rect 67766 25604 67772 25668
rect 67836 25666 67842 25668
rect 255957 25666 256023 25669
rect 67836 25664 256023 25666
rect 67836 25608 255962 25664
rect 256018 25608 256023 25664
rect 67836 25606 256023 25608
rect 67836 25604 67842 25606
rect 255957 25603 256023 25606
rect 20621 25530 20687 25533
rect 244038 25530 244044 25532
rect 20621 25528 244044 25530
rect 20621 25472 20626 25528
rect 20682 25472 244044 25528
rect 20621 25470 244044 25472
rect 20621 25467 20687 25470
rect 244038 25468 244044 25470
rect 244108 25468 244114 25532
rect 103421 24170 103487 24173
rect 236494 24170 236500 24172
rect 103421 24168 236500 24170
rect 103421 24112 103426 24168
rect 103482 24112 236500 24168
rect 103421 24110 236500 24112
rect 103421 24107 103487 24110
rect 236494 24108 236500 24110
rect 236564 24108 236570 24172
rect 254577 24170 254643 24173
rect 435030 24170 435036 24172
rect 254577 24168 435036 24170
rect 254577 24112 254582 24168
rect 254638 24112 435036 24168
rect 254577 24110 435036 24112
rect 254577 24107 254643 24110
rect 435030 24108 435036 24110
rect 435100 24108 435106 24172
rect 302877 23354 302943 23357
rect 303521 23354 303587 23357
rect 419022 23354 419028 23356
rect 302877 23352 419028 23354
rect 302877 23296 302882 23352
rect 302938 23296 303526 23352
rect 303582 23296 419028 23352
rect 302877 23294 419028 23296
rect 302877 23291 302943 23294
rect 303521 23291 303587 23294
rect 419022 23292 419028 23294
rect 419092 23292 419098 23356
rect 204897 22674 204963 22677
rect 277485 22674 277551 22677
rect 204897 22672 277551 22674
rect 204897 22616 204902 22672
rect 204958 22616 277490 22672
rect 277546 22616 277551 22672
rect 204897 22614 277551 22616
rect 204897 22611 204963 22614
rect 277485 22611 277551 22614
rect 4061 21314 4127 21317
rect 226926 21314 226932 21316
rect 4061 21312 226932 21314
rect 4061 21256 4066 21312
rect 4122 21256 226932 21312
rect 4061 21254 226932 21256
rect 4061 21251 4127 21254
rect 226926 21252 226932 21254
rect 226996 21252 227002 21316
rect 185577 20634 185643 20637
rect 284385 20634 284451 20637
rect 284937 20634 285003 20637
rect 185577 20632 285003 20634
rect 185577 20576 185582 20632
rect 185638 20576 284390 20632
rect 284446 20576 284942 20632
rect 284998 20576 285003 20632
rect 185577 20574 285003 20576
rect 185577 20571 185643 20574
rect 284385 20571 284451 20574
rect 284937 20571 285003 20574
rect 582557 19818 582623 19821
rect 583520 19818 584960 19908
rect 582557 19816 584960 19818
rect 582557 19760 582562 19816
rect 582618 19760 584960 19816
rect 582557 19758 584960 19760
rect 582557 19755 582623 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 3417 19410 3483 19413
rect -960 19408 3483 19410
rect -960 19352 3422 19408
rect 3478 19352 3483 19408
rect -960 19350 3483 19352
rect -960 19260 480 19350
rect 3417 19347 3483 19350
rect 175089 19274 175155 19277
rect 267733 19274 267799 19277
rect 268377 19274 268443 19277
rect 175089 19272 268443 19274
rect 175089 19216 175094 19272
rect 175150 19216 267738 19272
rect 267794 19216 268382 19272
rect 268438 19216 268443 19272
rect 175089 19214 268443 19216
rect 175089 19211 175155 19214
rect 267733 19211 267799 19214
rect 268377 19211 268443 19214
rect 98637 18594 98703 18597
rect 135253 18594 135319 18597
rect 98637 18592 135319 18594
rect 98637 18536 98642 18592
rect 98698 18536 135258 18592
rect 135314 18536 135319 18592
rect 98637 18534 135319 18536
rect 98637 18531 98703 18534
rect 135253 18531 135319 18534
rect 310513 17914 310579 17917
rect 427854 17914 427860 17916
rect 310513 17912 427860 17914
rect 310513 17856 310518 17912
rect 310574 17856 427860 17912
rect 310513 17854 427860 17856
rect 310513 17851 310579 17854
rect 427854 17852 427860 17854
rect 427924 17852 427930 17916
rect 57237 17234 57303 17237
rect 266854 17234 266860 17236
rect 57237 17232 266860 17234
rect 57237 17176 57242 17232
rect 57298 17176 266860 17232
rect 57237 17174 266860 17176
rect 57237 17171 57303 17174
rect 266854 17172 266860 17174
rect 266924 17172 266930 17236
rect 133137 15874 133203 15877
rect 172462 15874 172468 15876
rect 133137 15872 172468 15874
rect 133137 15816 133142 15872
rect 133198 15816 172468 15872
rect 133137 15814 172468 15816
rect 133137 15811 133203 15814
rect 172462 15812 172468 15814
rect 172532 15812 172538 15876
rect 177246 15812 177252 15876
rect 177316 15874 177322 15876
rect 253473 15874 253539 15877
rect 177316 15872 253539 15874
rect 177316 15816 253478 15872
rect 253534 15816 253539 15872
rect 177316 15814 253539 15816
rect 177316 15812 177322 15814
rect 253473 15811 253539 15814
rect 253473 15330 253539 15333
rect 254577 15330 254643 15333
rect 253473 15328 254643 15330
rect 253473 15272 253478 15328
rect 253534 15272 254582 15328
rect 254638 15272 254643 15328
rect 253473 15270 254643 15272
rect 253473 15267 253539 15270
rect 254577 15267 254643 15270
rect 59118 15132 59124 15196
rect 59188 15194 59194 15196
rect 250529 15194 250595 15197
rect 59188 15192 250595 15194
rect 59188 15136 250534 15192
rect 250590 15136 250595 15192
rect 59188 15134 250595 15136
rect 59188 15132 59194 15134
rect 250529 15131 250595 15134
rect 249977 13834 250043 13837
rect 250529 13834 250595 13837
rect 249977 13832 250595 13834
rect 249977 13776 249982 13832
rect 250038 13776 250534 13832
rect 250590 13776 250595 13832
rect 249977 13774 250595 13776
rect 249977 13771 250043 13774
rect 250529 13771 250595 13774
rect 295885 13700 295951 13701
rect 295885 13696 295932 13700
rect 295996 13698 296002 13700
rect 295885 13640 295890 13696
rect 295885 13636 295932 13640
rect 295996 13638 296042 13698
rect 295996 13636 296002 13638
rect 295885 13635 295951 13636
rect 299657 13156 299723 13157
rect 299606 13092 299612 13156
rect 299676 13154 299723 13156
rect 299676 13152 299768 13154
rect 299718 13096 299768 13152
rect 299676 13094 299768 13096
rect 299676 13092 299723 13094
rect 299657 13091 299723 13092
rect 252318 11732 252324 11796
rect 252388 11794 252394 11796
rect 253197 11794 253263 11797
rect 252388 11792 253263 11794
rect 252388 11736 253202 11792
rect 253258 11736 253263 11792
rect 252388 11734 253263 11736
rect 252388 11732 252394 11734
rect 253197 11731 253263 11734
rect 182766 11596 182772 11660
rect 182836 11658 182842 11660
rect 261753 11658 261819 11661
rect 182836 11656 261819 11658
rect 182836 11600 261758 11656
rect 261814 11600 261819 11656
rect 182836 11598 261819 11600
rect 182836 11596 182842 11598
rect 261753 11595 261819 11598
rect 180057 10298 180123 10301
rect 260097 10298 260163 10301
rect 180057 10296 260163 10298
rect 180057 10240 180062 10296
rect 180118 10240 260102 10296
rect 260158 10240 260163 10296
rect 180057 10238 260163 10240
rect 180057 10235 180123 10238
rect 260097 10235 260163 10238
rect 314009 9618 314075 9621
rect 439078 9618 439084 9620
rect 314009 9616 439084 9618
rect 314009 9560 314014 9616
rect 314070 9560 439084 9616
rect 314009 9558 439084 9560
rect 314009 9555 314075 9558
rect 439078 9556 439084 9558
rect 439148 9556 439154 9620
rect 297357 8258 297423 8261
rect 452653 8258 452719 8261
rect 297357 8256 452719 8258
rect 297357 8200 297362 8256
rect 297418 8200 452658 8256
rect 452714 8200 452719 8256
rect 297357 8198 452719 8200
rect 297357 8195 297423 8198
rect 452653 8195 452719 8198
rect 178718 7516 178724 7580
rect 178788 7578 178794 7580
rect 242893 7578 242959 7581
rect 178788 7576 242959 7578
rect 178788 7520 242898 7576
rect 242954 7520 242959 7576
rect 178788 7518 242959 7520
rect 178788 7516 178794 7518
rect 242893 7515 242959 7518
rect 13 6762 79 6765
rect 188337 6762 188403 6765
rect 289077 6762 289143 6765
rect 13 6760 122 6762
rect 13 6704 18 6760
rect 74 6704 122 6760
rect 13 6699 122 6704
rect 188337 6760 289143 6762
rect 188337 6704 188342 6760
rect 188398 6704 289082 6760
rect 289138 6704 289143 6760
rect 188337 6702 289143 6704
rect 188337 6699 188403 6702
rect 289077 6699 289143 6702
rect 62 6626 122 6699
rect 582465 6626 582531 6629
rect 583520 6626 584960 6716
rect 62 6580 674 6626
rect -960 6566 674 6580
rect -960 6490 480 6566
rect 614 6490 674 6566
rect 582465 6624 584960 6626
rect 582465 6568 582470 6624
rect 582526 6568 584960 6624
rect 582465 6566 584960 6568
rect 582465 6563 582531 6566
rect -960 6430 674 6490
rect 583520 6476 584960 6566
rect -960 6340 480 6430
rect 25313 6218 25379 6221
rect 186957 6218 187023 6221
rect 25313 6216 187023 6218
rect 25313 6160 25318 6216
rect 25374 6160 186962 6216
rect 187018 6160 187023 6216
rect 25313 6158 187023 6160
rect 25313 6155 25379 6158
rect 186957 6155 187023 6158
rect 287789 5674 287855 5677
rect 288341 5674 288407 5677
rect 287789 5672 288407 5674
rect 287789 5616 287794 5672
rect 287850 5616 288346 5672
rect 288402 5616 288407 5672
rect 287789 5614 288407 5616
rect 287789 5611 287855 5614
rect 288341 5611 288407 5614
rect 1669 4858 1735 4861
rect 227662 4858 227668 4860
rect 1669 4856 227668 4858
rect 1669 4800 1674 4856
rect 1730 4800 227668 4856
rect 1669 4798 227668 4800
rect 1669 4795 1735 4798
rect 227662 4796 227668 4798
rect 227732 4796 227738 4860
rect 195237 4042 195303 4045
rect 257061 4042 257127 4045
rect 257337 4042 257403 4045
rect 195237 4040 257403 4042
rect 195237 3984 195242 4040
rect 195298 3984 257066 4040
rect 257122 3984 257342 4040
rect 257398 3984 257403 4040
rect 195237 3982 257403 3984
rect 195237 3979 195303 3982
rect 257061 3979 257127 3982
rect 257337 3979 257403 3982
rect 326337 4042 326403 4045
rect 352557 4042 352623 4045
rect 326337 4040 352623 4042
rect 326337 3984 326342 4040
rect 326398 3984 352562 4040
rect 352618 3984 352623 4040
rect 326337 3982 352623 3984
rect 326337 3979 326403 3982
rect 352557 3979 352623 3982
rect 196617 3906 196683 3909
rect 246205 3906 246271 3909
rect 196617 3904 246271 3906
rect 196617 3848 196622 3904
rect 196678 3848 246210 3904
rect 246266 3848 246271 3904
rect 196617 3846 246271 3848
rect 196617 3843 196683 3846
rect 246205 3843 246271 3846
rect 295977 3906 296043 3909
rect 300117 3906 300183 3909
rect 295977 3904 300183 3906
rect 295977 3848 295982 3904
rect 296038 3848 300122 3904
rect 300178 3848 300183 3904
rect 295977 3846 300183 3848
rect 295977 3843 296043 3846
rect 300117 3843 300183 3846
rect 351637 3906 351703 3909
rect 376017 3906 376083 3909
rect 351637 3904 376083 3906
rect 351637 3848 351642 3904
rect 351698 3848 376022 3904
rect 376078 3848 376083 3904
rect 351637 3846 376083 3848
rect 351637 3843 351703 3846
rect 376017 3843 376083 3846
rect 322197 3770 322263 3773
rect 267690 3768 322263 3770
rect 267690 3712 322202 3768
rect 322258 3712 322263 3768
rect 267690 3710 322263 3712
rect 260097 3634 260163 3637
rect 260649 3634 260715 3637
rect 267690 3634 267750 3710
rect 322197 3707 322263 3710
rect 260097 3632 267750 3634
rect 260097 3576 260102 3632
rect 260158 3576 260654 3632
rect 260710 3576 267750 3632
rect 260097 3574 267750 3576
rect 260097 3571 260163 3574
rect 260649 3571 260715 3574
rect 132953 3498 133019 3501
rect 165654 3498 165660 3500
rect 132953 3496 165660 3498
rect 132953 3440 132958 3496
rect 133014 3440 165660 3496
rect 132953 3438 165660 3440
rect 132953 3435 133019 3438
rect 165654 3436 165660 3438
rect 165724 3436 165730 3500
rect 255865 3498 255931 3501
rect 256601 3498 256667 3501
rect 255865 3496 256667 3498
rect 255865 3440 255870 3496
rect 255926 3440 256606 3496
rect 256662 3440 256667 3496
rect 255865 3438 256667 3440
rect 255865 3435 255931 3438
rect 256601 3435 256667 3438
rect 290181 3498 290247 3501
rect 290590 3498 290596 3500
rect 290181 3496 290596 3498
rect 290181 3440 290186 3496
rect 290242 3440 290596 3496
rect 290181 3438 290596 3440
rect 290181 3435 290247 3438
rect 290590 3436 290596 3438
rect 290660 3436 290666 3500
rect 291694 3436 291700 3500
rect 291764 3498 291770 3500
rect 294873 3498 294939 3501
rect 291764 3496 294939 3498
rect 291764 3440 294878 3496
rect 294934 3440 294939 3496
rect 291764 3438 294939 3440
rect 291764 3436 291770 3438
rect 294873 3435 294939 3438
rect 299606 3436 299612 3500
rect 299676 3498 299682 3500
rect 300761 3498 300827 3501
rect 299676 3496 300827 3498
rect 299676 3440 300766 3496
rect 300822 3440 300827 3496
rect 299676 3438 300827 3440
rect 299676 3436 299682 3438
rect 300761 3435 300827 3438
rect 340965 3498 341031 3501
rect 344277 3498 344343 3501
rect 340965 3496 344343 3498
rect 340965 3440 340970 3496
rect 341026 3440 344282 3496
rect 344338 3440 344343 3496
rect 340965 3438 344343 3440
rect 340965 3435 341031 3438
rect 344277 3435 344343 3438
rect 2865 3362 2931 3365
rect 57145 3362 57211 3365
rect 2865 3360 57211 3362
rect 2865 3304 2870 3360
rect 2926 3304 57150 3360
rect 57206 3304 57211 3360
rect 2865 3302 57211 3304
rect 2865 3299 2931 3302
rect 57145 3299 57211 3302
rect 77385 3362 77451 3365
rect 196801 3362 196867 3365
rect 77385 3360 196867 3362
rect 77385 3304 77390 3360
rect 77446 3304 196806 3360
rect 196862 3304 196867 3360
rect 77385 3302 196867 3304
rect 77385 3299 77451 3302
rect 196801 3299 196867 3302
rect 256550 3300 256556 3364
rect 256620 3362 256626 3364
rect 266353 3362 266419 3365
rect 256620 3360 266419 3362
rect 256620 3304 266358 3360
rect 266414 3304 266419 3360
rect 256620 3302 266419 3304
rect 256620 3300 256626 3302
rect 266353 3299 266419 3302
rect 318517 3362 318583 3365
rect 329097 3362 329163 3365
rect 318517 3360 329163 3362
rect 318517 3304 318522 3360
rect 318578 3304 329102 3360
rect 329158 3304 329163 3360
rect 318517 3302 329163 3304
rect 318517 3299 318583 3302
rect 329097 3299 329163 3302
rect 346945 3362 347011 3365
rect 359457 3362 359523 3365
rect 346945 3360 359523 3362
rect 346945 3304 346950 3360
rect 347006 3304 359462 3360
rect 359518 3304 359523 3360
rect 346945 3302 359523 3304
rect 346945 3299 347011 3302
rect 359457 3299 359523 3302
rect 184197 2682 184263 2685
rect 278681 2682 278747 2685
rect 184197 2680 278747 2682
rect 184197 2624 184202 2680
rect 184258 2624 278686 2680
rect 278742 2624 278747 2680
rect 184197 2622 278747 2624
rect 184197 2619 184263 2622
rect 278681 2619 278747 2622
<< via3 >>
rect 69612 702476 69676 702540
rect 66116 590684 66180 590748
rect 88196 588508 88260 588572
rect 88196 585652 88260 585716
rect 69428 582252 69492 582316
rect 91140 578036 91204 578100
rect 178540 564436 178604 564500
rect 67404 556820 67468 556884
rect 66668 551380 66732 551444
rect 198596 551244 198660 551308
rect 184796 550700 184860 550764
rect 170260 546620 170324 546684
rect 358860 546484 358924 546548
rect 197860 542540 197924 542604
rect 69428 542268 69492 542332
rect 91140 542268 91204 542332
rect 353340 541316 353404 541380
rect 199332 541180 199396 541244
rect 185348 539684 185412 539748
rect 196572 538596 196636 538660
rect 194364 538324 194428 538388
rect 67404 537372 67468 537436
rect 69612 535528 69676 535532
rect 69612 535472 69626 535528
rect 69626 535472 69676 535528
rect 69612 535468 69676 535472
rect 71636 535468 71700 535532
rect 72372 535528 72436 535532
rect 72372 535472 72386 535528
rect 72386 535472 72436 535528
rect 72372 535468 72436 535472
rect 199516 535468 199580 535532
rect 200620 535468 200684 535532
rect 200068 532476 200132 532540
rect 97948 531448 98012 531452
rect 97948 531392 97998 531448
rect 97998 531392 98012 531448
rect 97948 531388 98012 531392
rect 197860 526356 197924 526420
rect 168972 523636 169036 523700
rect 199516 523636 199580 523700
rect 66668 522956 66732 523020
rect 66484 522820 66548 522884
rect 161980 518876 162044 518940
rect 191788 518060 191852 518124
rect 199332 513300 199396 513364
rect 188844 502420 188908 502484
rect 198596 500380 198660 500444
rect 356100 499836 356164 499900
rect 195100 490452 195164 490516
rect 361620 487188 361684 487252
rect 198412 483108 198476 483172
rect 122604 479436 122668 479500
rect 356652 475492 356716 475556
rect 106412 471140 106476 471204
rect 104940 469780 105004 469844
rect 115980 468420 116044 468484
rect 356284 467876 356348 467940
rect 91140 465700 91204 465764
rect 89668 464340 89732 464404
rect 107700 464340 107764 464404
rect 118004 464340 118068 464404
rect 92612 462844 92676 462908
rect 111748 460124 111812 460188
rect 93900 459580 93964 459644
rect 118740 458764 118804 458828
rect 198780 458356 198844 458420
rect 100708 457404 100772 457468
rect 108988 456996 109052 457060
rect 69796 456860 69860 456924
rect 98132 456044 98196 456108
rect 102180 456044 102244 456108
rect 96660 453188 96724 453252
rect 66116 450468 66180 450532
rect 160692 449924 160756 449988
rect 120212 449108 120276 449172
rect 72740 448624 72804 448628
rect 72740 448568 72754 448624
rect 72754 448568 72804 448624
rect 72740 448564 72804 448568
rect 95188 447748 95252 447812
rect 194548 446388 194612 446452
rect 96476 445708 96540 445772
rect 100524 445708 100588 445772
rect 115796 445708 115860 445772
rect 118556 445768 118620 445772
rect 118556 445712 118606 445768
rect 118606 445712 118620 445768
rect 118556 445708 118620 445712
rect 115796 444756 115860 444820
rect 124260 444756 124324 444820
rect 94452 444680 94516 444684
rect 94452 444624 94502 444680
rect 94502 444624 94516 444680
rect 94452 444620 94516 444624
rect 108804 444484 108868 444548
rect 111564 444544 111628 444548
rect 111564 444488 111578 444544
rect 111578 444488 111628 444544
rect 111564 444484 111628 444488
rect 114324 444544 114388 444548
rect 114324 444488 114374 444544
rect 114374 444488 114388 444544
rect 114324 444484 114388 444488
rect 67772 442172 67836 442236
rect 121684 435236 121748 435300
rect 120028 430612 120092 430676
rect 120212 425988 120276 426052
rect 198596 421636 198660 421700
rect 124260 420880 124324 420884
rect 124260 420824 124310 420880
rect 124310 420824 124324 420880
rect 124260 420820 124324 420824
rect 66668 419596 66732 419660
rect 198964 419596 199028 419660
rect 154620 411300 154684 411364
rect 69244 407764 69308 407828
rect 69244 407084 69308 407148
rect 186820 404500 186884 404564
rect 122604 403684 122668 403748
rect 177436 401644 177500 401708
rect 400260 393348 400324 393412
rect 119476 392124 119540 392188
rect 71820 391172 71884 391236
rect 92612 391036 92676 391100
rect 71820 390688 71884 390692
rect 71820 390632 71870 390688
rect 71870 390632 71884 390688
rect 71820 390628 71884 390632
rect 102180 390552 102244 390556
rect 102180 390496 102194 390552
rect 102194 390496 102244 390552
rect 102180 390492 102244 390496
rect 69612 390356 69676 390420
rect 89484 390356 89548 390420
rect 91140 390356 91204 390420
rect 93900 390356 93964 390420
rect 96660 390356 96724 390420
rect 98132 390356 98196 390420
rect 104940 390416 105004 390420
rect 104940 390360 104990 390416
rect 104990 390360 105004 390416
rect 104940 390356 105004 390360
rect 106412 390356 106476 390420
rect 107700 390356 107764 390420
rect 108988 390356 109052 390420
rect 115980 390416 116044 390420
rect 115980 390360 115994 390416
rect 115994 390360 116044 390416
rect 115980 390356 116044 390360
rect 118740 390416 118804 390420
rect 118740 390360 118790 390416
rect 118790 390360 118804 390416
rect 118740 390356 118804 390360
rect 100708 390280 100772 390284
rect 100708 390224 100758 390280
rect 100758 390224 100772 390280
rect 100708 390220 100772 390224
rect 95188 388996 95252 389060
rect 111748 388996 111812 389060
rect 118004 388996 118068 389060
rect 97948 388588 98012 388652
rect 96476 388452 96540 388516
rect 72372 388316 72436 388380
rect 95188 385596 95252 385660
rect 83964 384976 84028 384980
rect 83964 384920 83978 384976
rect 83978 384920 84028 384976
rect 83964 384916 84028 384920
rect 197308 384916 197372 384980
rect 197308 383692 197372 383756
rect 158668 380156 158732 380220
rect 124812 378796 124876 378860
rect 200620 378252 200684 378316
rect 194364 378116 194428 378180
rect 197308 377980 197372 378044
rect 120028 377300 120092 377364
rect 198964 376484 199028 376548
rect 114324 375260 114388 375324
rect 358860 375124 358924 375188
rect 166396 374580 166460 374644
rect 253060 374036 253124 374100
rect 119476 371860 119540 371924
rect 198780 369140 198844 369204
rect 154068 369004 154132 369068
rect 186820 368324 186884 368388
rect 69796 367644 69860 367708
rect 200620 367644 200684 367708
rect 287652 367508 287716 367572
rect 166212 367236 166276 367300
rect 194548 364924 194612 364988
rect 267596 364380 267660 364444
rect 108804 361720 108868 361724
rect 203012 361796 203076 361860
rect 108804 361664 108818 361720
rect 108818 361664 108868 361720
rect 108804 361660 108868 361664
rect 354444 360980 354508 361044
rect 356284 360844 356348 360908
rect 124812 360164 124876 360228
rect 166396 360028 166460 360092
rect 81020 359348 81084 359412
rect 356100 359348 356164 359412
rect 353340 357988 353404 358052
rect 111564 357580 111628 357644
rect 191236 357580 191300 357644
rect 69612 356084 69676 356148
rect 251220 355404 251284 355468
rect 100524 353500 100588 353564
rect 295932 350508 295996 350572
rect 67956 349692 68020 349756
rect 118556 349148 118620 349212
rect 121684 349012 121748 349076
rect 67772 348876 67836 348940
rect 208900 348468 208964 348532
rect 66668 346972 66732 347036
rect 94452 345748 94516 345812
rect 186820 345748 186884 345812
rect 248460 345536 248524 345540
rect 248460 345480 248510 345536
rect 248510 345480 248524 345536
rect 248460 345476 248524 345480
rect 198412 345068 198476 345132
rect 196572 344932 196636 344996
rect 156460 343844 156524 343908
rect 111748 342892 111812 342956
rect 230428 342348 230492 342412
rect 157748 341532 157812 341596
rect 219940 341396 220004 341460
rect 157748 340716 157812 340780
rect 158484 340716 158548 340780
rect 158852 340172 158916 340236
rect 115796 339900 115860 339964
rect 115796 339492 115860 339556
rect 67772 338812 67836 338876
rect 160876 337996 160940 338060
rect 213132 337452 213196 337516
rect 66116 337316 66180 337380
rect 169524 337316 169588 337380
rect 152596 333236 152660 333300
rect 69796 332556 69860 332620
rect 82676 331740 82740 331804
rect 177252 331740 177316 331804
rect 157748 331468 157812 331532
rect 141924 331332 141988 331396
rect 178724 331332 178788 331396
rect 75684 331196 75748 331260
rect 151860 329836 151924 329900
rect 157196 329700 157260 329764
rect 77156 329428 77220 329492
rect 142292 329156 142356 329220
rect 151676 329156 151740 329220
rect 152596 329216 152660 329220
rect 152596 329160 152646 329216
rect 152646 329160 152660 329216
rect 152596 329156 152660 329160
rect 259500 328536 259564 328540
rect 259500 328480 259550 328536
rect 259550 328480 259564 328536
rect 259500 328476 259564 328480
rect 69428 328340 69492 328404
rect 166212 328340 166276 328404
rect 198412 327116 198476 327180
rect 66116 325620 66180 325684
rect 157748 325348 157812 325412
rect 237420 324940 237484 325004
rect 255268 324940 255332 325004
rect 157748 324396 157812 324460
rect 69428 323988 69492 324052
rect 249748 323716 249812 323780
rect 158668 322144 158732 322148
rect 158668 322088 158718 322144
rect 158718 322088 158732 322144
rect 158668 322084 158732 322088
rect 244780 321736 244844 321740
rect 244780 321680 244794 321736
rect 244794 321680 244844 321736
rect 244780 321676 244844 321680
rect 227668 320860 227732 320924
rect 157196 320724 157260 320788
rect 210740 319500 210804 319564
rect 166396 319364 166460 319428
rect 173020 317324 173084 317388
rect 168972 316644 169036 316708
rect 187556 316644 187620 316708
rect 166212 314604 166276 314668
rect 206876 314060 206940 314124
rect 191052 313108 191116 313172
rect 156828 312564 156892 312628
rect 199332 312428 199396 312492
rect 240732 311884 240796 311948
rect 157196 310388 157260 310452
rect 173204 309844 173268 309908
rect 158852 309708 158916 309772
rect 188292 309708 188356 309772
rect 231900 306444 231964 306508
rect 159036 305764 159100 305828
rect 220860 305628 220924 305692
rect 169524 304132 169588 304196
rect 182772 304132 182836 304196
rect 248644 302500 248708 302564
rect 168420 302364 168484 302428
rect 197124 301412 197188 301476
rect 244228 300868 244292 300932
rect 226196 298692 226260 298756
rect 159036 298148 159100 298212
rect 202644 297468 202708 297532
rect 208164 297332 208228 297396
rect 67956 296244 68020 296308
rect 219204 296108 219268 296172
rect 242940 295972 243004 296036
rect 159956 295292 160020 295356
rect 267780 295292 267844 295356
rect 177436 294476 177500 294540
rect 217548 293116 217612 293180
rect 219940 292028 220004 292092
rect 211660 289852 211724 289916
rect 159220 288688 159284 288692
rect 159220 288632 159270 288688
rect 159270 288632 159284 288688
rect 159220 288628 159284 288632
rect 66668 287812 66732 287876
rect 69428 287676 69492 287740
rect 238524 287676 238588 287740
rect 233188 287132 233252 287196
rect 191236 286316 191300 286380
rect 438900 286316 438964 286380
rect 200252 285908 200316 285972
rect 232452 285908 232516 285972
rect 223620 285772 223684 285836
rect 222332 285636 222396 285700
rect 286180 285636 286244 285700
rect 425652 284956 425716 285020
rect 227852 284412 227916 284476
rect 243492 284412 243556 284476
rect 61884 284276 61948 284340
rect 214420 283928 214484 283932
rect 214420 283872 214470 283928
rect 214470 283872 214484 283928
rect 214420 283868 214484 283872
rect 216444 283928 216508 283932
rect 216444 283872 216458 283928
rect 216458 283872 216508 283928
rect 216444 283868 216508 283872
rect 218652 283868 218716 283932
rect 226932 283868 226996 283932
rect 227668 283868 227732 283932
rect 228220 283868 228284 283932
rect 229692 283868 229756 283932
rect 231716 283868 231780 283932
rect 236500 283868 236564 283932
rect 186820 283188 186884 283252
rect 198780 282916 198844 282980
rect 186820 281420 186884 281484
rect 243492 280740 243556 280804
rect 67772 280196 67836 280260
rect 244780 280196 244844 280260
rect 280292 280256 280356 280260
rect 280292 280200 280342 280256
rect 280342 280200 280356 280256
rect 280292 280196 280356 280200
rect 200068 279788 200132 279852
rect 248644 279380 248708 279444
rect 173204 278700 173268 278764
rect 158484 278020 158548 278084
rect 180012 278020 180076 278084
rect 158484 277748 158548 277812
rect 67956 277204 68020 277268
rect 160876 275164 160940 275228
rect 66116 273668 66180 273732
rect 195284 273260 195348 273324
rect 198780 273260 198844 273324
rect 185348 272444 185412 272508
rect 161980 271764 162044 271828
rect 198412 270948 198476 271012
rect 282132 270540 282196 270604
rect 244228 269044 244292 269108
rect 157932 268364 157996 268428
rect 67404 267412 67468 267476
rect 197124 267140 197188 267204
rect 244412 265780 244476 265844
rect 184612 265100 184676 265164
rect 197124 264964 197188 265028
rect 199332 264964 199396 265028
rect 186820 263604 186884 263668
rect 180196 262924 180260 262988
rect 195100 262924 195164 262988
rect 156828 262788 156892 262852
rect 245700 263060 245764 263124
rect 185348 261564 185412 261628
rect 195284 261564 195348 261628
rect 244228 261292 244292 261356
rect 195836 260884 195900 260948
rect 159956 260748 160020 260812
rect 161980 260612 162044 260676
rect 243492 259796 243556 259860
rect 251220 252452 251284 252516
rect 198596 251772 198660 251836
rect 172468 251228 172532 251292
rect 195100 249868 195164 249932
rect 67772 248916 67836 248980
rect 244780 248100 244844 248164
rect 59124 247012 59188 247076
rect 188292 247012 188356 247076
rect 197124 246468 197188 246532
rect 193812 245788 193876 245852
rect 197124 245788 197188 245852
rect 191788 245712 191852 245716
rect 191788 245656 191838 245712
rect 191838 245656 191852 245712
rect 191788 245652 191852 245656
rect 195836 245652 195900 245716
rect 156828 243476 156892 243540
rect 199332 243068 199396 243132
rect 259500 242932 259564 242996
rect 165660 242796 165724 242860
rect 81020 242040 81084 242044
rect 81020 241984 81034 242040
rect 81034 241984 81084 242040
rect 81020 241980 81084 241984
rect 154620 242040 154684 242044
rect 154620 241984 154670 242040
rect 154670 241984 154684 242040
rect 154620 241980 154684 241984
rect 196756 241708 196820 241772
rect 67404 241436 67468 241500
rect 83964 241436 84028 241500
rect 243492 241300 243556 241364
rect 160692 241164 160756 241228
rect 170260 241028 170324 241092
rect 155724 240136 155788 240140
rect 155724 240080 155738 240136
rect 155738 240080 155788 240136
rect 155724 240076 155788 240080
rect 157380 240076 157444 240140
rect 202644 240136 202708 240140
rect 202644 240080 202658 240136
rect 202658 240080 202708 240136
rect 202644 240076 202708 240080
rect 208164 240076 208228 240140
rect 208900 240076 208964 240140
rect 210740 240136 210804 240140
rect 210740 240080 210754 240136
rect 210754 240080 210804 240136
rect 210740 240076 210804 240080
rect 217548 240136 217612 240140
rect 217548 240080 217562 240136
rect 217562 240080 217612 240136
rect 217548 240076 217612 240080
rect 219204 240076 219268 240140
rect 226196 240076 226260 240140
rect 230428 240076 230492 240140
rect 231900 240076 231964 240140
rect 237420 240076 237484 240140
rect 203012 239940 203076 240004
rect 220860 239940 220924 240004
rect 226932 239396 226996 239460
rect 156644 238580 156708 238644
rect 206876 238580 206940 238644
rect 222332 238580 222396 238644
rect 244044 238580 244108 238644
rect 240732 237492 240796 237556
rect 154068 237356 154132 237420
rect 168236 237356 168300 237420
rect 196756 237356 196820 237420
rect 209820 237356 209884 237420
rect 227668 237356 227732 237420
rect 241652 237356 241716 237420
rect 72740 237220 72804 237284
rect 188844 237220 188908 237284
rect 195100 237220 195164 237284
rect 211660 237084 211724 237148
rect 199332 236948 199396 237012
rect 218652 235996 218716 236060
rect 224172 235996 224236 236060
rect 166212 235860 166276 235924
rect 156460 235724 156524 235788
rect 180196 235724 180260 235788
rect 213132 235452 213196 235516
rect 223620 234636 223684 234700
rect 242940 234500 243004 234564
rect 82676 234364 82740 234428
rect 184612 233140 184676 233204
rect 187556 233140 187620 233204
rect 168236 232868 168300 232932
rect 234660 231644 234724 231708
rect 168236 231100 168300 231164
rect 195652 231100 195716 231164
rect 185348 230284 185412 230348
rect 195836 229740 195900 229804
rect 180012 228924 180076 228988
rect 184796 228788 184860 228852
rect 184796 228244 184860 228308
rect 157932 227428 157996 227492
rect 242756 226884 242820 226948
rect 204852 226340 204916 226404
rect 283788 225524 283852 225588
rect 244412 225312 244476 225316
rect 244412 225256 244426 225312
rect 244426 225256 244476 225312
rect 244412 225252 244476 225256
rect 244780 225116 244844 225180
rect 196572 224980 196636 225044
rect 242756 224844 242820 224908
rect 178540 224300 178604 224364
rect 248644 222048 248708 222052
rect 248644 221992 248658 222048
rect 248658 221992 248708 222048
rect 248644 221988 248708 221992
rect 298140 217228 298204 217292
rect 442028 215868 442092 215932
rect 67956 215188 68020 215252
rect 252324 215188 252388 215252
rect 255268 215188 255332 215252
rect 173020 215052 173084 215116
rect 209820 215052 209884 215116
rect 237420 214644 237484 214708
rect 248460 213692 248524 213756
rect 216444 212604 216508 212668
rect 193812 212528 193876 212532
rect 193812 212472 193862 212528
rect 193862 212472 193876 212528
rect 193812 212468 193876 212472
rect 168420 212332 168484 212396
rect 230428 210428 230492 210492
rect 233372 208388 233436 208452
rect 159220 207572 159284 207636
rect 284524 207572 284588 207636
rect 290596 207572 290660 207636
rect 423996 207572 424060 207636
rect 227668 205728 227732 205732
rect 227668 205672 227718 205728
rect 227718 205672 227732 205728
rect 227668 205668 227732 205672
rect 214420 205592 214484 205596
rect 214420 205536 214470 205592
rect 214470 205536 214484 205592
rect 214420 205532 214484 205536
rect 195652 203628 195716 203692
rect 288572 201452 288636 201516
rect 204852 200636 204916 200700
rect 291700 199412 291764 199476
rect 288388 194440 288452 194444
rect 288388 194384 288438 194440
rect 288438 194384 288452 194440
rect 288388 194380 288452 194384
rect 240364 193836 240428 193900
rect 287100 193836 287164 193900
rect 256556 192476 256620 192540
rect 77156 191116 77220 191180
rect 277900 189892 277964 189956
rect 75684 189620 75748 189684
rect 237420 188532 237484 188596
rect 299612 188396 299676 188460
rect 69612 188260 69676 188324
rect 303660 187036 303724 187100
rect 155724 184316 155788 184380
rect 228220 183500 228284 183564
rect 228772 182956 228836 183020
rect 285628 182956 285692 183020
rect 280476 182820 280540 182884
rect 242940 182276 243004 182340
rect 169708 182004 169772 182068
rect 278820 181460 278884 181524
rect 169708 180780 169772 180844
rect 161980 180644 162044 180708
rect 281580 179964 281644 180028
rect 221228 179556 221292 179620
rect 282132 179420 282196 179484
rect 231900 179012 231964 179076
rect 237604 178876 237668 178940
rect 197308 178740 197372 178804
rect 232452 178060 232516 178124
rect 110644 177924 110708 177988
rect 118372 177924 118436 177988
rect 98316 177516 98380 177580
rect 100708 177516 100772 177580
rect 105676 177576 105740 177580
rect 105676 177520 105726 177576
rect 105726 177520 105740 177576
rect 105676 177516 105740 177520
rect 108068 177516 108132 177580
rect 109540 177516 109604 177580
rect 113220 177516 113284 177580
rect 115796 177576 115860 177580
rect 115796 177520 115846 177576
rect 115846 177520 115860 177576
rect 115796 177516 115860 177520
rect 116900 177516 116964 177580
rect 123156 177516 123220 177580
rect 133092 177516 133156 177580
rect 134380 177516 134444 177580
rect 148180 177576 148244 177580
rect 148180 177520 148230 177576
rect 148230 177520 148244 177576
rect 148180 177516 148244 177520
rect 112116 177380 112180 177444
rect 104572 177108 104636 177172
rect 279372 177108 279436 177172
rect 106964 177032 107028 177036
rect 106964 176976 107014 177032
rect 107014 176976 107028 177032
rect 106964 176972 107028 176976
rect 119476 176972 119540 177036
rect 127020 176972 127084 177036
rect 97028 176836 97092 176900
rect 120764 176836 120828 176900
rect 229324 176836 229388 176900
rect 101996 176760 102060 176764
rect 101996 176704 102046 176760
rect 102046 176704 102060 176760
rect 101996 176700 102060 176704
rect 124444 176700 124508 176764
rect 130700 176760 130764 176764
rect 130700 176704 130750 176760
rect 130750 176704 130764 176760
rect 130700 176700 130764 176704
rect 132356 176760 132420 176764
rect 132356 176704 132406 176760
rect 132406 176704 132420 176760
rect 132356 176700 132420 176704
rect 136036 176760 136100 176764
rect 136036 176704 136086 176760
rect 136086 176704 136100 176760
rect 136036 176700 136100 176704
rect 158852 176700 158916 176764
rect 232084 176700 232148 176764
rect 284340 176700 284404 176764
rect 99420 176428 99484 176492
rect 103284 176428 103348 176492
rect 128124 176428 128188 176492
rect 221228 175944 221292 175948
rect 221228 175888 221242 175944
rect 221242 175888 221292 175944
rect 221228 175884 221292 175888
rect 224172 175944 224236 175948
rect 224172 175888 224222 175944
rect 224222 175888 224236 175944
rect 224172 175884 224236 175888
rect 227668 175884 227732 175948
rect 125732 175748 125796 175812
rect 129412 175672 129476 175676
rect 129412 175616 129462 175672
rect 129462 175616 129476 175672
rect 129412 175612 129476 175616
rect 121868 175476 121932 175540
rect 114324 175340 114388 175404
rect 277900 175748 277964 175812
rect 229140 174388 229204 174452
rect 279372 170580 279436 170644
rect 236500 168540 236564 168604
rect 236684 168404 236748 168468
rect 244412 167588 244476 167652
rect 237604 165684 237668 165748
rect 242940 162012 243004 162076
rect 240364 161468 240428 161532
rect 286180 160652 286244 160716
rect 233372 160516 233436 160580
rect 233740 160108 233804 160172
rect 236684 160108 236748 160172
rect 240732 160108 240796 160172
rect 283788 157252 283852 157316
rect 233188 157116 233252 157180
rect 230428 156164 230492 156228
rect 281580 154940 281644 155004
rect 244228 153716 244292 153780
rect 282132 153716 282196 153780
rect 231900 151540 231964 151604
rect 170260 150996 170324 151060
rect 215892 150996 215956 151060
rect 233188 150996 233252 151060
rect 241652 150996 241716 151060
rect 232084 150588 232148 150652
rect 229140 150044 229204 150108
rect 233740 149092 233804 149156
rect 234108 148004 234172 148068
rect 298140 147732 298204 147796
rect 231164 146916 231228 146980
rect 409828 143440 409892 143444
rect 409828 143384 409878 143440
rect 409878 143384 409892 143440
rect 409828 143380 409892 143384
rect 417372 143380 417436 143444
rect 230980 142700 231044 142764
rect 233188 142428 233252 142492
rect 431908 142216 431972 142220
rect 431908 142160 431958 142216
rect 431958 142160 431972 142216
rect 431908 142156 431972 142160
rect 238708 142020 238772 142084
rect 248644 141068 248708 141132
rect 303660 140856 303724 140860
rect 303660 140800 303674 140856
rect 303674 140800 303724 140856
rect 303660 140796 303724 140800
rect 441660 140856 441724 140860
rect 441660 140800 441710 140856
rect 441710 140800 441724 140856
rect 441660 140796 441724 140800
rect 266860 140388 266924 140452
rect 231900 139708 231964 139772
rect 280108 139708 280172 139772
rect 419028 139708 419092 139772
rect 420684 139572 420748 139636
rect 421052 139436 421116 139500
rect 426388 139436 426452 139500
rect 427860 139436 427924 139500
rect 429148 139436 429212 139500
rect 435036 139496 435100 139500
rect 435036 139440 435050 139496
rect 435050 139440 435100 139496
rect 435036 139436 435100 139440
rect 439084 139496 439148 139500
rect 439084 139440 439098 139496
rect 439098 139440 439148 139496
rect 439084 139436 439148 139440
rect 234660 139164 234724 139228
rect 237420 138756 237484 138820
rect 441660 138620 441724 138684
rect 229692 137260 229756 137324
rect 236500 137260 236564 137324
rect 229876 137124 229940 137188
rect 400260 135084 400324 135148
rect 262812 134812 262876 134876
rect 231164 134404 231228 134468
rect 249012 133860 249076 133924
rect 230428 133588 230492 133652
rect 284524 133588 284588 133652
rect 282132 132092 282196 132156
rect 258580 130596 258644 130660
rect 242756 130188 242820 130252
rect 264100 130052 264164 130116
rect 232452 128964 232516 129028
rect 244044 127332 244108 127396
rect 260052 126380 260116 126444
rect 442212 125020 442276 125084
rect 244780 124612 244844 124676
rect 214420 123252 214484 123316
rect 230980 123116 231044 123180
rect 439268 120532 439332 120596
rect 439636 120532 439700 120596
rect 240732 119988 240796 120052
rect 361620 117132 361684 117196
rect 233740 113460 233804 113524
rect 439268 113052 439332 113116
rect 285628 111556 285692 111620
rect 168236 109652 168300 109716
rect 287100 109380 287164 109444
rect 267780 108836 267844 108900
rect 267964 107068 268028 107132
rect 234108 106116 234172 106180
rect 264100 105572 264164 105636
rect 280292 105436 280356 105500
rect 442028 105300 442092 105364
rect 197308 104756 197372 104820
rect 237972 102852 238036 102916
rect 398788 102716 398852 102780
rect 262996 102172 263060 102236
rect 284340 101628 284404 101692
rect 423996 100676 424060 100740
rect 425652 100676 425716 100740
rect 279372 100540 279436 100604
rect 262996 99996 263060 100060
rect 398788 99316 398852 99380
rect 267780 99180 267844 99244
rect 264100 97412 264164 97476
rect 229140 97004 229204 97068
rect 225092 95976 225156 95980
rect 225092 95920 225106 95976
rect 225106 95920 225156 95976
rect 225092 95916 225156 95920
rect 226380 95976 226444 95980
rect 226380 95920 226430 95976
rect 226430 95920 226444 95976
rect 226380 95916 226444 95920
rect 226932 95916 226996 95980
rect 242756 95644 242820 95708
rect 442212 95780 442276 95844
rect 113142 94752 113206 94756
rect 113142 94696 113178 94752
rect 113178 94696 113206 94752
rect 113142 94692 113206 94696
rect 130686 94692 130750 94756
rect 151492 94692 151556 94756
rect 151766 94692 151830 94756
rect 230428 94692 230492 94756
rect 267596 94556 267660 94620
rect 214420 94420 214484 94484
rect 100892 93876 100956 93940
rect 99236 93740 99300 93804
rect 118188 93604 118252 93668
rect 228772 93604 228836 93668
rect 110092 93468 110156 93532
rect 119660 93392 119724 93396
rect 119660 93336 119710 93392
rect 119710 93336 119724 93392
rect 119660 93332 119724 93336
rect 122972 93392 123036 93396
rect 122972 93336 123022 93392
rect 123022 93336 123036 93392
rect 122972 93332 123036 93336
rect 103284 93196 103348 93260
rect 74764 92440 74828 92444
rect 74764 92384 74814 92440
rect 74814 92384 74828 92440
rect 74764 92380 74828 92384
rect 97212 92380 97276 92444
rect 99972 92380 100036 92444
rect 102732 92380 102796 92444
rect 108068 92380 108132 92444
rect 116716 92440 116780 92444
rect 116716 92384 116766 92440
rect 116766 92384 116780 92440
rect 116716 92380 116780 92384
rect 124076 92440 124140 92444
rect 124076 92384 124126 92440
rect 124126 92384 124140 92440
rect 124076 92380 124140 92384
rect 134380 92440 134444 92444
rect 134380 92384 134430 92440
rect 134430 92384 134444 92440
rect 134380 92380 134444 92384
rect 151308 92440 151372 92444
rect 151308 92384 151358 92440
rect 151358 92384 151372 92440
rect 151308 92380 151372 92384
rect 106780 92244 106844 92308
rect 253060 92244 253124 92308
rect 88012 92168 88076 92172
rect 88012 92112 88062 92168
rect 88062 92112 88076 92168
rect 88012 92108 88076 92112
rect 133092 92108 133156 92172
rect 91324 91972 91388 92036
rect 109172 91700 109236 91764
rect 120580 91700 120644 91764
rect 136036 91700 136100 91764
rect 101996 91564 102060 91628
rect 126652 91488 126716 91492
rect 126652 91432 126702 91488
rect 126702 91432 126716 91488
rect 126652 91428 126716 91432
rect 85804 91292 85868 91356
rect 95004 91352 95068 91356
rect 95004 91296 95054 91352
rect 95054 91296 95068 91352
rect 95004 91292 95068 91296
rect 98500 91292 98564 91356
rect 110644 91292 110708 91356
rect 113220 91292 113284 91356
rect 115428 91352 115492 91356
rect 115428 91296 115478 91352
rect 115478 91296 115492 91352
rect 115428 91292 115492 91296
rect 115796 91352 115860 91356
rect 115796 91296 115810 91352
rect 115810 91296 115860 91352
rect 115796 91292 115860 91296
rect 124444 91292 124508 91356
rect 125732 91292 125796 91356
rect 151492 91352 151556 91356
rect 151492 91296 151542 91352
rect 151542 91296 151556 91352
rect 151492 91292 151556 91296
rect 84332 91156 84396 91220
rect 86724 91216 86788 91220
rect 86724 91160 86774 91216
rect 86774 91160 86788 91216
rect 86724 91156 86788 91160
rect 88932 91156 88996 91220
rect 90220 91156 90284 91220
rect 92612 91156 92676 91220
rect 93900 91156 93964 91220
rect 96292 91156 96356 91220
rect 96660 91156 96724 91220
rect 98132 91156 98196 91220
rect 100524 91216 100588 91220
rect 100524 91160 100574 91216
rect 100574 91160 100588 91216
rect 100524 91156 100588 91160
rect 101812 91156 101876 91220
rect 104204 91216 104268 91220
rect 104204 91160 104254 91216
rect 104254 91160 104268 91216
rect 104204 91156 104268 91160
rect 104572 91156 104636 91220
rect 105492 91216 105556 91220
rect 105492 91160 105542 91216
rect 105542 91160 105556 91216
rect 105492 91156 105556 91160
rect 105676 91156 105740 91220
rect 106412 91156 106476 91220
rect 107700 91156 107764 91220
rect 109540 91156 109604 91220
rect 111196 91156 111260 91220
rect 111932 91156 111996 91220
rect 112300 91156 112364 91220
rect 114324 91156 114388 91220
rect 114876 91156 114940 91220
rect 117084 91216 117148 91220
rect 117084 91160 117134 91216
rect 117134 91160 117148 91216
rect 117084 91156 117148 91160
rect 118004 91156 118068 91220
rect 119292 91156 119356 91220
rect 120212 91156 120276 91220
rect 121684 91156 121748 91220
rect 122052 91156 122116 91220
rect 123156 91156 123220 91220
rect 125364 91216 125428 91220
rect 125364 91160 125414 91216
rect 125414 91160 125428 91216
rect 125364 91156 125428 91160
rect 126468 91156 126532 91220
rect 127572 91156 127636 91220
rect 129412 91156 129476 91220
rect 132356 91216 132420 91220
rect 132356 91160 132406 91216
rect 132406 91160 132420 91216
rect 132356 91156 132420 91160
rect 151676 91216 151740 91220
rect 151676 91160 151726 91216
rect 151726 91160 151740 91216
rect 151676 91156 151740 91160
rect 152044 91156 152108 91220
rect 224724 91020 224788 91084
rect 420684 90340 420748 90404
rect 245700 89116 245764 89180
rect 291700 86940 291764 87004
rect 215892 86124 215956 86188
rect 191052 84764 191116 84828
rect 244780 80820 244844 80884
rect 264100 80684 264164 80748
rect 237972 79596 238036 79660
rect 229876 77964 229940 78028
rect 421052 73748 421116 73812
rect 258580 71028 258644 71092
rect 168236 67492 168300 67556
rect 431724 65452 431788 65516
rect 287652 64092 287716 64156
rect 267964 62732 268028 62796
rect 288572 62732 288636 62796
rect 249012 61372 249076 61436
rect 288388 60480 288452 60484
rect 288388 60424 288402 60480
rect 288402 60424 288452 60480
rect 288388 60420 288452 60424
rect 262812 59876 262876 59940
rect 409828 57156 409892 57220
rect 260052 55796 260116 55860
rect 233740 54436 233804 54500
rect 252508 53076 252572 53140
rect 429148 53076 429212 53140
rect 249748 50960 249812 50964
rect 249748 50904 249798 50960
rect 249798 50904 249812 50960
rect 249748 50900 249812 50904
rect 232452 42060 232516 42124
rect 226380 37980 226444 38044
rect 66116 37844 66180 37908
rect 267780 36484 267844 36548
rect 186820 35124 186884 35188
rect 61884 33764 61948 33828
rect 417372 33764 417436 33828
rect 426388 33084 426452 33148
rect 169524 26828 169588 26892
rect 67772 25604 67836 25668
rect 244044 25468 244108 25532
rect 236500 24108 236564 24172
rect 435036 24108 435100 24172
rect 419028 23292 419092 23356
rect 226932 21252 226996 21316
rect 427860 17852 427924 17916
rect 266860 17172 266924 17236
rect 172468 15812 172532 15876
rect 177252 15812 177316 15876
rect 59124 15132 59188 15196
rect 295932 13696 295996 13700
rect 295932 13640 295946 13696
rect 295946 13640 295996 13696
rect 295932 13636 295996 13640
rect 299612 13152 299676 13156
rect 299612 13096 299662 13152
rect 299662 13096 299676 13152
rect 299612 13092 299676 13096
rect 252324 11732 252388 11796
rect 182772 11596 182836 11660
rect 439084 9556 439148 9620
rect 178724 7516 178788 7580
rect 227668 4796 227732 4860
rect 165660 3436 165724 3500
rect 290596 3436 290660 3500
rect 291700 3436 291764 3500
rect 299612 3436 299676 3500
rect 256556 3300 256620 3364
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 680614 -8106 711002
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 -8106 680614
rect -8726 680294 -8106 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 -8106 680294
rect -8726 644614 -8106 680058
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 -8106 644614
rect -8726 644294 -8106 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 -8106 644294
rect -8726 608614 -8106 644058
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 -8106 608614
rect -8726 608294 -8106 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 -8106 608294
rect -8726 572614 -8106 608058
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 -8106 572614
rect -8726 572294 -8106 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 -8106 572294
rect -8726 536614 -8106 572058
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 -8106 536614
rect -8726 536294 -8106 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 -8106 536294
rect -8726 500614 -8106 536058
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 -8106 500614
rect -8726 500294 -8106 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 -8106 500294
rect -8726 464614 -8106 500058
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 -8106 464614
rect -8726 464294 -8106 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 -8106 464294
rect -8726 428614 -8106 464058
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 -8106 428614
rect -8726 428294 -8106 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 -8106 428294
rect -8726 392614 -8106 428058
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 -8106 392614
rect -8726 392294 -8106 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 -8106 392294
rect -8726 356614 -8106 392058
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 -8106 356614
rect -8726 356294 -8106 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 -8106 356294
rect -8726 320614 -8106 356058
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 -8106 320614
rect -8726 320294 -8106 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 -8106 320294
rect -8726 284614 -8106 320058
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 -8106 284614
rect -8726 284294 -8106 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 -8106 284294
rect -8726 248614 -8106 284058
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 -8106 248614
rect -8726 248294 -8106 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 -8106 248294
rect -8726 212614 -8106 248058
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 -8106 212614
rect -8726 212294 -8106 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 -8106 212294
rect -8726 176614 -8106 212058
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 -8106 176614
rect -8726 176294 -8106 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 -8106 176294
rect -8726 140614 -8106 176058
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 -8106 140614
rect -8726 140294 -8106 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 -8106 140294
rect -8726 104614 -8106 140058
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 -8106 104614
rect -8726 104294 -8106 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 -8106 104294
rect -8726 68614 -8106 104058
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 -8106 68614
rect -8726 68294 -8106 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 -8106 68294
rect -8726 32614 -8106 68058
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 -8106 32614
rect -8726 32294 -8106 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 -8106 32294
rect -8726 -7066 -8106 32058
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 698614 -7146 710042
rect 12954 710598 13574 711590
rect 12954 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 13574 710598
rect 12954 710278 13574 710362
rect 12954 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 13574 710278
rect -7766 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 -7146 698614
rect -7766 698294 -7146 698378
rect -7766 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 -7146 698294
rect -7766 662614 -7146 698058
rect -7766 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 -7146 662614
rect -7766 662294 -7146 662378
rect -7766 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 -7146 662294
rect -7766 626614 -7146 662058
rect -7766 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 -7146 626614
rect -7766 626294 -7146 626378
rect -7766 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 -7146 626294
rect -7766 590614 -7146 626058
rect -7766 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 -7146 590614
rect -7766 590294 -7146 590378
rect -7766 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 -7146 590294
rect -7766 554614 -7146 590058
rect -7766 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 -7146 554614
rect -7766 554294 -7146 554378
rect -7766 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 -7146 554294
rect -7766 518614 -7146 554058
rect -7766 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 -7146 518614
rect -7766 518294 -7146 518378
rect -7766 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 -7146 518294
rect -7766 482614 -7146 518058
rect -7766 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 -7146 482614
rect -7766 482294 -7146 482378
rect -7766 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 -7146 482294
rect -7766 446614 -7146 482058
rect -7766 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 -7146 446614
rect -7766 446294 -7146 446378
rect -7766 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 -7146 446294
rect -7766 410614 -7146 446058
rect -7766 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 -7146 410614
rect -7766 410294 -7146 410378
rect -7766 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 -7146 410294
rect -7766 374614 -7146 410058
rect -7766 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 -7146 374614
rect -7766 374294 -7146 374378
rect -7766 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 -7146 374294
rect -7766 338614 -7146 374058
rect -7766 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 -7146 338614
rect -7766 338294 -7146 338378
rect -7766 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 -7146 338294
rect -7766 302614 -7146 338058
rect -7766 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 -7146 302614
rect -7766 302294 -7146 302378
rect -7766 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 -7146 302294
rect -7766 266614 -7146 302058
rect -7766 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 -7146 266614
rect -7766 266294 -7146 266378
rect -7766 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 -7146 266294
rect -7766 230614 -7146 266058
rect -7766 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 -7146 230614
rect -7766 230294 -7146 230378
rect -7766 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 -7146 230294
rect -7766 194614 -7146 230058
rect -7766 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 -7146 194614
rect -7766 194294 -7146 194378
rect -7766 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 -7146 194294
rect -7766 158614 -7146 194058
rect -7766 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 -7146 158614
rect -7766 158294 -7146 158378
rect -7766 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 -7146 158294
rect -7766 122614 -7146 158058
rect -7766 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 -7146 122614
rect -7766 122294 -7146 122378
rect -7766 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 -7146 122294
rect -7766 86614 -7146 122058
rect -7766 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 -7146 86614
rect -7766 86294 -7146 86378
rect -7766 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 -7146 86294
rect -7766 50614 -7146 86058
rect -7766 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 -7146 50614
rect -7766 50294 -7146 50378
rect -7766 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 -7146 50294
rect -7766 14614 -7146 50058
rect -7766 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 -7146 14614
rect -7766 14294 -7146 14378
rect -7766 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 -7146 14294
rect -7766 -6106 -7146 14058
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 676894 -6186 709082
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 -6186 676894
rect -6806 676574 -6186 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 -6186 676574
rect -6806 640894 -6186 676338
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 -6186 640894
rect -6806 640574 -6186 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 -6186 640574
rect -6806 604894 -6186 640338
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 -6186 604894
rect -6806 604574 -6186 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 -6186 604574
rect -6806 568894 -6186 604338
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 -6186 568894
rect -6806 568574 -6186 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 -6186 568574
rect -6806 532894 -6186 568338
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 -6186 532894
rect -6806 532574 -6186 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 -6186 532574
rect -6806 496894 -6186 532338
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 -6186 496894
rect -6806 496574 -6186 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 -6186 496574
rect -6806 460894 -6186 496338
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 -6186 460894
rect -6806 460574 -6186 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 -6186 460574
rect -6806 424894 -6186 460338
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 -6186 424894
rect -6806 424574 -6186 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 -6186 424574
rect -6806 388894 -6186 424338
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 -6186 388894
rect -6806 388574 -6186 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 -6186 388574
rect -6806 352894 -6186 388338
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 -6186 352894
rect -6806 352574 -6186 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 -6186 352574
rect -6806 316894 -6186 352338
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 -6186 316894
rect -6806 316574 -6186 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 -6186 316574
rect -6806 280894 -6186 316338
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 -6186 280894
rect -6806 280574 -6186 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 -6186 280574
rect -6806 244894 -6186 280338
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 -6186 244894
rect -6806 244574 -6186 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 -6186 244574
rect -6806 208894 -6186 244338
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 -6186 208894
rect -6806 208574 -6186 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 -6186 208574
rect -6806 172894 -6186 208338
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 -6186 172894
rect -6806 172574 -6186 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 -6186 172574
rect -6806 136894 -6186 172338
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 -6186 136894
rect -6806 136574 -6186 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 -6186 136574
rect -6806 100894 -6186 136338
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 -6186 100894
rect -6806 100574 -6186 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 -6186 100574
rect -6806 64894 -6186 100338
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 -6186 64894
rect -6806 64574 -6186 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 -6186 64574
rect -6806 28894 -6186 64338
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 -6186 28894
rect -6806 28574 -6186 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 -6186 28574
rect -6806 -5146 -6186 28338
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 694894 -5226 708122
rect 9234 708678 9854 709670
rect 9234 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 9854 708678
rect 9234 708358 9854 708442
rect 9234 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 9854 708358
rect -5846 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 -5226 694894
rect -5846 694574 -5226 694658
rect -5846 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 -5226 694574
rect -5846 658894 -5226 694338
rect -5846 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 -5226 658894
rect -5846 658574 -5226 658658
rect -5846 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 -5226 658574
rect -5846 622894 -5226 658338
rect -5846 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 -5226 622894
rect -5846 622574 -5226 622658
rect -5846 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 -5226 622574
rect -5846 586894 -5226 622338
rect -5846 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 -5226 586894
rect -5846 586574 -5226 586658
rect -5846 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 -5226 586574
rect -5846 550894 -5226 586338
rect -5846 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 -5226 550894
rect -5846 550574 -5226 550658
rect -5846 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 -5226 550574
rect -5846 514894 -5226 550338
rect -5846 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 -5226 514894
rect -5846 514574 -5226 514658
rect -5846 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 -5226 514574
rect -5846 478894 -5226 514338
rect -5846 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 -5226 478894
rect -5846 478574 -5226 478658
rect -5846 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 -5226 478574
rect -5846 442894 -5226 478338
rect -5846 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 -5226 442894
rect -5846 442574 -5226 442658
rect -5846 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 -5226 442574
rect -5846 406894 -5226 442338
rect -5846 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 -5226 406894
rect -5846 406574 -5226 406658
rect -5846 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 -5226 406574
rect -5846 370894 -5226 406338
rect -5846 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 -5226 370894
rect -5846 370574 -5226 370658
rect -5846 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 -5226 370574
rect -5846 334894 -5226 370338
rect -5846 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 -5226 334894
rect -5846 334574 -5226 334658
rect -5846 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 -5226 334574
rect -5846 298894 -5226 334338
rect -5846 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 -5226 298894
rect -5846 298574 -5226 298658
rect -5846 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 -5226 298574
rect -5846 262894 -5226 298338
rect -5846 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 -5226 262894
rect -5846 262574 -5226 262658
rect -5846 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 -5226 262574
rect -5846 226894 -5226 262338
rect -5846 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 -5226 226894
rect -5846 226574 -5226 226658
rect -5846 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 -5226 226574
rect -5846 190894 -5226 226338
rect -5846 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 -5226 190894
rect -5846 190574 -5226 190658
rect -5846 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 -5226 190574
rect -5846 154894 -5226 190338
rect -5846 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 -5226 154894
rect -5846 154574 -5226 154658
rect -5846 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 -5226 154574
rect -5846 118894 -5226 154338
rect -5846 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 -5226 118894
rect -5846 118574 -5226 118658
rect -5846 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 -5226 118574
rect -5846 82894 -5226 118338
rect -5846 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 -5226 82894
rect -5846 82574 -5226 82658
rect -5846 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 -5226 82574
rect -5846 46894 -5226 82338
rect -5846 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 -5226 46894
rect -5846 46574 -5226 46658
rect -5846 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 -5226 46574
rect -5846 10894 -5226 46338
rect -5846 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 -5226 10894
rect -5846 10574 -5226 10658
rect -5846 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 -5226 10574
rect -5846 -4186 -5226 10338
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 673174 -4266 707162
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 -4266 673174
rect -4886 672854 -4266 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 -4266 672854
rect -4886 637174 -4266 672618
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 -4266 637174
rect -4886 636854 -4266 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 -4266 636854
rect -4886 601174 -4266 636618
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 -4266 601174
rect -4886 600854 -4266 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 -4266 600854
rect -4886 565174 -4266 600618
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 -4266 565174
rect -4886 564854 -4266 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 -4266 564854
rect -4886 529174 -4266 564618
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 -4266 529174
rect -4886 528854 -4266 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 -4266 528854
rect -4886 493174 -4266 528618
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 -4266 493174
rect -4886 492854 -4266 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 -4266 492854
rect -4886 457174 -4266 492618
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 -4266 457174
rect -4886 456854 -4266 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 -4266 456854
rect -4886 421174 -4266 456618
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 -4266 421174
rect -4886 420854 -4266 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 -4266 420854
rect -4886 385174 -4266 420618
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 -4266 385174
rect -4886 384854 -4266 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 -4266 384854
rect -4886 349174 -4266 384618
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 -4266 349174
rect -4886 348854 -4266 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 -4266 348854
rect -4886 313174 -4266 348618
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 -4266 313174
rect -4886 312854 -4266 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 -4266 312854
rect -4886 277174 -4266 312618
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 -4266 277174
rect -4886 276854 -4266 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 -4266 276854
rect -4886 241174 -4266 276618
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 -4266 241174
rect -4886 240854 -4266 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 -4266 240854
rect -4886 205174 -4266 240618
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 -4266 205174
rect -4886 204854 -4266 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 -4266 204854
rect -4886 169174 -4266 204618
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 -4266 169174
rect -4886 168854 -4266 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 -4266 168854
rect -4886 133174 -4266 168618
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 -4266 133174
rect -4886 132854 -4266 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 -4266 132854
rect -4886 97174 -4266 132618
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 -4266 97174
rect -4886 96854 -4266 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 -4266 96854
rect -4886 61174 -4266 96618
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 -4266 61174
rect -4886 60854 -4266 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 -4266 60854
rect -4886 25174 -4266 60618
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 -4266 25174
rect -4886 24854 -4266 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 -4266 24854
rect -4886 -3226 -4266 24618
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 691174 -3306 706202
rect 5514 706758 6134 707750
rect 5514 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 6134 706758
rect 5514 706438 6134 706522
rect 5514 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 6134 706438
rect -3926 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 -3306 691174
rect -3926 690854 -3306 690938
rect -3926 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 -3306 690854
rect -3926 655174 -3306 690618
rect -3926 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 -3306 655174
rect -3926 654854 -3306 654938
rect -3926 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 -3306 654854
rect -3926 619174 -3306 654618
rect -3926 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 -3306 619174
rect -3926 618854 -3306 618938
rect -3926 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 -3306 618854
rect -3926 583174 -3306 618618
rect -3926 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 -3306 583174
rect -3926 582854 -3306 582938
rect -3926 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 -3306 582854
rect -3926 547174 -3306 582618
rect -3926 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 -3306 547174
rect -3926 546854 -3306 546938
rect -3926 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 -3306 546854
rect -3926 511174 -3306 546618
rect -3926 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 -3306 511174
rect -3926 510854 -3306 510938
rect -3926 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 -3306 510854
rect -3926 475174 -3306 510618
rect -3926 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 -3306 475174
rect -3926 474854 -3306 474938
rect -3926 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 -3306 474854
rect -3926 439174 -3306 474618
rect -3926 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 -3306 439174
rect -3926 438854 -3306 438938
rect -3926 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 -3306 438854
rect -3926 403174 -3306 438618
rect -3926 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 -3306 403174
rect -3926 402854 -3306 402938
rect -3926 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 -3306 402854
rect -3926 367174 -3306 402618
rect -3926 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 -3306 367174
rect -3926 366854 -3306 366938
rect -3926 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 -3306 366854
rect -3926 331174 -3306 366618
rect -3926 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 -3306 331174
rect -3926 330854 -3306 330938
rect -3926 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 -3306 330854
rect -3926 295174 -3306 330618
rect -3926 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 -3306 295174
rect -3926 294854 -3306 294938
rect -3926 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 -3306 294854
rect -3926 259174 -3306 294618
rect -3926 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 -3306 259174
rect -3926 258854 -3306 258938
rect -3926 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 -3306 258854
rect -3926 223174 -3306 258618
rect -3926 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 -3306 223174
rect -3926 222854 -3306 222938
rect -3926 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 -3306 222854
rect -3926 187174 -3306 222618
rect -3926 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 -3306 187174
rect -3926 186854 -3306 186938
rect -3926 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 -3306 186854
rect -3926 151174 -3306 186618
rect -3926 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 -3306 151174
rect -3926 150854 -3306 150938
rect -3926 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 -3306 150854
rect -3926 115174 -3306 150618
rect -3926 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 -3306 115174
rect -3926 114854 -3306 114938
rect -3926 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 -3306 114854
rect -3926 79174 -3306 114618
rect -3926 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 -3306 79174
rect -3926 78854 -3306 78938
rect -3926 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 -3306 78854
rect -3926 43174 -3306 78618
rect -3926 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 -3306 43174
rect -3926 42854 -3306 42938
rect -3926 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 -3306 42854
rect -3926 7174 -3306 42618
rect -3926 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 -3306 7174
rect -3926 6854 -3306 6938
rect -3926 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 -3306 6854
rect -3926 -2266 -3306 6618
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 669454 -2346 705242
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 -2346 669454
rect -2966 669134 -2346 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 -2346 669134
rect -2966 633454 -2346 668898
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 -2346 633454
rect -2966 633134 -2346 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 -2346 633134
rect -2966 597454 -2346 632898
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 -2346 597454
rect -2966 597134 -2346 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 -2346 597134
rect -2966 561454 -2346 596898
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 -2346 561454
rect -2966 561134 -2346 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 -2346 561134
rect -2966 525454 -2346 560898
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 -2346 525454
rect -2966 525134 -2346 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 -2346 525134
rect -2966 489454 -2346 524898
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 -2346 489454
rect -2966 489134 -2346 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 -2346 489134
rect -2966 453454 -2346 488898
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 -2346 453454
rect -2966 453134 -2346 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 -2346 453134
rect -2966 417454 -2346 452898
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 -2346 417454
rect -2966 417134 -2346 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 -2346 417134
rect -2966 381454 -2346 416898
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 -2346 381454
rect -2966 381134 -2346 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 -2346 381134
rect -2966 345454 -2346 380898
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 -2346 345454
rect -2966 345134 -2346 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 -2346 345134
rect -2966 309454 -2346 344898
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 -2346 309454
rect -2966 309134 -2346 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 -2346 309134
rect -2966 273454 -2346 308898
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 -2346 273454
rect -2966 273134 -2346 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 -2346 273134
rect -2966 237454 -2346 272898
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 -2346 237454
rect -2966 237134 -2346 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 -2346 237134
rect -2966 201454 -2346 236898
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 -2346 201454
rect -2966 201134 -2346 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 -2346 201134
rect -2966 165454 -2346 200898
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 -2346 165454
rect -2966 165134 -2346 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 -2346 165134
rect -2966 129454 -2346 164898
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 -2346 129454
rect -2966 129134 -2346 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 -2346 129134
rect -2966 93454 -2346 128898
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 -2346 93454
rect -2966 93134 -2346 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 -2346 93134
rect -2966 57454 -2346 92898
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 -2346 57454
rect -2966 57134 -2346 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 -2346 57134
rect -2966 21454 -2346 56898
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 -2346 21454
rect -2966 21134 -2346 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 -2346 21134
rect -2966 -1306 -2346 20898
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 705830
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect 1794 -1894 2414 -902
rect 5514 691174 6134 706202
rect 5514 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 6134 691174
rect 5514 690854 6134 690938
rect 5514 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 6134 690854
rect 5514 655174 6134 690618
rect 5514 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 6134 655174
rect 5514 654854 6134 654938
rect 5514 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 6134 654854
rect 5514 619174 6134 654618
rect 5514 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 6134 619174
rect 5514 618854 6134 618938
rect 5514 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 6134 618854
rect 5514 583174 6134 618618
rect 5514 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 6134 583174
rect 5514 582854 6134 582938
rect 5514 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 6134 582854
rect 5514 547174 6134 582618
rect 5514 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 6134 547174
rect 5514 546854 6134 546938
rect 5514 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 6134 546854
rect 5514 511174 6134 546618
rect 5514 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 6134 511174
rect 5514 510854 6134 510938
rect 5514 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 6134 510854
rect 5514 475174 6134 510618
rect 5514 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 6134 475174
rect 5514 474854 6134 474938
rect 5514 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 6134 474854
rect 5514 439174 6134 474618
rect 5514 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 6134 439174
rect 5514 438854 6134 438938
rect 5514 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 6134 438854
rect 5514 403174 6134 438618
rect 5514 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 6134 403174
rect 5514 402854 6134 402938
rect 5514 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 6134 402854
rect 5514 367174 6134 402618
rect 5514 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 6134 367174
rect 5514 366854 6134 366938
rect 5514 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 6134 366854
rect 5514 331174 6134 366618
rect 5514 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 6134 331174
rect 5514 330854 6134 330938
rect 5514 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 6134 330854
rect 5514 295174 6134 330618
rect 5514 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 6134 295174
rect 5514 294854 6134 294938
rect 5514 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 6134 294854
rect 5514 259174 6134 294618
rect 5514 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 6134 259174
rect 5514 258854 6134 258938
rect 5514 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 6134 258854
rect 5514 223174 6134 258618
rect 5514 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 6134 223174
rect 5514 222854 6134 222938
rect 5514 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 6134 222854
rect 5514 187174 6134 222618
rect 5514 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 6134 187174
rect 5514 186854 6134 186938
rect 5514 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 6134 186854
rect 5514 151174 6134 186618
rect 5514 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 6134 151174
rect 5514 150854 6134 150938
rect 5514 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 6134 150854
rect 5514 115174 6134 150618
rect 5514 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 6134 115174
rect 5514 114854 6134 114938
rect 5514 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 6134 114854
rect 5514 79174 6134 114618
rect 5514 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 6134 79174
rect 5514 78854 6134 78938
rect 5514 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 6134 78854
rect 5514 43174 6134 78618
rect 5514 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 6134 43174
rect 5514 42854 6134 42938
rect 5514 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 6134 42854
rect 5514 7174 6134 42618
rect 5514 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 6134 7174
rect 5514 6854 6134 6938
rect 5514 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 6134 6854
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect 5514 -2266 6134 6618
rect 5514 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 6134 -2266
rect 5514 -2586 6134 -2502
rect 5514 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 6134 -2586
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect 5514 -3814 6134 -2822
rect 9234 694894 9854 708122
rect 9234 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 9854 694894
rect 9234 694574 9854 694658
rect 9234 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 9854 694574
rect 9234 658894 9854 694338
rect 9234 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 9854 658894
rect 9234 658574 9854 658658
rect 9234 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 9854 658574
rect 9234 622894 9854 658338
rect 9234 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 9854 622894
rect 9234 622574 9854 622658
rect 9234 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 9854 622574
rect 9234 586894 9854 622338
rect 9234 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 9854 586894
rect 9234 586574 9854 586658
rect 9234 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 9854 586574
rect 9234 550894 9854 586338
rect 9234 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 9854 550894
rect 9234 550574 9854 550658
rect 9234 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 9854 550574
rect 9234 514894 9854 550338
rect 9234 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 9854 514894
rect 9234 514574 9854 514658
rect 9234 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 9854 514574
rect 9234 478894 9854 514338
rect 9234 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 9854 478894
rect 9234 478574 9854 478658
rect 9234 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 9854 478574
rect 9234 442894 9854 478338
rect 9234 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 9854 442894
rect 9234 442574 9854 442658
rect 9234 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 9854 442574
rect 9234 406894 9854 442338
rect 9234 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 9854 406894
rect 9234 406574 9854 406658
rect 9234 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 9854 406574
rect 9234 370894 9854 406338
rect 9234 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 9854 370894
rect 9234 370574 9854 370658
rect 9234 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 9854 370574
rect 9234 334894 9854 370338
rect 9234 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 9854 334894
rect 9234 334574 9854 334658
rect 9234 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 9854 334574
rect 9234 298894 9854 334338
rect 9234 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 9854 298894
rect 9234 298574 9854 298658
rect 9234 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 9854 298574
rect 9234 262894 9854 298338
rect 9234 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 9854 262894
rect 9234 262574 9854 262658
rect 9234 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 9854 262574
rect 9234 226894 9854 262338
rect 9234 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 9854 226894
rect 9234 226574 9854 226658
rect 9234 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 9854 226574
rect 9234 190894 9854 226338
rect 9234 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 9854 190894
rect 9234 190574 9854 190658
rect 9234 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 9854 190574
rect 9234 154894 9854 190338
rect 9234 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 9854 154894
rect 9234 154574 9854 154658
rect 9234 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 9854 154574
rect 9234 118894 9854 154338
rect 9234 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 9854 118894
rect 9234 118574 9854 118658
rect 9234 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 9854 118574
rect 9234 82894 9854 118338
rect 9234 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 9854 82894
rect 9234 82574 9854 82658
rect 9234 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 9854 82574
rect 9234 46894 9854 82338
rect 9234 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 9854 46894
rect 9234 46574 9854 46658
rect 9234 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 9854 46574
rect 9234 10894 9854 46338
rect 9234 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 9854 10894
rect 9234 10574 9854 10658
rect 9234 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 9854 10574
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect 9234 -4186 9854 10338
rect 9234 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 9854 -4186
rect 9234 -4506 9854 -4422
rect 9234 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 9854 -4506
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect 9234 -5734 9854 -4742
rect 12954 698614 13574 710042
rect 30954 711558 31574 711590
rect 30954 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 31574 711558
rect 30954 711238 31574 711322
rect 30954 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 31574 711238
rect 27234 709638 27854 709670
rect 27234 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 27854 709638
rect 27234 709318 27854 709402
rect 27234 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 27854 709318
rect 23514 707718 24134 707750
rect 23514 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 24134 707718
rect 23514 707398 24134 707482
rect 23514 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 24134 707398
rect 12954 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 13574 698614
rect 12954 698294 13574 698378
rect 12954 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 13574 698294
rect 12954 662614 13574 698058
rect 12954 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 13574 662614
rect 12954 662294 13574 662378
rect 12954 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 13574 662294
rect 12954 626614 13574 662058
rect 12954 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 13574 626614
rect 12954 626294 13574 626378
rect 12954 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 13574 626294
rect 12954 590614 13574 626058
rect 12954 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 13574 590614
rect 12954 590294 13574 590378
rect 12954 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 13574 590294
rect 12954 554614 13574 590058
rect 12954 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 13574 554614
rect 12954 554294 13574 554378
rect 12954 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 13574 554294
rect 12954 518614 13574 554058
rect 12954 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 13574 518614
rect 12954 518294 13574 518378
rect 12954 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 13574 518294
rect 12954 482614 13574 518058
rect 12954 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 13574 482614
rect 12954 482294 13574 482378
rect 12954 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 13574 482294
rect 12954 446614 13574 482058
rect 12954 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 13574 446614
rect 12954 446294 13574 446378
rect 12954 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 13574 446294
rect 12954 410614 13574 446058
rect 12954 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 13574 410614
rect 12954 410294 13574 410378
rect 12954 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 13574 410294
rect 12954 374614 13574 410058
rect 12954 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 13574 374614
rect 12954 374294 13574 374378
rect 12954 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 13574 374294
rect 12954 338614 13574 374058
rect 12954 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 13574 338614
rect 12954 338294 13574 338378
rect 12954 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 13574 338294
rect 12954 302614 13574 338058
rect 12954 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 13574 302614
rect 12954 302294 13574 302378
rect 12954 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 13574 302294
rect 12954 266614 13574 302058
rect 12954 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 13574 266614
rect 12954 266294 13574 266378
rect 12954 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 13574 266294
rect 12954 230614 13574 266058
rect 12954 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 13574 230614
rect 12954 230294 13574 230378
rect 12954 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 13574 230294
rect 12954 194614 13574 230058
rect 12954 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 13574 194614
rect 12954 194294 13574 194378
rect 12954 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 13574 194294
rect 12954 158614 13574 194058
rect 12954 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 13574 158614
rect 12954 158294 13574 158378
rect 12954 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 13574 158294
rect 12954 122614 13574 158058
rect 12954 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 13574 122614
rect 12954 122294 13574 122378
rect 12954 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 13574 122294
rect 12954 86614 13574 122058
rect 12954 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 13574 86614
rect 12954 86294 13574 86378
rect 12954 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 13574 86294
rect 12954 50614 13574 86058
rect 12954 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 13574 50614
rect 12954 50294 13574 50378
rect 12954 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 13574 50294
rect 12954 14614 13574 50058
rect 12954 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 13574 14614
rect 12954 14294 13574 14378
rect 12954 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 13574 14294
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect 12954 -6106 13574 14058
rect 19794 705798 20414 705830
rect 19794 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 20414 705798
rect 19794 705478 20414 705562
rect 19794 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 20414 705478
rect 19794 669454 20414 705242
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -1306 20414 20898
rect 19794 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 20414 -1306
rect 19794 -1626 20414 -1542
rect 19794 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 20414 -1626
rect 19794 -1894 20414 -1862
rect 23514 673174 24134 707162
rect 23514 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 24134 673174
rect 23514 672854 24134 672938
rect 23514 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 24134 672854
rect 23514 637174 24134 672618
rect 23514 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 24134 637174
rect 23514 636854 24134 636938
rect 23514 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 24134 636854
rect 23514 601174 24134 636618
rect 23514 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 24134 601174
rect 23514 600854 24134 600938
rect 23514 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 24134 600854
rect 23514 565174 24134 600618
rect 23514 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 24134 565174
rect 23514 564854 24134 564938
rect 23514 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 24134 564854
rect 23514 529174 24134 564618
rect 23514 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 24134 529174
rect 23514 528854 24134 528938
rect 23514 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 24134 528854
rect 23514 493174 24134 528618
rect 23514 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 24134 493174
rect 23514 492854 24134 492938
rect 23514 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 24134 492854
rect 23514 457174 24134 492618
rect 23514 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 24134 457174
rect 23514 456854 24134 456938
rect 23514 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 24134 456854
rect 23514 421174 24134 456618
rect 23514 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 24134 421174
rect 23514 420854 24134 420938
rect 23514 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 24134 420854
rect 23514 385174 24134 420618
rect 23514 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 24134 385174
rect 23514 384854 24134 384938
rect 23514 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 24134 384854
rect 23514 349174 24134 384618
rect 23514 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 24134 349174
rect 23514 348854 24134 348938
rect 23514 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 24134 348854
rect 23514 313174 24134 348618
rect 23514 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 24134 313174
rect 23514 312854 24134 312938
rect 23514 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 24134 312854
rect 23514 277174 24134 312618
rect 23514 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 24134 277174
rect 23514 276854 24134 276938
rect 23514 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 24134 276854
rect 23514 241174 24134 276618
rect 23514 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 24134 241174
rect 23514 240854 24134 240938
rect 23514 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 24134 240854
rect 23514 205174 24134 240618
rect 23514 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 24134 205174
rect 23514 204854 24134 204938
rect 23514 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 24134 204854
rect 23514 169174 24134 204618
rect 23514 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 24134 169174
rect 23514 168854 24134 168938
rect 23514 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 24134 168854
rect 23514 133174 24134 168618
rect 23514 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 24134 133174
rect 23514 132854 24134 132938
rect 23514 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 24134 132854
rect 23514 97174 24134 132618
rect 23514 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 24134 97174
rect 23514 96854 24134 96938
rect 23514 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 24134 96854
rect 23514 61174 24134 96618
rect 23514 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 24134 61174
rect 23514 60854 24134 60938
rect 23514 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 24134 60854
rect 23514 25174 24134 60618
rect 23514 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 24134 25174
rect 23514 24854 24134 24938
rect 23514 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 24134 24854
rect 23514 -3226 24134 24618
rect 23514 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 24134 -3226
rect 23514 -3546 24134 -3462
rect 23514 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 24134 -3546
rect 23514 -3814 24134 -3782
rect 27234 676894 27854 709082
rect 27234 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 27854 676894
rect 27234 676574 27854 676658
rect 27234 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 27854 676574
rect 27234 640894 27854 676338
rect 27234 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 27854 640894
rect 27234 640574 27854 640658
rect 27234 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 27854 640574
rect 27234 604894 27854 640338
rect 27234 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 27854 604894
rect 27234 604574 27854 604658
rect 27234 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 27854 604574
rect 27234 568894 27854 604338
rect 27234 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 27854 568894
rect 27234 568574 27854 568658
rect 27234 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 27854 568574
rect 27234 532894 27854 568338
rect 27234 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 27854 532894
rect 27234 532574 27854 532658
rect 27234 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 27854 532574
rect 27234 496894 27854 532338
rect 27234 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 27854 496894
rect 27234 496574 27854 496658
rect 27234 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 27854 496574
rect 27234 460894 27854 496338
rect 27234 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 27854 460894
rect 27234 460574 27854 460658
rect 27234 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 27854 460574
rect 27234 424894 27854 460338
rect 27234 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 27854 424894
rect 27234 424574 27854 424658
rect 27234 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 27854 424574
rect 27234 388894 27854 424338
rect 27234 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 27854 388894
rect 27234 388574 27854 388658
rect 27234 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 27854 388574
rect 27234 352894 27854 388338
rect 27234 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 27854 352894
rect 27234 352574 27854 352658
rect 27234 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 27854 352574
rect 27234 316894 27854 352338
rect 27234 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 27854 316894
rect 27234 316574 27854 316658
rect 27234 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 27854 316574
rect 27234 280894 27854 316338
rect 27234 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 27854 280894
rect 27234 280574 27854 280658
rect 27234 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 27854 280574
rect 27234 244894 27854 280338
rect 27234 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 27854 244894
rect 27234 244574 27854 244658
rect 27234 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 27854 244574
rect 27234 208894 27854 244338
rect 27234 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 27854 208894
rect 27234 208574 27854 208658
rect 27234 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 27854 208574
rect 27234 172894 27854 208338
rect 27234 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 27854 172894
rect 27234 172574 27854 172658
rect 27234 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 27854 172574
rect 27234 136894 27854 172338
rect 27234 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 27854 136894
rect 27234 136574 27854 136658
rect 27234 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 27854 136574
rect 27234 100894 27854 136338
rect 27234 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 27854 100894
rect 27234 100574 27854 100658
rect 27234 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 27854 100574
rect 27234 64894 27854 100338
rect 27234 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 27854 64894
rect 27234 64574 27854 64658
rect 27234 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 27854 64574
rect 27234 28894 27854 64338
rect 27234 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 27854 28894
rect 27234 28574 27854 28658
rect 27234 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 27854 28574
rect 27234 -5146 27854 28338
rect 27234 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 27854 -5146
rect 27234 -5466 27854 -5382
rect 27234 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 27854 -5466
rect 27234 -5734 27854 -5702
rect 30954 680614 31574 711002
rect 48954 710598 49574 711590
rect 48954 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 49574 710598
rect 48954 710278 49574 710362
rect 48954 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 49574 710278
rect 45234 708678 45854 709670
rect 45234 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 45854 708678
rect 45234 708358 45854 708442
rect 45234 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 45854 708358
rect 41514 706758 42134 707750
rect 41514 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 42134 706758
rect 41514 706438 42134 706522
rect 41514 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 42134 706438
rect 30954 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 31574 680614
rect 30954 680294 31574 680378
rect 30954 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 31574 680294
rect 30954 644614 31574 680058
rect 30954 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 31574 644614
rect 30954 644294 31574 644378
rect 30954 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 31574 644294
rect 30954 608614 31574 644058
rect 30954 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 31574 608614
rect 30954 608294 31574 608378
rect 30954 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 31574 608294
rect 30954 572614 31574 608058
rect 30954 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 31574 572614
rect 30954 572294 31574 572378
rect 30954 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 31574 572294
rect 30954 536614 31574 572058
rect 30954 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 31574 536614
rect 30954 536294 31574 536378
rect 30954 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 31574 536294
rect 30954 500614 31574 536058
rect 30954 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 31574 500614
rect 30954 500294 31574 500378
rect 30954 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 31574 500294
rect 30954 464614 31574 500058
rect 30954 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 31574 464614
rect 30954 464294 31574 464378
rect 30954 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 31574 464294
rect 30954 428614 31574 464058
rect 30954 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 31574 428614
rect 30954 428294 31574 428378
rect 30954 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 31574 428294
rect 30954 392614 31574 428058
rect 30954 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 31574 392614
rect 30954 392294 31574 392378
rect 30954 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 31574 392294
rect 30954 356614 31574 392058
rect 30954 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 31574 356614
rect 30954 356294 31574 356378
rect 30954 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 31574 356294
rect 30954 320614 31574 356058
rect 30954 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 31574 320614
rect 30954 320294 31574 320378
rect 30954 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 31574 320294
rect 30954 284614 31574 320058
rect 30954 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 31574 284614
rect 30954 284294 31574 284378
rect 30954 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 31574 284294
rect 30954 248614 31574 284058
rect 30954 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 31574 248614
rect 30954 248294 31574 248378
rect 30954 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 31574 248294
rect 30954 212614 31574 248058
rect 30954 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 31574 212614
rect 30954 212294 31574 212378
rect 30954 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 31574 212294
rect 30954 176614 31574 212058
rect 30954 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 31574 176614
rect 30954 176294 31574 176378
rect 30954 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 31574 176294
rect 30954 140614 31574 176058
rect 30954 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 31574 140614
rect 30954 140294 31574 140378
rect 30954 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 31574 140294
rect 30954 104614 31574 140058
rect 30954 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 31574 104614
rect 30954 104294 31574 104378
rect 30954 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 31574 104294
rect 30954 68614 31574 104058
rect 30954 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 31574 68614
rect 30954 68294 31574 68378
rect 30954 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 31574 68294
rect 30954 32614 31574 68058
rect 30954 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 31574 32614
rect 30954 32294 31574 32378
rect 30954 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 31574 32294
rect 12954 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 13574 -6106
rect 12954 -6426 13574 -6342
rect 12954 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 13574 -6426
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 12954 -7654 13574 -6662
rect 30954 -7066 31574 32058
rect 37794 704838 38414 705830
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -1894 38414 -902
rect 41514 691174 42134 706202
rect 41514 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 42134 691174
rect 41514 690854 42134 690938
rect 41514 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 42134 690854
rect 41514 655174 42134 690618
rect 41514 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 42134 655174
rect 41514 654854 42134 654938
rect 41514 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 42134 654854
rect 41514 619174 42134 654618
rect 41514 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 42134 619174
rect 41514 618854 42134 618938
rect 41514 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 42134 618854
rect 41514 583174 42134 618618
rect 41514 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 42134 583174
rect 41514 582854 42134 582938
rect 41514 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 42134 582854
rect 41514 547174 42134 582618
rect 41514 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 42134 547174
rect 41514 546854 42134 546938
rect 41514 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 42134 546854
rect 41514 511174 42134 546618
rect 41514 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 42134 511174
rect 41514 510854 42134 510938
rect 41514 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 42134 510854
rect 41514 475174 42134 510618
rect 41514 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 42134 475174
rect 41514 474854 42134 474938
rect 41514 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 42134 474854
rect 41514 439174 42134 474618
rect 41514 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 42134 439174
rect 41514 438854 42134 438938
rect 41514 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 42134 438854
rect 41514 403174 42134 438618
rect 41514 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 42134 403174
rect 41514 402854 42134 402938
rect 41514 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 42134 402854
rect 41514 367174 42134 402618
rect 41514 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 42134 367174
rect 41514 366854 42134 366938
rect 41514 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 42134 366854
rect 41514 331174 42134 366618
rect 41514 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 42134 331174
rect 41514 330854 42134 330938
rect 41514 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 42134 330854
rect 41514 295174 42134 330618
rect 41514 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 42134 295174
rect 41514 294854 42134 294938
rect 41514 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 42134 294854
rect 41514 259174 42134 294618
rect 41514 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 42134 259174
rect 41514 258854 42134 258938
rect 41514 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 42134 258854
rect 41514 223174 42134 258618
rect 41514 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 42134 223174
rect 41514 222854 42134 222938
rect 41514 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 42134 222854
rect 41514 187174 42134 222618
rect 41514 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 42134 187174
rect 41514 186854 42134 186938
rect 41514 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 42134 186854
rect 41514 151174 42134 186618
rect 41514 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 42134 151174
rect 41514 150854 42134 150938
rect 41514 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 42134 150854
rect 41514 115174 42134 150618
rect 41514 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 42134 115174
rect 41514 114854 42134 114938
rect 41514 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 42134 114854
rect 41514 79174 42134 114618
rect 41514 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 42134 79174
rect 41514 78854 42134 78938
rect 41514 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 42134 78854
rect 41514 43174 42134 78618
rect 41514 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 42134 43174
rect 41514 42854 42134 42938
rect 41514 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 42134 42854
rect 41514 7174 42134 42618
rect 41514 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 42134 7174
rect 41514 6854 42134 6938
rect 41514 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 42134 6854
rect 41514 -2266 42134 6618
rect 41514 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 42134 -2266
rect 41514 -2586 42134 -2502
rect 41514 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 42134 -2586
rect 41514 -3814 42134 -2822
rect 45234 694894 45854 708122
rect 45234 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 45854 694894
rect 45234 694574 45854 694658
rect 45234 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 45854 694574
rect 45234 658894 45854 694338
rect 45234 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 45854 658894
rect 45234 658574 45854 658658
rect 45234 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 45854 658574
rect 45234 622894 45854 658338
rect 45234 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 45854 622894
rect 45234 622574 45854 622658
rect 45234 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 45854 622574
rect 45234 586894 45854 622338
rect 45234 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 45854 586894
rect 45234 586574 45854 586658
rect 45234 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 45854 586574
rect 45234 550894 45854 586338
rect 45234 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 45854 550894
rect 45234 550574 45854 550658
rect 45234 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 45854 550574
rect 45234 514894 45854 550338
rect 45234 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 45854 514894
rect 45234 514574 45854 514658
rect 45234 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 45854 514574
rect 45234 478894 45854 514338
rect 45234 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 45854 478894
rect 45234 478574 45854 478658
rect 45234 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 45854 478574
rect 45234 442894 45854 478338
rect 45234 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 45854 442894
rect 45234 442574 45854 442658
rect 45234 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 45854 442574
rect 45234 406894 45854 442338
rect 45234 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 45854 406894
rect 45234 406574 45854 406658
rect 45234 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 45854 406574
rect 45234 370894 45854 406338
rect 45234 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 45854 370894
rect 45234 370574 45854 370658
rect 45234 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 45854 370574
rect 45234 334894 45854 370338
rect 45234 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 45854 334894
rect 45234 334574 45854 334658
rect 45234 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 45854 334574
rect 45234 298894 45854 334338
rect 45234 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 45854 298894
rect 45234 298574 45854 298658
rect 45234 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 45854 298574
rect 45234 262894 45854 298338
rect 45234 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 45854 262894
rect 45234 262574 45854 262658
rect 45234 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 45854 262574
rect 45234 226894 45854 262338
rect 45234 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 45854 226894
rect 45234 226574 45854 226658
rect 45234 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 45854 226574
rect 45234 190894 45854 226338
rect 45234 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 45854 190894
rect 45234 190574 45854 190658
rect 45234 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 45854 190574
rect 45234 154894 45854 190338
rect 45234 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 45854 154894
rect 45234 154574 45854 154658
rect 45234 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 45854 154574
rect 45234 118894 45854 154338
rect 45234 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 45854 118894
rect 45234 118574 45854 118658
rect 45234 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 45854 118574
rect 45234 82894 45854 118338
rect 45234 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 45854 82894
rect 45234 82574 45854 82658
rect 45234 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 45854 82574
rect 45234 46894 45854 82338
rect 45234 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 45854 46894
rect 45234 46574 45854 46658
rect 45234 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 45854 46574
rect 45234 10894 45854 46338
rect 45234 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 45854 10894
rect 45234 10574 45854 10658
rect 45234 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 45854 10574
rect 45234 -4186 45854 10338
rect 45234 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 45854 -4186
rect 45234 -4506 45854 -4422
rect 45234 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 45854 -4506
rect 45234 -5734 45854 -4742
rect 48954 698614 49574 710042
rect 66954 711558 67574 711590
rect 66954 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 67574 711558
rect 66954 711238 67574 711322
rect 66954 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 67574 711238
rect 63234 709638 63854 709670
rect 63234 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 63854 709638
rect 63234 709318 63854 709402
rect 63234 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 63854 709318
rect 59514 707718 60134 707750
rect 59514 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 60134 707718
rect 59514 707398 60134 707482
rect 59514 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 60134 707398
rect 48954 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 49574 698614
rect 48954 698294 49574 698378
rect 48954 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 49574 698294
rect 48954 662614 49574 698058
rect 48954 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 49574 662614
rect 48954 662294 49574 662378
rect 48954 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 49574 662294
rect 48954 626614 49574 662058
rect 48954 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 49574 626614
rect 48954 626294 49574 626378
rect 48954 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 49574 626294
rect 48954 590614 49574 626058
rect 48954 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 49574 590614
rect 48954 590294 49574 590378
rect 48954 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 49574 590294
rect 48954 554614 49574 590058
rect 48954 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 49574 554614
rect 48954 554294 49574 554378
rect 48954 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 49574 554294
rect 48954 518614 49574 554058
rect 48954 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 49574 518614
rect 48954 518294 49574 518378
rect 48954 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 49574 518294
rect 48954 482614 49574 518058
rect 48954 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 49574 482614
rect 48954 482294 49574 482378
rect 48954 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 49574 482294
rect 48954 446614 49574 482058
rect 48954 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 49574 446614
rect 48954 446294 49574 446378
rect 48954 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 49574 446294
rect 48954 410614 49574 446058
rect 48954 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 49574 410614
rect 48954 410294 49574 410378
rect 48954 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 49574 410294
rect 48954 374614 49574 410058
rect 48954 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 49574 374614
rect 48954 374294 49574 374378
rect 48954 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 49574 374294
rect 48954 338614 49574 374058
rect 48954 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 49574 338614
rect 48954 338294 49574 338378
rect 48954 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 49574 338294
rect 48954 302614 49574 338058
rect 48954 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 49574 302614
rect 48954 302294 49574 302378
rect 48954 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 49574 302294
rect 48954 266614 49574 302058
rect 48954 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 49574 266614
rect 48954 266294 49574 266378
rect 48954 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 49574 266294
rect 48954 230614 49574 266058
rect 48954 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 49574 230614
rect 48954 230294 49574 230378
rect 48954 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 49574 230294
rect 48954 194614 49574 230058
rect 48954 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 49574 194614
rect 48954 194294 49574 194378
rect 48954 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 49574 194294
rect 48954 158614 49574 194058
rect 48954 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 49574 158614
rect 48954 158294 49574 158378
rect 48954 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 49574 158294
rect 48954 122614 49574 158058
rect 48954 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 49574 122614
rect 48954 122294 49574 122378
rect 48954 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 49574 122294
rect 48954 86614 49574 122058
rect 48954 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 49574 86614
rect 48954 86294 49574 86378
rect 48954 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 49574 86294
rect 48954 50614 49574 86058
rect 48954 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 49574 50614
rect 48954 50294 49574 50378
rect 48954 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 49574 50294
rect 48954 14614 49574 50058
rect 48954 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 49574 14614
rect 48954 14294 49574 14378
rect 48954 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 49574 14294
rect 30954 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 31574 -7066
rect 30954 -7386 31574 -7302
rect 30954 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 31574 -7386
rect 30954 -7654 31574 -7622
rect 48954 -6106 49574 14058
rect 55794 705798 56414 705830
rect 55794 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 56414 705798
rect 55794 705478 56414 705562
rect 55794 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 56414 705478
rect 55794 669454 56414 705242
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55794 525454 56414 560898
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55794 453454 56414 488898
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55794 417454 56414 452898
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55794 381454 56414 416898
rect 55794 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 56414 381454
rect 55794 381134 56414 381218
rect 55794 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 56414 381134
rect 55794 345454 56414 380898
rect 55794 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 56414 345454
rect 55794 345134 56414 345218
rect 55794 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 56414 345134
rect 55794 309454 56414 344898
rect 55794 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 56414 309454
rect 55794 309134 56414 309218
rect 55794 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 56414 309134
rect 55794 273454 56414 308898
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 55794 237454 56414 272898
rect 59514 673174 60134 707162
rect 59514 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 60134 673174
rect 59514 672854 60134 672938
rect 59514 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 60134 672854
rect 59514 637174 60134 672618
rect 59514 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 60134 637174
rect 59514 636854 60134 636938
rect 59514 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 60134 636854
rect 59514 601174 60134 636618
rect 59514 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 60134 601174
rect 59514 600854 60134 600938
rect 59514 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 60134 600854
rect 59514 565174 60134 600618
rect 59514 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 60134 565174
rect 59514 564854 60134 564938
rect 59514 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 60134 564854
rect 59514 529174 60134 564618
rect 59514 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 60134 529174
rect 59514 528854 60134 528938
rect 59514 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 60134 528854
rect 59514 493174 60134 528618
rect 59514 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 60134 493174
rect 59514 492854 60134 492938
rect 59514 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 60134 492854
rect 59514 457174 60134 492618
rect 59514 456938 59546 457174
rect 59782 456938 59866 457174
rect 60102 456938 60134 457174
rect 59514 456854 60134 456938
rect 59514 456618 59546 456854
rect 59782 456618 59866 456854
rect 60102 456618 60134 456854
rect 59514 421174 60134 456618
rect 59514 420938 59546 421174
rect 59782 420938 59866 421174
rect 60102 420938 60134 421174
rect 59514 420854 60134 420938
rect 59514 420618 59546 420854
rect 59782 420618 59866 420854
rect 60102 420618 60134 420854
rect 59514 385174 60134 420618
rect 59514 384938 59546 385174
rect 59782 384938 59866 385174
rect 60102 384938 60134 385174
rect 59514 384854 60134 384938
rect 59514 384618 59546 384854
rect 59782 384618 59866 384854
rect 60102 384618 60134 384854
rect 59514 349174 60134 384618
rect 59514 348938 59546 349174
rect 59782 348938 59866 349174
rect 60102 348938 60134 349174
rect 59514 348854 60134 348938
rect 59514 348618 59546 348854
rect 59782 348618 59866 348854
rect 60102 348618 60134 348854
rect 59514 313174 60134 348618
rect 59514 312938 59546 313174
rect 59782 312938 59866 313174
rect 60102 312938 60134 313174
rect 59514 312854 60134 312938
rect 59514 312618 59546 312854
rect 59782 312618 59866 312854
rect 60102 312618 60134 312854
rect 59514 277174 60134 312618
rect 63234 676894 63854 709082
rect 63234 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 63854 676894
rect 63234 676574 63854 676658
rect 63234 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 63854 676574
rect 63234 640894 63854 676338
rect 63234 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 63854 640894
rect 63234 640574 63854 640658
rect 63234 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 63854 640574
rect 63234 604894 63854 640338
rect 63234 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 63854 604894
rect 63234 604574 63854 604658
rect 63234 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 63854 604574
rect 63234 568894 63854 604338
rect 66954 680614 67574 711002
rect 84954 710598 85574 711590
rect 84954 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 85574 710598
rect 84954 710278 85574 710362
rect 84954 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 85574 710278
rect 81234 708678 81854 709670
rect 81234 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 81854 708678
rect 81234 708358 81854 708442
rect 81234 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 81854 708358
rect 77514 706758 78134 707750
rect 77514 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 78134 706758
rect 77514 706438 78134 706522
rect 77514 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 78134 706438
rect 73794 704838 74414 705830
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 69611 702540 69677 702541
rect 69611 702476 69612 702540
rect 69676 702476 69677 702540
rect 69611 702475 69677 702476
rect 66954 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 67574 680614
rect 66954 680294 67574 680378
rect 66954 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 67574 680294
rect 66954 644614 67574 680058
rect 66954 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 67574 644614
rect 66954 644294 67574 644378
rect 66954 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 67574 644294
rect 66954 608614 67574 644058
rect 66954 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 67574 608614
rect 66954 608294 67574 608378
rect 66954 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 67574 608294
rect 66954 591166 67574 608058
rect 66115 590748 66181 590749
rect 66115 590684 66116 590748
rect 66180 590684 66181 590748
rect 66115 590683 66181 590684
rect 63234 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 63854 568894
rect 63234 568574 63854 568658
rect 63234 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 63854 568574
rect 63234 532894 63854 568338
rect 63234 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 63854 532894
rect 63234 532574 63854 532658
rect 63234 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 63854 532574
rect 63234 496894 63854 532338
rect 63234 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 63854 496894
rect 63234 496574 63854 496658
rect 63234 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 63854 496574
rect 63234 460894 63854 496338
rect 63234 460658 63266 460894
rect 63502 460658 63586 460894
rect 63822 460658 63854 460894
rect 63234 460574 63854 460658
rect 63234 460338 63266 460574
rect 63502 460338 63586 460574
rect 63822 460338 63854 460574
rect 63234 424894 63854 460338
rect 66118 450533 66178 590683
rect 69614 586530 69674 702475
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73794 591166 74414 614898
rect 77514 691174 78134 706202
rect 77514 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 78134 691174
rect 77514 690854 78134 690938
rect 77514 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 78134 690854
rect 77514 655174 78134 690618
rect 77514 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 78134 655174
rect 77514 654854 78134 654938
rect 77514 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 78134 654854
rect 77514 619174 78134 654618
rect 77514 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 78134 619174
rect 77514 618854 78134 618938
rect 77514 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 78134 618854
rect 77514 591166 78134 618618
rect 81234 694894 81854 708122
rect 81234 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 81854 694894
rect 81234 694574 81854 694658
rect 81234 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 81854 694574
rect 81234 658894 81854 694338
rect 81234 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 81854 658894
rect 81234 658574 81854 658658
rect 81234 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 81854 658574
rect 81234 622894 81854 658338
rect 81234 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 81854 622894
rect 81234 622574 81854 622658
rect 81234 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 81854 622574
rect 81234 591166 81854 622338
rect 84954 698614 85574 710042
rect 102954 711558 103574 711590
rect 102954 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 103574 711558
rect 102954 711238 103574 711322
rect 102954 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 103574 711238
rect 99234 709638 99854 709670
rect 99234 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 99854 709638
rect 99234 709318 99854 709402
rect 99234 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 99854 709318
rect 95514 707718 96134 707750
rect 95514 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 96134 707718
rect 95514 707398 96134 707482
rect 95514 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 96134 707398
rect 84954 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 85574 698614
rect 84954 698294 85574 698378
rect 84954 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 85574 698294
rect 84954 662614 85574 698058
rect 84954 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 85574 662614
rect 84954 662294 85574 662378
rect 84954 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 85574 662294
rect 84954 626614 85574 662058
rect 84954 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 85574 626614
rect 84954 626294 85574 626378
rect 84954 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 85574 626294
rect 84954 591166 85574 626058
rect 91794 705798 92414 705830
rect 91794 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 92414 705798
rect 91794 705478 92414 705562
rect 91794 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 92414 705478
rect 91794 669454 92414 705242
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 633454 92414 668898
rect 91794 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 92414 633454
rect 91794 633134 92414 633218
rect 91794 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 92414 633134
rect 91794 597454 92414 632898
rect 91794 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 92414 597454
rect 91794 597134 92414 597218
rect 91794 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 92414 597134
rect 88195 588572 88261 588573
rect 88195 588508 88196 588572
rect 88260 588508 88261 588572
rect 88195 588507 88261 588508
rect 69430 586470 69674 586530
rect 69430 582317 69490 586470
rect 88198 585717 88258 588507
rect 88195 585716 88261 585717
rect 88195 585652 88196 585716
rect 88260 585652 88261 585716
rect 88195 585651 88261 585652
rect 69427 582316 69493 582317
rect 69427 582252 69428 582316
rect 69492 582252 69493 582316
rect 69427 582251 69493 582252
rect 72679 579454 72999 579486
rect 72679 579218 72721 579454
rect 72957 579218 72999 579454
rect 72679 579134 72999 579218
rect 72679 578898 72721 579134
rect 72957 578898 72999 579134
rect 72679 578866 72999 578898
rect 78609 579454 78929 579486
rect 78609 579218 78651 579454
rect 78887 579218 78929 579454
rect 78609 579134 78929 579218
rect 78609 578898 78651 579134
rect 78887 578898 78929 579134
rect 78609 578866 78929 578898
rect 84540 579454 84860 579486
rect 84540 579218 84582 579454
rect 84818 579218 84860 579454
rect 84540 579134 84860 579218
rect 84540 578898 84582 579134
rect 84818 578898 84860 579134
rect 84540 578866 84860 578898
rect 91139 578100 91205 578101
rect 91139 578036 91140 578100
rect 91204 578036 91205 578100
rect 91139 578035 91205 578036
rect 75644 561454 75964 561486
rect 75644 561218 75686 561454
rect 75922 561218 75964 561454
rect 75644 561134 75964 561218
rect 75644 560898 75686 561134
rect 75922 560898 75964 561134
rect 75644 560866 75964 560898
rect 81575 561454 81895 561486
rect 81575 561218 81617 561454
rect 81853 561218 81895 561454
rect 81575 561134 81895 561218
rect 81575 560898 81617 561134
rect 81853 560898 81895 561134
rect 81575 560866 81895 560898
rect 67403 556884 67469 556885
rect 67403 556820 67404 556884
rect 67468 556820 67469 556884
rect 67403 556819 67469 556820
rect 66667 551444 66733 551445
rect 66667 551380 66668 551444
rect 66732 551380 66733 551444
rect 66667 551379 66733 551380
rect 66670 528570 66730 551379
rect 67406 537437 67466 556819
rect 72679 543454 72999 543486
rect 72679 543218 72721 543454
rect 72957 543218 72999 543454
rect 72679 543134 72999 543218
rect 72679 542898 72721 543134
rect 72957 542898 72999 543134
rect 72679 542866 72999 542898
rect 78609 543454 78929 543486
rect 78609 543218 78651 543454
rect 78887 543218 78929 543454
rect 78609 543134 78929 543218
rect 78609 542898 78651 543134
rect 78887 542898 78929 543134
rect 78609 542866 78929 542898
rect 84540 543454 84860 543486
rect 84540 543218 84582 543454
rect 84818 543218 84860 543454
rect 84540 543134 84860 543218
rect 84540 542898 84582 543134
rect 84818 542898 84860 543134
rect 84540 542866 84860 542898
rect 91142 542333 91202 578035
rect 91794 561454 92414 596898
rect 91794 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 92414 561454
rect 91794 561134 92414 561218
rect 91794 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 92414 561134
rect 69427 542332 69493 542333
rect 69427 542268 69428 542332
rect 69492 542268 69493 542332
rect 69427 542267 69493 542268
rect 91139 542332 91205 542333
rect 91139 542268 91140 542332
rect 91204 542268 91205 542332
rect 91139 542267 91205 542268
rect 69430 538230 69490 542267
rect 69430 538170 69858 538230
rect 67403 537436 67469 537437
rect 67403 537372 67404 537436
rect 67468 537372 67469 537436
rect 67403 537371 67469 537372
rect 66486 528510 66730 528570
rect 66954 536614 67574 537166
rect 66954 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 67574 536614
rect 66954 536294 67574 536378
rect 66954 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 67574 536294
rect 66486 522885 66546 528510
rect 66667 523020 66733 523021
rect 66667 522956 66668 523020
rect 66732 522956 66733 523020
rect 66667 522955 66733 522956
rect 66483 522884 66549 522885
rect 66483 522820 66484 522884
rect 66548 522820 66549 522884
rect 66483 522819 66549 522820
rect 66115 450532 66181 450533
rect 66115 450468 66116 450532
rect 66180 450468 66181 450532
rect 66115 450467 66181 450468
rect 63234 424658 63266 424894
rect 63502 424658 63586 424894
rect 63822 424658 63854 424894
rect 63234 424574 63854 424658
rect 63234 424338 63266 424574
rect 63502 424338 63586 424574
rect 63822 424338 63854 424574
rect 63234 388894 63854 424338
rect 66670 419661 66730 522955
rect 66954 500614 67574 536058
rect 69611 535532 69677 535533
rect 69611 535468 69612 535532
rect 69676 535468 69677 535532
rect 69611 535467 69677 535468
rect 66954 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 67574 500614
rect 66954 500294 67574 500378
rect 66954 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 67574 500294
rect 66954 464614 67574 500058
rect 66954 464378 66986 464614
rect 67222 464378 67306 464614
rect 67542 464378 67574 464614
rect 66954 464294 67574 464378
rect 66954 464058 66986 464294
rect 67222 464058 67306 464294
rect 67542 464058 67574 464294
rect 66954 446407 67574 464058
rect 67771 442236 67837 442237
rect 67771 442172 67772 442236
rect 67836 442172 67837 442236
rect 67771 442171 67837 442172
rect 66667 419660 66733 419661
rect 66667 419596 66668 419660
rect 66732 419596 66733 419660
rect 66667 419595 66733 419596
rect 63234 388658 63266 388894
rect 63502 388658 63586 388894
rect 63822 388658 63854 388894
rect 63234 388574 63854 388658
rect 63234 388338 63266 388574
rect 63502 388338 63586 388574
rect 63822 388338 63854 388574
rect 63234 352894 63854 388338
rect 63234 352658 63266 352894
rect 63502 352658 63586 352894
rect 63822 352658 63854 352894
rect 63234 352574 63854 352658
rect 63234 352338 63266 352574
rect 63502 352338 63586 352574
rect 63822 352338 63854 352574
rect 63234 316894 63854 352338
rect 66954 356614 67574 388356
rect 66954 356378 66986 356614
rect 67222 356378 67306 356614
rect 67542 356378 67574 356614
rect 66954 356294 67574 356378
rect 66954 356058 66986 356294
rect 67222 356058 67306 356294
rect 67542 356058 67574 356294
rect 66667 347036 66733 347037
rect 66667 346972 66668 347036
rect 66732 346972 66733 347036
rect 66667 346971 66733 346972
rect 66115 337380 66181 337381
rect 66115 337316 66116 337380
rect 66180 337316 66181 337380
rect 66115 337315 66181 337316
rect 66118 325685 66178 337315
rect 66115 325684 66181 325685
rect 66115 325620 66116 325684
rect 66180 325620 66181 325684
rect 66115 325619 66181 325620
rect 63234 316658 63266 316894
rect 63502 316658 63586 316894
rect 63822 316658 63854 316894
rect 63234 316574 63854 316658
rect 63234 316338 63266 316574
rect 63502 316338 63586 316574
rect 63822 316338 63854 316574
rect 61883 284340 61949 284341
rect 61883 284276 61884 284340
rect 61948 284276 61949 284340
rect 61883 284275 61949 284276
rect 59514 276938 59546 277174
rect 59782 276938 59866 277174
rect 60102 276938 60134 277174
rect 59514 276854 60134 276938
rect 59514 276618 59546 276854
rect 59782 276618 59866 276854
rect 60102 276618 60134 276854
rect 59123 247076 59189 247077
rect 59123 247012 59124 247076
rect 59188 247012 59189 247076
rect 59123 247011 59189 247012
rect 55794 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 56414 237454
rect 55794 237134 56414 237218
rect 55794 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 56414 237134
rect 55794 201454 56414 236898
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 55794 165454 56414 200898
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 129454 56414 164898
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55794 57454 56414 92898
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55794 21454 56414 56898
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -1306 56414 20898
rect 59126 15197 59186 247011
rect 59514 241174 60134 276618
rect 59514 240938 59546 241174
rect 59782 240938 59866 241174
rect 60102 240938 60134 241174
rect 59514 240854 60134 240938
rect 59514 240618 59546 240854
rect 59782 240618 59866 240854
rect 60102 240618 60134 240854
rect 59514 205174 60134 240618
rect 59514 204938 59546 205174
rect 59782 204938 59866 205174
rect 60102 204938 60134 205174
rect 59514 204854 60134 204938
rect 59514 204618 59546 204854
rect 59782 204618 59866 204854
rect 60102 204618 60134 204854
rect 59514 169174 60134 204618
rect 59514 168938 59546 169174
rect 59782 168938 59866 169174
rect 60102 168938 60134 169174
rect 59514 168854 60134 168938
rect 59514 168618 59546 168854
rect 59782 168618 59866 168854
rect 60102 168618 60134 168854
rect 59514 133174 60134 168618
rect 59514 132938 59546 133174
rect 59782 132938 59866 133174
rect 60102 132938 60134 133174
rect 59514 132854 60134 132938
rect 59514 132618 59546 132854
rect 59782 132618 59866 132854
rect 60102 132618 60134 132854
rect 59514 97174 60134 132618
rect 59514 96938 59546 97174
rect 59782 96938 59866 97174
rect 60102 96938 60134 97174
rect 59514 96854 60134 96938
rect 59514 96618 59546 96854
rect 59782 96618 59866 96854
rect 60102 96618 60134 96854
rect 59514 61174 60134 96618
rect 59514 60938 59546 61174
rect 59782 60938 59866 61174
rect 60102 60938 60134 61174
rect 59514 60854 60134 60938
rect 59514 60618 59546 60854
rect 59782 60618 59866 60854
rect 60102 60618 60134 60854
rect 59514 25174 60134 60618
rect 61886 33829 61946 284275
rect 63234 280894 63854 316338
rect 66670 287877 66730 346971
rect 66954 331592 67574 356058
rect 67774 348941 67834 442171
rect 69614 414030 69674 535467
rect 69798 456925 69858 538170
rect 71635 535532 71701 535533
rect 71635 535468 71636 535532
rect 71700 535468 71701 535532
rect 71635 535467 71701 535468
rect 72371 535532 72437 535533
rect 72371 535468 72372 535532
rect 72436 535468 72437 535532
rect 72371 535467 72437 535468
rect 69795 456924 69861 456925
rect 69795 456860 69796 456924
rect 69860 456860 69861 456924
rect 69795 456859 69861 456860
rect 69062 413970 69674 414030
rect 69062 404370 69122 413970
rect 69243 407828 69309 407829
rect 69243 407764 69244 407828
rect 69308 407826 69309 407828
rect 69308 407766 69490 407826
rect 69308 407764 69309 407766
rect 69243 407763 69309 407764
rect 69246 407149 69306 407763
rect 69243 407148 69309 407149
rect 69243 407084 69244 407148
rect 69308 407084 69309 407148
rect 69243 407083 69309 407084
rect 69430 404370 69490 407766
rect 69062 404310 69306 404370
rect 69430 404310 69858 404370
rect 69246 396130 69306 404310
rect 69798 404290 69858 404310
rect 69798 404230 70042 404290
rect 69982 396130 70042 404230
rect 69246 396070 69674 396130
rect 69614 390421 69674 396070
rect 69798 396070 70042 396130
rect 69611 390420 69677 390421
rect 69611 390356 69612 390420
rect 69676 390356 69677 390420
rect 69611 390355 69677 390356
rect 69798 367709 69858 396070
rect 71638 391370 71698 535467
rect 71638 391310 71882 391370
rect 71638 390690 71698 391310
rect 71822 391237 71882 391310
rect 71819 391236 71885 391237
rect 71819 391172 71820 391236
rect 71884 391172 71885 391236
rect 71819 391171 71885 391172
rect 71819 390692 71885 390693
rect 71819 390690 71820 390692
rect 71638 390630 71820 390690
rect 71819 390628 71820 390630
rect 71884 390628 71885 390692
rect 71819 390627 71885 390628
rect 72374 388381 72434 535467
rect 73794 507454 74414 537166
rect 73794 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 74414 507454
rect 73794 507134 74414 507218
rect 73794 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 74414 507134
rect 73794 471454 74414 506898
rect 73794 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 74414 471454
rect 73794 471134 74414 471218
rect 73794 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 74414 471134
rect 72739 448628 72805 448629
rect 72739 448564 72740 448628
rect 72804 448564 72805 448628
rect 72739 448563 72805 448564
rect 72371 388380 72437 388381
rect 72371 388316 72372 388380
rect 72436 388316 72437 388380
rect 72371 388315 72437 388316
rect 69795 367708 69861 367709
rect 69795 367644 69796 367708
rect 69860 367644 69861 367708
rect 69795 367643 69861 367644
rect 69611 356148 69677 356149
rect 69611 356084 69612 356148
rect 69676 356084 69677 356148
rect 69611 356083 69677 356084
rect 67955 349756 68021 349757
rect 67955 349692 67956 349756
rect 68020 349692 68021 349756
rect 67955 349691 68021 349692
rect 67771 348940 67837 348941
rect 67771 348876 67772 348940
rect 67836 348876 67837 348940
rect 67771 348875 67837 348876
rect 67771 338876 67837 338877
rect 67771 338812 67772 338876
rect 67836 338812 67837 338876
rect 67771 338811 67837 338812
rect 66667 287876 66733 287877
rect 66667 287812 66668 287876
rect 66732 287812 66733 287876
rect 66667 287811 66733 287812
rect 63234 280658 63266 280894
rect 63502 280658 63586 280894
rect 63822 280658 63854 280894
rect 63234 280574 63854 280658
rect 63234 280338 63266 280574
rect 63502 280338 63586 280574
rect 63822 280338 63854 280574
rect 63234 244894 63854 280338
rect 67774 280261 67834 338811
rect 67958 296309 68018 349691
rect 69614 335370 69674 356083
rect 69430 335310 69674 335370
rect 69430 328405 69490 335310
rect 69795 332620 69861 332621
rect 69795 332556 69796 332620
rect 69860 332556 69861 332620
rect 69795 332555 69861 332556
rect 69427 328404 69493 328405
rect 69427 328340 69428 328404
rect 69492 328340 69493 328404
rect 69427 328339 69493 328340
rect 69798 325710 69858 332555
rect 69430 325650 69858 325710
rect 69430 324053 69490 325650
rect 69427 324052 69493 324053
rect 69427 323988 69428 324052
rect 69492 323988 69493 324052
rect 69427 323987 69493 323988
rect 67955 296308 68021 296309
rect 67955 296244 67956 296308
rect 68020 296244 68021 296308
rect 67955 296243 68021 296244
rect 69427 287740 69493 287741
rect 69427 287676 69428 287740
rect 69492 287676 69493 287740
rect 69427 287675 69493 287676
rect 69430 287070 69490 287675
rect 69430 287010 69674 287070
rect 67771 280260 67837 280261
rect 67771 280196 67772 280260
rect 67836 280196 67837 280260
rect 67771 280195 67837 280196
rect 67955 277268 68021 277269
rect 67955 277204 67956 277268
rect 68020 277204 68021 277268
rect 67955 277203 68021 277204
rect 66115 273732 66181 273733
rect 66115 273668 66116 273732
rect 66180 273668 66181 273732
rect 66115 273667 66181 273668
rect 63234 244658 63266 244894
rect 63502 244658 63586 244894
rect 63822 244658 63854 244894
rect 63234 244574 63854 244658
rect 63234 244338 63266 244574
rect 63502 244338 63586 244574
rect 63822 244338 63854 244574
rect 63234 208894 63854 244338
rect 63234 208658 63266 208894
rect 63502 208658 63586 208894
rect 63822 208658 63854 208894
rect 63234 208574 63854 208658
rect 63234 208338 63266 208574
rect 63502 208338 63586 208574
rect 63822 208338 63854 208574
rect 63234 172894 63854 208338
rect 63234 172658 63266 172894
rect 63502 172658 63586 172894
rect 63822 172658 63854 172894
rect 63234 172574 63854 172658
rect 63234 172338 63266 172574
rect 63502 172338 63586 172574
rect 63822 172338 63854 172574
rect 63234 136894 63854 172338
rect 63234 136658 63266 136894
rect 63502 136658 63586 136894
rect 63822 136658 63854 136894
rect 63234 136574 63854 136658
rect 63234 136338 63266 136574
rect 63502 136338 63586 136574
rect 63822 136338 63854 136574
rect 63234 100894 63854 136338
rect 63234 100658 63266 100894
rect 63502 100658 63586 100894
rect 63822 100658 63854 100894
rect 63234 100574 63854 100658
rect 63234 100338 63266 100574
rect 63502 100338 63586 100574
rect 63822 100338 63854 100574
rect 63234 64894 63854 100338
rect 63234 64658 63266 64894
rect 63502 64658 63586 64894
rect 63822 64658 63854 64894
rect 63234 64574 63854 64658
rect 63234 64338 63266 64574
rect 63502 64338 63586 64574
rect 63822 64338 63854 64574
rect 61883 33828 61949 33829
rect 61883 33764 61884 33828
rect 61948 33764 61949 33828
rect 61883 33763 61949 33764
rect 59514 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 60134 25174
rect 59514 24854 60134 24938
rect 59514 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 60134 24854
rect 59123 15196 59189 15197
rect 59123 15132 59124 15196
rect 59188 15132 59189 15196
rect 59123 15131 59189 15132
rect 55794 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 56414 -1306
rect 55794 -1626 56414 -1542
rect 55794 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 56414 -1626
rect 55794 -1894 56414 -1862
rect 59514 -3226 60134 24618
rect 59514 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 60134 -3226
rect 59514 -3546 60134 -3462
rect 59514 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 60134 -3546
rect 59514 -3814 60134 -3782
rect 63234 28894 63854 64338
rect 66118 37909 66178 273667
rect 67403 267476 67469 267477
rect 67403 267412 67404 267476
rect 67468 267412 67469 267476
rect 67403 267411 67469 267412
rect 67406 241501 67466 267411
rect 67771 248980 67837 248981
rect 67771 248916 67772 248980
rect 67836 248916 67837 248980
rect 67771 248915 67837 248916
rect 67403 241500 67469 241501
rect 67403 241436 67404 241500
rect 67468 241436 67469 241500
rect 67403 241435 67469 241436
rect 66954 212614 67574 239592
rect 66954 212378 66986 212614
rect 67222 212378 67306 212614
rect 67542 212378 67574 212614
rect 66954 212294 67574 212378
rect 66954 212058 66986 212294
rect 67222 212058 67306 212294
rect 67542 212058 67574 212294
rect 66954 176600 67574 212058
rect 66954 68614 67574 93100
rect 66954 68378 66986 68614
rect 67222 68378 67306 68614
rect 67542 68378 67574 68614
rect 66954 68294 67574 68378
rect 66954 68058 66986 68294
rect 67222 68058 67306 68294
rect 67542 68058 67574 68294
rect 66115 37908 66181 37909
rect 66115 37844 66116 37908
rect 66180 37844 66181 37908
rect 66115 37843 66181 37844
rect 63234 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 63854 28894
rect 63234 28574 63854 28658
rect 63234 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 63854 28574
rect 63234 -5146 63854 28338
rect 63234 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 63854 -5146
rect 63234 -5466 63854 -5382
rect 63234 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 63854 -5466
rect 63234 -5734 63854 -5702
rect 66954 32614 67574 68058
rect 66954 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 67574 32614
rect 66954 32294 67574 32378
rect 66954 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 67574 32294
rect 48954 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 49574 -6106
rect 48954 -6426 49574 -6342
rect 48954 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 49574 -6426
rect 48954 -7654 49574 -6662
rect 66954 -7066 67574 32058
rect 67774 25669 67834 248915
rect 67958 215253 68018 277203
rect 67955 215252 68021 215253
rect 67955 215188 67956 215252
rect 68020 215188 68021 215252
rect 67955 215187 68021 215188
rect 69614 188325 69674 287010
rect 72742 237285 72802 448563
rect 73794 446407 74414 470898
rect 77514 511174 78134 537166
rect 77514 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 78134 511174
rect 77514 510854 78134 510938
rect 77514 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 78134 510854
rect 77514 475174 78134 510618
rect 77514 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 78134 475174
rect 77514 474854 78134 474938
rect 77514 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 78134 474854
rect 77514 446407 78134 474618
rect 81234 514894 81854 537166
rect 81234 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 81854 514894
rect 81234 514574 81854 514658
rect 81234 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 81854 514574
rect 81234 478894 81854 514338
rect 81234 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 81854 478894
rect 81234 478574 81854 478658
rect 81234 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 81854 478574
rect 81234 446407 81854 478338
rect 84954 518614 85574 537166
rect 84954 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 85574 518614
rect 84954 518294 85574 518378
rect 84954 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 85574 518294
rect 84954 482614 85574 518058
rect 84954 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 85574 482614
rect 84954 482294 85574 482378
rect 84954 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 85574 482294
rect 84954 446407 85574 482058
rect 91794 525454 92414 560898
rect 91794 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 92414 525454
rect 91794 525134 92414 525218
rect 91794 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 92414 525134
rect 91794 489454 92414 524898
rect 91794 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 92414 489454
rect 91794 489134 92414 489218
rect 91794 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 92414 489134
rect 91139 465764 91205 465765
rect 91139 465700 91140 465764
rect 91204 465700 91205 465764
rect 91139 465699 91205 465700
rect 89667 464404 89733 464405
rect 89667 464340 89668 464404
rect 89732 464340 89733 464404
rect 89667 464339 89733 464340
rect 72978 435454 73298 435486
rect 72978 435218 73020 435454
rect 73256 435218 73298 435454
rect 72978 435134 73298 435218
rect 72978 434898 73020 435134
rect 73256 434898 73298 435134
rect 72978 434866 73298 434898
rect 88338 417454 88658 417486
rect 88338 417218 88380 417454
rect 88616 417218 88658 417454
rect 88338 417134 88658 417218
rect 88338 416898 88380 417134
rect 88616 416898 88658 417134
rect 88338 416866 88658 416898
rect 72978 399454 73298 399486
rect 72978 399218 73020 399454
rect 73256 399218 73298 399454
rect 72978 399134 73298 399218
rect 72978 398898 73020 399134
rect 73256 398898 73298 399134
rect 72978 398866 73298 398898
rect 89670 398850 89730 464339
rect 89486 398790 89730 398850
rect 89486 390421 89546 398790
rect 91142 390421 91202 465699
rect 91794 453454 92414 488898
rect 95514 673174 96134 707162
rect 95514 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 96134 673174
rect 95514 672854 96134 672938
rect 95514 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 96134 672854
rect 95514 637174 96134 672618
rect 95514 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 96134 637174
rect 95514 636854 96134 636938
rect 95514 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 96134 636854
rect 95514 601174 96134 636618
rect 95514 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 96134 601174
rect 95514 600854 96134 600938
rect 95514 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 96134 600854
rect 95514 565174 96134 600618
rect 95514 564938 95546 565174
rect 95782 564938 95866 565174
rect 96102 564938 96134 565174
rect 95514 564854 96134 564938
rect 95514 564618 95546 564854
rect 95782 564618 95866 564854
rect 96102 564618 96134 564854
rect 95514 529174 96134 564618
rect 99234 676894 99854 709082
rect 99234 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 99854 676894
rect 99234 676574 99854 676658
rect 99234 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 99854 676574
rect 99234 640894 99854 676338
rect 99234 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 99854 640894
rect 99234 640574 99854 640658
rect 99234 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 99854 640574
rect 99234 604894 99854 640338
rect 99234 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 99854 604894
rect 99234 604574 99854 604658
rect 99234 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 99854 604574
rect 99234 568894 99854 604338
rect 99234 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 99854 568894
rect 99234 568574 99854 568658
rect 99234 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 99854 568574
rect 99234 532894 99854 568338
rect 99234 532658 99266 532894
rect 99502 532658 99586 532894
rect 99822 532658 99854 532894
rect 99234 532574 99854 532658
rect 99234 532338 99266 532574
rect 99502 532338 99586 532574
rect 99822 532338 99854 532574
rect 97947 531452 98013 531453
rect 97947 531388 97948 531452
rect 98012 531388 98013 531452
rect 97947 531387 98013 531388
rect 95514 528938 95546 529174
rect 95782 528938 95866 529174
rect 96102 528938 96134 529174
rect 95514 528854 96134 528938
rect 95514 528618 95546 528854
rect 95782 528618 95866 528854
rect 96102 528618 96134 528854
rect 95514 493174 96134 528618
rect 95514 492938 95546 493174
rect 95782 492938 95866 493174
rect 96102 492938 96134 493174
rect 95514 492854 96134 492938
rect 95514 492618 95546 492854
rect 95782 492618 95866 492854
rect 96102 492618 96134 492854
rect 92611 462908 92677 462909
rect 92611 462844 92612 462908
rect 92676 462844 92677 462908
rect 92611 462843 92677 462844
rect 91794 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 92414 453454
rect 91794 453134 92414 453218
rect 91794 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 92414 453134
rect 91794 446407 92414 452898
rect 92614 391101 92674 462843
rect 93899 459644 93965 459645
rect 93899 459580 93900 459644
rect 93964 459580 93965 459644
rect 93899 459579 93965 459580
rect 92611 391100 92677 391101
rect 92611 391036 92612 391100
rect 92676 391036 92677 391100
rect 92611 391035 92677 391036
rect 93902 390421 93962 459579
rect 95514 457174 96134 492618
rect 95514 456938 95546 457174
rect 95782 456938 95866 457174
rect 96102 456938 96134 457174
rect 95514 456854 96134 456938
rect 95514 456618 95546 456854
rect 95782 456618 95866 456854
rect 96102 456618 96134 456854
rect 95187 447812 95253 447813
rect 95187 447748 95188 447812
rect 95252 447810 95253 447812
rect 95252 447750 95434 447810
rect 95252 447748 95253 447750
rect 95187 447747 95253 447748
rect 94451 444684 94517 444685
rect 94451 444620 94452 444684
rect 94516 444620 94517 444684
rect 94451 444619 94517 444620
rect 89483 390420 89549 390421
rect 89483 390356 89484 390420
rect 89548 390356 89549 390420
rect 89483 390355 89549 390356
rect 91139 390420 91205 390421
rect 91139 390356 91140 390420
rect 91204 390356 91205 390420
rect 91139 390355 91205 390356
rect 93899 390420 93965 390421
rect 93899 390356 93900 390420
rect 93964 390356 93965 390420
rect 93899 390355 93965 390356
rect 73794 363454 74414 388356
rect 73794 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 74414 363454
rect 73794 363134 74414 363218
rect 73794 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 74414 363134
rect 73794 331592 74414 362898
rect 77514 367174 78134 388356
rect 77514 366938 77546 367174
rect 77782 366938 77866 367174
rect 78102 366938 78134 367174
rect 77514 366854 78134 366938
rect 77514 366618 77546 366854
rect 77782 366618 77866 366854
rect 78102 366618 78134 366854
rect 77514 331592 78134 366618
rect 81234 370894 81854 388356
rect 83963 384980 84029 384981
rect 83963 384916 83964 384980
rect 84028 384916 84029 384980
rect 83963 384915 84029 384916
rect 81234 370658 81266 370894
rect 81502 370658 81586 370894
rect 81822 370658 81854 370894
rect 81234 370574 81854 370658
rect 81234 370338 81266 370574
rect 81502 370338 81586 370574
rect 81822 370338 81854 370574
rect 81019 359412 81085 359413
rect 81019 359348 81020 359412
rect 81084 359348 81085 359412
rect 81019 359347 81085 359348
rect 75683 331260 75749 331261
rect 75683 331196 75684 331260
rect 75748 331196 75749 331260
rect 75683 331195 75749 331196
rect 72978 291454 73298 291486
rect 72978 291218 73020 291454
rect 73256 291218 73298 291454
rect 72978 291134 73298 291218
rect 72978 290898 73020 291134
rect 73256 290898 73298 291134
rect 72978 290866 73298 290898
rect 72978 255454 73298 255486
rect 72978 255218 73020 255454
rect 73256 255218 73298 255454
rect 72978 255134 73298 255218
rect 72978 254898 73020 255134
rect 73256 254898 73298 255134
rect 72978 254866 73298 254898
rect 72739 237284 72805 237285
rect 72739 237220 72740 237284
rect 72804 237220 72805 237284
rect 72739 237219 72805 237220
rect 73794 219454 74414 239592
rect 73794 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 74414 219454
rect 73794 219134 74414 219218
rect 73794 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 74414 219134
rect 69611 188324 69677 188325
rect 69611 188260 69612 188324
rect 69676 188260 69677 188324
rect 69611 188259 69677 188260
rect 73794 183454 74414 218898
rect 75686 189685 75746 331195
rect 77155 329492 77221 329493
rect 77155 329428 77156 329492
rect 77220 329428 77221 329492
rect 77155 329427 77221 329428
rect 77158 191181 77218 329427
rect 81022 242045 81082 359347
rect 81234 334894 81854 370338
rect 81234 334658 81266 334894
rect 81502 334658 81586 334894
rect 81822 334658 81854 334894
rect 81234 334574 81854 334658
rect 81234 334338 81266 334574
rect 81502 334338 81586 334574
rect 81822 334338 81854 334574
rect 81234 331592 81854 334338
rect 82675 331804 82741 331805
rect 82675 331740 82676 331804
rect 82740 331740 82741 331804
rect 82675 331739 82741 331740
rect 81019 242044 81085 242045
rect 81019 241980 81020 242044
rect 81084 241980 81085 242044
rect 81019 241979 81085 241980
rect 77514 223174 78134 239592
rect 77514 222938 77546 223174
rect 77782 222938 77866 223174
rect 78102 222938 78134 223174
rect 77514 222854 78134 222938
rect 77514 222618 77546 222854
rect 77782 222618 77866 222854
rect 78102 222618 78134 222854
rect 77155 191180 77221 191181
rect 77155 191116 77156 191180
rect 77220 191116 77221 191180
rect 77155 191115 77221 191116
rect 75683 189684 75749 189685
rect 75683 189620 75684 189684
rect 75748 189620 75749 189684
rect 75683 189619 75749 189620
rect 73794 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 74414 183454
rect 73794 183134 74414 183218
rect 73794 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 74414 183134
rect 73794 176600 74414 182898
rect 77514 187174 78134 222618
rect 77514 186938 77546 187174
rect 77782 186938 77866 187174
rect 78102 186938 78134 187174
rect 77514 186854 78134 186938
rect 77514 186618 77546 186854
rect 77782 186618 77866 186854
rect 78102 186618 78134 186854
rect 77514 176600 78134 186618
rect 81234 226894 81854 239592
rect 82678 234429 82738 331739
rect 83966 241501 84026 384915
rect 84954 374614 85574 388356
rect 84954 374378 84986 374614
rect 85222 374378 85306 374614
rect 85542 374378 85574 374614
rect 84954 374294 85574 374378
rect 84954 374058 84986 374294
rect 85222 374058 85306 374294
rect 85542 374058 85574 374294
rect 84954 338614 85574 374058
rect 84954 338378 84986 338614
rect 85222 338378 85306 338614
rect 85542 338378 85574 338614
rect 84954 338294 85574 338378
rect 84954 338058 84986 338294
rect 85222 338058 85306 338294
rect 85542 338058 85574 338294
rect 84954 331592 85574 338058
rect 91794 381454 92414 388356
rect 91794 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 92414 381454
rect 91794 381134 92414 381218
rect 91794 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 92414 381134
rect 91794 345454 92414 380898
rect 94454 345813 94514 444619
rect 95374 393330 95434 447750
rect 95514 446407 96134 456618
rect 96659 453252 96725 453253
rect 96659 453188 96660 453252
rect 96724 453188 96725 453252
rect 96659 453187 96725 453188
rect 96475 445772 96541 445773
rect 96475 445708 96476 445772
rect 96540 445708 96541 445772
rect 96475 445707 96541 445708
rect 95190 393270 95434 393330
rect 95190 389061 95250 393270
rect 95187 389060 95253 389061
rect 95187 388996 95188 389060
rect 95252 388996 95253 389060
rect 95187 388995 95253 388996
rect 95190 385661 95250 388995
rect 96478 388517 96538 445707
rect 96662 390421 96722 453187
rect 96659 390420 96725 390421
rect 96659 390356 96660 390420
rect 96724 390356 96725 390420
rect 96659 390355 96725 390356
rect 97950 388653 98010 531387
rect 99234 496894 99854 532338
rect 99234 496658 99266 496894
rect 99502 496658 99586 496894
rect 99822 496658 99854 496894
rect 99234 496574 99854 496658
rect 99234 496338 99266 496574
rect 99502 496338 99586 496574
rect 99822 496338 99854 496574
rect 99234 460894 99854 496338
rect 99234 460658 99266 460894
rect 99502 460658 99586 460894
rect 99822 460658 99854 460894
rect 99234 460574 99854 460658
rect 99234 460338 99266 460574
rect 99502 460338 99586 460574
rect 99822 460338 99854 460574
rect 98131 456108 98197 456109
rect 98131 456044 98132 456108
rect 98196 456044 98197 456108
rect 98131 456043 98197 456044
rect 98134 390421 98194 456043
rect 99234 446407 99854 460338
rect 102954 680614 103574 711002
rect 120954 710598 121574 711590
rect 120954 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 121574 710598
rect 120954 710278 121574 710362
rect 120954 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 121574 710278
rect 117234 708678 117854 709670
rect 117234 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 117854 708678
rect 117234 708358 117854 708442
rect 117234 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 117854 708358
rect 113514 706758 114134 707750
rect 113514 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 114134 706758
rect 113514 706438 114134 706522
rect 113514 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 114134 706438
rect 102954 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 103574 680614
rect 102954 680294 103574 680378
rect 102954 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 103574 680294
rect 102954 644614 103574 680058
rect 102954 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 103574 644614
rect 102954 644294 103574 644378
rect 102954 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 103574 644294
rect 102954 608614 103574 644058
rect 102954 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 103574 608614
rect 102954 608294 103574 608378
rect 102954 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 103574 608294
rect 102954 572614 103574 608058
rect 102954 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 103574 572614
rect 102954 572294 103574 572378
rect 102954 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 103574 572294
rect 102954 536614 103574 572058
rect 102954 536378 102986 536614
rect 103222 536378 103306 536614
rect 103542 536378 103574 536614
rect 102954 536294 103574 536378
rect 102954 536058 102986 536294
rect 103222 536058 103306 536294
rect 103542 536058 103574 536294
rect 102954 500614 103574 536058
rect 102954 500378 102986 500614
rect 103222 500378 103306 500614
rect 103542 500378 103574 500614
rect 102954 500294 103574 500378
rect 102954 500058 102986 500294
rect 103222 500058 103306 500294
rect 103542 500058 103574 500294
rect 102954 464614 103574 500058
rect 109794 704838 110414 705830
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 615454 110414 650898
rect 109794 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 110414 615454
rect 109794 615134 110414 615218
rect 109794 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 110414 615134
rect 109794 579454 110414 614898
rect 109794 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 110414 579454
rect 109794 579134 110414 579218
rect 109794 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 110414 579134
rect 109794 543454 110414 578898
rect 109794 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 110414 543454
rect 109794 543134 110414 543218
rect 109794 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 110414 543134
rect 109794 507454 110414 542898
rect 109794 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 110414 507454
rect 109794 507134 110414 507218
rect 109794 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 110414 507134
rect 109794 471454 110414 506898
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 106411 471204 106477 471205
rect 106411 471140 106412 471204
rect 106476 471140 106477 471204
rect 106411 471139 106477 471140
rect 104939 469844 105005 469845
rect 104939 469780 104940 469844
rect 105004 469780 105005 469844
rect 104939 469779 105005 469780
rect 102954 464378 102986 464614
rect 103222 464378 103306 464614
rect 103542 464378 103574 464614
rect 102954 464294 103574 464378
rect 102954 464058 102986 464294
rect 103222 464058 103306 464294
rect 103542 464058 103574 464294
rect 100707 457468 100773 457469
rect 100707 457404 100708 457468
rect 100772 457404 100773 457468
rect 100707 457403 100773 457404
rect 100523 445772 100589 445773
rect 100523 445708 100524 445772
rect 100588 445708 100589 445772
rect 100523 445707 100589 445708
rect 98131 390420 98197 390421
rect 98131 390356 98132 390420
rect 98196 390356 98197 390420
rect 98131 390355 98197 390356
rect 97947 388652 98013 388653
rect 97947 388588 97948 388652
rect 98012 388588 98013 388652
rect 97947 388587 98013 388588
rect 96475 388516 96541 388517
rect 96475 388452 96476 388516
rect 96540 388452 96541 388516
rect 96475 388451 96541 388452
rect 95187 385660 95253 385661
rect 95187 385596 95188 385660
rect 95252 385596 95253 385660
rect 95187 385595 95253 385596
rect 95514 385174 96134 388356
rect 95514 384938 95546 385174
rect 95782 384938 95866 385174
rect 96102 384938 96134 385174
rect 95514 384854 96134 384938
rect 95514 384618 95546 384854
rect 95782 384618 95866 384854
rect 96102 384618 96134 384854
rect 95514 349174 96134 384618
rect 95514 348938 95546 349174
rect 95782 348938 95866 349174
rect 96102 348938 96134 349174
rect 95514 348854 96134 348938
rect 95514 348618 95546 348854
rect 95782 348618 95866 348854
rect 96102 348618 96134 348854
rect 94451 345812 94517 345813
rect 94451 345748 94452 345812
rect 94516 345748 94517 345812
rect 94451 345747 94517 345748
rect 91794 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 92414 345454
rect 91794 345134 92414 345218
rect 91794 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 92414 345134
rect 91794 331592 92414 344898
rect 95514 331592 96134 348618
rect 99234 352894 99854 388356
rect 100526 353565 100586 445707
rect 100710 390285 100770 457403
rect 102179 456108 102245 456109
rect 102179 456044 102180 456108
rect 102244 456044 102245 456108
rect 102179 456043 102245 456044
rect 102182 390557 102242 456043
rect 102954 446407 103574 464058
rect 103698 435454 104018 435486
rect 103698 435218 103740 435454
rect 103976 435218 104018 435454
rect 103698 435134 104018 435218
rect 103698 434898 103740 435134
rect 103976 434898 104018 435134
rect 103698 434866 104018 434898
rect 103698 399454 104018 399486
rect 103698 399218 103740 399454
rect 103976 399218 104018 399454
rect 103698 399134 104018 399218
rect 103698 398898 103740 399134
rect 103976 398898 104018 399134
rect 103698 398866 104018 398898
rect 102179 390556 102245 390557
rect 102179 390492 102180 390556
rect 102244 390492 102245 390556
rect 102179 390491 102245 390492
rect 104942 390421 105002 469779
rect 106414 390421 106474 471139
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 107699 464404 107765 464405
rect 107699 464340 107700 464404
rect 107764 464340 107765 464404
rect 107699 464339 107765 464340
rect 107702 390421 107762 464339
rect 108987 457060 109053 457061
rect 108987 456996 108988 457060
rect 109052 456996 109053 457060
rect 108987 456995 109053 456996
rect 108803 444548 108869 444549
rect 108803 444484 108804 444548
rect 108868 444484 108869 444548
rect 108803 444483 108869 444484
rect 104939 390420 105005 390421
rect 104939 390356 104940 390420
rect 105004 390356 105005 390420
rect 104939 390355 105005 390356
rect 106411 390420 106477 390421
rect 106411 390356 106412 390420
rect 106476 390356 106477 390420
rect 106411 390355 106477 390356
rect 107699 390420 107765 390421
rect 107699 390356 107700 390420
rect 107764 390356 107765 390420
rect 107699 390355 107765 390356
rect 100707 390284 100773 390285
rect 100707 390220 100708 390284
rect 100772 390220 100773 390284
rect 100707 390219 100773 390220
rect 102954 356614 103574 388356
rect 108806 361725 108866 444483
rect 108990 390421 109050 456995
rect 109794 446407 110414 470898
rect 113514 691174 114134 706202
rect 113514 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 114134 691174
rect 113514 690854 114134 690938
rect 113514 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 114134 690854
rect 113514 655174 114134 690618
rect 113514 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 114134 655174
rect 113514 654854 114134 654938
rect 113514 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 114134 654854
rect 113514 619174 114134 654618
rect 113514 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 114134 619174
rect 113514 618854 114134 618938
rect 113514 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 114134 618854
rect 113514 583174 114134 618618
rect 113514 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 114134 583174
rect 113514 582854 114134 582938
rect 113514 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 114134 582854
rect 113514 547174 114134 582618
rect 113514 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 114134 547174
rect 113514 546854 114134 546938
rect 113514 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 114134 546854
rect 113514 511174 114134 546618
rect 113514 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 114134 511174
rect 113514 510854 114134 510938
rect 113514 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 114134 510854
rect 113514 475174 114134 510618
rect 113514 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 114134 475174
rect 113514 474854 114134 474938
rect 113514 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 114134 474854
rect 111747 460188 111813 460189
rect 111747 460124 111748 460188
rect 111812 460124 111813 460188
rect 111747 460123 111813 460124
rect 111563 444548 111629 444549
rect 111563 444484 111564 444548
rect 111628 444484 111629 444548
rect 111563 444483 111629 444484
rect 108987 390420 109053 390421
rect 108987 390356 108988 390420
rect 109052 390356 109053 390420
rect 108987 390355 109053 390356
rect 109794 363454 110414 388356
rect 109794 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 110414 363454
rect 109794 363134 110414 363218
rect 109794 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 110414 363134
rect 108803 361724 108869 361725
rect 108803 361660 108804 361724
rect 108868 361660 108869 361724
rect 108803 361659 108869 361660
rect 102954 356378 102986 356614
rect 103222 356378 103306 356614
rect 103542 356378 103574 356614
rect 102954 356294 103574 356378
rect 102954 356058 102986 356294
rect 103222 356058 103306 356294
rect 103542 356058 103574 356294
rect 100523 353564 100589 353565
rect 100523 353500 100524 353564
rect 100588 353500 100589 353564
rect 100523 353499 100589 353500
rect 99234 352658 99266 352894
rect 99502 352658 99586 352894
rect 99822 352658 99854 352894
rect 99234 352574 99854 352658
rect 99234 352338 99266 352574
rect 99502 352338 99586 352574
rect 99822 352338 99854 352574
rect 99234 331592 99854 352338
rect 102954 331592 103574 356058
rect 109794 331592 110414 362898
rect 111566 357645 111626 444483
rect 111750 389061 111810 460123
rect 113514 446407 114134 474618
rect 117234 694894 117854 708122
rect 117234 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 117854 694894
rect 117234 694574 117854 694658
rect 117234 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 117854 694574
rect 117234 658894 117854 694338
rect 117234 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 117854 658894
rect 117234 658574 117854 658658
rect 117234 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 117854 658574
rect 117234 622894 117854 658338
rect 117234 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 117854 622894
rect 117234 622574 117854 622658
rect 117234 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 117854 622574
rect 117234 586894 117854 622338
rect 117234 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 117854 586894
rect 117234 586574 117854 586658
rect 117234 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 117854 586574
rect 117234 550894 117854 586338
rect 117234 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 117854 550894
rect 117234 550574 117854 550658
rect 117234 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 117854 550574
rect 117234 514894 117854 550338
rect 117234 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 117854 514894
rect 117234 514574 117854 514658
rect 117234 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 117854 514574
rect 117234 478894 117854 514338
rect 117234 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 117854 478894
rect 117234 478574 117854 478658
rect 117234 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 117854 478574
rect 115979 468484 116045 468485
rect 115979 468420 115980 468484
rect 116044 468420 116045 468484
rect 115979 468419 116045 468420
rect 115795 445772 115861 445773
rect 115795 445708 115796 445772
rect 115860 445708 115861 445772
rect 115795 445707 115861 445708
rect 115798 444821 115858 445707
rect 115795 444820 115861 444821
rect 115795 444756 115796 444820
rect 115860 444756 115861 444820
rect 115795 444755 115861 444756
rect 114323 444548 114389 444549
rect 114323 444484 114324 444548
rect 114388 444484 114389 444548
rect 114323 444483 114389 444484
rect 111747 389060 111813 389061
rect 111747 388996 111748 389060
rect 111812 388996 111813 389060
rect 111747 388995 111813 388996
rect 111563 357644 111629 357645
rect 111563 357580 111564 357644
rect 111628 357580 111629 357644
rect 111563 357579 111629 357580
rect 111750 342957 111810 388995
rect 113514 367174 114134 388356
rect 114326 375325 114386 444483
rect 114323 375324 114389 375325
rect 114323 375260 114324 375324
rect 114388 375260 114389 375324
rect 114323 375259 114389 375260
rect 113514 366938 113546 367174
rect 113782 366938 113866 367174
rect 114102 366938 114134 367174
rect 113514 366854 114134 366938
rect 113514 366618 113546 366854
rect 113782 366618 113866 366854
rect 114102 366618 114134 366854
rect 111747 342956 111813 342957
rect 111747 342892 111748 342956
rect 111812 342892 111813 342956
rect 111747 342891 111813 342892
rect 113514 331592 114134 366618
rect 115798 339965 115858 444755
rect 115982 390421 116042 468419
rect 117234 446407 117854 478338
rect 120954 698614 121574 710042
rect 138954 711558 139574 711590
rect 138954 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 139574 711558
rect 138954 711238 139574 711322
rect 138954 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 139574 711238
rect 135234 709638 135854 709670
rect 135234 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 135854 709638
rect 135234 709318 135854 709402
rect 135234 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 135854 709318
rect 131514 707718 132134 707750
rect 131514 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 132134 707718
rect 131514 707398 132134 707482
rect 131514 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 132134 707398
rect 120954 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 121574 698614
rect 120954 698294 121574 698378
rect 120954 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 121574 698294
rect 120954 662614 121574 698058
rect 120954 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 121574 662614
rect 120954 662294 121574 662378
rect 120954 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 121574 662294
rect 120954 626614 121574 662058
rect 120954 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 121574 626614
rect 120954 626294 121574 626378
rect 120954 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 121574 626294
rect 120954 590614 121574 626058
rect 120954 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 121574 590614
rect 120954 590294 121574 590378
rect 120954 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 121574 590294
rect 120954 554614 121574 590058
rect 120954 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 121574 554614
rect 120954 554294 121574 554378
rect 120954 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 121574 554294
rect 120954 518614 121574 554058
rect 120954 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 121574 518614
rect 120954 518294 121574 518378
rect 120954 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 121574 518294
rect 120954 482614 121574 518058
rect 120954 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 121574 482614
rect 120954 482294 121574 482378
rect 120954 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 121574 482294
rect 118003 464404 118069 464405
rect 118003 464340 118004 464404
rect 118068 464340 118069 464404
rect 118003 464339 118069 464340
rect 115979 390420 116045 390421
rect 115979 390356 115980 390420
rect 116044 390356 116045 390420
rect 115979 390355 116045 390356
rect 118006 389061 118066 464339
rect 118739 458828 118805 458829
rect 118739 458764 118740 458828
rect 118804 458764 118805 458828
rect 118739 458763 118805 458764
rect 118555 445772 118621 445773
rect 118555 445708 118556 445772
rect 118620 445708 118621 445772
rect 118555 445707 118621 445708
rect 118003 389060 118069 389061
rect 118003 388996 118004 389060
rect 118068 388996 118069 389060
rect 118003 388995 118069 388996
rect 117234 370894 117854 388356
rect 117234 370658 117266 370894
rect 117502 370658 117586 370894
rect 117822 370658 117854 370894
rect 117234 370574 117854 370658
rect 117234 370338 117266 370574
rect 117502 370338 117586 370574
rect 117822 370338 117854 370574
rect 115795 339964 115861 339965
rect 115795 339900 115796 339964
rect 115860 339900 115861 339964
rect 115795 339899 115861 339900
rect 115798 339557 115858 339899
rect 115795 339556 115861 339557
rect 115795 339492 115796 339556
rect 115860 339492 115861 339556
rect 115795 339491 115861 339492
rect 117234 334894 117854 370338
rect 118558 349213 118618 445707
rect 118742 390421 118802 458763
rect 120211 449172 120277 449173
rect 120211 449108 120212 449172
rect 120276 449108 120277 449172
rect 120211 449107 120277 449108
rect 120027 430676 120093 430677
rect 120027 430612 120028 430676
rect 120092 430612 120093 430676
rect 120027 430611 120093 430612
rect 119058 417454 119378 417486
rect 119058 417218 119100 417454
rect 119336 417218 119378 417454
rect 119058 417134 119378 417218
rect 119058 416898 119100 417134
rect 119336 416898 119378 417134
rect 119058 416866 119378 416898
rect 119475 392188 119541 392189
rect 119475 392124 119476 392188
rect 119540 392124 119541 392188
rect 119475 392123 119541 392124
rect 118739 390420 118805 390421
rect 118739 390356 118740 390420
rect 118804 390356 118805 390420
rect 118739 390355 118805 390356
rect 119478 371925 119538 392123
rect 120030 377365 120090 430611
rect 120214 426053 120274 449107
rect 120954 446407 121574 482058
rect 127794 705798 128414 705830
rect 127794 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 128414 705798
rect 127794 705478 128414 705562
rect 127794 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 128414 705478
rect 127794 669454 128414 705242
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 633454 128414 668898
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 127794 597454 128414 632898
rect 127794 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 128414 597454
rect 127794 597134 128414 597218
rect 127794 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 128414 597134
rect 127794 561454 128414 596898
rect 127794 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 128414 561454
rect 127794 561134 128414 561218
rect 127794 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 128414 561134
rect 127794 525454 128414 560898
rect 127794 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 128414 525454
rect 127794 525134 128414 525218
rect 127794 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 128414 525134
rect 127794 489454 128414 524898
rect 127794 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 128414 489454
rect 127794 489134 128414 489218
rect 127794 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 128414 489134
rect 122603 479500 122669 479501
rect 122603 479436 122604 479500
rect 122668 479436 122669 479500
rect 122603 479435 122669 479436
rect 121683 435300 121749 435301
rect 121683 435236 121684 435300
rect 121748 435236 121749 435300
rect 121683 435235 121749 435236
rect 120211 426052 120277 426053
rect 120211 425988 120212 426052
rect 120276 425988 120277 426052
rect 120211 425987 120277 425988
rect 120027 377364 120093 377365
rect 120027 377300 120028 377364
rect 120092 377300 120093 377364
rect 120027 377299 120093 377300
rect 120954 374614 121574 388356
rect 120954 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 121574 374614
rect 120954 374294 121574 374378
rect 120954 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 121574 374294
rect 119475 371924 119541 371925
rect 119475 371860 119476 371924
rect 119540 371860 119541 371924
rect 119475 371859 119541 371860
rect 118555 349212 118621 349213
rect 118555 349148 118556 349212
rect 118620 349148 118621 349212
rect 118555 349147 118621 349148
rect 117234 334658 117266 334894
rect 117502 334658 117586 334894
rect 117822 334658 117854 334894
rect 117234 334574 117854 334658
rect 117234 334338 117266 334574
rect 117502 334338 117586 334574
rect 117822 334338 117854 334574
rect 117234 331592 117854 334338
rect 120954 338614 121574 374058
rect 121686 349077 121746 435235
rect 122606 403749 122666 479435
rect 127794 453454 128414 488898
rect 127794 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 128414 453454
rect 127794 453134 128414 453218
rect 127794 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 128414 453134
rect 124259 444820 124325 444821
rect 124259 444756 124260 444820
rect 124324 444756 124325 444820
rect 124259 444755 124325 444756
rect 124262 420885 124322 444755
rect 124259 420884 124325 420885
rect 124259 420820 124260 420884
rect 124324 420820 124325 420884
rect 124259 420819 124325 420820
rect 127794 417454 128414 452898
rect 127794 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 128414 417454
rect 127794 417134 128414 417218
rect 127794 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 128414 417134
rect 122603 403748 122669 403749
rect 122603 403684 122604 403748
rect 122668 403684 122669 403748
rect 122603 403683 122669 403684
rect 127794 381454 128414 416898
rect 127794 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 128414 381454
rect 127794 381134 128414 381218
rect 127794 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 128414 381134
rect 124811 378860 124877 378861
rect 124811 378796 124812 378860
rect 124876 378796 124877 378860
rect 124811 378795 124877 378796
rect 124814 360229 124874 378795
rect 124811 360228 124877 360229
rect 124811 360164 124812 360228
rect 124876 360164 124877 360228
rect 124811 360163 124877 360164
rect 121683 349076 121749 349077
rect 121683 349012 121684 349076
rect 121748 349012 121749 349076
rect 121683 349011 121749 349012
rect 120954 338378 120986 338614
rect 121222 338378 121306 338614
rect 121542 338378 121574 338614
rect 120954 338294 121574 338378
rect 120954 338058 120986 338294
rect 121222 338058 121306 338294
rect 121542 338058 121574 338294
rect 120954 331592 121574 338058
rect 127794 345454 128414 380898
rect 127794 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 128414 345454
rect 127794 345134 128414 345218
rect 127794 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 128414 345134
rect 127794 331592 128414 344898
rect 131514 673174 132134 707162
rect 131514 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 132134 673174
rect 131514 672854 132134 672938
rect 131514 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 132134 672854
rect 131514 637174 132134 672618
rect 131514 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 132134 637174
rect 131514 636854 132134 636938
rect 131514 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 132134 636854
rect 131514 601174 132134 636618
rect 131514 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 132134 601174
rect 131514 600854 132134 600938
rect 131514 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 132134 600854
rect 131514 565174 132134 600618
rect 131514 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 132134 565174
rect 131514 564854 132134 564938
rect 131514 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 132134 564854
rect 131514 529174 132134 564618
rect 131514 528938 131546 529174
rect 131782 528938 131866 529174
rect 132102 528938 132134 529174
rect 131514 528854 132134 528938
rect 131514 528618 131546 528854
rect 131782 528618 131866 528854
rect 132102 528618 132134 528854
rect 131514 493174 132134 528618
rect 131514 492938 131546 493174
rect 131782 492938 131866 493174
rect 132102 492938 132134 493174
rect 131514 492854 132134 492938
rect 131514 492618 131546 492854
rect 131782 492618 131866 492854
rect 132102 492618 132134 492854
rect 131514 457174 132134 492618
rect 131514 456938 131546 457174
rect 131782 456938 131866 457174
rect 132102 456938 132134 457174
rect 131514 456854 132134 456938
rect 131514 456618 131546 456854
rect 131782 456618 131866 456854
rect 132102 456618 132134 456854
rect 131514 421174 132134 456618
rect 131514 420938 131546 421174
rect 131782 420938 131866 421174
rect 132102 420938 132134 421174
rect 131514 420854 132134 420938
rect 131514 420618 131546 420854
rect 131782 420618 131866 420854
rect 132102 420618 132134 420854
rect 131514 385174 132134 420618
rect 131514 384938 131546 385174
rect 131782 384938 131866 385174
rect 132102 384938 132134 385174
rect 131514 384854 132134 384938
rect 131514 384618 131546 384854
rect 131782 384618 131866 384854
rect 132102 384618 132134 384854
rect 131514 349174 132134 384618
rect 131514 348938 131546 349174
rect 131782 348938 131866 349174
rect 132102 348938 132134 349174
rect 131514 348854 132134 348938
rect 131514 348618 131546 348854
rect 131782 348618 131866 348854
rect 132102 348618 132134 348854
rect 131514 331592 132134 348618
rect 135234 676894 135854 709082
rect 135234 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 135854 676894
rect 135234 676574 135854 676658
rect 135234 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 135854 676574
rect 135234 640894 135854 676338
rect 135234 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 135854 640894
rect 135234 640574 135854 640658
rect 135234 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 135854 640574
rect 135234 604894 135854 640338
rect 135234 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 135854 604894
rect 135234 604574 135854 604658
rect 135234 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 135854 604574
rect 135234 568894 135854 604338
rect 135234 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 135854 568894
rect 135234 568574 135854 568658
rect 135234 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 135854 568574
rect 135234 532894 135854 568338
rect 135234 532658 135266 532894
rect 135502 532658 135586 532894
rect 135822 532658 135854 532894
rect 135234 532574 135854 532658
rect 135234 532338 135266 532574
rect 135502 532338 135586 532574
rect 135822 532338 135854 532574
rect 135234 496894 135854 532338
rect 135234 496658 135266 496894
rect 135502 496658 135586 496894
rect 135822 496658 135854 496894
rect 135234 496574 135854 496658
rect 135234 496338 135266 496574
rect 135502 496338 135586 496574
rect 135822 496338 135854 496574
rect 135234 460894 135854 496338
rect 135234 460658 135266 460894
rect 135502 460658 135586 460894
rect 135822 460658 135854 460894
rect 135234 460574 135854 460658
rect 135234 460338 135266 460574
rect 135502 460338 135586 460574
rect 135822 460338 135854 460574
rect 135234 424894 135854 460338
rect 135234 424658 135266 424894
rect 135502 424658 135586 424894
rect 135822 424658 135854 424894
rect 135234 424574 135854 424658
rect 135234 424338 135266 424574
rect 135502 424338 135586 424574
rect 135822 424338 135854 424574
rect 135234 388894 135854 424338
rect 135234 388658 135266 388894
rect 135502 388658 135586 388894
rect 135822 388658 135854 388894
rect 135234 388574 135854 388658
rect 135234 388338 135266 388574
rect 135502 388338 135586 388574
rect 135822 388338 135854 388574
rect 135234 352894 135854 388338
rect 135234 352658 135266 352894
rect 135502 352658 135586 352894
rect 135822 352658 135854 352894
rect 135234 352574 135854 352658
rect 135234 352338 135266 352574
rect 135502 352338 135586 352574
rect 135822 352338 135854 352574
rect 135234 331592 135854 352338
rect 138954 680614 139574 711002
rect 156954 710598 157574 711590
rect 156954 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 157574 710598
rect 156954 710278 157574 710362
rect 156954 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 157574 710278
rect 153234 708678 153854 709670
rect 153234 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 153854 708678
rect 153234 708358 153854 708442
rect 153234 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 153854 708358
rect 149514 706758 150134 707750
rect 149514 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 150134 706758
rect 149514 706438 150134 706522
rect 149514 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 150134 706438
rect 138954 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 139574 680614
rect 138954 680294 139574 680378
rect 138954 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 139574 680294
rect 138954 644614 139574 680058
rect 138954 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 139574 644614
rect 138954 644294 139574 644378
rect 138954 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 139574 644294
rect 138954 608614 139574 644058
rect 138954 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 139574 608614
rect 138954 608294 139574 608378
rect 138954 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 139574 608294
rect 138954 572614 139574 608058
rect 138954 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 139574 572614
rect 138954 572294 139574 572378
rect 138954 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 139574 572294
rect 138954 536614 139574 572058
rect 138954 536378 138986 536614
rect 139222 536378 139306 536614
rect 139542 536378 139574 536614
rect 138954 536294 139574 536378
rect 138954 536058 138986 536294
rect 139222 536058 139306 536294
rect 139542 536058 139574 536294
rect 138954 500614 139574 536058
rect 138954 500378 138986 500614
rect 139222 500378 139306 500614
rect 139542 500378 139574 500614
rect 138954 500294 139574 500378
rect 138954 500058 138986 500294
rect 139222 500058 139306 500294
rect 139542 500058 139574 500294
rect 138954 464614 139574 500058
rect 138954 464378 138986 464614
rect 139222 464378 139306 464614
rect 139542 464378 139574 464614
rect 138954 464294 139574 464378
rect 138954 464058 138986 464294
rect 139222 464058 139306 464294
rect 139542 464058 139574 464294
rect 138954 428614 139574 464058
rect 138954 428378 138986 428614
rect 139222 428378 139306 428614
rect 139542 428378 139574 428614
rect 138954 428294 139574 428378
rect 138954 428058 138986 428294
rect 139222 428058 139306 428294
rect 139542 428058 139574 428294
rect 138954 392614 139574 428058
rect 138954 392378 138986 392614
rect 139222 392378 139306 392614
rect 139542 392378 139574 392614
rect 138954 392294 139574 392378
rect 138954 392058 138986 392294
rect 139222 392058 139306 392294
rect 139542 392058 139574 392294
rect 138954 356614 139574 392058
rect 138954 356378 138986 356614
rect 139222 356378 139306 356614
rect 139542 356378 139574 356614
rect 138954 356294 139574 356378
rect 138954 356058 138986 356294
rect 139222 356058 139306 356294
rect 139542 356058 139574 356294
rect 138954 331592 139574 356058
rect 145794 704838 146414 705830
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 579454 146414 614898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 543454 146414 578898
rect 145794 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 146414 543454
rect 145794 543134 146414 543218
rect 145794 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 146414 543134
rect 145794 507454 146414 542898
rect 145794 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 146414 507454
rect 145794 507134 146414 507218
rect 145794 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 146414 507134
rect 145794 471454 146414 506898
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 145794 435454 146414 470898
rect 145794 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 146414 435454
rect 145794 435134 146414 435218
rect 145794 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 146414 435134
rect 145794 399454 146414 434898
rect 145794 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 146414 399454
rect 145794 399134 146414 399218
rect 145794 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 146414 399134
rect 145794 363454 146414 398898
rect 145794 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 146414 363454
rect 145794 363134 146414 363218
rect 145794 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 146414 363134
rect 145794 331592 146414 362898
rect 149514 691174 150134 706202
rect 149514 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 150134 691174
rect 149514 690854 150134 690938
rect 149514 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 150134 690854
rect 149514 655174 150134 690618
rect 149514 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 150134 655174
rect 149514 654854 150134 654938
rect 149514 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 150134 654854
rect 149514 619174 150134 654618
rect 149514 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 150134 619174
rect 149514 618854 150134 618938
rect 149514 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 150134 618854
rect 149514 583174 150134 618618
rect 149514 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 150134 583174
rect 149514 582854 150134 582938
rect 149514 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 150134 582854
rect 149514 547174 150134 582618
rect 149514 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 150134 547174
rect 149514 546854 150134 546938
rect 149514 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 150134 546854
rect 149514 511174 150134 546618
rect 149514 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 150134 511174
rect 149514 510854 150134 510938
rect 149514 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 150134 510854
rect 149514 475174 150134 510618
rect 149514 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 150134 475174
rect 149514 474854 150134 474938
rect 149514 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 150134 474854
rect 149514 439174 150134 474618
rect 149514 438938 149546 439174
rect 149782 438938 149866 439174
rect 150102 438938 150134 439174
rect 149514 438854 150134 438938
rect 149514 438618 149546 438854
rect 149782 438618 149866 438854
rect 150102 438618 150134 438854
rect 149514 403174 150134 438618
rect 149514 402938 149546 403174
rect 149782 402938 149866 403174
rect 150102 402938 150134 403174
rect 149514 402854 150134 402938
rect 149514 402618 149546 402854
rect 149782 402618 149866 402854
rect 150102 402618 150134 402854
rect 149514 367174 150134 402618
rect 149514 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 150134 367174
rect 149514 366854 150134 366938
rect 149514 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 150134 366854
rect 149514 331592 150134 366618
rect 153234 694894 153854 708122
rect 153234 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 153854 694894
rect 153234 694574 153854 694658
rect 153234 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 153854 694574
rect 153234 658894 153854 694338
rect 153234 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 153854 658894
rect 153234 658574 153854 658658
rect 153234 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 153854 658574
rect 153234 622894 153854 658338
rect 153234 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 153854 622894
rect 153234 622574 153854 622658
rect 153234 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 153854 622574
rect 153234 586894 153854 622338
rect 153234 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 153854 586894
rect 153234 586574 153854 586658
rect 153234 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 153854 586574
rect 153234 550894 153854 586338
rect 153234 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 153854 550894
rect 153234 550574 153854 550658
rect 153234 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 153854 550574
rect 153234 514894 153854 550338
rect 153234 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 153854 514894
rect 153234 514574 153854 514658
rect 153234 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 153854 514574
rect 153234 478894 153854 514338
rect 153234 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 153854 478894
rect 153234 478574 153854 478658
rect 153234 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 153854 478574
rect 153234 442894 153854 478338
rect 153234 442658 153266 442894
rect 153502 442658 153586 442894
rect 153822 442658 153854 442894
rect 153234 442574 153854 442658
rect 153234 442338 153266 442574
rect 153502 442338 153586 442574
rect 153822 442338 153854 442574
rect 153234 406894 153854 442338
rect 156954 698614 157574 710042
rect 174954 711558 175574 711590
rect 174954 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 175574 711558
rect 174954 711238 175574 711322
rect 174954 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 175574 711238
rect 171234 709638 171854 709670
rect 171234 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 171854 709638
rect 171234 709318 171854 709402
rect 171234 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 171854 709318
rect 167514 707718 168134 707750
rect 167514 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 168134 707718
rect 167514 707398 168134 707482
rect 167514 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 168134 707398
rect 156954 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 157574 698614
rect 156954 698294 157574 698378
rect 156954 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 157574 698294
rect 156954 662614 157574 698058
rect 156954 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 157574 662614
rect 156954 662294 157574 662378
rect 156954 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 157574 662294
rect 156954 626614 157574 662058
rect 156954 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 157574 626614
rect 156954 626294 157574 626378
rect 156954 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 157574 626294
rect 156954 590614 157574 626058
rect 156954 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 157574 590614
rect 156954 590294 157574 590378
rect 156954 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 157574 590294
rect 156954 554614 157574 590058
rect 156954 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 157574 554614
rect 156954 554294 157574 554378
rect 156954 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 157574 554294
rect 156954 518614 157574 554058
rect 163794 705798 164414 705830
rect 163794 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 164414 705798
rect 163794 705478 164414 705562
rect 163794 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 164414 705478
rect 163794 669454 164414 705242
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 633454 164414 668898
rect 163794 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 164414 633454
rect 163794 633134 164414 633218
rect 163794 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 164414 633134
rect 163794 597454 164414 632898
rect 163794 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 164414 597454
rect 163794 597134 164414 597218
rect 163794 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 164414 597134
rect 163794 561454 164414 596898
rect 163794 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 164414 561454
rect 163794 561134 164414 561218
rect 163794 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 164414 561134
rect 163794 525454 164414 560898
rect 163794 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 164414 525454
rect 163794 525134 164414 525218
rect 163794 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 164414 525134
rect 161979 518940 162045 518941
rect 161979 518876 161980 518940
rect 162044 518876 162045 518940
rect 161979 518875 162045 518876
rect 156954 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 157574 518614
rect 156954 518294 157574 518378
rect 156954 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 157574 518294
rect 156954 482614 157574 518058
rect 156954 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 157574 482614
rect 156954 482294 157574 482378
rect 156954 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 157574 482294
rect 156954 446614 157574 482058
rect 160691 449988 160757 449989
rect 160691 449924 160692 449988
rect 160756 449924 160757 449988
rect 160691 449923 160757 449924
rect 156954 446378 156986 446614
rect 157222 446378 157306 446614
rect 157542 446378 157574 446614
rect 156954 446294 157574 446378
rect 156954 446058 156986 446294
rect 157222 446058 157306 446294
rect 157542 446058 157574 446294
rect 154619 411364 154685 411365
rect 154619 411300 154620 411364
rect 154684 411300 154685 411364
rect 154619 411299 154685 411300
rect 153234 406658 153266 406894
rect 153502 406658 153586 406894
rect 153822 406658 153854 406894
rect 153234 406574 153854 406658
rect 153234 406338 153266 406574
rect 153502 406338 153586 406574
rect 153822 406338 153854 406574
rect 153234 370894 153854 406338
rect 153234 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 153854 370894
rect 153234 370574 153854 370658
rect 153234 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 153854 370574
rect 153234 334894 153854 370338
rect 154067 369068 154133 369069
rect 154067 369004 154068 369068
rect 154132 369004 154133 369068
rect 154067 369003 154133 369004
rect 153234 334658 153266 334894
rect 153502 334658 153586 334894
rect 153822 334658 153854 334894
rect 153234 334574 153854 334658
rect 153234 334338 153266 334574
rect 153502 334338 153586 334574
rect 153822 334338 153854 334574
rect 152595 333300 152661 333301
rect 152595 333236 152596 333300
rect 152660 333236 152661 333300
rect 152595 333235 152661 333236
rect 141923 331396 141989 331397
rect 141923 331332 141924 331396
rect 141988 331332 141989 331396
rect 141923 331331 141989 331332
rect 141926 328130 141986 331331
rect 151859 329900 151925 329901
rect 151859 329836 151860 329900
rect 151924 329836 151925 329900
rect 151859 329835 151925 329836
rect 142291 329220 142357 329221
rect 142291 329156 142292 329220
rect 142356 329156 142357 329220
rect 142291 329155 142357 329156
rect 151675 329220 151741 329221
rect 151675 329156 151676 329220
rect 151740 329156 151741 329220
rect 151675 329155 151741 329156
rect 142294 328130 142354 329155
rect 141926 328070 142354 328130
rect 151678 328130 151738 329155
rect 151862 328130 151922 329835
rect 152598 329221 152658 333235
rect 153234 331592 153854 334338
rect 152595 329220 152661 329221
rect 152595 329156 152596 329220
rect 152660 329156 152661 329220
rect 152595 329155 152661 329156
rect 151678 328070 151922 328130
rect 88338 309454 88658 309486
rect 88338 309218 88380 309454
rect 88616 309218 88658 309454
rect 88338 309134 88658 309218
rect 88338 308898 88380 309134
rect 88616 308898 88658 309134
rect 88338 308866 88658 308898
rect 119058 309454 119378 309486
rect 119058 309218 119100 309454
rect 119336 309218 119378 309454
rect 119058 309134 119378 309218
rect 119058 308898 119100 309134
rect 119336 308898 119378 309134
rect 119058 308866 119378 308898
rect 149778 309454 150098 309486
rect 149778 309218 149820 309454
rect 150056 309218 150098 309454
rect 149778 309134 150098 309218
rect 149778 308898 149820 309134
rect 150056 308898 150098 309134
rect 149778 308866 150098 308898
rect 103698 291454 104018 291486
rect 103698 291218 103740 291454
rect 103976 291218 104018 291454
rect 103698 291134 104018 291218
rect 103698 290898 103740 291134
rect 103976 290898 104018 291134
rect 103698 290866 104018 290898
rect 134418 291454 134738 291486
rect 134418 291218 134460 291454
rect 134696 291218 134738 291454
rect 134418 291134 134738 291218
rect 134418 290898 134460 291134
rect 134696 290898 134738 291134
rect 134418 290866 134738 290898
rect 88338 273454 88658 273486
rect 88338 273218 88380 273454
rect 88616 273218 88658 273454
rect 88338 273134 88658 273218
rect 88338 272898 88380 273134
rect 88616 272898 88658 273134
rect 88338 272866 88658 272898
rect 119058 273454 119378 273486
rect 119058 273218 119100 273454
rect 119336 273218 119378 273454
rect 119058 273134 119378 273218
rect 119058 272898 119100 273134
rect 119336 272898 119378 273134
rect 119058 272866 119378 272898
rect 149778 273454 150098 273486
rect 149778 273218 149820 273454
rect 150056 273218 150098 273454
rect 149778 273134 150098 273218
rect 149778 272898 149820 273134
rect 150056 272898 150098 273134
rect 149778 272866 150098 272898
rect 103698 255454 104018 255486
rect 103698 255218 103740 255454
rect 103976 255218 104018 255454
rect 103698 255134 104018 255218
rect 103698 254898 103740 255134
rect 103976 254898 104018 255134
rect 103698 254866 104018 254898
rect 134418 255454 134738 255486
rect 134418 255218 134460 255454
rect 134696 255218 134738 255454
rect 134418 255134 134738 255218
rect 134418 254898 134460 255134
rect 134696 254898 134738 255134
rect 134418 254866 134738 254898
rect 83963 241500 84029 241501
rect 83963 241436 83964 241500
rect 84028 241436 84029 241500
rect 83963 241435 84029 241436
rect 82675 234428 82741 234429
rect 82675 234364 82676 234428
rect 82740 234364 82741 234428
rect 82675 234363 82741 234364
rect 81234 226658 81266 226894
rect 81502 226658 81586 226894
rect 81822 226658 81854 226894
rect 81234 226574 81854 226658
rect 81234 226338 81266 226574
rect 81502 226338 81586 226574
rect 81822 226338 81854 226574
rect 81234 190894 81854 226338
rect 81234 190658 81266 190894
rect 81502 190658 81586 190894
rect 81822 190658 81854 190894
rect 81234 190574 81854 190658
rect 81234 190338 81266 190574
rect 81502 190338 81586 190574
rect 81822 190338 81854 190574
rect 81234 176600 81854 190338
rect 84954 230614 85574 239592
rect 84954 230378 84986 230614
rect 85222 230378 85306 230614
rect 85542 230378 85574 230614
rect 84954 230294 85574 230378
rect 84954 230058 84986 230294
rect 85222 230058 85306 230294
rect 85542 230058 85574 230294
rect 84954 194614 85574 230058
rect 84954 194378 84986 194614
rect 85222 194378 85306 194614
rect 85542 194378 85574 194614
rect 84954 194294 85574 194378
rect 84954 194058 84986 194294
rect 85222 194058 85306 194294
rect 85542 194058 85574 194294
rect 84954 176600 85574 194058
rect 91794 237454 92414 239592
rect 91794 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 92414 237454
rect 91794 237134 92414 237218
rect 91794 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 92414 237134
rect 91794 201454 92414 236898
rect 91794 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 92414 201454
rect 91794 201134 92414 201218
rect 91794 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 92414 201134
rect 91794 176600 92414 200898
rect 95514 205174 96134 239592
rect 95514 204938 95546 205174
rect 95782 204938 95866 205174
rect 96102 204938 96134 205174
rect 95514 204854 96134 204938
rect 95514 204618 95546 204854
rect 95782 204618 95866 204854
rect 96102 204618 96134 204854
rect 95514 176600 96134 204618
rect 99234 208894 99854 239592
rect 99234 208658 99266 208894
rect 99502 208658 99586 208894
rect 99822 208658 99854 208894
rect 99234 208574 99854 208658
rect 99234 208338 99266 208574
rect 99502 208338 99586 208574
rect 99822 208338 99854 208574
rect 98315 177580 98381 177581
rect 98315 177516 98316 177580
rect 98380 177516 98381 177580
rect 98315 177515 98381 177516
rect 97027 176900 97093 176901
rect 97027 176836 97028 176900
rect 97092 176836 97093 176900
rect 97027 176835 97093 176836
rect 97030 175130 97090 176835
rect 96960 175070 97090 175130
rect 98318 175130 98378 177515
rect 99234 176600 99854 208338
rect 102954 212614 103574 239592
rect 102954 212378 102986 212614
rect 103222 212378 103306 212614
rect 103542 212378 103574 212614
rect 102954 212294 103574 212378
rect 102954 212058 102986 212294
rect 103222 212058 103306 212294
rect 103542 212058 103574 212294
rect 100707 177580 100773 177581
rect 100707 177516 100708 177580
rect 100772 177516 100773 177580
rect 100707 177515 100773 177516
rect 99419 176492 99485 176493
rect 99419 176428 99420 176492
rect 99484 176428 99485 176492
rect 99419 176427 99485 176428
rect 99422 175130 99482 176427
rect 98318 175070 98380 175130
rect 96960 174494 97020 175070
rect 98320 174494 98380 175070
rect 99408 175070 99482 175130
rect 100710 175130 100770 177515
rect 101995 176764 102061 176765
rect 101995 176700 101996 176764
rect 102060 176700 102061 176764
rect 101995 176699 102061 176700
rect 101998 175130 102058 176699
rect 102954 176600 103574 212058
rect 109794 219454 110414 239592
rect 109794 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 110414 219454
rect 109794 219134 110414 219218
rect 109794 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 110414 219134
rect 109794 183454 110414 218898
rect 109794 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 110414 183454
rect 109794 183134 110414 183218
rect 109794 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 110414 183134
rect 105675 177580 105741 177581
rect 105675 177516 105676 177580
rect 105740 177516 105741 177580
rect 105675 177515 105741 177516
rect 108067 177580 108133 177581
rect 108067 177516 108068 177580
rect 108132 177516 108133 177580
rect 108067 177515 108133 177516
rect 109539 177580 109605 177581
rect 109539 177516 109540 177580
rect 109604 177516 109605 177580
rect 109539 177515 109605 177516
rect 104571 177172 104637 177173
rect 104571 177108 104572 177172
rect 104636 177108 104637 177172
rect 104571 177107 104637 177108
rect 103283 176492 103349 176493
rect 103283 176428 103284 176492
rect 103348 176428 103349 176492
rect 103283 176427 103349 176428
rect 100710 175070 100828 175130
rect 99408 174494 99468 175070
rect 100768 174494 100828 175070
rect 101992 175070 102058 175130
rect 103286 175130 103346 176427
rect 104574 175130 104634 177107
rect 105678 175130 105738 177515
rect 106963 177036 107029 177037
rect 106963 176972 106964 177036
rect 107028 176972 107029 177036
rect 106963 176971 107029 176972
rect 103286 175070 103412 175130
rect 104574 175070 104636 175130
rect 101992 174494 102052 175070
rect 103352 174494 103412 175070
rect 104576 174494 104636 175070
rect 105664 175070 105738 175130
rect 106966 175130 107026 176971
rect 108070 175130 108130 177515
rect 109542 175130 109602 177515
rect 109794 176600 110414 182898
rect 113514 223174 114134 239592
rect 113514 222938 113546 223174
rect 113782 222938 113866 223174
rect 114102 222938 114134 223174
rect 113514 222854 114134 222938
rect 113514 222618 113546 222854
rect 113782 222618 113866 222854
rect 114102 222618 114134 222854
rect 113514 187174 114134 222618
rect 113514 186938 113546 187174
rect 113782 186938 113866 187174
rect 114102 186938 114134 187174
rect 113514 186854 114134 186938
rect 113514 186618 113546 186854
rect 113782 186618 113866 186854
rect 114102 186618 114134 186854
rect 110643 177988 110709 177989
rect 110643 177924 110644 177988
rect 110708 177924 110709 177988
rect 110643 177923 110709 177924
rect 106966 175070 107084 175130
rect 108070 175070 108172 175130
rect 105664 174494 105724 175070
rect 107024 174494 107084 175070
rect 108112 174494 108172 175070
rect 109472 175070 109602 175130
rect 110646 175130 110706 177923
rect 113219 177580 113285 177581
rect 113219 177516 113220 177580
rect 113284 177516 113285 177580
rect 113219 177515 113285 177516
rect 112115 177444 112181 177445
rect 112115 177380 112116 177444
rect 112180 177380 112181 177444
rect 112115 177379 112181 177380
rect 112118 175130 112178 177379
rect 113222 175130 113282 177515
rect 113514 176600 114134 186618
rect 117234 226894 117854 239592
rect 117234 226658 117266 226894
rect 117502 226658 117586 226894
rect 117822 226658 117854 226894
rect 117234 226574 117854 226658
rect 117234 226338 117266 226574
rect 117502 226338 117586 226574
rect 117822 226338 117854 226574
rect 117234 190894 117854 226338
rect 117234 190658 117266 190894
rect 117502 190658 117586 190894
rect 117822 190658 117854 190894
rect 117234 190574 117854 190658
rect 117234 190338 117266 190574
rect 117502 190338 117586 190574
rect 117822 190338 117854 190574
rect 115795 177580 115861 177581
rect 115795 177516 115796 177580
rect 115860 177516 115861 177580
rect 115795 177515 115861 177516
rect 116899 177580 116965 177581
rect 116899 177516 116900 177580
rect 116964 177516 116965 177580
rect 116899 177515 116965 177516
rect 114323 175404 114389 175405
rect 114323 175340 114324 175404
rect 114388 175340 114389 175404
rect 114323 175339 114389 175340
rect 110646 175070 110756 175130
rect 109472 174494 109532 175070
rect 110696 174494 110756 175070
rect 112056 175070 112178 175130
rect 113144 175070 113282 175130
rect 114326 175130 114386 175339
rect 115798 175130 115858 177515
rect 114326 175070 114428 175130
rect 112056 174494 112116 175070
rect 113144 174494 113204 175070
rect 114368 174494 114428 175070
rect 115728 175070 115858 175130
rect 116902 175130 116962 177515
rect 117234 176600 117854 190338
rect 120954 230614 121574 239592
rect 120954 230378 120986 230614
rect 121222 230378 121306 230614
rect 121542 230378 121574 230614
rect 120954 230294 121574 230378
rect 120954 230058 120986 230294
rect 121222 230058 121306 230294
rect 121542 230058 121574 230294
rect 120954 194614 121574 230058
rect 120954 194378 120986 194614
rect 121222 194378 121306 194614
rect 121542 194378 121574 194614
rect 120954 194294 121574 194378
rect 120954 194058 120986 194294
rect 121222 194058 121306 194294
rect 121542 194058 121574 194294
rect 118371 177988 118437 177989
rect 118371 177924 118372 177988
rect 118436 177924 118437 177988
rect 118371 177923 118437 177924
rect 118374 175130 118434 177923
rect 119475 177036 119541 177037
rect 119475 176972 119476 177036
rect 119540 176972 119541 177036
rect 119475 176971 119541 176972
rect 119478 175130 119538 176971
rect 120763 176900 120829 176901
rect 120763 176836 120764 176900
rect 120828 176836 120829 176900
rect 120763 176835 120829 176836
rect 120766 175130 120826 176835
rect 120954 176600 121574 194058
rect 127794 237454 128414 239592
rect 127794 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 128414 237454
rect 127794 237134 128414 237218
rect 127794 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 128414 237134
rect 127794 201454 128414 236898
rect 127794 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 128414 201454
rect 127794 201134 128414 201218
rect 127794 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 128414 201134
rect 123155 177580 123221 177581
rect 123155 177516 123156 177580
rect 123220 177516 123221 177580
rect 123155 177515 123221 177516
rect 121867 175540 121933 175541
rect 121867 175476 121868 175540
rect 121932 175476 121933 175540
rect 121867 175475 121933 175476
rect 121870 175130 121930 175475
rect 123158 175130 123218 177515
rect 127019 177036 127085 177037
rect 127019 176972 127020 177036
rect 127084 176972 127085 177036
rect 127019 176971 127085 176972
rect 124443 176764 124509 176765
rect 124443 176700 124444 176764
rect 124508 176700 124509 176764
rect 124443 176699 124509 176700
rect 124446 175130 124506 176699
rect 125731 175812 125797 175813
rect 125731 175748 125732 175812
rect 125796 175748 125797 175812
rect 125731 175747 125797 175748
rect 125734 175130 125794 175747
rect 127022 175130 127082 176971
rect 127794 176600 128414 200898
rect 131514 205174 132134 239592
rect 131514 204938 131546 205174
rect 131782 204938 131866 205174
rect 132102 204938 132134 205174
rect 131514 204854 132134 204938
rect 131514 204618 131546 204854
rect 131782 204618 131866 204854
rect 132102 204618 132134 204854
rect 130699 176764 130765 176765
rect 130699 176700 130700 176764
rect 130764 176700 130765 176764
rect 130699 176699 130765 176700
rect 128123 176492 128189 176493
rect 128123 176428 128124 176492
rect 128188 176428 128189 176492
rect 128123 176427 128189 176428
rect 128126 175130 128186 176427
rect 129411 175676 129477 175677
rect 129411 175612 129412 175676
rect 129476 175612 129477 175676
rect 129411 175611 129477 175612
rect 116902 175070 117012 175130
rect 115728 174494 115788 175070
rect 116952 174494 117012 175070
rect 118312 175070 118434 175130
rect 119400 175070 119538 175130
rect 120760 175070 120826 175130
rect 121848 175070 121930 175130
rect 123072 175070 123218 175130
rect 124432 175070 124506 175130
rect 125656 175070 125794 175130
rect 127016 175070 127082 175130
rect 128104 175070 128186 175130
rect 129414 175130 129474 175611
rect 130702 175130 130762 176699
rect 131514 176600 132134 204618
rect 135234 208894 135854 239592
rect 135234 208658 135266 208894
rect 135502 208658 135586 208894
rect 135822 208658 135854 208894
rect 135234 208574 135854 208658
rect 135234 208338 135266 208574
rect 135502 208338 135586 208574
rect 135822 208338 135854 208574
rect 133091 177580 133157 177581
rect 133091 177516 133092 177580
rect 133156 177516 133157 177580
rect 133091 177515 133157 177516
rect 134379 177580 134445 177581
rect 134379 177516 134380 177580
rect 134444 177516 134445 177580
rect 134379 177515 134445 177516
rect 132355 176764 132421 176765
rect 132355 176700 132356 176764
rect 132420 176700 132421 176764
rect 132355 176699 132421 176700
rect 132358 175130 132418 176699
rect 129414 175070 129524 175130
rect 118312 174494 118372 175070
rect 119400 174494 119460 175070
rect 120760 174494 120820 175070
rect 121848 174494 121908 175070
rect 123072 174494 123132 175070
rect 124432 174494 124492 175070
rect 125656 174494 125716 175070
rect 127016 174494 127076 175070
rect 128104 174494 128164 175070
rect 129464 174494 129524 175070
rect 130688 175070 130762 175130
rect 132048 175070 132418 175130
rect 133094 175130 133154 177515
rect 134382 175130 134442 177515
rect 135234 176600 135854 208338
rect 138954 212614 139574 239592
rect 138954 212378 138986 212614
rect 139222 212378 139306 212614
rect 139542 212378 139574 212614
rect 138954 212294 139574 212378
rect 138954 212058 138986 212294
rect 139222 212058 139306 212294
rect 139542 212058 139574 212294
rect 136035 176764 136101 176765
rect 136035 176700 136036 176764
rect 136100 176700 136101 176764
rect 136035 176699 136101 176700
rect 136038 175130 136098 176699
rect 138954 176600 139574 212058
rect 145794 219454 146414 239592
rect 145794 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 146414 219454
rect 145794 219134 146414 219218
rect 145794 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 146414 219134
rect 145794 183454 146414 218898
rect 145794 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 146414 183454
rect 145794 183134 146414 183218
rect 145794 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 146414 183134
rect 145794 176600 146414 182898
rect 149514 223174 150134 239592
rect 149514 222938 149546 223174
rect 149782 222938 149866 223174
rect 150102 222938 150134 223174
rect 149514 222854 150134 222938
rect 149514 222618 149546 222854
rect 149782 222618 149866 222854
rect 150102 222618 150134 222854
rect 149514 187174 150134 222618
rect 149514 186938 149546 187174
rect 149782 186938 149866 187174
rect 150102 186938 150134 187174
rect 149514 186854 150134 186938
rect 149514 186618 149546 186854
rect 149782 186618 149866 186854
rect 150102 186618 150134 186854
rect 148179 177580 148245 177581
rect 148179 177516 148180 177580
rect 148244 177516 148245 177580
rect 148179 177515 148245 177516
rect 133094 175070 133196 175130
rect 130688 174494 130748 175070
rect 132048 174494 132108 175070
rect 133136 174494 133196 175070
rect 134360 175070 134442 175130
rect 135720 175070 136098 175130
rect 148182 175130 148242 177515
rect 149514 176600 150134 186618
rect 153234 226894 153854 239592
rect 154070 237421 154130 369003
rect 154622 242045 154682 411299
rect 156954 410614 157574 446058
rect 156954 410378 156986 410614
rect 157222 410378 157306 410614
rect 157542 410378 157574 410614
rect 156954 410294 157574 410378
rect 156954 410058 156986 410294
rect 157222 410058 157306 410294
rect 157542 410058 157574 410294
rect 156954 374614 157574 410058
rect 158667 380220 158733 380221
rect 158667 380156 158668 380220
rect 158732 380156 158733 380220
rect 158667 380155 158733 380156
rect 156954 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 157574 374614
rect 156954 374294 157574 374378
rect 156954 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 157574 374294
rect 156459 343908 156525 343909
rect 156459 343844 156460 343908
rect 156524 343844 156525 343908
rect 156459 343843 156525 343844
rect 156462 325710 156522 343843
rect 156954 338614 157574 374058
rect 157747 341596 157813 341597
rect 157747 341532 157748 341596
rect 157812 341532 157813 341596
rect 157747 341531 157813 341532
rect 157750 340781 157810 341531
rect 157747 340780 157813 340781
rect 157747 340716 157748 340780
rect 157812 340716 157813 340780
rect 157747 340715 157813 340716
rect 158483 340780 158549 340781
rect 158483 340716 158484 340780
rect 158548 340716 158549 340780
rect 158483 340715 158549 340716
rect 156954 338378 156986 338614
rect 157222 338378 157306 338614
rect 157542 338378 157574 338614
rect 156954 338294 157574 338378
rect 156954 338058 156986 338294
rect 157222 338058 157306 338294
rect 157542 338058 157574 338294
rect 156954 331592 157574 338058
rect 157747 331532 157813 331533
rect 157747 331468 157748 331532
rect 157812 331468 157813 331532
rect 157747 331467 157813 331468
rect 157195 329764 157261 329765
rect 157195 329700 157196 329764
rect 157260 329700 157261 329764
rect 157195 329699 157261 329700
rect 156462 325650 156890 325710
rect 156830 312629 156890 325650
rect 157198 320789 157258 329699
rect 157750 325413 157810 331467
rect 157747 325412 157813 325413
rect 157747 325348 157748 325412
rect 157812 325348 157813 325412
rect 157747 325347 157813 325348
rect 157750 324461 157810 325347
rect 157747 324460 157813 324461
rect 157747 324396 157748 324460
rect 157812 324396 157813 324460
rect 157747 324395 157813 324396
rect 157195 320788 157261 320789
rect 157195 320724 157196 320788
rect 157260 320724 157261 320788
rect 157195 320723 157261 320724
rect 156827 312628 156893 312629
rect 156827 312564 156828 312628
rect 156892 312564 156893 312628
rect 156827 312563 156893 312564
rect 157195 310452 157261 310453
rect 157195 310388 157196 310452
rect 157260 310388 157261 310452
rect 157195 310387 157261 310388
rect 157198 273730 157258 310387
rect 158486 278085 158546 340715
rect 158670 322149 158730 380155
rect 158851 340236 158917 340237
rect 158851 340172 158852 340236
rect 158916 340172 158917 340236
rect 158851 340171 158917 340172
rect 158667 322148 158733 322149
rect 158667 322084 158668 322148
rect 158732 322084 158733 322148
rect 158667 322083 158733 322084
rect 158854 309773 158914 340171
rect 158851 309772 158917 309773
rect 158851 309708 158852 309772
rect 158916 309708 158917 309772
rect 158851 309707 158917 309708
rect 159035 305828 159101 305829
rect 159035 305764 159036 305828
rect 159100 305764 159101 305828
rect 159035 305763 159101 305764
rect 159038 298213 159098 305763
rect 159035 298212 159101 298213
rect 159035 298148 159036 298212
rect 159100 298148 159101 298212
rect 159035 298147 159101 298148
rect 159955 295356 160021 295357
rect 159955 295292 159956 295356
rect 160020 295292 160021 295356
rect 159955 295291 160021 295292
rect 159219 288692 159285 288693
rect 159219 288628 159220 288692
rect 159284 288628 159285 288692
rect 159219 288627 159285 288628
rect 158483 278084 158549 278085
rect 158483 278020 158484 278084
rect 158548 278020 158549 278084
rect 158483 278019 158549 278020
rect 158486 277813 158546 278019
rect 158483 277812 158549 277813
rect 158483 277748 158484 277812
rect 158548 277748 158549 277812
rect 158483 277747 158549 277748
rect 157198 273670 157442 273730
rect 156827 262852 156893 262853
rect 156827 262788 156828 262852
rect 156892 262788 156893 262852
rect 156827 262787 156893 262788
rect 156830 258090 156890 262787
rect 156462 258030 156890 258090
rect 154619 242044 154685 242045
rect 154619 241980 154620 242044
rect 154684 241980 154685 242044
rect 154619 241979 154685 241980
rect 155723 240140 155789 240141
rect 155723 240076 155724 240140
rect 155788 240076 155789 240140
rect 155723 240075 155789 240076
rect 154067 237420 154133 237421
rect 154067 237356 154068 237420
rect 154132 237356 154133 237420
rect 154067 237355 154133 237356
rect 153234 226658 153266 226894
rect 153502 226658 153586 226894
rect 153822 226658 153854 226894
rect 153234 226574 153854 226658
rect 153234 226338 153266 226574
rect 153502 226338 153586 226574
rect 153822 226338 153854 226574
rect 153234 190894 153854 226338
rect 153234 190658 153266 190894
rect 153502 190658 153586 190894
rect 153822 190658 153854 190894
rect 153234 190574 153854 190658
rect 153234 190338 153266 190574
rect 153502 190338 153586 190574
rect 153822 190338 153854 190574
rect 153234 176600 153854 190338
rect 155726 184381 155786 240075
rect 156462 235789 156522 258030
rect 156827 243540 156893 243541
rect 156827 243476 156828 243540
rect 156892 243476 156893 243540
rect 156827 243475 156893 243476
rect 156830 241090 156890 243475
rect 156646 241030 156890 241090
rect 156646 238645 156706 241030
rect 157382 240141 157442 273670
rect 157931 268428 157997 268429
rect 157931 268364 157932 268428
rect 157996 268364 157997 268428
rect 157931 268363 157997 268364
rect 157379 240140 157445 240141
rect 157379 240076 157380 240140
rect 157444 240076 157445 240140
rect 157379 240075 157445 240076
rect 156643 238644 156709 238645
rect 156643 238580 156644 238644
rect 156708 238580 156709 238644
rect 156643 238579 156709 238580
rect 156459 235788 156525 235789
rect 156459 235724 156460 235788
rect 156524 235724 156525 235788
rect 156459 235723 156525 235724
rect 156954 230614 157574 239592
rect 156954 230378 156986 230614
rect 157222 230378 157306 230614
rect 157542 230378 157574 230614
rect 156954 230294 157574 230378
rect 156954 230058 156986 230294
rect 157222 230058 157306 230294
rect 157542 230058 157574 230294
rect 156954 194614 157574 230058
rect 157934 227493 157994 268363
rect 157931 227492 157997 227493
rect 157931 227428 157932 227492
rect 157996 227428 157997 227492
rect 157931 227427 157997 227428
rect 159222 207637 159282 288627
rect 159958 260813 160018 295291
rect 159955 260812 160021 260813
rect 159955 260748 159956 260812
rect 160020 260748 160021 260812
rect 159955 260747 160021 260748
rect 160694 241229 160754 449923
rect 160875 338060 160941 338061
rect 160875 337996 160876 338060
rect 160940 337996 160941 338060
rect 160875 337995 160941 337996
rect 160878 275229 160938 337995
rect 160875 275228 160941 275229
rect 160875 275164 160876 275228
rect 160940 275164 160941 275228
rect 160875 275163 160941 275164
rect 161982 271829 162042 518875
rect 163794 489454 164414 524898
rect 163794 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 164414 489454
rect 163794 489134 164414 489218
rect 163794 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 164414 489134
rect 163794 453454 164414 488898
rect 163794 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 164414 453454
rect 163794 453134 164414 453218
rect 163794 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 164414 453134
rect 163794 417454 164414 452898
rect 163794 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 164414 417454
rect 163794 417134 164414 417218
rect 163794 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 164414 417134
rect 163794 381454 164414 416898
rect 163794 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 164414 381454
rect 163794 381134 164414 381218
rect 163794 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 164414 381134
rect 163794 345454 164414 380898
rect 167514 673174 168134 707162
rect 167514 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 168134 673174
rect 167514 672854 168134 672938
rect 167514 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 168134 672854
rect 167514 637174 168134 672618
rect 167514 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 168134 637174
rect 167514 636854 168134 636938
rect 167514 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 168134 636854
rect 167514 601174 168134 636618
rect 167514 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 168134 601174
rect 167514 600854 168134 600938
rect 167514 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 168134 600854
rect 167514 565174 168134 600618
rect 167514 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 168134 565174
rect 167514 564854 168134 564938
rect 167514 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 168134 564854
rect 167514 529174 168134 564618
rect 171234 676894 171854 709082
rect 171234 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 171854 676894
rect 171234 676574 171854 676658
rect 171234 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 171854 676574
rect 171234 640894 171854 676338
rect 171234 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 171854 640894
rect 171234 640574 171854 640658
rect 171234 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 171854 640574
rect 171234 604894 171854 640338
rect 171234 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 171854 604894
rect 171234 604574 171854 604658
rect 171234 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 171854 604574
rect 171234 568894 171854 604338
rect 171234 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 171854 568894
rect 171234 568574 171854 568658
rect 171234 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 171854 568574
rect 170259 546684 170325 546685
rect 170259 546620 170260 546684
rect 170324 546620 170325 546684
rect 170259 546619 170325 546620
rect 167514 528938 167546 529174
rect 167782 528938 167866 529174
rect 168102 528938 168134 529174
rect 167514 528854 168134 528938
rect 167514 528618 167546 528854
rect 167782 528618 167866 528854
rect 168102 528618 168134 528854
rect 167514 493174 168134 528618
rect 168971 523700 169037 523701
rect 168971 523636 168972 523700
rect 169036 523636 169037 523700
rect 168971 523635 169037 523636
rect 167514 492938 167546 493174
rect 167782 492938 167866 493174
rect 168102 492938 168134 493174
rect 167514 492854 168134 492938
rect 167514 492618 167546 492854
rect 167782 492618 167866 492854
rect 168102 492618 168134 492854
rect 167514 457174 168134 492618
rect 167514 456938 167546 457174
rect 167782 456938 167866 457174
rect 168102 456938 168134 457174
rect 167514 456854 168134 456938
rect 167514 456618 167546 456854
rect 167782 456618 167866 456854
rect 168102 456618 168134 456854
rect 167514 421174 168134 456618
rect 167514 420938 167546 421174
rect 167782 420938 167866 421174
rect 168102 420938 168134 421174
rect 167514 420854 168134 420938
rect 167514 420618 167546 420854
rect 167782 420618 167866 420854
rect 168102 420618 168134 420854
rect 167514 385174 168134 420618
rect 167514 384938 167546 385174
rect 167782 384938 167866 385174
rect 168102 384938 168134 385174
rect 167514 384854 168134 384938
rect 167514 384618 167546 384854
rect 167782 384618 167866 384854
rect 168102 384618 168134 384854
rect 166395 374644 166461 374645
rect 166395 374580 166396 374644
rect 166460 374580 166461 374644
rect 166395 374579 166461 374580
rect 166211 367300 166277 367301
rect 166211 367236 166212 367300
rect 166276 367236 166277 367300
rect 166211 367235 166277 367236
rect 163794 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 164414 345454
rect 163794 345134 164414 345218
rect 163794 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 164414 345134
rect 163794 309454 164414 344898
rect 166214 328405 166274 367235
rect 166398 360093 166458 374579
rect 166395 360092 166461 360093
rect 166395 360028 166396 360092
rect 166460 360028 166461 360092
rect 166395 360027 166461 360028
rect 166211 328404 166277 328405
rect 166211 328340 166212 328404
rect 166276 328340 166277 328404
rect 166211 328339 166277 328340
rect 166398 319429 166458 360027
rect 167514 349174 168134 384618
rect 167514 348938 167546 349174
rect 167782 348938 167866 349174
rect 168102 348938 168134 349174
rect 167514 348854 168134 348938
rect 167514 348618 167546 348854
rect 167782 348618 167866 348854
rect 168102 348618 168134 348854
rect 166395 319428 166461 319429
rect 166395 319364 166396 319428
rect 166460 319364 166461 319428
rect 166395 319363 166461 319364
rect 166211 314668 166277 314669
rect 166211 314604 166212 314668
rect 166276 314604 166277 314668
rect 166211 314603 166277 314604
rect 163794 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 164414 309454
rect 163794 309134 164414 309218
rect 163794 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 164414 309134
rect 163794 273454 164414 308898
rect 163794 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 164414 273454
rect 163794 273134 164414 273218
rect 163794 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 164414 273134
rect 161979 271828 162045 271829
rect 161979 271764 161980 271828
rect 162044 271764 162045 271828
rect 161979 271763 162045 271764
rect 161979 260676 162045 260677
rect 161979 260612 161980 260676
rect 162044 260612 162045 260676
rect 161979 260611 162045 260612
rect 160691 241228 160757 241229
rect 160691 241164 160692 241228
rect 160756 241164 160757 241228
rect 160691 241163 160757 241164
rect 159219 207636 159285 207637
rect 159219 207572 159220 207636
rect 159284 207572 159285 207636
rect 159219 207571 159285 207572
rect 156954 194378 156986 194614
rect 157222 194378 157306 194614
rect 157542 194378 157574 194614
rect 156954 194294 157574 194378
rect 156954 194058 156986 194294
rect 157222 194058 157306 194294
rect 157542 194058 157574 194294
rect 155723 184380 155789 184381
rect 155723 184316 155724 184380
rect 155788 184316 155789 184380
rect 155723 184315 155789 184316
rect 156954 176600 157574 194058
rect 161982 180709 162042 260611
rect 163794 237454 164414 272898
rect 165659 242860 165725 242861
rect 165659 242796 165660 242860
rect 165724 242796 165725 242860
rect 165659 242795 165725 242796
rect 163794 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 164414 237454
rect 163794 237134 164414 237218
rect 163794 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 164414 237134
rect 163794 201454 164414 236898
rect 163794 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 164414 201454
rect 163794 201134 164414 201218
rect 163794 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 164414 201134
rect 161979 180708 162045 180709
rect 161979 180644 161980 180708
rect 162044 180644 162045 180708
rect 161979 180643 162045 180644
rect 158851 176764 158917 176765
rect 158851 176700 158852 176764
rect 158916 176700 158917 176764
rect 158851 176699 158917 176700
rect 158854 175130 158914 176699
rect 163794 176600 164414 200898
rect 148182 175070 148292 175130
rect 134360 174494 134420 175070
rect 135720 174494 135780 175070
rect 148232 174494 148292 175070
rect 158840 175070 158914 175130
rect 158840 174494 158900 175070
rect 69072 165454 69420 165486
rect 69072 165218 69128 165454
rect 69364 165218 69420 165454
rect 69072 165134 69420 165218
rect 69072 164898 69128 165134
rect 69364 164898 69420 165134
rect 69072 164866 69420 164898
rect 164136 165454 164484 165486
rect 164136 165218 164192 165454
rect 164428 165218 164484 165454
rect 164136 165134 164484 165218
rect 164136 164898 164192 165134
rect 164428 164898 164484 165134
rect 164136 164866 164484 164898
rect 69752 147454 70100 147486
rect 69752 147218 69808 147454
rect 70044 147218 70100 147454
rect 69752 147134 70100 147218
rect 69752 146898 69808 147134
rect 70044 146898 70100 147134
rect 69752 146866 70100 146898
rect 163456 147454 163804 147486
rect 163456 147218 163512 147454
rect 163748 147218 163804 147454
rect 163456 147134 163804 147218
rect 163456 146898 163512 147134
rect 163748 146898 163804 147134
rect 163456 146866 163804 146898
rect 69072 129454 69420 129486
rect 69072 129218 69128 129454
rect 69364 129218 69420 129454
rect 69072 129134 69420 129218
rect 69072 128898 69128 129134
rect 69364 128898 69420 129134
rect 69072 128866 69420 128898
rect 164136 129454 164484 129486
rect 164136 129218 164192 129454
rect 164428 129218 164484 129454
rect 164136 129134 164484 129218
rect 164136 128898 164192 129134
rect 164428 128898 164484 129134
rect 164136 128866 164484 128898
rect 69752 111454 70100 111486
rect 69752 111218 69808 111454
rect 70044 111218 70100 111454
rect 69752 111134 70100 111218
rect 69752 110898 69808 111134
rect 70044 110898 70100 111134
rect 69752 110866 70100 110898
rect 163456 111454 163804 111486
rect 163456 111218 163512 111454
rect 163748 111218 163804 111454
rect 163456 111134 163804 111218
rect 163456 110898 163512 111134
rect 163748 110898 163804 111134
rect 163456 110866 163804 110898
rect 74656 94890 74716 95200
rect 84312 94890 84372 95200
rect 85536 94890 85596 95200
rect 86624 94890 86684 95200
rect 87984 94890 88044 95200
rect 88936 94890 88996 95200
rect 74656 94830 74826 94890
rect 84312 94830 84394 94890
rect 85536 94830 85866 94890
rect 86624 94830 86786 94890
rect 87984 94830 88074 94890
rect 73794 75454 74414 93100
rect 74766 92445 74826 94830
rect 74763 92444 74829 92445
rect 74763 92380 74764 92444
rect 74828 92380 74829 92444
rect 74763 92379 74829 92380
rect 73794 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 74414 75454
rect 73794 75134 74414 75218
rect 73794 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 74414 75134
rect 73794 39454 74414 74898
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 67771 25668 67837 25669
rect 67771 25604 67772 25668
rect 67836 25604 67837 25668
rect 67771 25603 67837 25604
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -1894 74414 -902
rect 77514 79174 78134 93100
rect 77514 78938 77546 79174
rect 77782 78938 77866 79174
rect 78102 78938 78134 79174
rect 77514 78854 78134 78938
rect 77514 78618 77546 78854
rect 77782 78618 77866 78854
rect 78102 78618 78134 78854
rect 77514 43174 78134 78618
rect 77514 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 78134 43174
rect 77514 42854 78134 42938
rect 77514 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 78134 42854
rect 77514 7174 78134 42618
rect 77514 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 78134 7174
rect 77514 6854 78134 6938
rect 77514 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 78134 6854
rect 77514 -2266 78134 6618
rect 77514 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 78134 -2266
rect 77514 -2586 78134 -2502
rect 77514 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 78134 -2586
rect 77514 -3814 78134 -2822
rect 81234 82894 81854 93100
rect 84334 91221 84394 94830
rect 84331 91220 84397 91221
rect 84331 91156 84332 91220
rect 84396 91156 84397 91220
rect 84331 91155 84397 91156
rect 81234 82658 81266 82894
rect 81502 82658 81586 82894
rect 81822 82658 81854 82894
rect 81234 82574 81854 82658
rect 81234 82338 81266 82574
rect 81502 82338 81586 82574
rect 81822 82338 81854 82574
rect 81234 46894 81854 82338
rect 81234 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 81854 46894
rect 81234 46574 81854 46658
rect 81234 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 81854 46574
rect 81234 10894 81854 46338
rect 81234 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 81854 10894
rect 81234 10574 81854 10658
rect 81234 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 81854 10574
rect 81234 -4186 81854 10338
rect 81234 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 81854 -4186
rect 81234 -4506 81854 -4422
rect 81234 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 81854 -4506
rect 81234 -5734 81854 -4742
rect 84954 86614 85574 93100
rect 85806 91357 85866 94830
rect 85803 91356 85869 91357
rect 85803 91292 85804 91356
rect 85868 91292 85869 91356
rect 85803 91291 85869 91292
rect 86726 91221 86786 94830
rect 88014 92173 88074 94830
rect 88934 94830 88996 94890
rect 90160 94890 90220 95200
rect 91384 94890 91444 95200
rect 90160 94830 90282 94890
rect 88011 92172 88077 92173
rect 88011 92108 88012 92172
rect 88076 92108 88077 92172
rect 88011 92107 88077 92108
rect 88934 91221 88994 94830
rect 90222 91221 90282 94830
rect 91326 94830 91444 94890
rect 92472 94890 92532 95200
rect 93832 94890 93892 95200
rect 94920 94890 94980 95200
rect 96008 94890 96068 95200
rect 96688 94890 96748 95200
rect 92472 94830 92674 94890
rect 93832 94830 93962 94890
rect 94920 94830 95066 94890
rect 96008 94830 96354 94890
rect 91326 92037 91386 94830
rect 91323 92036 91389 92037
rect 91323 91972 91324 92036
rect 91388 91972 91389 92036
rect 91323 91971 91389 91972
rect 86723 91220 86789 91221
rect 86723 91156 86724 91220
rect 86788 91156 86789 91220
rect 86723 91155 86789 91156
rect 88931 91220 88997 91221
rect 88931 91156 88932 91220
rect 88996 91156 88997 91220
rect 88931 91155 88997 91156
rect 90219 91220 90285 91221
rect 90219 91156 90220 91220
rect 90284 91156 90285 91220
rect 90219 91155 90285 91156
rect 84954 86378 84986 86614
rect 85222 86378 85306 86614
rect 85542 86378 85574 86614
rect 84954 86294 85574 86378
rect 84954 86058 84986 86294
rect 85222 86058 85306 86294
rect 85542 86058 85574 86294
rect 84954 50614 85574 86058
rect 84954 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 85574 50614
rect 84954 50294 85574 50378
rect 84954 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 85574 50294
rect 84954 14614 85574 50058
rect 84954 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 85574 14614
rect 84954 14294 85574 14378
rect 84954 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 85574 14294
rect 66954 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 67574 -7066
rect 66954 -7386 67574 -7302
rect 66954 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 67574 -7386
rect 66954 -7654 67574 -7622
rect 84954 -6106 85574 14058
rect 91794 57454 92414 93100
rect 92614 91221 92674 94830
rect 93902 91221 93962 94830
rect 95006 91357 95066 94830
rect 95003 91356 95069 91357
rect 95003 91292 95004 91356
rect 95068 91292 95069 91356
rect 95003 91291 95069 91292
rect 92611 91220 92677 91221
rect 92611 91156 92612 91220
rect 92676 91156 92677 91220
rect 92611 91155 92677 91156
rect 93899 91220 93965 91221
rect 93899 91156 93900 91220
rect 93964 91156 93965 91220
rect 93899 91155 93965 91156
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -1306 92414 20898
rect 91794 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 92414 -1306
rect 91794 -1626 92414 -1542
rect 91794 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 92414 -1626
rect 91794 -1894 92414 -1862
rect 95514 61174 96134 93100
rect 96294 91221 96354 94830
rect 96662 94830 96748 94890
rect 97096 94890 97156 95200
rect 98048 94890 98108 95200
rect 98456 94890 98516 95200
rect 99136 94890 99196 95200
rect 99544 94890 99604 95200
rect 100632 94890 100692 95200
rect 97096 94830 97274 94890
rect 98048 94830 98194 94890
rect 98456 94830 98562 94890
rect 99136 94830 99298 94890
rect 99544 94830 100034 94890
rect 96662 91221 96722 94830
rect 97214 92445 97274 94830
rect 97211 92444 97277 92445
rect 97211 92380 97212 92444
rect 97276 92380 97277 92444
rect 97211 92379 97277 92380
rect 98134 91221 98194 94830
rect 98502 91357 98562 94830
rect 99238 93805 99298 94830
rect 99235 93804 99301 93805
rect 99235 93740 99236 93804
rect 99300 93740 99301 93804
rect 99235 93739 99301 93740
rect 98499 91356 98565 91357
rect 98499 91292 98500 91356
rect 98564 91292 98565 91356
rect 98499 91291 98565 91292
rect 96291 91220 96357 91221
rect 96291 91156 96292 91220
rect 96356 91156 96357 91220
rect 96291 91155 96357 91156
rect 96659 91220 96725 91221
rect 96659 91156 96660 91220
rect 96724 91156 96725 91220
rect 96659 91155 96725 91156
rect 98131 91220 98197 91221
rect 98131 91156 98132 91220
rect 98196 91156 98197 91220
rect 98131 91155 98197 91156
rect 95514 60938 95546 61174
rect 95782 60938 95866 61174
rect 96102 60938 96134 61174
rect 95514 60854 96134 60938
rect 95514 60618 95546 60854
rect 95782 60618 95866 60854
rect 96102 60618 96134 60854
rect 95514 25174 96134 60618
rect 95514 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 96134 25174
rect 95514 24854 96134 24938
rect 95514 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 96134 24854
rect 95514 -3226 96134 24618
rect 95514 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 96134 -3226
rect 95514 -3546 96134 -3462
rect 95514 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 96134 -3546
rect 95514 -3814 96134 -3782
rect 99234 64894 99854 93100
rect 99974 92445 100034 94830
rect 100526 94830 100692 94890
rect 100768 94890 100828 95200
rect 101856 94890 101916 95200
rect 100768 94830 100954 94890
rect 99971 92444 100037 92445
rect 99971 92380 99972 92444
rect 100036 92380 100037 92444
rect 99971 92379 100037 92380
rect 100526 91221 100586 94830
rect 100894 93941 100954 94830
rect 101814 94830 101916 94890
rect 101992 94890 102052 95200
rect 102944 94890 103004 95200
rect 101992 94830 102058 94890
rect 100891 93940 100957 93941
rect 100891 93876 100892 93940
rect 100956 93876 100957 93940
rect 100891 93875 100957 93876
rect 101814 91221 101874 94830
rect 101998 91629 102058 94830
rect 102918 94830 103004 94890
rect 103216 94890 103276 95200
rect 103216 94830 103346 94890
rect 102918 93870 102978 94830
rect 102734 93810 102978 93870
rect 102734 92445 102794 93810
rect 103286 93261 103346 94830
rect 104304 94754 104364 95200
rect 104206 94694 104364 94754
rect 104440 94754 104500 95200
rect 105392 94754 105452 95200
rect 105664 94754 105724 95200
rect 106480 94754 106540 95200
rect 104440 94694 104634 94754
rect 105392 94694 105554 94754
rect 105664 94694 105738 94754
rect 103283 93260 103349 93261
rect 103283 93196 103284 93260
rect 103348 93196 103349 93260
rect 103283 93195 103349 93196
rect 102731 92444 102797 92445
rect 102731 92380 102732 92444
rect 102796 92380 102797 92444
rect 102731 92379 102797 92380
rect 101995 91628 102061 91629
rect 101995 91564 101996 91628
rect 102060 91564 102061 91628
rect 101995 91563 102061 91564
rect 100523 91220 100589 91221
rect 100523 91156 100524 91220
rect 100588 91156 100589 91220
rect 100523 91155 100589 91156
rect 101811 91220 101877 91221
rect 101811 91156 101812 91220
rect 101876 91156 101877 91220
rect 101811 91155 101877 91156
rect 99234 64658 99266 64894
rect 99502 64658 99586 64894
rect 99822 64658 99854 64894
rect 99234 64574 99854 64658
rect 99234 64338 99266 64574
rect 99502 64338 99586 64574
rect 99822 64338 99854 64574
rect 99234 28894 99854 64338
rect 99234 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 99854 28894
rect 99234 28574 99854 28658
rect 99234 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 99854 28574
rect 99234 -5146 99854 28338
rect 99234 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 99854 -5146
rect 99234 -5466 99854 -5382
rect 99234 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 99854 -5466
rect 99234 -5734 99854 -5702
rect 102954 68614 103574 93100
rect 104206 91221 104266 94694
rect 104574 91221 104634 94694
rect 105494 91221 105554 94694
rect 105678 91221 105738 94694
rect 106414 94694 106540 94754
rect 106616 94754 106676 95200
rect 107704 94754 107764 95200
rect 108112 94754 108172 95200
rect 106616 94694 106842 94754
rect 106414 91221 106474 94694
rect 106782 92309 106842 94694
rect 107702 94694 107764 94754
rect 108070 94694 108172 94754
rect 109064 94754 109124 95200
rect 109472 94754 109532 95200
rect 110152 94754 110212 95200
rect 110696 94754 110756 95200
rect 111240 94754 111300 95200
rect 109064 94694 109234 94754
rect 109472 94694 109602 94754
rect 106779 92308 106845 92309
rect 106779 92244 106780 92308
rect 106844 92244 106845 92308
rect 106779 92243 106845 92244
rect 107702 91221 107762 94694
rect 108070 92445 108130 94694
rect 108067 92444 108133 92445
rect 108067 92380 108068 92444
rect 108132 92380 108133 92444
rect 108067 92379 108133 92380
rect 109174 91765 109234 94694
rect 109171 91764 109237 91765
rect 109171 91700 109172 91764
rect 109236 91700 109237 91764
rect 109171 91699 109237 91700
rect 109542 91221 109602 94694
rect 110094 94694 110212 94754
rect 110646 94694 110756 94754
rect 111198 94694 111300 94754
rect 111920 94754 111980 95200
rect 112328 94754 112388 95200
rect 113144 94757 113204 95200
rect 113688 94890 113748 95200
rect 114368 94890 114428 95200
rect 113406 94830 113748 94890
rect 114326 94830 114428 94890
rect 114776 94890 114836 95200
rect 115456 94890 115516 95200
rect 115864 94890 115924 95200
rect 114776 94830 114938 94890
rect 111920 94694 111994 94754
rect 110094 93533 110154 94694
rect 110091 93532 110157 93533
rect 110091 93468 110092 93532
rect 110156 93468 110157 93532
rect 110091 93467 110157 93468
rect 104203 91220 104269 91221
rect 104203 91156 104204 91220
rect 104268 91156 104269 91220
rect 104203 91155 104269 91156
rect 104571 91220 104637 91221
rect 104571 91156 104572 91220
rect 104636 91156 104637 91220
rect 104571 91155 104637 91156
rect 105491 91220 105557 91221
rect 105491 91156 105492 91220
rect 105556 91156 105557 91220
rect 105491 91155 105557 91156
rect 105675 91220 105741 91221
rect 105675 91156 105676 91220
rect 105740 91156 105741 91220
rect 105675 91155 105741 91156
rect 106411 91220 106477 91221
rect 106411 91156 106412 91220
rect 106476 91156 106477 91220
rect 106411 91155 106477 91156
rect 107699 91220 107765 91221
rect 107699 91156 107700 91220
rect 107764 91156 107765 91220
rect 107699 91155 107765 91156
rect 109539 91220 109605 91221
rect 109539 91156 109540 91220
rect 109604 91156 109605 91220
rect 109539 91155 109605 91156
rect 102954 68378 102986 68614
rect 103222 68378 103306 68614
rect 103542 68378 103574 68614
rect 102954 68294 103574 68378
rect 102954 68058 102986 68294
rect 103222 68058 103306 68294
rect 103542 68058 103574 68294
rect 102954 32614 103574 68058
rect 102954 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 103574 32614
rect 102954 32294 103574 32378
rect 102954 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 103574 32294
rect 84954 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 85574 -6106
rect 84954 -6426 85574 -6342
rect 84954 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 85574 -6426
rect 84954 -7654 85574 -6662
rect 102954 -7066 103574 32058
rect 109794 75454 110414 93100
rect 110646 91357 110706 94694
rect 110643 91356 110709 91357
rect 110643 91292 110644 91356
rect 110708 91292 110709 91356
rect 110643 91291 110709 91292
rect 111198 91221 111258 94694
rect 111934 91221 111994 94694
rect 112302 94694 112388 94754
rect 113141 94756 113207 94757
rect 112302 91221 112362 94694
rect 113141 94692 113142 94756
rect 113206 94692 113207 94756
rect 113141 94691 113207 94692
rect 113406 93870 113466 94830
rect 113222 93810 113466 93870
rect 113222 91357 113282 93810
rect 113219 91356 113285 91357
rect 113219 91292 113220 91356
rect 113284 91292 113285 91356
rect 113219 91291 113285 91292
rect 111195 91220 111261 91221
rect 111195 91156 111196 91220
rect 111260 91156 111261 91220
rect 111195 91155 111261 91156
rect 111931 91220 111997 91221
rect 111931 91156 111932 91220
rect 111996 91156 111997 91220
rect 111931 91155 111997 91156
rect 112299 91220 112365 91221
rect 112299 91156 112300 91220
rect 112364 91156 112365 91220
rect 112299 91155 112365 91156
rect 109794 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 110414 75454
rect 109794 75134 110414 75218
rect 109794 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 110414 75134
rect 109794 39454 110414 74898
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -1894 110414 -902
rect 113514 79174 114134 93100
rect 114326 91221 114386 94830
rect 114878 91221 114938 94830
rect 115430 94830 115516 94890
rect 115798 94830 115924 94890
rect 116680 94890 116740 95200
rect 117088 94890 117148 95200
rect 116680 94830 116778 94890
rect 115430 91357 115490 94830
rect 115798 91357 115858 94830
rect 116718 92445 116778 94830
rect 117086 94830 117148 94890
rect 117904 94890 117964 95200
rect 118176 94890 118236 95200
rect 119400 94890 119460 95200
rect 117904 94830 118066 94890
rect 118176 94830 118250 94890
rect 116715 92444 116781 92445
rect 116715 92380 116716 92444
rect 116780 92380 116781 92444
rect 116715 92379 116781 92380
rect 115427 91356 115493 91357
rect 115427 91292 115428 91356
rect 115492 91292 115493 91356
rect 115427 91291 115493 91292
rect 115795 91356 115861 91357
rect 115795 91292 115796 91356
rect 115860 91292 115861 91356
rect 115795 91291 115861 91292
rect 117086 91221 117146 94830
rect 114323 91220 114389 91221
rect 114323 91156 114324 91220
rect 114388 91156 114389 91220
rect 114323 91155 114389 91156
rect 114875 91220 114941 91221
rect 114875 91156 114876 91220
rect 114940 91156 114941 91220
rect 114875 91155 114941 91156
rect 117083 91220 117149 91221
rect 117083 91156 117084 91220
rect 117148 91156 117149 91220
rect 117083 91155 117149 91156
rect 113514 78938 113546 79174
rect 113782 78938 113866 79174
rect 114102 78938 114134 79174
rect 113514 78854 114134 78938
rect 113514 78618 113546 78854
rect 113782 78618 113866 78854
rect 114102 78618 114134 78854
rect 113514 43174 114134 78618
rect 113514 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 114134 43174
rect 113514 42854 114134 42938
rect 113514 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 114134 42854
rect 113514 7174 114134 42618
rect 113514 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 114134 7174
rect 113514 6854 114134 6938
rect 113514 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 114134 6854
rect 113514 -2266 114134 6618
rect 113514 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 114134 -2266
rect 113514 -2586 114134 -2502
rect 113514 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 114134 -2586
rect 113514 -3814 114134 -2822
rect 117234 82894 117854 93100
rect 118006 91221 118066 94830
rect 118190 93669 118250 94830
rect 119294 94830 119460 94890
rect 119536 94890 119596 95200
rect 120216 94890 120276 95200
rect 120624 94890 120684 95200
rect 121712 94890 121772 95200
rect 119536 94830 119722 94890
rect 118187 93668 118253 93669
rect 118187 93604 118188 93668
rect 118252 93604 118253 93668
rect 118187 93603 118253 93604
rect 119294 91221 119354 94830
rect 119662 93397 119722 94830
rect 120214 94830 120276 94890
rect 120582 94830 120684 94890
rect 121686 94830 121772 94890
rect 121984 94890 122044 95200
rect 122800 94890 122860 95200
rect 123208 94890 123268 95200
rect 121984 94830 122114 94890
rect 122800 94830 123034 94890
rect 119659 93396 119725 93397
rect 119659 93332 119660 93396
rect 119724 93332 119725 93396
rect 119659 93331 119725 93332
rect 120214 91221 120274 94830
rect 120582 91765 120642 94830
rect 120579 91764 120645 91765
rect 120579 91700 120580 91764
rect 120644 91700 120645 91764
rect 120579 91699 120645 91700
rect 118003 91220 118069 91221
rect 118003 91156 118004 91220
rect 118068 91156 118069 91220
rect 118003 91155 118069 91156
rect 119291 91220 119357 91221
rect 119291 91156 119292 91220
rect 119356 91156 119357 91220
rect 119291 91155 119357 91156
rect 120211 91220 120277 91221
rect 120211 91156 120212 91220
rect 120276 91156 120277 91220
rect 120211 91155 120277 91156
rect 117234 82658 117266 82894
rect 117502 82658 117586 82894
rect 117822 82658 117854 82894
rect 117234 82574 117854 82658
rect 117234 82338 117266 82574
rect 117502 82338 117586 82574
rect 117822 82338 117854 82574
rect 117234 46894 117854 82338
rect 117234 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 117854 46894
rect 117234 46574 117854 46658
rect 117234 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 117854 46574
rect 117234 10894 117854 46338
rect 117234 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 117854 10894
rect 117234 10574 117854 10658
rect 117234 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 117854 10574
rect 117234 -4186 117854 10338
rect 117234 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 117854 -4186
rect 117234 -4506 117854 -4422
rect 117234 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 117854 -4506
rect 117234 -5734 117854 -4742
rect 120954 86614 121574 93100
rect 121686 91221 121746 94830
rect 122054 91221 122114 94830
rect 122974 93397 123034 94830
rect 123158 94830 123268 94890
rect 124024 94890 124084 95200
rect 124432 94890 124492 95200
rect 125384 94890 125444 95200
rect 124024 94830 124138 94890
rect 124432 94830 124506 94890
rect 122971 93396 123037 93397
rect 122971 93332 122972 93396
rect 123036 93332 123037 93396
rect 122971 93331 123037 93332
rect 123158 91221 123218 94830
rect 124078 92445 124138 94830
rect 124075 92444 124141 92445
rect 124075 92380 124076 92444
rect 124140 92380 124141 92444
rect 124075 92379 124141 92380
rect 124446 91357 124506 94830
rect 125366 94830 125444 94890
rect 125656 94890 125716 95200
rect 126472 94890 126532 95200
rect 125656 94830 125794 94890
rect 124443 91356 124509 91357
rect 124443 91292 124444 91356
rect 124508 91292 124509 91356
rect 124443 91291 124509 91292
rect 125366 91221 125426 94830
rect 125734 91357 125794 94830
rect 126470 94830 126532 94890
rect 126608 94890 126668 95200
rect 128104 94890 128164 95200
rect 126608 94830 126714 94890
rect 125731 91356 125797 91357
rect 125731 91292 125732 91356
rect 125796 91292 125797 91356
rect 125731 91291 125797 91292
rect 126470 91221 126530 94830
rect 126654 91493 126714 94830
rect 127574 94830 128164 94890
rect 129328 94890 129388 95200
rect 129328 94830 129474 94890
rect 126651 91492 126717 91493
rect 126651 91428 126652 91492
rect 126716 91428 126717 91492
rect 126651 91427 126717 91428
rect 127574 91221 127634 94830
rect 121683 91220 121749 91221
rect 121683 91156 121684 91220
rect 121748 91156 121749 91220
rect 121683 91155 121749 91156
rect 122051 91220 122117 91221
rect 122051 91156 122052 91220
rect 122116 91156 122117 91220
rect 122051 91155 122117 91156
rect 123155 91220 123221 91221
rect 123155 91156 123156 91220
rect 123220 91156 123221 91220
rect 123155 91155 123221 91156
rect 125363 91220 125429 91221
rect 125363 91156 125364 91220
rect 125428 91156 125429 91220
rect 125363 91155 125429 91156
rect 126467 91220 126533 91221
rect 126467 91156 126468 91220
rect 126532 91156 126533 91220
rect 126467 91155 126533 91156
rect 127571 91220 127637 91221
rect 127571 91156 127572 91220
rect 127636 91156 127637 91220
rect 127571 91155 127637 91156
rect 120954 86378 120986 86614
rect 121222 86378 121306 86614
rect 121542 86378 121574 86614
rect 120954 86294 121574 86378
rect 120954 86058 120986 86294
rect 121222 86058 121306 86294
rect 121542 86058 121574 86294
rect 120954 50614 121574 86058
rect 120954 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 121574 50614
rect 120954 50294 121574 50378
rect 120954 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 121574 50294
rect 120954 14614 121574 50058
rect 120954 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 121574 14614
rect 120954 14294 121574 14378
rect 120954 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 121574 14294
rect 102954 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 103574 -7066
rect 102954 -7386 103574 -7302
rect 102954 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 103574 -7386
rect 102954 -7654 103574 -7622
rect 120954 -6106 121574 14058
rect 127794 57454 128414 93100
rect 129414 91221 129474 94830
rect 130688 94757 130748 95200
rect 131912 94890 131972 95200
rect 133136 94890 133196 95200
rect 131912 94830 132418 94890
rect 130685 94756 130751 94757
rect 130685 94692 130686 94756
rect 130750 94692 130751 94756
rect 130685 94691 130751 94692
rect 129411 91220 129477 91221
rect 129411 91156 129412 91220
rect 129476 91156 129477 91220
rect 129411 91155 129477 91156
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -1306 128414 20898
rect 127794 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 128414 -1306
rect 127794 -1626 128414 -1542
rect 127794 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 128414 -1626
rect 127794 -1894 128414 -1862
rect 131514 61174 132134 93100
rect 132358 91221 132418 94830
rect 133094 94830 133196 94890
rect 134360 94890 134420 95200
rect 135584 94890 135644 95200
rect 151496 94890 151556 95200
rect 134360 94830 134442 94890
rect 135584 94830 136098 94890
rect 133094 92173 133154 94830
rect 134382 92445 134442 94830
rect 134379 92444 134445 92445
rect 134379 92380 134380 92444
rect 134444 92380 134445 92444
rect 134379 92379 134445 92380
rect 133091 92172 133157 92173
rect 133091 92108 133092 92172
rect 133156 92108 133157 92172
rect 133091 92107 133157 92108
rect 132355 91220 132421 91221
rect 132355 91156 132356 91220
rect 132420 91156 132421 91220
rect 132355 91155 132421 91156
rect 131514 60938 131546 61174
rect 131782 60938 131866 61174
rect 132102 60938 132134 61174
rect 131514 60854 132134 60938
rect 131514 60618 131546 60854
rect 131782 60618 131866 60854
rect 132102 60618 132134 60854
rect 131514 25174 132134 60618
rect 131514 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 132134 25174
rect 131514 24854 132134 24938
rect 131514 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 132134 24854
rect 131514 -3226 132134 24618
rect 131514 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 132134 -3226
rect 131514 -3546 132134 -3462
rect 131514 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 132134 -3546
rect 131514 -3814 132134 -3782
rect 135234 64894 135854 93100
rect 136038 91765 136098 94830
rect 151310 94830 151556 94890
rect 136035 91764 136101 91765
rect 136035 91700 136036 91764
rect 136100 91700 136101 91764
rect 136035 91699 136101 91700
rect 135234 64658 135266 64894
rect 135502 64658 135586 64894
rect 135822 64658 135854 64894
rect 135234 64574 135854 64658
rect 135234 64338 135266 64574
rect 135502 64338 135586 64574
rect 135822 64338 135854 64574
rect 135234 28894 135854 64338
rect 135234 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 135854 28894
rect 135234 28574 135854 28658
rect 135234 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 135854 28574
rect 135234 -5146 135854 28338
rect 135234 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 135854 -5146
rect 135234 -5466 135854 -5382
rect 135234 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 135854 -5466
rect 135234 -5734 135854 -5702
rect 138954 68614 139574 93100
rect 138954 68378 138986 68614
rect 139222 68378 139306 68614
rect 139542 68378 139574 68614
rect 138954 68294 139574 68378
rect 138954 68058 138986 68294
rect 139222 68058 139306 68294
rect 139542 68058 139574 68294
rect 138954 32614 139574 68058
rect 138954 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 139574 32614
rect 138954 32294 139574 32378
rect 138954 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 139574 32294
rect 120954 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 121574 -6106
rect 120954 -6426 121574 -6342
rect 120954 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 121574 -6426
rect 120954 -7654 121574 -6662
rect 138954 -7066 139574 32058
rect 145794 75454 146414 93100
rect 145794 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 146414 75454
rect 145794 75134 146414 75218
rect 145794 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 146414 75134
rect 145794 39454 146414 74898
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -1894 146414 -902
rect 149514 79174 150134 93100
rect 151310 92445 151370 94830
rect 151491 94756 151557 94757
rect 151491 94692 151492 94756
rect 151556 94692 151557 94756
rect 151491 94691 151557 94692
rect 151307 92444 151373 92445
rect 151307 92380 151308 92444
rect 151372 92380 151373 92444
rect 151307 92379 151373 92380
rect 151494 91357 151554 94691
rect 151632 94210 151692 95200
rect 151768 94757 151828 95200
rect 151904 94890 151964 95200
rect 151904 94830 152106 94890
rect 151765 94756 151831 94757
rect 151765 94692 151766 94756
rect 151830 94692 151831 94756
rect 151765 94691 151831 94692
rect 151632 94150 151738 94210
rect 151491 91356 151557 91357
rect 151491 91292 151492 91356
rect 151556 91292 151557 91356
rect 151491 91291 151557 91292
rect 151678 91221 151738 94150
rect 152046 91221 152106 94830
rect 151675 91220 151741 91221
rect 151675 91156 151676 91220
rect 151740 91156 151741 91220
rect 151675 91155 151741 91156
rect 152043 91220 152109 91221
rect 152043 91156 152044 91220
rect 152108 91156 152109 91220
rect 152043 91155 152109 91156
rect 149514 78938 149546 79174
rect 149782 78938 149866 79174
rect 150102 78938 150134 79174
rect 149514 78854 150134 78938
rect 149514 78618 149546 78854
rect 149782 78618 149866 78854
rect 150102 78618 150134 78854
rect 149514 43174 150134 78618
rect 149514 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 150134 43174
rect 149514 42854 150134 42938
rect 149514 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 150134 42854
rect 149514 7174 150134 42618
rect 149514 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 150134 7174
rect 149514 6854 150134 6938
rect 149514 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 150134 6854
rect 149514 -2266 150134 6618
rect 149514 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 150134 -2266
rect 149514 -2586 150134 -2502
rect 149514 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 150134 -2586
rect 149514 -3814 150134 -2822
rect 153234 82894 153854 93100
rect 153234 82658 153266 82894
rect 153502 82658 153586 82894
rect 153822 82658 153854 82894
rect 153234 82574 153854 82658
rect 153234 82338 153266 82574
rect 153502 82338 153586 82574
rect 153822 82338 153854 82574
rect 153234 46894 153854 82338
rect 153234 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 153854 46894
rect 153234 46574 153854 46658
rect 153234 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 153854 46574
rect 153234 10894 153854 46338
rect 153234 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 153854 10894
rect 153234 10574 153854 10658
rect 153234 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 153854 10574
rect 153234 -4186 153854 10338
rect 153234 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 153854 -4186
rect 153234 -4506 153854 -4422
rect 153234 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 153854 -4506
rect 153234 -5734 153854 -4742
rect 156954 86614 157574 93100
rect 156954 86378 156986 86614
rect 157222 86378 157306 86614
rect 157542 86378 157574 86614
rect 156954 86294 157574 86378
rect 156954 86058 156986 86294
rect 157222 86058 157306 86294
rect 157542 86058 157574 86294
rect 156954 50614 157574 86058
rect 156954 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 157574 50614
rect 156954 50294 157574 50378
rect 156954 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 157574 50294
rect 156954 14614 157574 50058
rect 156954 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 157574 14614
rect 156954 14294 157574 14378
rect 156954 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 157574 14294
rect 138954 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 139574 -7066
rect 138954 -7386 139574 -7302
rect 138954 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 139574 -7386
rect 138954 -7654 139574 -7622
rect 156954 -6106 157574 14058
rect 163794 57454 164414 93100
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163794 21454 164414 56898
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -1306 164414 20898
rect 165662 3501 165722 242795
rect 166214 235925 166274 314603
rect 167514 313174 168134 348618
rect 168974 316709 169034 523635
rect 169523 337380 169589 337381
rect 169523 337316 169524 337380
rect 169588 337316 169589 337380
rect 169523 337315 169589 337316
rect 168971 316708 169037 316709
rect 168971 316644 168972 316708
rect 169036 316644 169037 316708
rect 168971 316643 169037 316644
rect 167514 312938 167546 313174
rect 167782 312938 167866 313174
rect 168102 312938 168134 313174
rect 167514 312854 168134 312938
rect 167514 312618 167546 312854
rect 167782 312618 167866 312854
rect 168102 312618 168134 312854
rect 167514 277174 168134 312618
rect 169526 304197 169586 337315
rect 169523 304196 169589 304197
rect 169523 304132 169524 304196
rect 169588 304132 169589 304196
rect 169523 304131 169589 304132
rect 168419 302428 168485 302429
rect 168419 302364 168420 302428
rect 168484 302364 168485 302428
rect 168419 302363 168485 302364
rect 167514 276938 167546 277174
rect 167782 276938 167866 277174
rect 168102 276938 168134 277174
rect 167514 276854 168134 276938
rect 167514 276618 167546 276854
rect 167782 276618 167866 276854
rect 168102 276618 168134 276854
rect 167514 241174 168134 276618
rect 167514 240938 167546 241174
rect 167782 240938 167866 241174
rect 168102 240938 168134 241174
rect 167514 240854 168134 240938
rect 167514 240618 167546 240854
rect 167782 240618 167866 240854
rect 168102 240618 168134 240854
rect 166211 235924 166277 235925
rect 166211 235860 166212 235924
rect 166276 235860 166277 235924
rect 166211 235859 166277 235860
rect 167514 205174 168134 240618
rect 168235 237420 168301 237421
rect 168235 237356 168236 237420
rect 168300 237356 168301 237420
rect 168235 237355 168301 237356
rect 168238 232933 168298 237355
rect 168235 232932 168301 232933
rect 168235 232868 168236 232932
rect 168300 232868 168301 232932
rect 168235 232867 168301 232868
rect 168238 231165 168298 232867
rect 168235 231164 168301 231165
rect 168235 231100 168236 231164
rect 168300 231100 168301 231164
rect 168235 231099 168301 231100
rect 168422 212397 168482 302363
rect 170262 241093 170322 546619
rect 171234 532894 171854 568338
rect 171234 532658 171266 532894
rect 171502 532658 171586 532894
rect 171822 532658 171854 532894
rect 171234 532574 171854 532658
rect 171234 532338 171266 532574
rect 171502 532338 171586 532574
rect 171822 532338 171854 532574
rect 171234 496894 171854 532338
rect 171234 496658 171266 496894
rect 171502 496658 171586 496894
rect 171822 496658 171854 496894
rect 171234 496574 171854 496658
rect 171234 496338 171266 496574
rect 171502 496338 171586 496574
rect 171822 496338 171854 496574
rect 171234 460894 171854 496338
rect 171234 460658 171266 460894
rect 171502 460658 171586 460894
rect 171822 460658 171854 460894
rect 171234 460574 171854 460658
rect 171234 460338 171266 460574
rect 171502 460338 171586 460574
rect 171822 460338 171854 460574
rect 171234 424894 171854 460338
rect 171234 424658 171266 424894
rect 171502 424658 171586 424894
rect 171822 424658 171854 424894
rect 171234 424574 171854 424658
rect 171234 424338 171266 424574
rect 171502 424338 171586 424574
rect 171822 424338 171854 424574
rect 171234 388894 171854 424338
rect 171234 388658 171266 388894
rect 171502 388658 171586 388894
rect 171822 388658 171854 388894
rect 171234 388574 171854 388658
rect 171234 388338 171266 388574
rect 171502 388338 171586 388574
rect 171822 388338 171854 388574
rect 171234 352894 171854 388338
rect 171234 352658 171266 352894
rect 171502 352658 171586 352894
rect 171822 352658 171854 352894
rect 171234 352574 171854 352658
rect 171234 352338 171266 352574
rect 171502 352338 171586 352574
rect 171822 352338 171854 352574
rect 171234 316894 171854 352338
rect 174954 680614 175574 711002
rect 192954 710598 193574 711590
rect 192954 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 193574 710598
rect 192954 710278 193574 710362
rect 192954 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 193574 710278
rect 189234 708678 189854 709670
rect 189234 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 189854 708678
rect 189234 708358 189854 708442
rect 189234 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 189854 708358
rect 185514 706758 186134 707750
rect 185514 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 186134 706758
rect 185514 706438 186134 706522
rect 185514 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 186134 706438
rect 174954 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 175574 680614
rect 174954 680294 175574 680378
rect 174954 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 175574 680294
rect 174954 644614 175574 680058
rect 174954 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 175574 644614
rect 174954 644294 175574 644378
rect 174954 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 175574 644294
rect 174954 608614 175574 644058
rect 174954 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 175574 608614
rect 174954 608294 175574 608378
rect 174954 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 175574 608294
rect 174954 572614 175574 608058
rect 174954 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 175574 572614
rect 174954 572294 175574 572378
rect 174954 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 175574 572294
rect 174954 536614 175574 572058
rect 181794 704838 182414 705830
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 178539 564500 178605 564501
rect 178539 564436 178540 564500
rect 178604 564436 178605 564500
rect 178539 564435 178605 564436
rect 174954 536378 174986 536614
rect 175222 536378 175306 536614
rect 175542 536378 175574 536614
rect 174954 536294 175574 536378
rect 174954 536058 174986 536294
rect 175222 536058 175306 536294
rect 175542 536058 175574 536294
rect 174954 500614 175574 536058
rect 174954 500378 174986 500614
rect 175222 500378 175306 500614
rect 175542 500378 175574 500614
rect 174954 500294 175574 500378
rect 174954 500058 174986 500294
rect 175222 500058 175306 500294
rect 175542 500058 175574 500294
rect 174954 464614 175574 500058
rect 174954 464378 174986 464614
rect 175222 464378 175306 464614
rect 175542 464378 175574 464614
rect 174954 464294 175574 464378
rect 174954 464058 174986 464294
rect 175222 464058 175306 464294
rect 175542 464058 175574 464294
rect 174954 428614 175574 464058
rect 174954 428378 174986 428614
rect 175222 428378 175306 428614
rect 175542 428378 175574 428614
rect 174954 428294 175574 428378
rect 174954 428058 174986 428294
rect 175222 428058 175306 428294
rect 175542 428058 175574 428294
rect 174954 392614 175574 428058
rect 177435 401708 177501 401709
rect 177435 401644 177436 401708
rect 177500 401644 177501 401708
rect 177435 401643 177501 401644
rect 174954 392378 174986 392614
rect 175222 392378 175306 392614
rect 175542 392378 175574 392614
rect 174954 392294 175574 392378
rect 174954 392058 174986 392294
rect 175222 392058 175306 392294
rect 175542 392058 175574 392294
rect 174954 356614 175574 392058
rect 174954 356378 174986 356614
rect 175222 356378 175306 356614
rect 175542 356378 175574 356614
rect 174954 356294 175574 356378
rect 174954 356058 174986 356294
rect 175222 356058 175306 356294
rect 175542 356058 175574 356294
rect 174954 320614 175574 356058
rect 177251 331804 177317 331805
rect 177251 331740 177252 331804
rect 177316 331740 177317 331804
rect 177251 331739 177317 331740
rect 174954 320378 174986 320614
rect 175222 320378 175306 320614
rect 175542 320378 175574 320614
rect 174954 320294 175574 320378
rect 174954 320058 174986 320294
rect 175222 320058 175306 320294
rect 175542 320058 175574 320294
rect 173019 317388 173085 317389
rect 173019 317324 173020 317388
rect 173084 317324 173085 317388
rect 173019 317323 173085 317324
rect 171234 316658 171266 316894
rect 171502 316658 171586 316894
rect 171822 316658 171854 316894
rect 171234 316574 171854 316658
rect 171234 316338 171266 316574
rect 171502 316338 171586 316574
rect 171822 316338 171854 316574
rect 171234 280894 171854 316338
rect 171234 280658 171266 280894
rect 171502 280658 171586 280894
rect 171822 280658 171854 280894
rect 171234 280574 171854 280658
rect 171234 280338 171266 280574
rect 171502 280338 171586 280574
rect 171822 280338 171854 280574
rect 171234 244894 171854 280338
rect 172467 251292 172533 251293
rect 172467 251228 172468 251292
rect 172532 251228 172533 251292
rect 172467 251227 172533 251228
rect 171234 244658 171266 244894
rect 171502 244658 171586 244894
rect 171822 244658 171854 244894
rect 171234 244574 171854 244658
rect 171234 244338 171266 244574
rect 171502 244338 171586 244574
rect 171822 244338 171854 244574
rect 170259 241092 170325 241093
rect 170259 241028 170260 241092
rect 170324 241028 170325 241092
rect 170259 241027 170325 241028
rect 168419 212396 168485 212397
rect 168419 212332 168420 212396
rect 168484 212332 168485 212396
rect 168419 212331 168485 212332
rect 167514 204938 167546 205174
rect 167782 204938 167866 205174
rect 168102 204938 168134 205174
rect 167514 204854 168134 204938
rect 167514 204618 167546 204854
rect 167782 204618 167866 204854
rect 168102 204618 168134 204854
rect 167514 169174 168134 204618
rect 169707 182068 169773 182069
rect 169707 182004 169708 182068
rect 169772 182004 169773 182068
rect 169707 182003 169773 182004
rect 169710 180845 169770 182003
rect 169707 180844 169773 180845
rect 169707 180780 169708 180844
rect 169772 180780 169773 180844
rect 169707 180779 169773 180780
rect 167514 168938 167546 169174
rect 167782 168938 167866 169174
rect 168102 168938 168134 169174
rect 167514 168854 168134 168938
rect 167514 168618 167546 168854
rect 167782 168618 167866 168854
rect 168102 168618 168134 168854
rect 167514 133174 168134 168618
rect 169710 161490 169770 180779
rect 167514 132938 167546 133174
rect 167782 132938 167866 133174
rect 168102 132938 168134 133174
rect 167514 132854 168134 132938
rect 167514 132618 167546 132854
rect 167782 132618 167866 132854
rect 168102 132618 168134 132854
rect 167514 97174 168134 132618
rect 169526 161430 169770 161490
rect 168235 109716 168301 109717
rect 168235 109652 168236 109716
rect 168300 109652 168301 109716
rect 168235 109651 168301 109652
rect 167514 96938 167546 97174
rect 167782 96938 167866 97174
rect 168102 96938 168134 97174
rect 167514 96854 168134 96938
rect 167514 96618 167546 96854
rect 167782 96618 167866 96854
rect 168102 96618 168134 96854
rect 167514 61174 168134 96618
rect 168238 67557 168298 109651
rect 168235 67556 168301 67557
rect 168235 67492 168236 67556
rect 168300 67492 168301 67556
rect 168235 67491 168301 67492
rect 167514 60938 167546 61174
rect 167782 60938 167866 61174
rect 168102 60938 168134 61174
rect 167514 60854 168134 60938
rect 167514 60618 167546 60854
rect 167782 60618 167866 60854
rect 168102 60618 168134 60854
rect 167514 25174 168134 60618
rect 169526 26893 169586 161430
rect 170262 151061 170322 241027
rect 171234 208894 171854 244338
rect 171234 208658 171266 208894
rect 171502 208658 171586 208894
rect 171822 208658 171854 208894
rect 171234 208574 171854 208658
rect 171234 208338 171266 208574
rect 171502 208338 171586 208574
rect 171822 208338 171854 208574
rect 171234 172894 171854 208338
rect 171234 172658 171266 172894
rect 171502 172658 171586 172894
rect 171822 172658 171854 172894
rect 171234 172574 171854 172658
rect 171234 172338 171266 172574
rect 171502 172338 171586 172574
rect 171822 172338 171854 172574
rect 170259 151060 170325 151061
rect 170259 150996 170260 151060
rect 170324 150996 170325 151060
rect 170259 150995 170325 150996
rect 171234 136894 171854 172338
rect 171234 136658 171266 136894
rect 171502 136658 171586 136894
rect 171822 136658 171854 136894
rect 171234 136574 171854 136658
rect 171234 136338 171266 136574
rect 171502 136338 171586 136574
rect 171822 136338 171854 136574
rect 171234 100894 171854 136338
rect 171234 100658 171266 100894
rect 171502 100658 171586 100894
rect 171822 100658 171854 100894
rect 171234 100574 171854 100658
rect 171234 100338 171266 100574
rect 171502 100338 171586 100574
rect 171822 100338 171854 100574
rect 171234 64894 171854 100338
rect 171234 64658 171266 64894
rect 171502 64658 171586 64894
rect 171822 64658 171854 64894
rect 171234 64574 171854 64658
rect 171234 64338 171266 64574
rect 171502 64338 171586 64574
rect 171822 64338 171854 64574
rect 171234 28894 171854 64338
rect 171234 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 171854 28894
rect 171234 28574 171854 28658
rect 171234 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 171854 28574
rect 169523 26892 169589 26893
rect 169523 26828 169524 26892
rect 169588 26828 169589 26892
rect 169523 26827 169589 26828
rect 167514 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 168134 25174
rect 167514 24854 168134 24938
rect 167514 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 168134 24854
rect 165659 3500 165725 3501
rect 165659 3436 165660 3500
rect 165724 3436 165725 3500
rect 165659 3435 165725 3436
rect 163794 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 164414 -1306
rect 163794 -1626 164414 -1542
rect 163794 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 164414 -1626
rect 163794 -1894 164414 -1862
rect 167514 -3226 168134 24618
rect 167514 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 168134 -3226
rect 167514 -3546 168134 -3462
rect 167514 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 168134 -3546
rect 167514 -3814 168134 -3782
rect 171234 -5146 171854 28338
rect 172470 15877 172530 251227
rect 173022 215117 173082 317323
rect 173203 309908 173269 309909
rect 173203 309844 173204 309908
rect 173268 309844 173269 309908
rect 173203 309843 173269 309844
rect 173206 278765 173266 309843
rect 174954 284614 175574 320058
rect 174954 284378 174986 284614
rect 175222 284378 175306 284614
rect 175542 284378 175574 284614
rect 174954 284294 175574 284378
rect 174954 284058 174986 284294
rect 175222 284058 175306 284294
rect 175542 284058 175574 284294
rect 173203 278764 173269 278765
rect 173203 278700 173204 278764
rect 173268 278700 173269 278764
rect 173203 278699 173269 278700
rect 174954 248614 175574 284058
rect 174954 248378 174986 248614
rect 175222 248378 175306 248614
rect 175542 248378 175574 248614
rect 174954 248294 175574 248378
rect 174954 248058 174986 248294
rect 175222 248058 175306 248294
rect 175542 248058 175574 248294
rect 173019 215116 173085 215117
rect 173019 215052 173020 215116
rect 173084 215052 173085 215116
rect 173019 215051 173085 215052
rect 174954 212614 175574 248058
rect 174954 212378 174986 212614
rect 175222 212378 175306 212614
rect 175542 212378 175574 212614
rect 174954 212294 175574 212378
rect 174954 212058 174986 212294
rect 175222 212058 175306 212294
rect 175542 212058 175574 212294
rect 174954 176614 175574 212058
rect 174954 176378 174986 176614
rect 175222 176378 175306 176614
rect 175542 176378 175574 176614
rect 174954 176294 175574 176378
rect 174954 176058 174986 176294
rect 175222 176058 175306 176294
rect 175542 176058 175574 176294
rect 174954 140614 175574 176058
rect 174954 140378 174986 140614
rect 175222 140378 175306 140614
rect 175542 140378 175574 140614
rect 174954 140294 175574 140378
rect 174954 140058 174986 140294
rect 175222 140058 175306 140294
rect 175542 140058 175574 140294
rect 174954 104614 175574 140058
rect 174954 104378 174986 104614
rect 175222 104378 175306 104614
rect 175542 104378 175574 104614
rect 174954 104294 175574 104378
rect 174954 104058 174986 104294
rect 175222 104058 175306 104294
rect 175542 104058 175574 104294
rect 174954 68614 175574 104058
rect 174954 68378 174986 68614
rect 175222 68378 175306 68614
rect 175542 68378 175574 68614
rect 174954 68294 175574 68378
rect 174954 68058 174986 68294
rect 175222 68058 175306 68294
rect 175542 68058 175574 68294
rect 174954 32614 175574 68058
rect 174954 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 175574 32614
rect 174954 32294 175574 32378
rect 174954 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 175574 32294
rect 172467 15876 172533 15877
rect 172467 15812 172468 15876
rect 172532 15812 172533 15876
rect 172467 15811 172533 15812
rect 171234 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 171854 -5146
rect 171234 -5466 171854 -5382
rect 171234 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 171854 -5466
rect 171234 -5734 171854 -5702
rect 156954 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 157574 -6106
rect 156954 -6426 157574 -6342
rect 156954 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 157574 -6426
rect 156954 -7654 157574 -6662
rect 174954 -7066 175574 32058
rect 177254 15877 177314 331739
rect 177438 294541 177498 401643
rect 177435 294540 177501 294541
rect 177435 294476 177436 294540
rect 177500 294476 177501 294540
rect 177435 294475 177501 294476
rect 178542 224365 178602 564435
rect 181794 543454 182414 578898
rect 185514 691174 186134 706202
rect 185514 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 186134 691174
rect 185514 690854 186134 690938
rect 185514 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 186134 690854
rect 185514 655174 186134 690618
rect 185514 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 186134 655174
rect 185514 654854 186134 654938
rect 185514 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 186134 654854
rect 185514 619174 186134 654618
rect 185514 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 186134 619174
rect 185514 618854 186134 618938
rect 185514 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 186134 618854
rect 185514 583174 186134 618618
rect 185514 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 186134 583174
rect 185514 582854 186134 582938
rect 185514 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 186134 582854
rect 184795 550764 184861 550765
rect 184795 550700 184796 550764
rect 184860 550700 184861 550764
rect 184795 550699 184861 550700
rect 181794 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 182414 543454
rect 181794 543134 182414 543218
rect 181794 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 182414 543134
rect 181794 507454 182414 542898
rect 181794 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 182414 507454
rect 181794 507134 182414 507218
rect 181794 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 182414 507134
rect 181794 471454 182414 506898
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 181794 435454 182414 470898
rect 181794 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 182414 435454
rect 181794 435134 182414 435218
rect 181794 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 182414 435134
rect 181794 399454 182414 434898
rect 181794 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 182414 399454
rect 181794 399134 182414 399218
rect 181794 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 182414 399134
rect 181794 363454 182414 398898
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 178723 331396 178789 331397
rect 178723 331332 178724 331396
rect 178788 331332 178789 331396
rect 178723 331331 178789 331332
rect 178539 224364 178605 224365
rect 178539 224300 178540 224364
rect 178604 224300 178605 224364
rect 178539 224299 178605 224300
rect 177251 15876 177317 15877
rect 177251 15812 177252 15876
rect 177316 15812 177317 15876
rect 177251 15811 177317 15812
rect 178726 7581 178786 331331
rect 181794 327454 182414 362898
rect 181794 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 182414 327454
rect 181794 327134 182414 327218
rect 181794 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 182414 327134
rect 181794 291454 182414 326898
rect 182771 304196 182837 304197
rect 182771 304132 182772 304196
rect 182836 304132 182837 304196
rect 182771 304131 182837 304132
rect 181794 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 182414 291454
rect 181794 291134 182414 291218
rect 181794 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 182414 291134
rect 180011 278084 180077 278085
rect 180011 278020 180012 278084
rect 180076 278020 180077 278084
rect 180011 278019 180077 278020
rect 180014 228989 180074 278019
rect 180195 262988 180261 262989
rect 180195 262924 180196 262988
rect 180260 262924 180261 262988
rect 180195 262923 180261 262924
rect 180198 235789 180258 262923
rect 181794 255454 182414 290898
rect 181794 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 182414 255454
rect 181794 255134 182414 255218
rect 181794 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 182414 255134
rect 180195 235788 180261 235789
rect 180195 235724 180196 235788
rect 180260 235724 180261 235788
rect 180195 235723 180261 235724
rect 180011 228988 180077 228989
rect 180011 228924 180012 228988
rect 180076 228924 180077 228988
rect 180011 228923 180077 228924
rect 181794 219454 182414 254898
rect 181794 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 182414 219454
rect 181794 219134 182414 219218
rect 181794 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 182414 219134
rect 181794 183454 182414 218898
rect 181794 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 182414 183454
rect 181794 183134 182414 183218
rect 181794 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 182414 183134
rect 181794 147454 182414 182898
rect 181794 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 182414 147454
rect 181794 147134 182414 147218
rect 181794 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 182414 147134
rect 181794 111454 182414 146898
rect 181794 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 182414 111454
rect 181794 111134 182414 111218
rect 181794 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 182414 111134
rect 181794 75454 182414 110898
rect 181794 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 182414 75454
rect 181794 75134 182414 75218
rect 181794 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 182414 75134
rect 181794 39454 182414 74898
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 178723 7580 178789 7581
rect 178723 7516 178724 7580
rect 178788 7516 178789 7580
rect 178723 7515 178789 7516
rect 181794 3454 182414 38898
rect 182774 11661 182834 304131
rect 184611 265164 184677 265165
rect 184611 265100 184612 265164
rect 184676 265100 184677 265164
rect 184611 265099 184677 265100
rect 184614 233205 184674 265099
rect 184611 233204 184677 233205
rect 184611 233140 184612 233204
rect 184676 233140 184677 233204
rect 184611 233139 184677 233140
rect 184798 228853 184858 550699
rect 185514 547174 186134 582618
rect 185514 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 186134 547174
rect 185514 546854 186134 546938
rect 185514 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 186134 546854
rect 185347 539748 185413 539749
rect 185347 539684 185348 539748
rect 185412 539684 185413 539748
rect 185347 539683 185413 539684
rect 185350 272509 185410 539683
rect 185514 511174 186134 546618
rect 185514 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 186134 511174
rect 185514 510854 186134 510938
rect 185514 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 186134 510854
rect 185514 475174 186134 510618
rect 189234 694894 189854 708122
rect 189234 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 189854 694894
rect 189234 694574 189854 694658
rect 189234 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 189854 694574
rect 189234 658894 189854 694338
rect 189234 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 189854 658894
rect 189234 658574 189854 658658
rect 189234 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 189854 658574
rect 189234 622894 189854 658338
rect 189234 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 189854 622894
rect 189234 622574 189854 622658
rect 189234 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 189854 622574
rect 189234 586894 189854 622338
rect 189234 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 189854 586894
rect 189234 586574 189854 586658
rect 189234 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 189854 586574
rect 189234 550894 189854 586338
rect 189234 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 189854 550894
rect 189234 550574 189854 550658
rect 189234 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 189854 550574
rect 189234 514894 189854 550338
rect 192954 698614 193574 710042
rect 210954 711558 211574 711590
rect 210954 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 211574 711558
rect 210954 711238 211574 711322
rect 210954 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 211574 711238
rect 207234 709638 207854 709670
rect 207234 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 207854 709638
rect 207234 709318 207854 709402
rect 207234 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 207854 709318
rect 203514 707718 204134 707750
rect 203514 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 204134 707718
rect 203514 707398 204134 707482
rect 203514 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 204134 707398
rect 192954 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 193574 698614
rect 192954 698294 193574 698378
rect 192954 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 193574 698294
rect 192954 662614 193574 698058
rect 192954 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 193574 662614
rect 192954 662294 193574 662378
rect 192954 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 193574 662294
rect 192954 626614 193574 662058
rect 192954 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 193574 626614
rect 192954 626294 193574 626378
rect 192954 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 193574 626294
rect 192954 590614 193574 626058
rect 192954 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 193574 590614
rect 192954 590294 193574 590378
rect 192954 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 193574 590294
rect 192954 554614 193574 590058
rect 192954 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 193574 554614
rect 192954 554294 193574 554378
rect 192954 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 193574 554294
rect 192954 518614 193574 554058
rect 199794 705798 200414 705830
rect 199794 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 200414 705798
rect 199794 705478 200414 705562
rect 199794 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 200414 705478
rect 199794 669454 200414 705242
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 633454 200414 668898
rect 199794 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 200414 633454
rect 199794 633134 200414 633218
rect 199794 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 200414 633134
rect 199794 597454 200414 632898
rect 199794 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 200414 597454
rect 199794 597134 200414 597218
rect 199794 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 200414 597134
rect 199794 561454 200414 596898
rect 199794 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 200414 561454
rect 199794 561134 200414 561218
rect 199794 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 200414 561134
rect 198595 551308 198661 551309
rect 198595 551244 198596 551308
rect 198660 551244 198661 551308
rect 198595 551243 198661 551244
rect 197859 542604 197925 542605
rect 197859 542540 197860 542604
rect 197924 542540 197925 542604
rect 197859 542539 197925 542540
rect 196571 538660 196637 538661
rect 196571 538596 196572 538660
rect 196636 538596 196637 538660
rect 196571 538595 196637 538596
rect 194363 538388 194429 538389
rect 194363 538324 194364 538388
rect 194428 538324 194429 538388
rect 194363 538323 194429 538324
rect 192954 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 193574 518614
rect 192954 518294 193574 518378
rect 191787 518124 191853 518125
rect 191787 518060 191788 518124
rect 191852 518060 191853 518124
rect 191787 518059 191853 518060
rect 189234 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 189854 514894
rect 189234 514574 189854 514658
rect 189234 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 189854 514574
rect 188843 502484 188909 502485
rect 188843 502420 188844 502484
rect 188908 502420 188909 502484
rect 188843 502419 188909 502420
rect 185514 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 186134 475174
rect 185514 474854 186134 474938
rect 185514 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 186134 474854
rect 185514 439174 186134 474618
rect 185514 438938 185546 439174
rect 185782 438938 185866 439174
rect 186102 438938 186134 439174
rect 185514 438854 186134 438938
rect 185514 438618 185546 438854
rect 185782 438618 185866 438854
rect 186102 438618 186134 438854
rect 185514 403174 186134 438618
rect 186819 404564 186885 404565
rect 186819 404500 186820 404564
rect 186884 404500 186885 404564
rect 186819 404499 186885 404500
rect 185514 402938 185546 403174
rect 185782 402938 185866 403174
rect 186102 402938 186134 403174
rect 185514 402854 186134 402938
rect 185514 402618 185546 402854
rect 185782 402618 185866 402854
rect 186102 402618 186134 402854
rect 185514 367174 186134 402618
rect 186822 368389 186882 404499
rect 186819 368388 186885 368389
rect 186819 368324 186820 368388
rect 186884 368324 186885 368388
rect 186819 368323 186885 368324
rect 185514 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 186134 367174
rect 185514 366854 186134 366938
rect 185514 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 186134 366854
rect 185514 331174 186134 366618
rect 186819 345812 186885 345813
rect 186819 345748 186820 345812
rect 186884 345748 186885 345812
rect 186819 345747 186885 345748
rect 185514 330938 185546 331174
rect 185782 330938 185866 331174
rect 186102 330938 186134 331174
rect 185514 330854 186134 330938
rect 185514 330618 185546 330854
rect 185782 330618 185866 330854
rect 186102 330618 186134 330854
rect 185514 295174 186134 330618
rect 185514 294938 185546 295174
rect 185782 294938 185866 295174
rect 186102 294938 186134 295174
rect 185514 294854 186134 294938
rect 185514 294618 185546 294854
rect 185782 294618 185866 294854
rect 186102 294618 186134 294854
rect 185347 272508 185413 272509
rect 185347 272444 185348 272508
rect 185412 272444 185413 272508
rect 185347 272443 185413 272444
rect 185347 261628 185413 261629
rect 185347 261564 185348 261628
rect 185412 261564 185413 261628
rect 185347 261563 185413 261564
rect 185350 230349 185410 261563
rect 185514 259174 186134 294618
rect 186822 283253 186882 345747
rect 187555 316708 187621 316709
rect 187555 316644 187556 316708
rect 187620 316644 187621 316708
rect 187555 316643 187621 316644
rect 186819 283252 186885 283253
rect 186819 283188 186820 283252
rect 186884 283188 186885 283252
rect 186819 283187 186885 283188
rect 186822 281485 186882 283187
rect 186819 281484 186885 281485
rect 186819 281420 186820 281484
rect 186884 281420 186885 281484
rect 186819 281419 186885 281420
rect 186819 263668 186885 263669
rect 186819 263604 186820 263668
rect 186884 263604 186885 263668
rect 186819 263603 186885 263604
rect 185514 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 186134 259174
rect 185514 258854 186134 258938
rect 185514 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 186134 258854
rect 185347 230348 185413 230349
rect 185347 230284 185348 230348
rect 185412 230284 185413 230348
rect 185347 230283 185413 230284
rect 184795 228852 184861 228853
rect 184795 228788 184796 228852
rect 184860 228788 184861 228852
rect 184795 228787 184861 228788
rect 184798 228309 184858 228787
rect 184795 228308 184861 228309
rect 184795 228244 184796 228308
rect 184860 228244 184861 228308
rect 184795 228243 184861 228244
rect 185514 223174 186134 258618
rect 185514 222938 185546 223174
rect 185782 222938 185866 223174
rect 186102 222938 186134 223174
rect 185514 222854 186134 222938
rect 185514 222618 185546 222854
rect 185782 222618 185866 222854
rect 186102 222618 186134 222854
rect 185514 187174 186134 222618
rect 185514 186938 185546 187174
rect 185782 186938 185866 187174
rect 186102 186938 186134 187174
rect 185514 186854 186134 186938
rect 185514 186618 185546 186854
rect 185782 186618 185866 186854
rect 186102 186618 186134 186854
rect 185514 151174 186134 186618
rect 185514 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 186134 151174
rect 185514 150854 186134 150938
rect 185514 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 186134 150854
rect 185514 115174 186134 150618
rect 185514 114938 185546 115174
rect 185782 114938 185866 115174
rect 186102 114938 186134 115174
rect 185514 114854 186134 114938
rect 185514 114618 185546 114854
rect 185782 114618 185866 114854
rect 186102 114618 186134 114854
rect 185514 79174 186134 114618
rect 185514 78938 185546 79174
rect 185782 78938 185866 79174
rect 186102 78938 186134 79174
rect 185514 78854 186134 78938
rect 185514 78618 185546 78854
rect 185782 78618 185866 78854
rect 186102 78618 186134 78854
rect 185514 43174 186134 78618
rect 185514 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 186134 43174
rect 185514 42854 186134 42938
rect 185514 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 186134 42854
rect 182771 11660 182837 11661
rect 182771 11596 182772 11660
rect 182836 11596 182837 11660
rect 182771 11595 182837 11596
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -1894 182414 -902
rect 185514 7174 186134 42618
rect 186822 35189 186882 263603
rect 187558 233205 187618 316643
rect 188291 309772 188357 309773
rect 188291 309708 188292 309772
rect 188356 309708 188357 309772
rect 188291 309707 188357 309708
rect 188294 247077 188354 309707
rect 188291 247076 188357 247077
rect 188291 247012 188292 247076
rect 188356 247012 188357 247076
rect 188291 247011 188357 247012
rect 188846 237285 188906 502419
rect 189234 478894 189854 514338
rect 189234 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 189854 478894
rect 189234 478574 189854 478658
rect 189234 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 189854 478574
rect 189234 442894 189854 478338
rect 189234 442658 189266 442894
rect 189502 442658 189586 442894
rect 189822 442658 189854 442894
rect 189234 442574 189854 442658
rect 189234 442338 189266 442574
rect 189502 442338 189586 442574
rect 189822 442338 189854 442574
rect 189234 406894 189854 442338
rect 189234 406658 189266 406894
rect 189502 406658 189586 406894
rect 189822 406658 189854 406894
rect 189234 406574 189854 406658
rect 189234 406338 189266 406574
rect 189502 406338 189586 406574
rect 189822 406338 189854 406574
rect 189234 370894 189854 406338
rect 189234 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 189854 370894
rect 189234 370574 189854 370658
rect 189234 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 189854 370574
rect 189234 334894 189854 370338
rect 191235 357644 191301 357645
rect 191235 357580 191236 357644
rect 191300 357580 191301 357644
rect 191235 357579 191301 357580
rect 189234 334658 189266 334894
rect 189502 334658 189586 334894
rect 189822 334658 189854 334894
rect 189234 334574 189854 334658
rect 189234 334338 189266 334574
rect 189502 334338 189586 334574
rect 189822 334338 189854 334574
rect 189234 298894 189854 334338
rect 191051 313172 191117 313173
rect 191051 313108 191052 313172
rect 191116 313108 191117 313172
rect 191051 313107 191117 313108
rect 189234 298658 189266 298894
rect 189502 298658 189586 298894
rect 189822 298658 189854 298894
rect 189234 298574 189854 298658
rect 189234 298338 189266 298574
rect 189502 298338 189586 298574
rect 189822 298338 189854 298574
rect 189234 262894 189854 298338
rect 189234 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 189854 262894
rect 189234 262574 189854 262658
rect 189234 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 189854 262574
rect 188843 237284 188909 237285
rect 188843 237220 188844 237284
rect 188908 237220 188909 237284
rect 188843 237219 188909 237220
rect 187555 233204 187621 233205
rect 187555 233140 187556 233204
rect 187620 233140 187621 233204
rect 187555 233139 187621 233140
rect 189234 226894 189854 262338
rect 189234 226658 189266 226894
rect 189502 226658 189586 226894
rect 189822 226658 189854 226894
rect 189234 226574 189854 226658
rect 189234 226338 189266 226574
rect 189502 226338 189586 226574
rect 189822 226338 189854 226574
rect 189234 190894 189854 226338
rect 189234 190658 189266 190894
rect 189502 190658 189586 190894
rect 189822 190658 189854 190894
rect 189234 190574 189854 190658
rect 189234 190338 189266 190574
rect 189502 190338 189586 190574
rect 189822 190338 189854 190574
rect 189234 154894 189854 190338
rect 189234 154658 189266 154894
rect 189502 154658 189586 154894
rect 189822 154658 189854 154894
rect 189234 154574 189854 154658
rect 189234 154338 189266 154574
rect 189502 154338 189586 154574
rect 189822 154338 189854 154574
rect 189234 118894 189854 154338
rect 189234 118658 189266 118894
rect 189502 118658 189586 118894
rect 189822 118658 189854 118894
rect 189234 118574 189854 118658
rect 189234 118338 189266 118574
rect 189502 118338 189586 118574
rect 189822 118338 189854 118574
rect 189234 82894 189854 118338
rect 191054 84829 191114 313107
rect 191238 286381 191298 357579
rect 191235 286380 191301 286381
rect 191235 286316 191236 286380
rect 191300 286316 191301 286380
rect 191235 286315 191301 286316
rect 191790 245717 191850 518059
rect 192954 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 193574 518294
rect 192954 482614 193574 518058
rect 192954 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 193574 482614
rect 192954 482294 193574 482378
rect 192954 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 193574 482294
rect 192954 446614 193574 482058
rect 192954 446378 192986 446614
rect 193222 446378 193306 446614
rect 193542 446378 193574 446614
rect 192954 446294 193574 446378
rect 192954 446058 192986 446294
rect 193222 446058 193306 446294
rect 193542 446058 193574 446294
rect 192954 410614 193574 446058
rect 192954 410378 192986 410614
rect 193222 410378 193306 410614
rect 193542 410378 193574 410614
rect 192954 410294 193574 410378
rect 192954 410058 192986 410294
rect 193222 410058 193306 410294
rect 193542 410058 193574 410294
rect 192954 374614 193574 410058
rect 194366 378181 194426 538323
rect 195099 490516 195165 490517
rect 195099 490452 195100 490516
rect 195164 490452 195165 490516
rect 195099 490451 195165 490452
rect 194547 446452 194613 446453
rect 194547 446388 194548 446452
rect 194612 446388 194613 446452
rect 194547 446387 194613 446388
rect 194363 378180 194429 378181
rect 194363 378116 194364 378180
rect 194428 378116 194429 378180
rect 194363 378115 194429 378116
rect 192954 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 193574 374614
rect 192954 374294 193574 374378
rect 192954 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 193574 374294
rect 192954 338614 193574 374058
rect 194550 364989 194610 446387
rect 194547 364988 194613 364989
rect 194547 364924 194548 364988
rect 194612 364924 194613 364988
rect 194547 364923 194613 364924
rect 192954 338378 192986 338614
rect 193222 338378 193306 338614
rect 193542 338378 193574 338614
rect 192954 338294 193574 338378
rect 192954 338058 192986 338294
rect 193222 338058 193306 338294
rect 193542 338058 193574 338294
rect 192954 302614 193574 338058
rect 192954 302378 192986 302614
rect 193222 302378 193306 302614
rect 193542 302378 193574 302614
rect 192954 302294 193574 302378
rect 192954 302058 192986 302294
rect 193222 302058 193306 302294
rect 193542 302058 193574 302294
rect 192954 266614 193574 302058
rect 192954 266378 192986 266614
rect 193222 266378 193306 266614
rect 193542 266378 193574 266614
rect 192954 266294 193574 266378
rect 192954 266058 192986 266294
rect 193222 266058 193306 266294
rect 193542 266058 193574 266294
rect 191787 245716 191853 245717
rect 191787 245652 191788 245716
rect 191852 245652 191853 245716
rect 191787 245651 191853 245652
rect 192954 230614 193574 266058
rect 195102 262989 195162 490451
rect 196574 344997 196634 538595
rect 197862 526421 197922 542539
rect 197859 526420 197925 526421
rect 197859 526356 197860 526420
rect 197924 526356 197925 526420
rect 197859 526355 197925 526356
rect 198598 500445 198658 551243
rect 199331 541244 199397 541245
rect 199331 541180 199332 541244
rect 199396 541180 199397 541244
rect 199331 541179 199397 541180
rect 199334 513365 199394 541179
rect 199794 537993 200414 560898
rect 203514 673174 204134 707162
rect 203514 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 204134 673174
rect 203514 672854 204134 672938
rect 203514 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 204134 672854
rect 203514 637174 204134 672618
rect 203514 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 204134 637174
rect 203514 636854 204134 636938
rect 203514 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 204134 636854
rect 203514 601174 204134 636618
rect 203514 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 204134 601174
rect 203514 600854 204134 600938
rect 203514 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 204134 600854
rect 203514 565174 204134 600618
rect 203514 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 204134 565174
rect 203514 564854 204134 564938
rect 203514 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 204134 564854
rect 203514 537993 204134 564618
rect 207234 676894 207854 709082
rect 207234 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 207854 676894
rect 207234 676574 207854 676658
rect 207234 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 207854 676574
rect 207234 640894 207854 676338
rect 207234 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 207854 640894
rect 207234 640574 207854 640658
rect 207234 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 207854 640574
rect 207234 604894 207854 640338
rect 207234 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 207854 604894
rect 207234 604574 207854 604658
rect 207234 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 207854 604574
rect 207234 568894 207854 604338
rect 207234 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 207854 568894
rect 207234 568574 207854 568658
rect 207234 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 207854 568574
rect 207234 537993 207854 568338
rect 210954 680614 211574 711002
rect 228954 710598 229574 711590
rect 228954 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 229574 710598
rect 228954 710278 229574 710362
rect 228954 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 229574 710278
rect 225234 708678 225854 709670
rect 225234 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 225854 708678
rect 225234 708358 225854 708442
rect 225234 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 225854 708358
rect 221514 706758 222134 707750
rect 221514 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 222134 706758
rect 221514 706438 222134 706522
rect 221514 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 222134 706438
rect 210954 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 211574 680614
rect 210954 680294 211574 680378
rect 210954 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 211574 680294
rect 210954 644614 211574 680058
rect 210954 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 211574 644614
rect 210954 644294 211574 644378
rect 210954 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 211574 644294
rect 210954 608614 211574 644058
rect 210954 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 211574 608614
rect 210954 608294 211574 608378
rect 210954 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 211574 608294
rect 210954 572614 211574 608058
rect 210954 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 211574 572614
rect 210954 572294 211574 572378
rect 210954 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 211574 572294
rect 210954 537993 211574 572058
rect 217794 704838 218414 705830
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 579454 218414 614898
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 217794 543454 218414 578898
rect 217794 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 218414 543454
rect 217794 543134 218414 543218
rect 217794 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 218414 543134
rect 217794 537993 218414 542898
rect 221514 691174 222134 706202
rect 221514 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 222134 691174
rect 221514 690854 222134 690938
rect 221514 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 222134 690854
rect 221514 655174 222134 690618
rect 221514 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 222134 655174
rect 221514 654854 222134 654938
rect 221514 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 222134 654854
rect 221514 619174 222134 654618
rect 221514 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 222134 619174
rect 221514 618854 222134 618938
rect 221514 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 222134 618854
rect 221514 583174 222134 618618
rect 221514 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 222134 583174
rect 221514 582854 222134 582938
rect 221514 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 222134 582854
rect 221514 547174 222134 582618
rect 221514 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 222134 547174
rect 221514 546854 222134 546938
rect 221514 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 222134 546854
rect 221514 537993 222134 546618
rect 225234 694894 225854 708122
rect 225234 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 225854 694894
rect 225234 694574 225854 694658
rect 225234 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 225854 694574
rect 225234 658894 225854 694338
rect 225234 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 225854 658894
rect 225234 658574 225854 658658
rect 225234 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 225854 658574
rect 225234 622894 225854 658338
rect 225234 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 225854 622894
rect 225234 622574 225854 622658
rect 225234 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 225854 622574
rect 225234 586894 225854 622338
rect 225234 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 225854 586894
rect 225234 586574 225854 586658
rect 225234 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 225854 586574
rect 225234 550894 225854 586338
rect 225234 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 225854 550894
rect 225234 550574 225854 550658
rect 225234 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 225854 550574
rect 225234 537993 225854 550338
rect 228954 698614 229574 710042
rect 246954 711558 247574 711590
rect 246954 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 247574 711558
rect 246954 711238 247574 711322
rect 246954 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 247574 711238
rect 243234 709638 243854 709670
rect 243234 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 243854 709638
rect 243234 709318 243854 709402
rect 243234 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 243854 709318
rect 239514 707718 240134 707750
rect 239514 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 240134 707718
rect 239514 707398 240134 707482
rect 239514 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 240134 707398
rect 228954 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 229574 698614
rect 228954 698294 229574 698378
rect 228954 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 229574 698294
rect 228954 662614 229574 698058
rect 228954 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 229574 662614
rect 228954 662294 229574 662378
rect 228954 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 229574 662294
rect 228954 626614 229574 662058
rect 228954 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 229574 626614
rect 228954 626294 229574 626378
rect 228954 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 229574 626294
rect 228954 590614 229574 626058
rect 228954 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 229574 590614
rect 228954 590294 229574 590378
rect 228954 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 229574 590294
rect 228954 554614 229574 590058
rect 228954 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 229574 554614
rect 228954 554294 229574 554378
rect 228954 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 229574 554294
rect 228954 537993 229574 554058
rect 235794 705798 236414 705830
rect 235794 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 236414 705798
rect 235794 705478 236414 705562
rect 235794 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 236414 705478
rect 235794 669454 236414 705242
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 633454 236414 668898
rect 235794 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 236414 633454
rect 235794 633134 236414 633218
rect 235794 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 236414 633134
rect 235794 597454 236414 632898
rect 235794 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 236414 597454
rect 235794 597134 236414 597218
rect 235794 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 236414 597134
rect 235794 561454 236414 596898
rect 235794 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 236414 561454
rect 235794 561134 236414 561218
rect 235794 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 236414 561134
rect 235794 537993 236414 560898
rect 239514 673174 240134 707162
rect 239514 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 240134 673174
rect 239514 672854 240134 672938
rect 239514 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 240134 672854
rect 239514 637174 240134 672618
rect 239514 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 240134 637174
rect 239514 636854 240134 636938
rect 239514 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 240134 636854
rect 239514 601174 240134 636618
rect 239514 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 240134 601174
rect 239514 600854 240134 600938
rect 239514 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 240134 600854
rect 239514 565174 240134 600618
rect 239514 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 240134 565174
rect 239514 564854 240134 564938
rect 239514 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 240134 564854
rect 239514 537993 240134 564618
rect 243234 676894 243854 709082
rect 243234 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 243854 676894
rect 243234 676574 243854 676658
rect 243234 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 243854 676574
rect 243234 640894 243854 676338
rect 243234 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 243854 640894
rect 243234 640574 243854 640658
rect 243234 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 243854 640574
rect 243234 604894 243854 640338
rect 243234 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 243854 604894
rect 243234 604574 243854 604658
rect 243234 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 243854 604574
rect 243234 568894 243854 604338
rect 243234 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 243854 568894
rect 243234 568574 243854 568658
rect 243234 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 243854 568574
rect 243234 537993 243854 568338
rect 246954 680614 247574 711002
rect 264954 710598 265574 711590
rect 264954 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 265574 710598
rect 264954 710278 265574 710362
rect 264954 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 265574 710278
rect 261234 708678 261854 709670
rect 261234 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 261854 708678
rect 261234 708358 261854 708442
rect 261234 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 261854 708358
rect 257514 706758 258134 707750
rect 257514 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 258134 706758
rect 257514 706438 258134 706522
rect 257514 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 258134 706438
rect 246954 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 247574 680614
rect 246954 680294 247574 680378
rect 246954 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 247574 680294
rect 246954 644614 247574 680058
rect 246954 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 247574 644614
rect 246954 644294 247574 644378
rect 246954 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 247574 644294
rect 246954 608614 247574 644058
rect 246954 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 247574 608614
rect 246954 608294 247574 608378
rect 246954 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 247574 608294
rect 246954 572614 247574 608058
rect 246954 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 247574 572614
rect 246954 572294 247574 572378
rect 246954 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 247574 572294
rect 246954 537993 247574 572058
rect 253794 704838 254414 705830
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 615454 254414 650898
rect 253794 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 254414 615454
rect 253794 615134 254414 615218
rect 253794 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 254414 615134
rect 253794 579454 254414 614898
rect 253794 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 254414 579454
rect 253794 579134 254414 579218
rect 253794 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 254414 579134
rect 253794 543454 254414 578898
rect 253794 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 254414 543454
rect 253794 543134 254414 543218
rect 253794 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 254414 543134
rect 253794 537993 254414 542898
rect 257514 691174 258134 706202
rect 257514 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 258134 691174
rect 257514 690854 258134 690938
rect 257514 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 258134 690854
rect 257514 655174 258134 690618
rect 257514 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 258134 655174
rect 257514 654854 258134 654938
rect 257514 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 258134 654854
rect 257514 619174 258134 654618
rect 257514 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 258134 619174
rect 257514 618854 258134 618938
rect 257514 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 258134 618854
rect 257514 583174 258134 618618
rect 257514 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 258134 583174
rect 257514 582854 258134 582938
rect 257514 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 258134 582854
rect 257514 547174 258134 582618
rect 257514 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 258134 547174
rect 257514 546854 258134 546938
rect 257514 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 258134 546854
rect 257514 537993 258134 546618
rect 261234 694894 261854 708122
rect 261234 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 261854 694894
rect 261234 694574 261854 694658
rect 261234 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 261854 694574
rect 261234 658894 261854 694338
rect 261234 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 261854 658894
rect 261234 658574 261854 658658
rect 261234 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 261854 658574
rect 261234 622894 261854 658338
rect 261234 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 261854 622894
rect 261234 622574 261854 622658
rect 261234 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 261854 622574
rect 261234 586894 261854 622338
rect 261234 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 261854 586894
rect 261234 586574 261854 586658
rect 261234 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 261854 586574
rect 261234 550894 261854 586338
rect 261234 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 261854 550894
rect 261234 550574 261854 550658
rect 261234 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 261854 550574
rect 261234 537993 261854 550338
rect 264954 698614 265574 710042
rect 282954 711558 283574 711590
rect 282954 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 283574 711558
rect 282954 711238 283574 711322
rect 282954 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 283574 711238
rect 279234 709638 279854 709670
rect 279234 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 279854 709638
rect 279234 709318 279854 709402
rect 279234 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 279854 709318
rect 275514 707718 276134 707750
rect 275514 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 276134 707718
rect 275514 707398 276134 707482
rect 275514 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 276134 707398
rect 264954 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 265574 698614
rect 264954 698294 265574 698378
rect 264954 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 265574 698294
rect 264954 662614 265574 698058
rect 264954 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 265574 662614
rect 264954 662294 265574 662378
rect 264954 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 265574 662294
rect 264954 626614 265574 662058
rect 264954 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 265574 626614
rect 264954 626294 265574 626378
rect 264954 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 265574 626294
rect 264954 590614 265574 626058
rect 264954 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 265574 590614
rect 264954 590294 265574 590378
rect 264954 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 265574 590294
rect 264954 554614 265574 590058
rect 264954 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 265574 554614
rect 264954 554294 265574 554378
rect 264954 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 265574 554294
rect 264954 537993 265574 554058
rect 271794 705798 272414 705830
rect 271794 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 272414 705798
rect 271794 705478 272414 705562
rect 271794 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 272414 705478
rect 271794 669454 272414 705242
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 633454 272414 668898
rect 271794 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 272414 633454
rect 271794 633134 272414 633218
rect 271794 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 272414 633134
rect 271794 597454 272414 632898
rect 271794 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 272414 597454
rect 271794 597134 272414 597218
rect 271794 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 272414 597134
rect 271794 561454 272414 596898
rect 271794 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 272414 561454
rect 271794 561134 272414 561218
rect 271794 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 272414 561134
rect 271794 537993 272414 560898
rect 275514 673174 276134 707162
rect 275514 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 276134 673174
rect 275514 672854 276134 672938
rect 275514 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 276134 672854
rect 275514 637174 276134 672618
rect 275514 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 276134 637174
rect 275514 636854 276134 636938
rect 275514 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 276134 636854
rect 275514 601174 276134 636618
rect 275514 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 276134 601174
rect 275514 600854 276134 600938
rect 275514 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 276134 600854
rect 275514 565174 276134 600618
rect 275514 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 276134 565174
rect 275514 564854 276134 564938
rect 275514 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 276134 564854
rect 275514 537993 276134 564618
rect 279234 676894 279854 709082
rect 279234 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 279854 676894
rect 279234 676574 279854 676658
rect 279234 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 279854 676574
rect 279234 640894 279854 676338
rect 279234 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 279854 640894
rect 279234 640574 279854 640658
rect 279234 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 279854 640574
rect 279234 604894 279854 640338
rect 279234 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 279854 604894
rect 279234 604574 279854 604658
rect 279234 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 279854 604574
rect 279234 568894 279854 604338
rect 279234 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 279854 568894
rect 279234 568574 279854 568658
rect 279234 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 279854 568574
rect 279234 537993 279854 568338
rect 282954 680614 283574 711002
rect 300954 710598 301574 711590
rect 300954 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 301574 710598
rect 300954 710278 301574 710362
rect 300954 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 301574 710278
rect 297234 708678 297854 709670
rect 297234 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 297854 708678
rect 297234 708358 297854 708442
rect 297234 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 297854 708358
rect 293514 706758 294134 707750
rect 293514 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 294134 706758
rect 293514 706438 294134 706522
rect 293514 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 294134 706438
rect 282954 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 283574 680614
rect 282954 680294 283574 680378
rect 282954 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 283574 680294
rect 282954 644614 283574 680058
rect 282954 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 283574 644614
rect 282954 644294 283574 644378
rect 282954 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 283574 644294
rect 282954 608614 283574 644058
rect 282954 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 283574 608614
rect 282954 608294 283574 608378
rect 282954 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 283574 608294
rect 282954 572614 283574 608058
rect 282954 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 283574 572614
rect 282954 572294 283574 572378
rect 282954 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 283574 572294
rect 282954 537993 283574 572058
rect 289794 704838 290414 705830
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 543454 290414 578898
rect 289794 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 290414 543454
rect 289794 543134 290414 543218
rect 289794 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 290414 543134
rect 289794 537993 290414 542898
rect 293514 691174 294134 706202
rect 293514 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 294134 691174
rect 293514 690854 294134 690938
rect 293514 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 294134 690854
rect 293514 655174 294134 690618
rect 293514 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 294134 655174
rect 293514 654854 294134 654938
rect 293514 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 294134 654854
rect 293514 619174 294134 654618
rect 293514 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 294134 619174
rect 293514 618854 294134 618938
rect 293514 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 294134 618854
rect 293514 583174 294134 618618
rect 293514 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 294134 583174
rect 293514 582854 294134 582938
rect 293514 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 294134 582854
rect 293514 547174 294134 582618
rect 293514 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 294134 547174
rect 293514 546854 294134 546938
rect 293514 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 294134 546854
rect 293514 537993 294134 546618
rect 297234 694894 297854 708122
rect 297234 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 297854 694894
rect 297234 694574 297854 694658
rect 297234 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 297854 694574
rect 297234 658894 297854 694338
rect 297234 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 297854 658894
rect 297234 658574 297854 658658
rect 297234 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 297854 658574
rect 297234 622894 297854 658338
rect 297234 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 297854 622894
rect 297234 622574 297854 622658
rect 297234 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 297854 622574
rect 297234 586894 297854 622338
rect 297234 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 297854 586894
rect 297234 586574 297854 586658
rect 297234 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 297854 586574
rect 297234 550894 297854 586338
rect 297234 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 297854 550894
rect 297234 550574 297854 550658
rect 297234 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 297854 550574
rect 297234 537993 297854 550338
rect 300954 698614 301574 710042
rect 318954 711558 319574 711590
rect 318954 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 319574 711558
rect 318954 711238 319574 711322
rect 318954 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 319574 711238
rect 315234 709638 315854 709670
rect 315234 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 315854 709638
rect 315234 709318 315854 709402
rect 315234 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 315854 709318
rect 311514 707718 312134 707750
rect 311514 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 312134 707718
rect 311514 707398 312134 707482
rect 311514 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 312134 707398
rect 300954 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 301574 698614
rect 300954 698294 301574 698378
rect 300954 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 301574 698294
rect 300954 662614 301574 698058
rect 300954 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 301574 662614
rect 300954 662294 301574 662378
rect 300954 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 301574 662294
rect 300954 626614 301574 662058
rect 300954 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 301574 626614
rect 300954 626294 301574 626378
rect 300954 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 301574 626294
rect 300954 590614 301574 626058
rect 300954 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 301574 590614
rect 300954 590294 301574 590378
rect 300954 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 301574 590294
rect 300954 554614 301574 590058
rect 300954 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 301574 554614
rect 300954 554294 301574 554378
rect 300954 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 301574 554294
rect 300954 537993 301574 554058
rect 307794 705798 308414 705830
rect 307794 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 308414 705798
rect 307794 705478 308414 705562
rect 307794 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 308414 705478
rect 307794 669454 308414 705242
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 633454 308414 668898
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 307794 597454 308414 632898
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 307794 561454 308414 596898
rect 307794 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 308414 561454
rect 307794 561134 308414 561218
rect 307794 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 308414 561134
rect 307794 537993 308414 560898
rect 311514 673174 312134 707162
rect 311514 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 312134 673174
rect 311514 672854 312134 672938
rect 311514 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 312134 672854
rect 311514 637174 312134 672618
rect 311514 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 312134 637174
rect 311514 636854 312134 636938
rect 311514 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 312134 636854
rect 311514 601174 312134 636618
rect 311514 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 312134 601174
rect 311514 600854 312134 600938
rect 311514 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 312134 600854
rect 311514 565174 312134 600618
rect 311514 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 312134 565174
rect 311514 564854 312134 564938
rect 311514 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 312134 564854
rect 311514 537993 312134 564618
rect 315234 676894 315854 709082
rect 315234 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 315854 676894
rect 315234 676574 315854 676658
rect 315234 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 315854 676574
rect 315234 640894 315854 676338
rect 315234 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 315854 640894
rect 315234 640574 315854 640658
rect 315234 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 315854 640574
rect 315234 604894 315854 640338
rect 315234 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 315854 604894
rect 315234 604574 315854 604658
rect 315234 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 315854 604574
rect 315234 568894 315854 604338
rect 315234 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 315854 568894
rect 315234 568574 315854 568658
rect 315234 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 315854 568574
rect 315234 537993 315854 568338
rect 318954 680614 319574 711002
rect 336954 710598 337574 711590
rect 336954 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 337574 710598
rect 336954 710278 337574 710362
rect 336954 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 337574 710278
rect 333234 708678 333854 709670
rect 333234 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 333854 708678
rect 333234 708358 333854 708442
rect 333234 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 333854 708358
rect 329514 706758 330134 707750
rect 329514 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 330134 706758
rect 329514 706438 330134 706522
rect 329514 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 330134 706438
rect 318954 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 319574 680614
rect 318954 680294 319574 680378
rect 318954 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 319574 680294
rect 318954 644614 319574 680058
rect 318954 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 319574 644614
rect 318954 644294 319574 644378
rect 318954 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 319574 644294
rect 318954 608614 319574 644058
rect 318954 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 319574 608614
rect 318954 608294 319574 608378
rect 318954 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 319574 608294
rect 318954 572614 319574 608058
rect 318954 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 319574 572614
rect 318954 572294 319574 572378
rect 318954 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 319574 572294
rect 318954 537993 319574 572058
rect 325794 704838 326414 705830
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 543454 326414 578898
rect 325794 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 326414 543454
rect 325794 543134 326414 543218
rect 325794 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 326414 543134
rect 325794 537993 326414 542898
rect 329514 691174 330134 706202
rect 329514 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 330134 691174
rect 329514 690854 330134 690938
rect 329514 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 330134 690854
rect 329514 655174 330134 690618
rect 329514 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 330134 655174
rect 329514 654854 330134 654938
rect 329514 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 330134 654854
rect 329514 619174 330134 654618
rect 329514 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 330134 619174
rect 329514 618854 330134 618938
rect 329514 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 330134 618854
rect 329514 583174 330134 618618
rect 329514 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 330134 583174
rect 329514 582854 330134 582938
rect 329514 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 330134 582854
rect 329514 547174 330134 582618
rect 329514 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 330134 547174
rect 329514 546854 330134 546938
rect 329514 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 330134 546854
rect 329514 537993 330134 546618
rect 333234 694894 333854 708122
rect 333234 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 333854 694894
rect 333234 694574 333854 694658
rect 333234 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 333854 694574
rect 333234 658894 333854 694338
rect 333234 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 333854 658894
rect 333234 658574 333854 658658
rect 333234 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 333854 658574
rect 333234 622894 333854 658338
rect 333234 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 333854 622894
rect 333234 622574 333854 622658
rect 333234 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 333854 622574
rect 333234 586894 333854 622338
rect 333234 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 333854 586894
rect 333234 586574 333854 586658
rect 333234 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 333854 586574
rect 333234 550894 333854 586338
rect 333234 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 333854 550894
rect 333234 550574 333854 550658
rect 333234 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 333854 550574
rect 333234 537993 333854 550338
rect 336954 698614 337574 710042
rect 354954 711558 355574 711590
rect 354954 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 355574 711558
rect 354954 711238 355574 711322
rect 354954 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 355574 711238
rect 351234 709638 351854 709670
rect 351234 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 351854 709638
rect 351234 709318 351854 709402
rect 351234 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 351854 709318
rect 347514 707718 348134 707750
rect 347514 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 348134 707718
rect 347514 707398 348134 707482
rect 347514 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 348134 707398
rect 336954 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 337574 698614
rect 336954 698294 337574 698378
rect 336954 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 337574 698294
rect 336954 662614 337574 698058
rect 336954 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 337574 662614
rect 336954 662294 337574 662378
rect 336954 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 337574 662294
rect 336954 626614 337574 662058
rect 336954 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 337574 626614
rect 336954 626294 337574 626378
rect 336954 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 337574 626294
rect 336954 590614 337574 626058
rect 336954 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 337574 590614
rect 336954 590294 337574 590378
rect 336954 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 337574 590294
rect 336954 554614 337574 590058
rect 336954 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 337574 554614
rect 336954 554294 337574 554378
rect 336954 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 337574 554294
rect 336954 537993 337574 554058
rect 343794 705798 344414 705830
rect 343794 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 344414 705798
rect 343794 705478 344414 705562
rect 343794 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 344414 705478
rect 343794 669454 344414 705242
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 633454 344414 668898
rect 343794 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 344414 633454
rect 343794 633134 344414 633218
rect 343794 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 344414 633134
rect 343794 597454 344414 632898
rect 343794 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 344414 597454
rect 343794 597134 344414 597218
rect 343794 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 344414 597134
rect 343794 561454 344414 596898
rect 343794 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 344414 561454
rect 343794 561134 344414 561218
rect 343794 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 344414 561134
rect 343794 537993 344414 560898
rect 347514 673174 348134 707162
rect 347514 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 348134 673174
rect 347514 672854 348134 672938
rect 347514 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 348134 672854
rect 347514 637174 348134 672618
rect 347514 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 348134 637174
rect 347514 636854 348134 636938
rect 347514 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 348134 636854
rect 347514 601174 348134 636618
rect 347514 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 348134 601174
rect 347514 600854 348134 600938
rect 347514 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 348134 600854
rect 347514 565174 348134 600618
rect 347514 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 348134 565174
rect 347514 564854 348134 564938
rect 347514 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 348134 564854
rect 347514 537993 348134 564618
rect 351234 676894 351854 709082
rect 351234 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 351854 676894
rect 351234 676574 351854 676658
rect 351234 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 351854 676574
rect 351234 640894 351854 676338
rect 351234 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 351854 640894
rect 351234 640574 351854 640658
rect 351234 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 351854 640574
rect 351234 604894 351854 640338
rect 351234 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 351854 604894
rect 351234 604574 351854 604658
rect 351234 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 351854 604574
rect 351234 568894 351854 604338
rect 351234 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 351854 568894
rect 351234 568574 351854 568658
rect 351234 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 351854 568574
rect 351234 537993 351854 568338
rect 354954 680614 355574 711002
rect 372954 710598 373574 711590
rect 372954 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 373574 710598
rect 372954 710278 373574 710362
rect 372954 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 373574 710278
rect 369234 708678 369854 709670
rect 369234 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 369854 708678
rect 369234 708358 369854 708442
rect 369234 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 369854 708358
rect 365514 706758 366134 707750
rect 365514 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 366134 706758
rect 365514 706438 366134 706522
rect 365514 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 366134 706438
rect 354954 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 355574 680614
rect 354954 680294 355574 680378
rect 354954 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 355574 680294
rect 354954 644614 355574 680058
rect 354954 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 355574 644614
rect 354954 644294 355574 644378
rect 354954 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 355574 644294
rect 354954 608614 355574 644058
rect 354954 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 355574 608614
rect 354954 608294 355574 608378
rect 354954 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 355574 608294
rect 354954 572614 355574 608058
rect 354954 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 355574 572614
rect 354954 572294 355574 572378
rect 354954 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 355574 572294
rect 353339 541380 353405 541381
rect 353339 541316 353340 541380
rect 353404 541316 353405 541380
rect 353339 541315 353405 541316
rect 199515 535532 199581 535533
rect 199515 535468 199516 535532
rect 199580 535468 199581 535532
rect 200619 535532 200685 535533
rect 200619 535530 200620 535532
rect 199515 535467 199581 535468
rect 200254 535470 200620 535530
rect 199518 523701 199578 535467
rect 200254 532810 200314 535470
rect 200619 535468 200620 535470
rect 200684 535468 200685 535532
rect 200619 535467 200685 535468
rect 200070 532750 200314 532810
rect 200070 532541 200130 532750
rect 200067 532540 200133 532541
rect 200067 532476 200068 532540
rect 200132 532476 200133 532540
rect 200067 532475 200133 532476
rect 219568 525454 219888 525486
rect 219568 525218 219610 525454
rect 219846 525218 219888 525454
rect 219568 525134 219888 525218
rect 219568 524898 219610 525134
rect 219846 524898 219888 525134
rect 219568 524866 219888 524898
rect 250288 525454 250608 525486
rect 250288 525218 250330 525454
rect 250566 525218 250608 525454
rect 250288 525134 250608 525218
rect 250288 524898 250330 525134
rect 250566 524898 250608 525134
rect 250288 524866 250608 524898
rect 281008 525454 281328 525486
rect 281008 525218 281050 525454
rect 281286 525218 281328 525454
rect 281008 525134 281328 525218
rect 281008 524898 281050 525134
rect 281286 524898 281328 525134
rect 281008 524866 281328 524898
rect 311728 525454 312048 525486
rect 311728 525218 311770 525454
rect 312006 525218 312048 525454
rect 311728 525134 312048 525218
rect 311728 524898 311770 525134
rect 312006 524898 312048 525134
rect 311728 524866 312048 524898
rect 342448 525454 342768 525486
rect 342448 525218 342490 525454
rect 342726 525218 342768 525454
rect 342448 525134 342768 525218
rect 342448 524898 342490 525134
rect 342726 524898 342768 525134
rect 342448 524866 342768 524898
rect 199515 523700 199581 523701
rect 199515 523636 199516 523700
rect 199580 523636 199581 523700
rect 199515 523635 199581 523636
rect 199331 513364 199397 513365
rect 199331 513300 199332 513364
rect 199396 513300 199397 513364
rect 199331 513299 199397 513300
rect 204208 507454 204528 507486
rect 204208 507218 204250 507454
rect 204486 507218 204528 507454
rect 204208 507134 204528 507218
rect 204208 506898 204250 507134
rect 204486 506898 204528 507134
rect 204208 506866 204528 506898
rect 234928 507454 235248 507486
rect 234928 507218 234970 507454
rect 235206 507218 235248 507454
rect 234928 507134 235248 507218
rect 234928 506898 234970 507134
rect 235206 506898 235248 507134
rect 234928 506866 235248 506898
rect 265648 507454 265968 507486
rect 265648 507218 265690 507454
rect 265926 507218 265968 507454
rect 265648 507134 265968 507218
rect 265648 506898 265690 507134
rect 265926 506898 265968 507134
rect 265648 506866 265968 506898
rect 296368 507454 296688 507486
rect 296368 507218 296410 507454
rect 296646 507218 296688 507454
rect 296368 507134 296688 507218
rect 296368 506898 296410 507134
rect 296646 506898 296688 507134
rect 296368 506866 296688 506898
rect 327088 507454 327408 507486
rect 327088 507218 327130 507454
rect 327366 507218 327408 507454
rect 327088 507134 327408 507218
rect 327088 506898 327130 507134
rect 327366 506898 327408 507134
rect 327088 506866 327408 506898
rect 198595 500444 198661 500445
rect 198595 500380 198596 500444
rect 198660 500380 198661 500444
rect 198595 500379 198661 500380
rect 219568 489454 219888 489486
rect 219568 489218 219610 489454
rect 219846 489218 219888 489454
rect 219568 489134 219888 489218
rect 219568 488898 219610 489134
rect 219846 488898 219888 489134
rect 219568 488866 219888 488898
rect 250288 489454 250608 489486
rect 250288 489218 250330 489454
rect 250566 489218 250608 489454
rect 250288 489134 250608 489218
rect 250288 488898 250330 489134
rect 250566 488898 250608 489134
rect 250288 488866 250608 488898
rect 281008 489454 281328 489486
rect 281008 489218 281050 489454
rect 281286 489218 281328 489454
rect 281008 489134 281328 489218
rect 281008 488898 281050 489134
rect 281286 488898 281328 489134
rect 281008 488866 281328 488898
rect 311728 489454 312048 489486
rect 311728 489218 311770 489454
rect 312006 489218 312048 489454
rect 311728 489134 312048 489218
rect 311728 488898 311770 489134
rect 312006 488898 312048 489134
rect 311728 488866 312048 488898
rect 342448 489454 342768 489486
rect 342448 489218 342490 489454
rect 342726 489218 342768 489454
rect 342448 489134 342768 489218
rect 342448 488898 342490 489134
rect 342726 488898 342768 489134
rect 342448 488866 342768 488898
rect 198411 483172 198477 483173
rect 198411 483108 198412 483172
rect 198476 483108 198477 483172
rect 198411 483107 198477 483108
rect 197307 384980 197373 384981
rect 197307 384916 197308 384980
rect 197372 384916 197373 384980
rect 197307 384915 197373 384916
rect 197310 383757 197370 384915
rect 197307 383756 197373 383757
rect 197307 383692 197308 383756
rect 197372 383692 197373 383756
rect 197307 383691 197373 383692
rect 197310 378045 197370 383691
rect 197307 378044 197373 378045
rect 197307 377980 197308 378044
rect 197372 377980 197373 378044
rect 197307 377979 197373 377980
rect 198414 345133 198474 483107
rect 204208 471454 204528 471486
rect 204208 471218 204250 471454
rect 204486 471218 204528 471454
rect 204208 471134 204528 471218
rect 204208 470898 204250 471134
rect 204486 470898 204528 471134
rect 204208 470866 204528 470898
rect 234928 471454 235248 471486
rect 234928 471218 234970 471454
rect 235206 471218 235248 471454
rect 234928 471134 235248 471218
rect 234928 470898 234970 471134
rect 235206 470898 235248 471134
rect 234928 470866 235248 470898
rect 265648 471454 265968 471486
rect 265648 471218 265690 471454
rect 265926 471218 265968 471454
rect 265648 471134 265968 471218
rect 265648 470898 265690 471134
rect 265926 470898 265968 471134
rect 265648 470866 265968 470898
rect 296368 471454 296688 471486
rect 296368 471218 296410 471454
rect 296646 471218 296688 471454
rect 296368 471134 296688 471218
rect 296368 470898 296410 471134
rect 296646 470898 296688 471134
rect 296368 470866 296688 470898
rect 327088 471454 327408 471486
rect 327088 471218 327130 471454
rect 327366 471218 327408 471454
rect 327088 471134 327408 471218
rect 327088 470898 327130 471134
rect 327366 470898 327408 471134
rect 327088 470866 327408 470898
rect 198779 458420 198845 458421
rect 198779 458356 198780 458420
rect 198844 458356 198845 458420
rect 198779 458355 198845 458356
rect 198595 421700 198661 421701
rect 198595 421636 198596 421700
rect 198660 421636 198661 421700
rect 198595 421635 198661 421636
rect 198411 345132 198477 345133
rect 198411 345068 198412 345132
rect 198476 345068 198477 345132
rect 198411 345067 198477 345068
rect 196571 344996 196637 344997
rect 196571 344932 196572 344996
rect 196636 344932 196637 344996
rect 196571 344931 196637 344932
rect 198414 327181 198474 345067
rect 198411 327180 198477 327181
rect 198411 327116 198412 327180
rect 198476 327116 198477 327180
rect 198411 327115 198477 327116
rect 197123 301476 197189 301477
rect 197123 301412 197124 301476
rect 197188 301412 197189 301476
rect 197123 301411 197189 301412
rect 195283 273324 195349 273325
rect 195283 273260 195284 273324
rect 195348 273260 195349 273324
rect 195283 273259 195349 273260
rect 195099 262988 195165 262989
rect 195099 262924 195100 262988
rect 195164 262924 195165 262988
rect 195099 262923 195165 262924
rect 195286 261629 195346 273259
rect 197126 267205 197186 301411
rect 198414 271013 198474 327115
rect 198411 271012 198477 271013
rect 198411 270948 198412 271012
rect 198476 270948 198477 271012
rect 198411 270947 198477 270948
rect 197123 267204 197189 267205
rect 197123 267140 197124 267204
rect 197188 267140 197189 267204
rect 197123 267139 197189 267140
rect 197123 265028 197189 265029
rect 197123 264964 197124 265028
rect 197188 264964 197189 265028
rect 197123 264963 197189 264964
rect 195283 261628 195349 261629
rect 195283 261564 195284 261628
rect 195348 261564 195349 261628
rect 195283 261563 195349 261564
rect 195835 260948 195901 260949
rect 195835 260884 195836 260948
rect 195900 260884 195901 260948
rect 195835 260883 195901 260884
rect 195099 249932 195165 249933
rect 195099 249868 195100 249932
rect 195164 249868 195165 249932
rect 195099 249867 195165 249868
rect 193811 245852 193877 245853
rect 193811 245788 193812 245852
rect 193876 245788 193877 245852
rect 193811 245787 193877 245788
rect 192954 230378 192986 230614
rect 193222 230378 193306 230614
rect 193542 230378 193574 230614
rect 192954 230294 193574 230378
rect 192954 230058 192986 230294
rect 193222 230058 193306 230294
rect 193542 230058 193574 230294
rect 192954 194614 193574 230058
rect 193814 212533 193874 245787
rect 195102 237285 195162 249867
rect 195838 248430 195898 260883
rect 195838 248370 196634 248430
rect 195835 245716 195901 245717
rect 195835 245652 195836 245716
rect 195900 245652 195901 245716
rect 195835 245651 195901 245652
rect 195099 237284 195165 237285
rect 195099 237220 195100 237284
rect 195164 237220 195165 237284
rect 195099 237219 195165 237220
rect 195651 231164 195717 231165
rect 195651 231100 195652 231164
rect 195716 231100 195717 231164
rect 195651 231099 195717 231100
rect 193811 212532 193877 212533
rect 193811 212468 193812 212532
rect 193876 212468 193877 212532
rect 193811 212467 193877 212468
rect 195654 203693 195714 231099
rect 195838 229805 195898 245651
rect 195835 229804 195901 229805
rect 195835 229740 195836 229804
rect 195900 229740 195901 229804
rect 195835 229739 195901 229740
rect 196574 225045 196634 248370
rect 197126 246533 197186 264963
rect 198598 251837 198658 421635
rect 198782 369205 198842 458355
rect 219568 453454 219888 453486
rect 219568 453218 219610 453454
rect 219846 453218 219888 453454
rect 219568 453134 219888 453218
rect 219568 452898 219610 453134
rect 219846 452898 219888 453134
rect 219568 452866 219888 452898
rect 250288 453454 250608 453486
rect 250288 453218 250330 453454
rect 250566 453218 250608 453454
rect 250288 453134 250608 453218
rect 250288 452898 250330 453134
rect 250566 452898 250608 453134
rect 250288 452866 250608 452898
rect 281008 453454 281328 453486
rect 281008 453218 281050 453454
rect 281286 453218 281328 453454
rect 281008 453134 281328 453218
rect 281008 452898 281050 453134
rect 281286 452898 281328 453134
rect 281008 452866 281328 452898
rect 311728 453454 312048 453486
rect 311728 453218 311770 453454
rect 312006 453218 312048 453454
rect 311728 453134 312048 453218
rect 311728 452898 311770 453134
rect 312006 452898 312048 453134
rect 311728 452866 312048 452898
rect 342448 453454 342768 453486
rect 342448 453218 342490 453454
rect 342726 453218 342768 453454
rect 342448 453134 342768 453218
rect 342448 452898 342490 453134
rect 342726 452898 342768 453134
rect 342448 452866 342768 452898
rect 204208 435454 204528 435486
rect 204208 435218 204250 435454
rect 204486 435218 204528 435454
rect 204208 435134 204528 435218
rect 204208 434898 204250 435134
rect 204486 434898 204528 435134
rect 204208 434866 204528 434898
rect 234928 435454 235248 435486
rect 234928 435218 234970 435454
rect 235206 435218 235248 435454
rect 234928 435134 235248 435218
rect 234928 434898 234970 435134
rect 235206 434898 235248 435134
rect 234928 434866 235248 434898
rect 265648 435454 265968 435486
rect 265648 435218 265690 435454
rect 265926 435218 265968 435454
rect 265648 435134 265968 435218
rect 265648 434898 265690 435134
rect 265926 434898 265968 435134
rect 265648 434866 265968 434898
rect 296368 435454 296688 435486
rect 296368 435218 296410 435454
rect 296646 435218 296688 435454
rect 296368 435134 296688 435218
rect 296368 434898 296410 435134
rect 296646 434898 296688 435134
rect 296368 434866 296688 434898
rect 327088 435454 327408 435486
rect 327088 435218 327130 435454
rect 327366 435218 327408 435454
rect 327088 435134 327408 435218
rect 327088 434898 327130 435134
rect 327366 434898 327408 435134
rect 327088 434866 327408 434898
rect 198963 419660 199029 419661
rect 198963 419596 198964 419660
rect 199028 419596 199029 419660
rect 198963 419595 199029 419596
rect 198966 376549 199026 419595
rect 219568 417454 219888 417486
rect 219568 417218 219610 417454
rect 219846 417218 219888 417454
rect 219568 417134 219888 417218
rect 219568 416898 219610 417134
rect 219846 416898 219888 417134
rect 219568 416866 219888 416898
rect 250288 417454 250608 417486
rect 250288 417218 250330 417454
rect 250566 417218 250608 417454
rect 250288 417134 250608 417218
rect 250288 416898 250330 417134
rect 250566 416898 250608 417134
rect 250288 416866 250608 416898
rect 281008 417454 281328 417486
rect 281008 417218 281050 417454
rect 281286 417218 281328 417454
rect 281008 417134 281328 417218
rect 281008 416898 281050 417134
rect 281286 416898 281328 417134
rect 281008 416866 281328 416898
rect 311728 417454 312048 417486
rect 311728 417218 311770 417454
rect 312006 417218 312048 417454
rect 311728 417134 312048 417218
rect 311728 416898 311770 417134
rect 312006 416898 312048 417134
rect 311728 416866 312048 416898
rect 342448 417454 342768 417486
rect 342448 417218 342490 417454
rect 342726 417218 342768 417454
rect 342448 417134 342768 417218
rect 342448 416898 342490 417134
rect 342726 416898 342768 417134
rect 342448 416866 342768 416898
rect 204208 399454 204528 399486
rect 204208 399218 204250 399454
rect 204486 399218 204528 399454
rect 204208 399134 204528 399218
rect 204208 398898 204250 399134
rect 204486 398898 204528 399134
rect 204208 398866 204528 398898
rect 234928 399454 235248 399486
rect 234928 399218 234970 399454
rect 235206 399218 235248 399454
rect 234928 399134 235248 399218
rect 234928 398898 234970 399134
rect 235206 398898 235248 399134
rect 234928 398866 235248 398898
rect 265648 399454 265968 399486
rect 265648 399218 265690 399454
rect 265926 399218 265968 399454
rect 265648 399134 265968 399218
rect 265648 398898 265690 399134
rect 265926 398898 265968 399134
rect 265648 398866 265968 398898
rect 296368 399454 296688 399486
rect 296368 399218 296410 399454
rect 296646 399218 296688 399454
rect 296368 399134 296688 399218
rect 296368 398898 296410 399134
rect 296646 398898 296688 399134
rect 296368 398866 296688 398898
rect 327088 399454 327408 399486
rect 327088 399218 327130 399454
rect 327366 399218 327408 399454
rect 327088 399134 327408 399218
rect 327088 398898 327130 399134
rect 327366 398898 327408 399134
rect 327088 398866 327408 398898
rect 219568 381454 219888 381486
rect 219568 381218 219610 381454
rect 219846 381218 219888 381454
rect 219568 381134 219888 381218
rect 219568 380898 219610 381134
rect 219846 380898 219888 381134
rect 219568 380866 219888 380898
rect 250288 381454 250608 381486
rect 250288 381218 250330 381454
rect 250566 381218 250608 381454
rect 250288 381134 250608 381218
rect 250288 380898 250330 381134
rect 250566 380898 250608 381134
rect 250288 380866 250608 380898
rect 281008 381454 281328 381486
rect 281008 381218 281050 381454
rect 281286 381218 281328 381454
rect 281008 381134 281328 381218
rect 281008 380898 281050 381134
rect 281286 380898 281328 381134
rect 281008 380866 281328 380898
rect 311728 381454 312048 381486
rect 311728 381218 311770 381454
rect 312006 381218 312048 381454
rect 311728 381134 312048 381218
rect 311728 380898 311770 381134
rect 312006 380898 312048 381134
rect 311728 380866 312048 380898
rect 342448 381454 342768 381486
rect 342448 381218 342490 381454
rect 342726 381218 342768 381454
rect 342448 381134 342768 381218
rect 342448 380898 342490 381134
rect 342726 380898 342768 381134
rect 342448 380866 342768 380898
rect 200619 378316 200685 378317
rect 200619 378252 200620 378316
rect 200684 378252 200685 378316
rect 200619 378251 200685 378252
rect 198963 376548 199029 376549
rect 198963 376484 198964 376548
rect 199028 376484 199029 376548
rect 198963 376483 199029 376484
rect 198779 369204 198845 369205
rect 198779 369140 198780 369204
rect 198844 369140 198845 369204
rect 198779 369139 198845 369140
rect 199794 345454 200414 375600
rect 200622 367709 200682 378251
rect 200619 367708 200685 367709
rect 200619 367644 200620 367708
rect 200684 367644 200685 367708
rect 200619 367643 200685 367644
rect 203011 361860 203077 361861
rect 203011 361796 203012 361860
rect 203076 361796 203077 361860
rect 203011 361795 203077 361796
rect 199794 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 200414 345454
rect 199794 345134 200414 345218
rect 199794 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 200414 345134
rect 199331 312492 199397 312493
rect 199331 312428 199332 312492
rect 199396 312428 199397 312492
rect 199331 312427 199397 312428
rect 198779 282980 198845 282981
rect 198779 282916 198780 282980
rect 198844 282916 198845 282980
rect 198779 282915 198845 282916
rect 198782 273325 198842 282915
rect 198779 273324 198845 273325
rect 198779 273260 198780 273324
rect 198844 273260 198845 273324
rect 198779 273259 198845 273260
rect 199334 265029 199394 312427
rect 199794 309454 200414 344898
rect 199794 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 200414 309454
rect 199794 309134 200414 309218
rect 199794 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 200414 309134
rect 199794 286182 200414 308898
rect 202643 297532 202709 297533
rect 202643 297468 202644 297532
rect 202708 297468 202709 297532
rect 202643 297467 202709 297468
rect 200251 285972 200317 285973
rect 200251 285908 200252 285972
rect 200316 285908 200317 285972
rect 200251 285907 200317 285908
rect 200067 279852 200133 279853
rect 200067 279788 200068 279852
rect 200132 279850 200133 279852
rect 200254 279850 200314 285907
rect 200132 279790 200314 279850
rect 200132 279788 200133 279790
rect 200067 279787 200133 279788
rect 199331 265028 199397 265029
rect 199331 264964 199332 265028
rect 199396 264964 199397 265028
rect 199331 264963 199397 264964
rect 198595 251836 198661 251837
rect 198595 251772 198596 251836
rect 198660 251772 198661 251836
rect 198595 251771 198661 251772
rect 197123 246532 197189 246533
rect 197123 246468 197124 246532
rect 197188 246468 197189 246532
rect 197123 246467 197189 246468
rect 197126 245853 197186 246467
rect 197123 245852 197189 245853
rect 197123 245788 197124 245852
rect 197188 245788 197189 245852
rect 197123 245787 197189 245788
rect 199331 243132 199397 243133
rect 199331 243068 199332 243132
rect 199396 243068 199397 243132
rect 199331 243067 199397 243068
rect 196755 241772 196821 241773
rect 196755 241708 196756 241772
rect 196820 241708 196821 241772
rect 196755 241707 196821 241708
rect 196758 237421 196818 241707
rect 196755 237420 196821 237421
rect 196755 237356 196756 237420
rect 196820 237356 196821 237420
rect 196755 237355 196821 237356
rect 199334 237013 199394 243067
rect 202646 240141 202706 297467
rect 202643 240140 202709 240141
rect 202643 240076 202644 240140
rect 202708 240076 202709 240140
rect 202643 240075 202709 240076
rect 203014 240005 203074 361795
rect 203514 349174 204134 375600
rect 203514 348938 203546 349174
rect 203782 348938 203866 349174
rect 204102 348938 204134 349174
rect 203514 348854 204134 348938
rect 203514 348618 203546 348854
rect 203782 348618 203866 348854
rect 204102 348618 204134 348854
rect 203514 313174 204134 348618
rect 207234 352894 207854 375600
rect 207234 352658 207266 352894
rect 207502 352658 207586 352894
rect 207822 352658 207854 352894
rect 207234 352574 207854 352658
rect 207234 352338 207266 352574
rect 207502 352338 207586 352574
rect 207822 352338 207854 352574
rect 207234 316894 207854 352338
rect 210954 356614 211574 375600
rect 210954 356378 210986 356614
rect 211222 356378 211306 356614
rect 211542 356378 211574 356614
rect 210954 356294 211574 356378
rect 210954 356058 210986 356294
rect 211222 356058 211306 356294
rect 211542 356058 211574 356294
rect 208899 348532 208965 348533
rect 208899 348468 208900 348532
rect 208964 348468 208965 348532
rect 208899 348467 208965 348468
rect 207234 316658 207266 316894
rect 207502 316658 207586 316894
rect 207822 316658 207854 316894
rect 207234 316574 207854 316658
rect 207234 316338 207266 316574
rect 207502 316338 207586 316574
rect 207822 316338 207854 316574
rect 206875 314124 206941 314125
rect 206875 314060 206876 314124
rect 206940 314060 206941 314124
rect 206875 314059 206941 314060
rect 203514 312938 203546 313174
rect 203782 312938 203866 313174
rect 204102 312938 204134 313174
rect 203514 312854 204134 312938
rect 203514 312618 203546 312854
rect 203782 312618 203866 312854
rect 204102 312618 204134 312854
rect 203514 286182 204134 312618
rect 204408 255454 204728 255486
rect 204408 255218 204450 255454
rect 204686 255218 204728 255454
rect 204408 255134 204728 255218
rect 204408 254898 204450 255134
rect 204686 254898 204728 255134
rect 204408 254866 204728 254898
rect 203011 240004 203077 240005
rect 203011 239940 203012 240004
rect 203076 239940 203077 240004
rect 203011 239939 203077 239940
rect 206878 238645 206938 314059
rect 207234 286182 207854 316338
rect 208163 297396 208229 297397
rect 208163 297332 208164 297396
rect 208228 297332 208229 297396
rect 208163 297331 208229 297332
rect 208166 240141 208226 297331
rect 208902 240141 208962 348467
rect 210954 320614 211574 356058
rect 217794 363454 218414 375600
rect 217794 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 218414 363454
rect 217794 363134 218414 363218
rect 217794 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 218414 363134
rect 213131 337516 213197 337517
rect 213131 337452 213132 337516
rect 213196 337452 213197 337516
rect 213131 337451 213197 337452
rect 210954 320378 210986 320614
rect 211222 320378 211306 320614
rect 211542 320378 211574 320614
rect 210954 320294 211574 320378
rect 210954 320058 210986 320294
rect 211222 320058 211306 320294
rect 211542 320058 211574 320294
rect 210739 319564 210805 319565
rect 210739 319500 210740 319564
rect 210804 319500 210805 319564
rect 210739 319499 210805 319500
rect 210742 240141 210802 319499
rect 210954 286182 211574 320058
rect 211659 289916 211725 289917
rect 211659 289852 211660 289916
rect 211724 289852 211725 289916
rect 211659 289851 211725 289852
rect 208163 240140 208229 240141
rect 208163 240076 208164 240140
rect 208228 240076 208229 240140
rect 208163 240075 208229 240076
rect 208899 240140 208965 240141
rect 208899 240076 208900 240140
rect 208964 240076 208965 240140
rect 208899 240075 208965 240076
rect 210739 240140 210805 240141
rect 210739 240076 210740 240140
rect 210804 240076 210805 240140
rect 210739 240075 210805 240076
rect 206875 238644 206941 238645
rect 206875 238580 206876 238644
rect 206940 238580 206941 238644
rect 206875 238579 206941 238580
rect 199794 237454 200414 238182
rect 199794 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 200414 237454
rect 199794 237134 200414 237218
rect 199331 237012 199397 237013
rect 199331 236948 199332 237012
rect 199396 236948 199397 237012
rect 199331 236947 199397 236948
rect 199794 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 200414 237134
rect 196571 225044 196637 225045
rect 196571 224980 196572 225044
rect 196636 224980 196637 225044
rect 196571 224979 196637 224980
rect 195651 203692 195717 203693
rect 195651 203628 195652 203692
rect 195716 203628 195717 203692
rect 195651 203627 195717 203628
rect 192954 194378 192986 194614
rect 193222 194378 193306 194614
rect 193542 194378 193574 194614
rect 192954 194294 193574 194378
rect 192954 194058 192986 194294
rect 193222 194058 193306 194294
rect 193542 194058 193574 194294
rect 192954 158614 193574 194058
rect 199794 201454 200414 236898
rect 199794 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 200414 201454
rect 199794 201134 200414 201218
rect 199794 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 200414 201134
rect 197307 178804 197373 178805
rect 197307 178740 197308 178804
rect 197372 178740 197373 178804
rect 197307 178739 197373 178740
rect 192954 158378 192986 158614
rect 193222 158378 193306 158614
rect 193542 158378 193574 158614
rect 192954 158294 193574 158378
rect 192954 158058 192986 158294
rect 193222 158058 193306 158294
rect 193542 158058 193574 158294
rect 192954 122614 193574 158058
rect 192954 122378 192986 122614
rect 193222 122378 193306 122614
rect 193542 122378 193574 122614
rect 192954 122294 193574 122378
rect 192954 122058 192986 122294
rect 193222 122058 193306 122294
rect 193542 122058 193574 122294
rect 192954 86614 193574 122058
rect 197310 104821 197370 178739
rect 199794 165454 200414 200898
rect 199794 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 200414 165454
rect 199794 165134 200414 165218
rect 199794 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 200414 165134
rect 199794 129454 200414 164898
rect 199794 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 200414 129454
rect 199794 129134 200414 129218
rect 199794 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 200414 129134
rect 197307 104820 197373 104821
rect 197307 104756 197308 104820
rect 197372 104756 197373 104820
rect 197307 104755 197373 104756
rect 192954 86378 192986 86614
rect 193222 86378 193306 86614
rect 193542 86378 193574 86614
rect 192954 86294 193574 86378
rect 192954 86058 192986 86294
rect 193222 86058 193306 86294
rect 193542 86058 193574 86294
rect 191051 84828 191117 84829
rect 191051 84764 191052 84828
rect 191116 84764 191117 84828
rect 191051 84763 191117 84764
rect 189234 82658 189266 82894
rect 189502 82658 189586 82894
rect 189822 82658 189854 82894
rect 189234 82574 189854 82658
rect 189234 82338 189266 82574
rect 189502 82338 189586 82574
rect 189822 82338 189854 82574
rect 189234 46894 189854 82338
rect 189234 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 189854 46894
rect 189234 46574 189854 46658
rect 189234 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 189854 46574
rect 186819 35188 186885 35189
rect 186819 35124 186820 35188
rect 186884 35124 186885 35188
rect 186819 35123 186885 35124
rect 185514 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 186134 7174
rect 185514 6854 186134 6938
rect 185514 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 186134 6854
rect 185514 -2266 186134 6618
rect 185514 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 186134 -2266
rect 185514 -2586 186134 -2502
rect 185514 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 186134 -2586
rect 185514 -3814 186134 -2822
rect 189234 10894 189854 46338
rect 189234 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 189854 10894
rect 189234 10574 189854 10658
rect 189234 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 189854 10574
rect 189234 -4186 189854 10338
rect 189234 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 189854 -4186
rect 189234 -4506 189854 -4422
rect 189234 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 189854 -4506
rect 189234 -5734 189854 -4742
rect 192954 50614 193574 86058
rect 192954 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 193574 50614
rect 192954 50294 193574 50378
rect 192954 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 193574 50294
rect 192954 14614 193574 50058
rect 192954 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 193574 14614
rect 192954 14294 193574 14378
rect 192954 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 193574 14294
rect 174954 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 175574 -7066
rect 174954 -7386 175574 -7302
rect 174954 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 175574 -7386
rect 174954 -7654 175574 -7622
rect 192954 -6106 193574 14058
rect 199794 93454 200414 128898
rect 199794 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 200414 93454
rect 199794 93134 200414 93218
rect 199794 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 200414 93134
rect 199794 57454 200414 92898
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 199794 57134 200414 57218
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 199794 21454 200414 56898
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -1306 200414 20898
rect 199794 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 200414 -1306
rect 199794 -1626 200414 -1542
rect 199794 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 200414 -1626
rect 199794 -1894 200414 -1862
rect 203514 205174 204134 238182
rect 204851 226404 204917 226405
rect 204851 226340 204852 226404
rect 204916 226340 204917 226404
rect 204851 226339 204917 226340
rect 203514 204938 203546 205174
rect 203782 204938 203866 205174
rect 204102 204938 204134 205174
rect 203514 204854 204134 204938
rect 203514 204618 203546 204854
rect 203782 204618 203866 204854
rect 204102 204618 204134 204854
rect 203514 169174 204134 204618
rect 204854 200701 204914 226339
rect 207234 208894 207854 238182
rect 209819 237420 209885 237421
rect 209819 237356 209820 237420
rect 209884 237356 209885 237420
rect 209819 237355 209885 237356
rect 209822 215117 209882 237355
rect 209819 215116 209885 215117
rect 209819 215052 209820 215116
rect 209884 215052 209885 215116
rect 209819 215051 209885 215052
rect 207234 208658 207266 208894
rect 207502 208658 207586 208894
rect 207822 208658 207854 208894
rect 207234 208574 207854 208658
rect 207234 208338 207266 208574
rect 207502 208338 207586 208574
rect 207822 208338 207854 208574
rect 204851 200700 204917 200701
rect 204851 200636 204852 200700
rect 204916 200636 204917 200700
rect 204851 200635 204917 200636
rect 203514 168938 203546 169174
rect 203782 168938 203866 169174
rect 204102 168938 204134 169174
rect 203514 168854 204134 168938
rect 203514 168618 203546 168854
rect 203782 168618 203866 168854
rect 204102 168618 204134 168854
rect 203514 133174 204134 168618
rect 203514 132938 203546 133174
rect 203782 132938 203866 133174
rect 204102 132938 204134 133174
rect 203514 132854 204134 132938
rect 203514 132618 203546 132854
rect 203782 132618 203866 132854
rect 204102 132618 204134 132854
rect 203514 97174 204134 132618
rect 203514 96938 203546 97174
rect 203782 96938 203866 97174
rect 204102 96938 204134 97174
rect 203514 96854 204134 96938
rect 203514 96618 203546 96854
rect 203782 96618 203866 96854
rect 204102 96618 204134 96854
rect 203514 61174 204134 96618
rect 203514 60938 203546 61174
rect 203782 60938 203866 61174
rect 204102 60938 204134 61174
rect 203514 60854 204134 60938
rect 203514 60618 203546 60854
rect 203782 60618 203866 60854
rect 204102 60618 204134 60854
rect 203514 25174 204134 60618
rect 203514 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 204134 25174
rect 203514 24854 204134 24938
rect 203514 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 204134 24854
rect 203514 -3226 204134 24618
rect 203514 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 204134 -3226
rect 203514 -3546 204134 -3462
rect 203514 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 204134 -3546
rect 203514 -3814 204134 -3782
rect 207234 172894 207854 208338
rect 207234 172658 207266 172894
rect 207502 172658 207586 172894
rect 207822 172658 207854 172894
rect 207234 172574 207854 172658
rect 207234 172338 207266 172574
rect 207502 172338 207586 172574
rect 207822 172338 207854 172574
rect 207234 136894 207854 172338
rect 207234 136658 207266 136894
rect 207502 136658 207586 136894
rect 207822 136658 207854 136894
rect 207234 136574 207854 136658
rect 207234 136338 207266 136574
rect 207502 136338 207586 136574
rect 207822 136338 207854 136574
rect 207234 100894 207854 136338
rect 207234 100658 207266 100894
rect 207502 100658 207586 100894
rect 207822 100658 207854 100894
rect 207234 100574 207854 100658
rect 207234 100338 207266 100574
rect 207502 100338 207586 100574
rect 207822 100338 207854 100574
rect 207234 64894 207854 100338
rect 207234 64658 207266 64894
rect 207502 64658 207586 64894
rect 207822 64658 207854 64894
rect 207234 64574 207854 64658
rect 207234 64338 207266 64574
rect 207502 64338 207586 64574
rect 207822 64338 207854 64574
rect 207234 28894 207854 64338
rect 207234 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 207854 28894
rect 207234 28574 207854 28658
rect 207234 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 207854 28574
rect 207234 -5146 207854 28338
rect 207234 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 207854 -5146
rect 207234 -5466 207854 -5382
rect 207234 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 207854 -5466
rect 207234 -5734 207854 -5702
rect 210954 212614 211574 238182
rect 211662 237149 211722 289851
rect 211659 237148 211725 237149
rect 211659 237084 211660 237148
rect 211724 237084 211725 237148
rect 211659 237083 211725 237084
rect 213134 235517 213194 337451
rect 217794 327454 218414 362898
rect 221514 367174 222134 375600
rect 221514 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 222134 367174
rect 221514 366854 222134 366938
rect 221514 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 222134 366854
rect 219939 341460 220005 341461
rect 219939 341396 219940 341460
rect 220004 341396 220005 341460
rect 219939 341395 220005 341396
rect 217794 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 218414 327454
rect 217794 327134 218414 327218
rect 217794 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 218414 327134
rect 217547 293180 217613 293181
rect 217547 293116 217548 293180
rect 217612 293116 217613 293180
rect 217547 293115 217613 293116
rect 214419 283932 214485 283933
rect 214419 283868 214420 283932
rect 214484 283868 214485 283932
rect 214419 283867 214485 283868
rect 216443 283932 216509 283933
rect 216443 283868 216444 283932
rect 216508 283868 216509 283932
rect 216443 283867 216509 283868
rect 213131 235516 213197 235517
rect 213131 235452 213132 235516
rect 213196 235452 213197 235516
rect 213131 235451 213197 235452
rect 210954 212378 210986 212614
rect 211222 212378 211306 212614
rect 211542 212378 211574 212614
rect 210954 212294 211574 212378
rect 210954 212058 210986 212294
rect 211222 212058 211306 212294
rect 211542 212058 211574 212294
rect 210954 176614 211574 212058
rect 214422 205597 214482 283867
rect 216446 212669 216506 283867
rect 217550 240141 217610 293115
rect 217794 291454 218414 326898
rect 219203 296172 219269 296173
rect 219203 296108 219204 296172
rect 219268 296108 219269 296172
rect 219203 296107 219269 296108
rect 217794 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 218414 291454
rect 217794 291134 218414 291218
rect 217794 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 218414 291134
rect 217794 286182 218414 290898
rect 218651 283932 218717 283933
rect 218651 283868 218652 283932
rect 218716 283868 218717 283932
rect 218651 283867 218717 283868
rect 217547 240140 217613 240141
rect 217547 240076 217548 240140
rect 217612 240076 217613 240140
rect 217547 240075 217613 240076
rect 217794 219454 218414 238182
rect 218654 236061 218714 283867
rect 219206 240141 219266 296107
rect 219942 292093 220002 341395
rect 221514 331174 222134 366618
rect 221514 330938 221546 331174
rect 221782 330938 221866 331174
rect 222102 330938 222134 331174
rect 221514 330854 222134 330938
rect 221514 330618 221546 330854
rect 221782 330618 221866 330854
rect 222102 330618 222134 330854
rect 220859 305692 220925 305693
rect 220859 305628 220860 305692
rect 220924 305628 220925 305692
rect 220859 305627 220925 305628
rect 219939 292092 220005 292093
rect 219939 292028 219940 292092
rect 220004 292028 220005 292092
rect 219939 292027 220005 292028
rect 219768 273454 220088 273486
rect 219768 273218 219810 273454
rect 220046 273218 220088 273454
rect 219768 273134 220088 273218
rect 219768 272898 219810 273134
rect 220046 272898 220088 273134
rect 219768 272866 220088 272898
rect 219203 240140 219269 240141
rect 219203 240076 219204 240140
rect 219268 240076 219269 240140
rect 219203 240075 219269 240076
rect 220862 240005 220922 305627
rect 221514 295174 222134 330618
rect 221514 294938 221546 295174
rect 221782 294938 221866 295174
rect 222102 294938 222134 295174
rect 221514 294854 222134 294938
rect 221514 294618 221546 294854
rect 221782 294618 221866 294854
rect 222102 294618 222134 294854
rect 221514 286182 222134 294618
rect 225234 370894 225854 375600
rect 225234 370658 225266 370894
rect 225502 370658 225586 370894
rect 225822 370658 225854 370894
rect 225234 370574 225854 370658
rect 225234 370338 225266 370574
rect 225502 370338 225586 370574
rect 225822 370338 225854 370574
rect 225234 334894 225854 370338
rect 225234 334658 225266 334894
rect 225502 334658 225586 334894
rect 225822 334658 225854 334894
rect 225234 334574 225854 334658
rect 225234 334338 225266 334574
rect 225502 334338 225586 334574
rect 225822 334338 225854 334574
rect 225234 298894 225854 334338
rect 228954 374614 229574 375600
rect 228954 374378 228986 374614
rect 229222 374378 229306 374614
rect 229542 374378 229574 374614
rect 228954 374294 229574 374378
rect 228954 374058 228986 374294
rect 229222 374058 229306 374294
rect 229542 374058 229574 374294
rect 228954 338614 229574 374058
rect 235794 345454 236414 375600
rect 235794 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 236414 345454
rect 235794 345134 236414 345218
rect 235794 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 236414 345134
rect 230427 342412 230493 342413
rect 230427 342348 230428 342412
rect 230492 342348 230493 342412
rect 230427 342347 230493 342348
rect 228954 338378 228986 338614
rect 229222 338378 229306 338614
rect 229542 338378 229574 338614
rect 228954 338294 229574 338378
rect 228954 338058 228986 338294
rect 229222 338058 229306 338294
rect 229542 338058 229574 338294
rect 227667 320924 227733 320925
rect 227667 320860 227668 320924
rect 227732 320860 227733 320924
rect 227667 320859 227733 320860
rect 225234 298658 225266 298894
rect 225502 298658 225586 298894
rect 225822 298658 225854 298894
rect 226195 298756 226261 298757
rect 226195 298692 226196 298756
rect 226260 298692 226261 298756
rect 226195 298691 226261 298692
rect 225234 298574 225854 298658
rect 225234 298338 225266 298574
rect 225502 298338 225586 298574
rect 225822 298338 225854 298574
rect 225234 286182 225854 298338
rect 223619 285836 223685 285837
rect 223619 285772 223620 285836
rect 223684 285772 223685 285836
rect 223619 285771 223685 285772
rect 222331 285700 222397 285701
rect 222331 285636 222332 285700
rect 222396 285636 222397 285700
rect 222331 285635 222397 285636
rect 220859 240004 220925 240005
rect 220859 239940 220860 240004
rect 220924 239940 220925 240004
rect 220859 239939 220925 239940
rect 222334 238645 222394 285635
rect 222331 238644 222397 238645
rect 222331 238580 222332 238644
rect 222396 238580 222397 238644
rect 222331 238579 222397 238580
rect 218651 236060 218717 236061
rect 218651 235996 218652 236060
rect 218716 235996 218717 236060
rect 218651 235995 218717 235996
rect 217794 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 218414 219454
rect 217794 219134 218414 219218
rect 217794 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 218414 219134
rect 216443 212668 216509 212669
rect 216443 212604 216444 212668
rect 216508 212604 216509 212668
rect 216443 212603 216509 212604
rect 214419 205596 214485 205597
rect 214419 205532 214420 205596
rect 214484 205532 214485 205596
rect 214419 205531 214485 205532
rect 217794 183454 218414 218898
rect 217794 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 218414 183454
rect 217794 183134 218414 183218
rect 217794 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 218414 183134
rect 217794 178000 218414 182898
rect 221514 223174 222134 238182
rect 223622 234701 223682 285771
rect 226198 240141 226258 298691
rect 227670 283933 227730 320859
rect 228954 302614 229574 338058
rect 228954 302378 228986 302614
rect 229222 302378 229306 302614
rect 229542 302378 229574 302614
rect 228954 302294 229574 302378
rect 228954 302058 228986 302294
rect 229222 302058 229306 302294
rect 229542 302058 229574 302294
rect 228954 286182 229574 302058
rect 227851 284476 227917 284477
rect 227851 284412 227852 284476
rect 227916 284412 227917 284476
rect 227851 284411 227917 284412
rect 226931 283932 226997 283933
rect 226931 283868 226932 283932
rect 226996 283868 226997 283932
rect 226931 283867 226997 283868
rect 227667 283932 227733 283933
rect 227667 283868 227668 283932
rect 227732 283868 227733 283932
rect 227667 283867 227733 283868
rect 226195 240140 226261 240141
rect 226195 240076 226196 240140
rect 226260 240076 226261 240140
rect 226195 240075 226261 240076
rect 226934 239461 226994 283867
rect 227854 277410 227914 284411
rect 228219 283932 228285 283933
rect 228219 283868 228220 283932
rect 228284 283868 228285 283932
rect 228219 283867 228285 283868
rect 229691 283932 229757 283933
rect 229691 283868 229692 283932
rect 229756 283868 229757 283932
rect 229691 283867 229757 283868
rect 227670 277350 227914 277410
rect 226931 239460 226997 239461
rect 226931 239396 226932 239460
rect 226996 239396 226997 239460
rect 226931 239395 226997 239396
rect 224171 236060 224237 236061
rect 224171 235996 224172 236060
rect 224236 235996 224237 236060
rect 224171 235995 224237 235996
rect 223619 234700 223685 234701
rect 223619 234636 223620 234700
rect 223684 234636 223685 234700
rect 223619 234635 223685 234636
rect 221514 222938 221546 223174
rect 221782 222938 221866 223174
rect 222102 222938 222134 223174
rect 221514 222854 222134 222938
rect 221514 222618 221546 222854
rect 221782 222618 221866 222854
rect 222102 222618 222134 222854
rect 221514 187174 222134 222618
rect 221514 186938 221546 187174
rect 221782 186938 221866 187174
rect 222102 186938 222134 187174
rect 221514 186854 222134 186938
rect 221514 186618 221546 186854
rect 221782 186618 221866 186854
rect 222102 186618 222134 186854
rect 221227 179620 221293 179621
rect 221227 179556 221228 179620
rect 221292 179556 221293 179620
rect 221227 179555 221293 179556
rect 210954 176378 210986 176614
rect 211222 176378 211306 176614
rect 211542 176378 211574 176614
rect 210954 176294 211574 176378
rect 210954 176058 210986 176294
rect 211222 176058 211306 176294
rect 211542 176058 211574 176294
rect 210954 140614 211574 176058
rect 221230 175949 221290 179555
rect 221514 178000 222134 186618
rect 224174 175949 224234 235995
rect 225234 226894 225854 238182
rect 227670 237421 227730 277350
rect 227667 237420 227733 237421
rect 227667 237356 227668 237420
rect 227732 237356 227733 237420
rect 227667 237355 227733 237356
rect 225234 226658 225266 226894
rect 225502 226658 225586 226894
rect 225822 226658 225854 226894
rect 225234 226574 225854 226658
rect 225234 226338 225266 226574
rect 225502 226338 225586 226574
rect 225822 226338 225854 226574
rect 225234 190894 225854 226338
rect 227667 205732 227733 205733
rect 227667 205668 227668 205732
rect 227732 205668 227733 205732
rect 227667 205667 227733 205668
rect 225234 190658 225266 190894
rect 225502 190658 225586 190894
rect 225822 190658 225854 190894
rect 225234 190574 225854 190658
rect 225234 190338 225266 190574
rect 225502 190338 225586 190574
rect 225822 190338 225854 190574
rect 225234 178000 225854 190338
rect 227670 175949 227730 205667
rect 228222 183565 228282 283867
rect 228954 230614 229574 238182
rect 228954 230378 228986 230614
rect 229222 230378 229306 230614
rect 229542 230378 229574 230614
rect 228954 230294 229574 230378
rect 228954 230058 228986 230294
rect 229222 230058 229306 230294
rect 229542 230058 229574 230294
rect 228954 194614 229574 230058
rect 228954 194378 228986 194614
rect 229222 194378 229306 194614
rect 229542 194378 229574 194614
rect 228954 194294 229574 194378
rect 228954 194058 228986 194294
rect 229222 194058 229306 194294
rect 229542 194058 229574 194294
rect 228219 183564 228285 183565
rect 228219 183500 228220 183564
rect 228284 183500 228285 183564
rect 228219 183499 228285 183500
rect 228771 183020 228837 183021
rect 228771 182956 228772 183020
rect 228836 182956 228837 183020
rect 228771 182955 228837 182956
rect 221227 175948 221293 175949
rect 221227 175884 221228 175948
rect 221292 175884 221293 175948
rect 221227 175883 221293 175884
rect 224171 175948 224237 175949
rect 224171 175884 224172 175948
rect 224236 175884 224237 175948
rect 224171 175883 224237 175884
rect 227667 175948 227733 175949
rect 227667 175884 227668 175948
rect 227732 175884 227733 175948
rect 227667 175883 227733 175884
rect 228774 174450 228834 182955
rect 228954 178000 229574 194058
rect 229323 176900 229389 176901
rect 229323 176836 229324 176900
rect 229388 176836 229389 176900
rect 229323 176835 229389 176836
rect 229139 174452 229205 174453
rect 229139 174450 229140 174452
rect 228774 174390 229140 174450
rect 229139 174388 229140 174390
rect 229204 174388 229205 174452
rect 229139 174387 229205 174388
rect 221207 165454 221527 165486
rect 221207 165218 221249 165454
rect 221485 165218 221527 165454
rect 221207 165134 221527 165218
rect 221207 164898 221249 165134
rect 221485 164898 221527 165134
rect 221207 164866 221527 164898
rect 224471 165454 224791 165486
rect 224471 165218 224513 165454
rect 224749 165218 224791 165454
rect 224471 165134 224791 165218
rect 224471 164898 224513 165134
rect 224749 164898 224791 165134
rect 224471 164866 224791 164898
rect 229326 161490 229386 176835
rect 229142 161430 229386 161490
rect 215891 151060 215957 151061
rect 215891 150996 215892 151060
rect 215956 150996 215957 151060
rect 215891 150995 215957 150996
rect 210954 140378 210986 140614
rect 211222 140378 211306 140614
rect 211542 140378 211574 140614
rect 210954 140294 211574 140378
rect 210954 140058 210986 140294
rect 211222 140058 211306 140294
rect 211542 140058 211574 140294
rect 210954 104614 211574 140058
rect 214419 123316 214485 123317
rect 214419 123252 214420 123316
rect 214484 123252 214485 123316
rect 214419 123251 214485 123252
rect 210954 104378 210986 104614
rect 211222 104378 211306 104614
rect 211542 104378 211574 104614
rect 210954 104294 211574 104378
rect 210954 104058 210986 104294
rect 211222 104058 211306 104294
rect 211542 104058 211574 104294
rect 210954 68614 211574 104058
rect 214422 94485 214482 123251
rect 214419 94484 214485 94485
rect 214419 94420 214420 94484
rect 214484 94420 214485 94484
rect 214419 94419 214485 94420
rect 215894 86189 215954 150995
rect 229142 150109 229202 161430
rect 229139 150108 229205 150109
rect 229139 150044 229140 150108
rect 229204 150044 229205 150108
rect 229139 150043 229205 150044
rect 219575 147454 219895 147486
rect 219575 147218 219617 147454
rect 219853 147218 219895 147454
rect 219575 147134 219895 147218
rect 219575 146898 219617 147134
rect 219853 146898 219895 147134
rect 219575 146866 219895 146898
rect 222839 147454 223159 147486
rect 222839 147218 222881 147454
rect 223117 147218 223159 147454
rect 222839 147134 223159 147218
rect 222839 146898 222881 147134
rect 223117 146898 223159 147134
rect 222839 146866 223159 146898
rect 226103 147454 226423 147486
rect 226103 147218 226145 147454
rect 226381 147218 226423 147454
rect 226103 147134 226423 147218
rect 226103 146898 226145 147134
rect 226381 146898 226423 147134
rect 226103 146866 226423 146898
rect 229694 137325 229754 283867
rect 230430 240141 230490 342347
rect 235794 309454 236414 344898
rect 239514 349174 240134 375600
rect 239514 348938 239546 349174
rect 239782 348938 239866 349174
rect 240102 348938 240134 349174
rect 239514 348854 240134 348938
rect 239514 348618 239546 348854
rect 239782 348618 239866 348854
rect 240102 348618 240134 348854
rect 237419 325004 237485 325005
rect 237419 324940 237420 325004
rect 237484 324940 237485 325004
rect 237419 324939 237485 324940
rect 235794 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 236414 309454
rect 235794 309134 236414 309218
rect 235794 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 236414 309134
rect 231899 306508 231965 306509
rect 231899 306444 231900 306508
rect 231964 306444 231965 306508
rect 231899 306443 231965 306444
rect 231715 283932 231781 283933
rect 231715 283868 231716 283932
rect 231780 283868 231781 283932
rect 231715 283867 231781 283868
rect 230427 240140 230493 240141
rect 230427 240076 230428 240140
rect 230492 240076 230493 240140
rect 230427 240075 230493 240076
rect 230427 210492 230493 210493
rect 230427 210428 230428 210492
rect 230492 210428 230493 210492
rect 230427 210427 230493 210428
rect 230430 156229 230490 210427
rect 230427 156228 230493 156229
rect 230427 156164 230428 156228
rect 230492 156164 230493 156228
rect 230427 156163 230493 156164
rect 231718 147250 231778 283867
rect 231902 240141 231962 306443
rect 233187 287196 233253 287197
rect 233187 287132 233188 287196
rect 233252 287132 233253 287196
rect 233187 287131 233253 287132
rect 232451 285972 232517 285973
rect 232451 285908 232452 285972
rect 232516 285908 232517 285972
rect 232451 285907 232517 285908
rect 231899 240140 231965 240141
rect 231899 240076 231900 240140
rect 231964 240076 231965 240140
rect 231899 240075 231965 240076
rect 231899 179076 231965 179077
rect 231899 179012 231900 179076
rect 231964 179012 231965 179076
rect 231899 179011 231965 179012
rect 231902 151605 231962 179011
rect 232454 178125 232514 285907
rect 232451 178124 232517 178125
rect 232451 178060 232452 178124
rect 232516 178060 232517 178124
rect 232451 178059 232517 178060
rect 232083 176764 232149 176765
rect 232083 176700 232084 176764
rect 232148 176700 232149 176764
rect 232083 176699 232149 176700
rect 231899 151604 231965 151605
rect 231899 151540 231900 151604
rect 231964 151540 231965 151604
rect 231899 151539 231965 151540
rect 232086 150653 232146 176699
rect 233190 157181 233250 287131
rect 235794 286182 236414 308898
rect 236499 283932 236565 283933
rect 236499 283868 236500 283932
rect 236564 283868 236565 283932
rect 236499 283867 236565 283868
rect 235128 255454 235448 255486
rect 235128 255218 235170 255454
rect 235406 255218 235448 255454
rect 235128 255134 235448 255218
rect 235128 254898 235170 255134
rect 235406 254898 235448 255134
rect 235128 254866 235448 254898
rect 235794 237454 236414 238182
rect 235794 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 236414 237454
rect 235794 237134 236414 237218
rect 235794 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 236414 237134
rect 234659 231708 234725 231709
rect 234659 231644 234660 231708
rect 234724 231644 234725 231708
rect 234659 231643 234725 231644
rect 233371 208452 233437 208453
rect 233371 208388 233372 208452
rect 233436 208388 233437 208452
rect 233371 208387 233437 208388
rect 233374 160581 233434 208387
rect 233371 160580 233437 160581
rect 233371 160516 233372 160580
rect 233436 160516 233437 160580
rect 233371 160515 233437 160516
rect 233739 160172 233805 160173
rect 233739 160108 233740 160172
rect 233804 160108 233805 160172
rect 233739 160107 233805 160108
rect 233187 157180 233253 157181
rect 233187 157116 233188 157180
rect 233252 157116 233253 157180
rect 233187 157115 233253 157116
rect 233187 151060 233253 151061
rect 233187 150996 233188 151060
rect 233252 150996 233253 151060
rect 233187 150995 233253 150996
rect 232083 150652 232149 150653
rect 232083 150588 232084 150652
rect 232148 150588 232149 150652
rect 232083 150587 232149 150588
rect 231718 147190 231962 147250
rect 231163 146980 231229 146981
rect 231163 146916 231164 146980
rect 231228 146916 231229 146980
rect 231163 146915 231229 146916
rect 230979 142764 231045 142765
rect 230979 142700 230980 142764
rect 231044 142700 231045 142764
rect 230979 142699 231045 142700
rect 229691 137324 229757 137325
rect 229691 137260 229692 137324
rect 229756 137260 229757 137324
rect 229691 137259 229757 137260
rect 229875 137188 229941 137189
rect 229875 137124 229876 137188
rect 229940 137124 229941 137188
rect 229875 137123 229941 137124
rect 221207 129454 221527 129486
rect 221207 129218 221249 129454
rect 221485 129218 221527 129454
rect 221207 129134 221527 129218
rect 221207 128898 221249 129134
rect 221485 128898 221527 129134
rect 221207 128866 221527 128898
rect 224471 129454 224791 129486
rect 224471 129218 224513 129454
rect 224749 129218 224791 129454
rect 224471 129134 224791 129218
rect 224471 128898 224513 129134
rect 224749 128898 224791 129134
rect 224471 128866 224791 128898
rect 219575 111454 219895 111486
rect 219575 111218 219617 111454
rect 219853 111218 219895 111454
rect 219575 111134 219895 111218
rect 219575 110898 219617 111134
rect 219853 110898 219895 111134
rect 219575 110866 219895 110898
rect 222839 111454 223159 111486
rect 222839 111218 222881 111454
rect 223117 111218 223159 111454
rect 222839 111134 223159 111218
rect 222839 110898 222881 111134
rect 223117 110898 223159 111134
rect 222839 110866 223159 110898
rect 226103 111454 226423 111486
rect 226103 111218 226145 111454
rect 226381 111218 226423 111454
rect 226103 111134 226423 111218
rect 226103 110898 226145 111134
rect 226381 110898 226423 111134
rect 226103 110866 226423 110898
rect 224726 97550 225154 97610
rect 215891 86188 215957 86189
rect 215891 86124 215892 86188
rect 215956 86124 215957 86188
rect 215891 86123 215957 86124
rect 210954 68378 210986 68614
rect 211222 68378 211306 68614
rect 211542 68378 211574 68614
rect 210954 68294 211574 68378
rect 210954 68058 210986 68294
rect 211222 68058 211306 68294
rect 211542 68058 211574 68294
rect 210954 32614 211574 68058
rect 210954 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 211574 32614
rect 210954 32294 211574 32378
rect 210954 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 211574 32294
rect 192954 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 193574 -6106
rect 192954 -6426 193574 -6342
rect 192954 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 193574 -6426
rect 192954 -7654 193574 -6662
rect 210954 -7066 211574 32058
rect 217794 75454 218414 94000
rect 217794 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 218414 75454
rect 217794 75134 218414 75218
rect 217794 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 218414 75134
rect 217794 39454 218414 74898
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -1894 218414 -902
rect 221514 79174 222134 94000
rect 224726 91085 224786 97550
rect 225094 95981 225154 97550
rect 229139 97068 229205 97069
rect 229139 97004 229140 97068
rect 229204 97004 229205 97068
rect 229139 97003 229205 97004
rect 229142 96930 229202 97003
rect 228958 96870 229202 96930
rect 225091 95980 225157 95981
rect 225091 95916 225092 95980
rect 225156 95916 225157 95980
rect 225091 95915 225157 95916
rect 226379 95980 226445 95981
rect 226379 95916 226380 95980
rect 226444 95916 226445 95980
rect 226379 95915 226445 95916
rect 226931 95980 226997 95981
rect 226931 95916 226932 95980
rect 226996 95916 226997 95980
rect 226931 95915 226997 95916
rect 224723 91084 224789 91085
rect 224723 91020 224724 91084
rect 224788 91020 224789 91084
rect 224723 91019 224789 91020
rect 221514 78938 221546 79174
rect 221782 78938 221866 79174
rect 222102 78938 222134 79174
rect 221514 78854 222134 78938
rect 221514 78618 221546 78854
rect 221782 78618 221866 78854
rect 222102 78618 222134 78854
rect 221514 43174 222134 78618
rect 221514 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 222134 43174
rect 221514 42854 222134 42938
rect 221514 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 222134 42854
rect 221514 7174 222134 42618
rect 221514 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 222134 7174
rect 221514 6854 222134 6938
rect 221514 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 222134 6854
rect 221514 -2266 222134 6618
rect 221514 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 222134 -2266
rect 221514 -2586 222134 -2502
rect 221514 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 222134 -2586
rect 221514 -3814 222134 -2822
rect 225234 82894 225854 94000
rect 225234 82658 225266 82894
rect 225502 82658 225586 82894
rect 225822 82658 225854 82894
rect 225234 82574 225854 82658
rect 225234 82338 225266 82574
rect 225502 82338 225586 82574
rect 225822 82338 225854 82574
rect 225234 46894 225854 82338
rect 225234 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 225854 46894
rect 225234 46574 225854 46658
rect 225234 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 225854 46574
rect 225234 10894 225854 46338
rect 226382 38045 226442 95915
rect 226379 38044 226445 38045
rect 226379 37980 226380 38044
rect 226444 37980 226445 38044
rect 226379 37979 226445 37980
rect 226934 21317 226994 95915
rect 228958 94210 229018 96870
rect 228774 94150 229018 94210
rect 228774 93669 228834 94150
rect 228771 93668 228837 93669
rect 228771 93604 228772 93668
rect 228836 93604 228837 93668
rect 228771 93603 228837 93604
rect 228774 89730 228834 93603
rect 227670 89670 228834 89730
rect 226931 21316 226997 21317
rect 226931 21252 226932 21316
rect 226996 21252 226997 21316
rect 226931 21251 226997 21252
rect 225234 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 225854 10894
rect 225234 10574 225854 10658
rect 225234 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 225854 10574
rect 225234 -4186 225854 10338
rect 227670 4861 227730 89670
rect 228954 86614 229574 94000
rect 228954 86378 228986 86614
rect 229222 86378 229306 86614
rect 229542 86378 229574 86614
rect 228954 86294 229574 86378
rect 228954 86058 228986 86294
rect 229222 86058 229306 86294
rect 229542 86058 229574 86294
rect 228954 50614 229574 86058
rect 229878 78029 229938 137123
rect 230427 133652 230493 133653
rect 230427 133588 230428 133652
rect 230492 133588 230493 133652
rect 230427 133587 230493 133588
rect 230430 94757 230490 133587
rect 230982 123181 231042 142699
rect 231166 134469 231226 146915
rect 231902 139773 231962 147190
rect 233190 142493 233250 150995
rect 233742 149157 233802 160107
rect 233739 149156 233805 149157
rect 233739 149092 233740 149156
rect 233804 149092 233805 149156
rect 233739 149091 233805 149092
rect 234107 148068 234173 148069
rect 234107 148004 234108 148068
rect 234172 148004 234173 148068
rect 234107 148003 234173 148004
rect 233187 142492 233253 142493
rect 233187 142428 233188 142492
rect 233252 142428 233253 142492
rect 233187 142427 233253 142428
rect 231899 139772 231965 139773
rect 231899 139708 231900 139772
rect 231964 139708 231965 139772
rect 231899 139707 231965 139708
rect 231163 134468 231229 134469
rect 231163 134404 231164 134468
rect 231228 134404 231229 134468
rect 231163 134403 231229 134404
rect 232451 129028 232517 129029
rect 232451 128964 232452 129028
rect 232516 128964 232517 129028
rect 232451 128963 232517 128964
rect 230979 123180 231045 123181
rect 230979 123116 230980 123180
rect 231044 123116 231045 123180
rect 230979 123115 231045 123116
rect 230427 94756 230493 94757
rect 230427 94692 230428 94756
rect 230492 94692 230493 94756
rect 230427 94691 230493 94692
rect 229875 78028 229941 78029
rect 229875 77964 229876 78028
rect 229940 77964 229941 78028
rect 229875 77963 229941 77964
rect 228954 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 229574 50614
rect 228954 50294 229574 50378
rect 228954 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 229574 50294
rect 228954 14614 229574 50058
rect 232454 42125 232514 128963
rect 233739 113524 233805 113525
rect 233739 113460 233740 113524
rect 233804 113460 233805 113524
rect 233739 113459 233805 113460
rect 233742 54501 233802 113459
rect 234110 106181 234170 148003
rect 234662 139229 234722 231643
rect 235794 201454 236414 236898
rect 235794 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 236414 201454
rect 235794 201134 236414 201218
rect 235794 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 236414 201134
rect 235794 165454 236414 200898
rect 236502 168605 236562 283867
rect 237422 240141 237482 324939
rect 239514 313174 240134 348618
rect 239514 312938 239546 313174
rect 239782 312938 239866 313174
rect 240102 312938 240134 313174
rect 239514 312854 240134 312938
rect 239514 312618 239546 312854
rect 239782 312618 239866 312854
rect 240102 312618 240134 312854
rect 238523 287740 238589 287741
rect 238523 287676 238524 287740
rect 238588 287676 238589 287740
rect 238523 287675 238589 287676
rect 237419 240140 237485 240141
rect 237419 240076 237420 240140
rect 237484 240076 237485 240140
rect 237419 240075 237485 240076
rect 237422 214709 237482 240075
rect 237419 214708 237485 214709
rect 237419 214644 237420 214708
rect 237484 214644 237485 214708
rect 237419 214643 237485 214644
rect 237419 188596 237485 188597
rect 237419 188532 237420 188596
rect 237484 188532 237485 188596
rect 237419 188531 237485 188532
rect 236499 168604 236565 168605
rect 236499 168540 236500 168604
rect 236564 168540 236565 168604
rect 236499 168539 236565 168540
rect 236683 168468 236749 168469
rect 236683 168404 236684 168468
rect 236748 168404 236749 168468
rect 236683 168403 236749 168404
rect 235794 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 236414 165454
rect 235794 165134 236414 165218
rect 235794 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 236414 165134
rect 234659 139228 234725 139229
rect 234659 139164 234660 139228
rect 234724 139164 234725 139228
rect 234659 139163 234725 139164
rect 235794 129454 236414 164898
rect 236686 160173 236746 168403
rect 236683 160172 236749 160173
rect 236683 160108 236684 160172
rect 236748 160108 236749 160172
rect 236683 160107 236749 160108
rect 237422 138821 237482 188531
rect 237603 178940 237669 178941
rect 237603 178876 237604 178940
rect 237668 178876 237669 178940
rect 237603 178875 237669 178876
rect 237606 165749 237666 178875
rect 237603 165748 237669 165749
rect 237603 165684 237604 165748
rect 237668 165684 237669 165748
rect 237603 165683 237669 165684
rect 238526 142490 238586 287675
rect 239514 286182 240134 312618
rect 243234 352894 243854 375600
rect 243234 352658 243266 352894
rect 243502 352658 243586 352894
rect 243822 352658 243854 352894
rect 243234 352574 243854 352658
rect 243234 352338 243266 352574
rect 243502 352338 243586 352574
rect 243822 352338 243854 352574
rect 243234 316894 243854 352338
rect 246954 356614 247574 375600
rect 253059 374100 253125 374101
rect 253059 374036 253060 374100
rect 253124 374036 253125 374100
rect 253059 374035 253125 374036
rect 246954 356378 246986 356614
rect 247222 356378 247306 356614
rect 247542 356378 247574 356614
rect 246954 356294 247574 356378
rect 246954 356058 246986 356294
rect 247222 356058 247306 356294
rect 247542 356058 247574 356294
rect 244779 321740 244845 321741
rect 244779 321676 244780 321740
rect 244844 321676 244845 321740
rect 244779 321675 244845 321676
rect 243234 316658 243266 316894
rect 243502 316658 243586 316894
rect 243822 316658 243854 316894
rect 243234 316574 243854 316658
rect 243234 316338 243266 316574
rect 243502 316338 243586 316574
rect 243822 316338 243854 316574
rect 240731 311948 240797 311949
rect 240731 311884 240732 311948
rect 240796 311884 240797 311948
rect 240731 311883 240797 311884
rect 239514 205174 240134 238182
rect 240734 237557 240794 311883
rect 242939 296036 243005 296037
rect 242939 295972 242940 296036
rect 243004 295972 243005 296036
rect 242939 295971 243005 295972
rect 242942 267750 243002 295971
rect 243234 286182 243854 316338
rect 244227 300932 244293 300933
rect 244227 300868 244228 300932
rect 244292 300868 244293 300932
rect 244227 300867 244293 300868
rect 243491 284476 243557 284477
rect 243491 284412 243492 284476
rect 243556 284412 243557 284476
rect 243491 284411 243557 284412
rect 243494 280805 243554 284411
rect 243491 280804 243557 280805
rect 243491 280740 243492 280804
rect 243556 280740 243557 280804
rect 243491 280739 243557 280740
rect 244230 269109 244290 300867
rect 244782 280261 244842 321675
rect 246954 320614 247574 356058
rect 251219 355468 251285 355469
rect 251219 355404 251220 355468
rect 251284 355404 251285 355468
rect 251219 355403 251285 355404
rect 248459 345540 248525 345541
rect 248459 345476 248460 345540
rect 248524 345476 248525 345540
rect 248459 345475 248525 345476
rect 246954 320378 246986 320614
rect 247222 320378 247306 320614
rect 247542 320378 247574 320614
rect 246954 320294 247574 320378
rect 246954 320058 246986 320294
rect 247222 320058 247306 320294
rect 247542 320058 247574 320294
rect 246954 284614 247574 320058
rect 246954 284378 246986 284614
rect 247222 284378 247306 284614
rect 247542 284378 247574 284614
rect 246954 284294 247574 284378
rect 246954 284058 246986 284294
rect 247222 284058 247306 284294
rect 247542 284058 247574 284294
rect 244779 280260 244845 280261
rect 244779 280196 244780 280260
rect 244844 280196 244845 280260
rect 244779 280195 244845 280196
rect 244227 269108 244293 269109
rect 244227 269044 244228 269108
rect 244292 269044 244293 269108
rect 244227 269043 244293 269044
rect 242942 267690 243554 267750
rect 243494 259861 243554 267690
rect 244411 265844 244477 265845
rect 244411 265780 244412 265844
rect 244476 265780 244477 265844
rect 244411 265779 244477 265780
rect 244227 261356 244293 261357
rect 244227 261292 244228 261356
rect 244292 261292 244293 261356
rect 244227 261291 244293 261292
rect 243491 259860 243557 259861
rect 243491 259796 243492 259860
rect 243556 259796 243557 259860
rect 243491 259795 243557 259796
rect 244230 259450 244290 261291
rect 244046 259390 244290 259450
rect 243491 241364 243557 241365
rect 243491 241300 243492 241364
rect 243556 241300 243557 241364
rect 243491 241299 243557 241300
rect 243494 238770 243554 241299
rect 242942 238710 243554 238770
rect 240731 237556 240797 237557
rect 240731 237492 240732 237556
rect 240796 237492 240797 237556
rect 240731 237491 240797 237492
rect 241651 237420 241717 237421
rect 241651 237356 241652 237420
rect 241716 237356 241717 237420
rect 241651 237355 241717 237356
rect 239514 204938 239546 205174
rect 239782 204938 239866 205174
rect 240102 204938 240134 205174
rect 239514 204854 240134 204938
rect 239514 204618 239546 204854
rect 239782 204618 239866 204854
rect 240102 204618 240134 204854
rect 239514 169174 240134 204618
rect 240363 193900 240429 193901
rect 240363 193836 240364 193900
rect 240428 193836 240429 193900
rect 240363 193835 240429 193836
rect 239514 168938 239546 169174
rect 239782 168938 239866 169174
rect 240102 168938 240134 169174
rect 239514 168854 240134 168938
rect 239514 168618 239546 168854
rect 239782 168618 239866 168854
rect 240102 168618 240134 168854
rect 238526 142430 238770 142490
rect 238710 142085 238770 142430
rect 238707 142084 238773 142085
rect 238707 142020 238708 142084
rect 238772 142020 238773 142084
rect 238707 142019 238773 142020
rect 237419 138820 237485 138821
rect 237419 138756 237420 138820
rect 237484 138756 237485 138820
rect 237419 138755 237485 138756
rect 236499 137324 236565 137325
rect 236499 137260 236500 137324
rect 236564 137260 236565 137324
rect 236499 137259 236565 137260
rect 235794 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 236414 129454
rect 235794 129134 236414 129218
rect 235794 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 236414 129134
rect 234107 106180 234173 106181
rect 234107 106116 234108 106180
rect 234172 106116 234173 106180
rect 234107 106115 234173 106116
rect 235794 93454 236414 128898
rect 235794 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 236414 93454
rect 235794 93134 236414 93218
rect 235794 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 236414 93134
rect 235794 57454 236414 92898
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 233739 54500 233805 54501
rect 233739 54436 233740 54500
rect 233804 54436 233805 54500
rect 233739 54435 233805 54436
rect 232451 42124 232517 42125
rect 232451 42060 232452 42124
rect 232516 42060 232517 42124
rect 232451 42059 232517 42060
rect 228954 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 229574 14614
rect 228954 14294 229574 14378
rect 228954 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 229574 14294
rect 227667 4860 227733 4861
rect 227667 4796 227668 4860
rect 227732 4796 227733 4860
rect 227667 4795 227733 4796
rect 225234 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 225854 -4186
rect 225234 -4506 225854 -4422
rect 225234 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 225854 -4506
rect 225234 -5734 225854 -4742
rect 210954 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 211574 -7066
rect 210954 -7386 211574 -7302
rect 210954 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 211574 -7386
rect 210954 -7654 211574 -7622
rect 228954 -6106 229574 14058
rect 235794 21454 236414 56898
rect 236502 24173 236562 137259
rect 239514 133174 240134 168618
rect 240366 161533 240426 193835
rect 240363 161532 240429 161533
rect 240363 161468 240364 161532
rect 240428 161468 240429 161532
rect 240363 161467 240429 161468
rect 240731 160172 240797 160173
rect 240731 160108 240732 160172
rect 240796 160108 240797 160172
rect 240731 160107 240797 160108
rect 239514 132938 239546 133174
rect 239782 132938 239866 133174
rect 240102 132938 240134 133174
rect 239514 132854 240134 132938
rect 239514 132618 239546 132854
rect 239782 132618 239866 132854
rect 240102 132618 240134 132854
rect 237971 102916 238037 102917
rect 237971 102852 237972 102916
rect 238036 102852 238037 102916
rect 237971 102851 238037 102852
rect 237974 79661 238034 102851
rect 239514 97174 240134 132618
rect 240734 120053 240794 160107
rect 241654 151061 241714 237355
rect 242942 234565 243002 238710
rect 244046 238645 244106 259390
rect 244414 258090 244474 265779
rect 245699 263124 245765 263125
rect 245699 263060 245700 263124
rect 245764 263060 245765 263124
rect 245699 263059 245765 263060
rect 244230 258030 244474 258090
rect 244043 238644 244109 238645
rect 244043 238580 244044 238644
rect 244108 238580 244109 238644
rect 244043 238579 244109 238580
rect 242939 234564 243005 234565
rect 242939 234500 242940 234564
rect 243004 234500 243005 234564
rect 242939 234499 243005 234500
rect 242755 226948 242821 226949
rect 242755 226884 242756 226948
rect 242820 226884 242821 226948
rect 242755 226883 242821 226884
rect 242758 224909 242818 226883
rect 242755 224908 242821 224909
rect 242755 224844 242756 224908
rect 242820 224844 242821 224908
rect 242755 224843 242821 224844
rect 243234 208894 243854 238182
rect 243234 208658 243266 208894
rect 243502 208658 243586 208894
rect 243822 208658 243854 208894
rect 243234 208574 243854 208658
rect 243234 208338 243266 208574
rect 243502 208338 243586 208574
rect 243822 208338 243854 208574
rect 242939 182340 243005 182341
rect 242939 182276 242940 182340
rect 243004 182276 243005 182340
rect 242939 182275 243005 182276
rect 242942 162077 243002 182275
rect 243234 172894 243854 208338
rect 243234 172658 243266 172894
rect 243502 172658 243586 172894
rect 243822 172658 243854 172894
rect 243234 172574 243854 172658
rect 243234 172338 243266 172574
rect 243502 172338 243586 172574
rect 243822 172338 243854 172574
rect 242939 162076 243005 162077
rect 242939 162012 242940 162076
rect 243004 162012 243005 162076
rect 242939 162011 243005 162012
rect 241651 151060 241717 151061
rect 241651 150996 241652 151060
rect 241716 150996 241717 151060
rect 241651 150995 241717 150996
rect 243234 136894 243854 172338
rect 244230 153781 244290 258030
rect 244779 248164 244845 248165
rect 244779 248100 244780 248164
rect 244844 248100 244845 248164
rect 244779 248099 244845 248100
rect 244411 225316 244477 225317
rect 244411 225252 244412 225316
rect 244476 225252 244477 225316
rect 244411 225251 244477 225252
rect 244414 167653 244474 225251
rect 244782 225181 244842 248099
rect 244779 225180 244845 225181
rect 244779 225116 244780 225180
rect 244844 225116 244845 225180
rect 244779 225115 244845 225116
rect 244411 167652 244477 167653
rect 244411 167588 244412 167652
rect 244476 167588 244477 167652
rect 244411 167587 244477 167588
rect 244227 153780 244293 153781
rect 244227 153716 244228 153780
rect 244292 153716 244293 153780
rect 244227 153715 244293 153716
rect 243234 136658 243266 136894
rect 243502 136658 243586 136894
rect 243822 136658 243854 136894
rect 243234 136574 243854 136658
rect 243234 136338 243266 136574
rect 243502 136338 243586 136574
rect 243822 136338 243854 136574
rect 242755 130252 242821 130253
rect 242755 130188 242756 130252
rect 242820 130188 242821 130252
rect 242755 130187 242821 130188
rect 240731 120052 240797 120053
rect 240731 119988 240732 120052
rect 240796 119988 240797 120052
rect 240731 119987 240797 119988
rect 239514 96938 239546 97174
rect 239782 96938 239866 97174
rect 240102 96938 240134 97174
rect 239514 96854 240134 96938
rect 239514 96618 239546 96854
rect 239782 96618 239866 96854
rect 240102 96618 240134 96854
rect 237971 79660 238037 79661
rect 237971 79596 237972 79660
rect 238036 79596 238037 79660
rect 237971 79595 238037 79596
rect 239514 61174 240134 96618
rect 242758 95709 242818 130187
rect 243234 100894 243854 136338
rect 244043 127396 244109 127397
rect 244043 127332 244044 127396
rect 244108 127332 244109 127396
rect 244043 127331 244109 127332
rect 243234 100658 243266 100894
rect 243502 100658 243586 100894
rect 243822 100658 243854 100894
rect 243234 100574 243854 100658
rect 243234 100338 243266 100574
rect 243502 100338 243586 100574
rect 243822 100338 243854 100574
rect 242755 95708 242821 95709
rect 242755 95644 242756 95708
rect 242820 95644 242821 95708
rect 242755 95643 242821 95644
rect 239514 60938 239546 61174
rect 239782 60938 239866 61174
rect 240102 60938 240134 61174
rect 239514 60854 240134 60938
rect 239514 60618 239546 60854
rect 239782 60618 239866 60854
rect 240102 60618 240134 60854
rect 239514 25174 240134 60618
rect 239514 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 240134 25174
rect 239514 24854 240134 24938
rect 239514 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 240134 24854
rect 236499 24172 236565 24173
rect 236499 24108 236500 24172
rect 236564 24108 236565 24172
rect 236499 24107 236565 24108
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -1306 236414 20898
rect 235794 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 236414 -1306
rect 235794 -1626 236414 -1542
rect 235794 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 236414 -1626
rect 235794 -1894 236414 -1862
rect 239514 -3226 240134 24618
rect 239514 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 240134 -3226
rect 239514 -3546 240134 -3462
rect 239514 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 240134 -3546
rect 239514 -3814 240134 -3782
rect 243234 64894 243854 100338
rect 243234 64658 243266 64894
rect 243502 64658 243586 64894
rect 243822 64658 243854 64894
rect 243234 64574 243854 64658
rect 243234 64338 243266 64574
rect 243502 64338 243586 64574
rect 243822 64338 243854 64574
rect 243234 28894 243854 64338
rect 243234 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 243854 28894
rect 243234 28574 243854 28658
rect 243234 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 243854 28574
rect 243234 -5146 243854 28338
rect 244046 25533 244106 127331
rect 244779 124676 244845 124677
rect 244779 124612 244780 124676
rect 244844 124612 244845 124676
rect 244779 124611 244845 124612
rect 244782 80885 244842 124611
rect 245702 89181 245762 263059
rect 246954 248614 247574 284058
rect 246954 248378 246986 248614
rect 247222 248378 247306 248614
rect 247542 248378 247574 248614
rect 246954 248294 247574 248378
rect 246954 248058 246986 248294
rect 247222 248058 247306 248294
rect 247542 248058 247574 248294
rect 246954 212614 247574 248058
rect 248462 213757 248522 345475
rect 249747 323780 249813 323781
rect 249747 323716 249748 323780
rect 249812 323716 249813 323780
rect 249747 323715 249813 323716
rect 248643 302564 248709 302565
rect 248643 302500 248644 302564
rect 248708 302500 248709 302564
rect 248643 302499 248709 302500
rect 248646 279445 248706 302499
rect 248643 279444 248709 279445
rect 248643 279380 248644 279444
rect 248708 279380 248709 279444
rect 248643 279379 248709 279380
rect 248643 222052 248709 222053
rect 248643 221988 248644 222052
rect 248708 221988 248709 222052
rect 248643 221987 248709 221988
rect 248459 213756 248525 213757
rect 248459 213692 248460 213756
rect 248524 213692 248525 213756
rect 248459 213691 248525 213692
rect 246954 212378 246986 212614
rect 247222 212378 247306 212614
rect 247542 212378 247574 212614
rect 246954 212294 247574 212378
rect 246954 212058 246986 212294
rect 247222 212058 247306 212294
rect 247542 212058 247574 212294
rect 246954 176614 247574 212058
rect 246954 176378 246986 176614
rect 247222 176378 247306 176614
rect 247542 176378 247574 176614
rect 246954 176294 247574 176378
rect 246954 176058 246986 176294
rect 247222 176058 247306 176294
rect 247542 176058 247574 176294
rect 246954 140614 247574 176058
rect 248646 141133 248706 221987
rect 248643 141132 248709 141133
rect 248643 141068 248644 141132
rect 248708 141068 248709 141132
rect 248643 141067 248709 141068
rect 246954 140378 246986 140614
rect 247222 140378 247306 140614
rect 247542 140378 247574 140614
rect 246954 140294 247574 140378
rect 246954 140058 246986 140294
rect 247222 140058 247306 140294
rect 247542 140058 247574 140294
rect 246954 104614 247574 140058
rect 249011 133924 249077 133925
rect 249011 133860 249012 133924
rect 249076 133860 249077 133924
rect 249011 133859 249077 133860
rect 246954 104378 246986 104614
rect 247222 104378 247306 104614
rect 247542 104378 247574 104614
rect 246954 104294 247574 104378
rect 246954 104058 246986 104294
rect 247222 104058 247306 104294
rect 247542 104058 247574 104294
rect 245699 89180 245765 89181
rect 245699 89116 245700 89180
rect 245764 89116 245765 89180
rect 245699 89115 245765 89116
rect 244779 80884 244845 80885
rect 244779 80820 244780 80884
rect 244844 80820 244845 80884
rect 244779 80819 244845 80820
rect 246954 68614 247574 104058
rect 246954 68378 246986 68614
rect 247222 68378 247306 68614
rect 247542 68378 247574 68614
rect 246954 68294 247574 68378
rect 246954 68058 246986 68294
rect 247222 68058 247306 68294
rect 247542 68058 247574 68294
rect 246954 32614 247574 68058
rect 249014 61437 249074 133859
rect 249011 61436 249077 61437
rect 249011 61372 249012 61436
rect 249076 61372 249077 61436
rect 249011 61371 249077 61372
rect 249750 50965 249810 323715
rect 251222 252517 251282 355403
rect 251219 252516 251285 252517
rect 251219 252452 251220 252516
rect 251284 252452 251285 252516
rect 251219 252451 251285 252452
rect 252323 215252 252389 215253
rect 252323 215188 252324 215252
rect 252388 215188 252389 215252
rect 252323 215187 252389 215188
rect 252326 53410 252386 215187
rect 253062 92309 253122 374035
rect 253794 363454 254414 375600
rect 253794 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 254414 363454
rect 253794 363134 254414 363218
rect 253794 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 254414 363134
rect 253794 327454 254414 362898
rect 253794 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 254414 327454
rect 253794 327134 254414 327218
rect 253794 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 254414 327134
rect 253794 291454 254414 326898
rect 257514 367174 258134 375600
rect 257514 366938 257546 367174
rect 257782 366938 257866 367174
rect 258102 366938 258134 367174
rect 257514 366854 258134 366938
rect 257514 366618 257546 366854
rect 257782 366618 257866 366854
rect 258102 366618 258134 366854
rect 257514 331174 258134 366618
rect 257514 330938 257546 331174
rect 257782 330938 257866 331174
rect 258102 330938 258134 331174
rect 257514 330854 258134 330938
rect 257514 330618 257546 330854
rect 257782 330618 257866 330854
rect 258102 330618 258134 330854
rect 255267 325004 255333 325005
rect 255267 324940 255268 325004
rect 255332 324940 255333 325004
rect 255267 324939 255333 324940
rect 253794 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 254414 291454
rect 253794 291134 254414 291218
rect 253794 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 254414 291134
rect 253794 255454 254414 290898
rect 253794 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 254414 255454
rect 253794 255134 254414 255218
rect 253794 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 254414 255134
rect 253794 219454 254414 254898
rect 253794 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 254414 219454
rect 253794 219134 254414 219218
rect 253794 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 254414 219134
rect 253794 183454 254414 218898
rect 255270 215253 255330 324939
rect 257514 295174 258134 330618
rect 261234 370894 261854 375600
rect 261234 370658 261266 370894
rect 261502 370658 261586 370894
rect 261822 370658 261854 370894
rect 261234 370574 261854 370658
rect 261234 370338 261266 370574
rect 261502 370338 261586 370574
rect 261822 370338 261854 370574
rect 261234 334894 261854 370338
rect 261234 334658 261266 334894
rect 261502 334658 261586 334894
rect 261822 334658 261854 334894
rect 261234 334574 261854 334658
rect 261234 334338 261266 334574
rect 261502 334338 261586 334574
rect 261822 334338 261854 334574
rect 259499 328540 259565 328541
rect 259499 328476 259500 328540
rect 259564 328476 259565 328540
rect 259499 328475 259565 328476
rect 257514 294938 257546 295174
rect 257782 294938 257866 295174
rect 258102 294938 258134 295174
rect 257514 294854 258134 294938
rect 257514 294618 257546 294854
rect 257782 294618 257866 294854
rect 258102 294618 258134 294854
rect 257514 259174 258134 294618
rect 257514 258938 257546 259174
rect 257782 258938 257866 259174
rect 258102 258938 258134 259174
rect 257514 258854 258134 258938
rect 257514 258618 257546 258854
rect 257782 258618 257866 258854
rect 258102 258618 258134 258854
rect 257514 223174 258134 258618
rect 259502 242997 259562 328475
rect 261234 298894 261854 334338
rect 261234 298658 261266 298894
rect 261502 298658 261586 298894
rect 261822 298658 261854 298894
rect 261234 298574 261854 298658
rect 261234 298338 261266 298574
rect 261502 298338 261586 298574
rect 261822 298338 261854 298574
rect 261234 262894 261854 298338
rect 261234 262658 261266 262894
rect 261502 262658 261586 262894
rect 261822 262658 261854 262894
rect 261234 262574 261854 262658
rect 261234 262338 261266 262574
rect 261502 262338 261586 262574
rect 261822 262338 261854 262574
rect 259499 242996 259565 242997
rect 259499 242932 259500 242996
rect 259564 242932 259565 242996
rect 259499 242931 259565 242932
rect 257514 222938 257546 223174
rect 257782 222938 257866 223174
rect 258102 222938 258134 223174
rect 257514 222854 258134 222938
rect 257514 222618 257546 222854
rect 257782 222618 257866 222854
rect 258102 222618 258134 222854
rect 255267 215252 255333 215253
rect 255267 215188 255268 215252
rect 255332 215188 255333 215252
rect 255267 215187 255333 215188
rect 256555 192540 256621 192541
rect 256555 192476 256556 192540
rect 256620 192476 256621 192540
rect 256555 192475 256621 192476
rect 253794 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 254414 183454
rect 253794 183134 254414 183218
rect 253794 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 254414 183134
rect 253794 147454 254414 182898
rect 253794 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 254414 147454
rect 253794 147134 254414 147218
rect 253794 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 254414 147134
rect 253794 111454 254414 146898
rect 253794 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 254414 111454
rect 253794 111134 254414 111218
rect 253794 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 254414 111134
rect 253059 92308 253125 92309
rect 253059 92244 253060 92308
rect 253124 92244 253125 92308
rect 253059 92243 253125 92244
rect 253794 75454 254414 110898
rect 253794 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 254414 75454
rect 253794 75134 254414 75218
rect 253794 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 254414 75134
rect 252326 53350 252570 53410
rect 249747 50964 249813 50965
rect 249747 50900 249748 50964
rect 249812 50900 249813 50964
rect 249747 50899 249813 50900
rect 246954 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 247574 32614
rect 246954 32294 247574 32378
rect 246954 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 247574 32294
rect 244043 25532 244109 25533
rect 244043 25468 244044 25532
rect 244108 25468 244109 25532
rect 244043 25467 244109 25468
rect 243234 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 243854 -5146
rect 243234 -5466 243854 -5382
rect 243234 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 243854 -5466
rect 243234 -5734 243854 -5702
rect 228954 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 229574 -6106
rect 228954 -6426 229574 -6342
rect 228954 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 229574 -6426
rect 228954 -7654 229574 -6662
rect 246954 -7066 247574 32058
rect 252326 11797 252386 53350
rect 252510 53141 252570 53350
rect 252507 53140 252573 53141
rect 252507 53076 252508 53140
rect 252572 53076 252573 53140
rect 252507 53075 252573 53076
rect 253794 39454 254414 74898
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 252323 11796 252389 11797
rect 252323 11732 252324 11796
rect 252388 11732 252389 11796
rect 252323 11731 252389 11732
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 256558 3365 256618 192475
rect 257514 187174 258134 222618
rect 257514 186938 257546 187174
rect 257782 186938 257866 187174
rect 258102 186938 258134 187174
rect 257514 186854 258134 186938
rect 257514 186618 257546 186854
rect 257782 186618 257866 186854
rect 258102 186618 258134 186854
rect 257514 151174 258134 186618
rect 257514 150938 257546 151174
rect 257782 150938 257866 151174
rect 258102 150938 258134 151174
rect 257514 150854 258134 150938
rect 257514 150618 257546 150854
rect 257782 150618 257866 150854
rect 258102 150618 258134 150854
rect 257514 115174 258134 150618
rect 261234 226894 261854 262338
rect 261234 226658 261266 226894
rect 261502 226658 261586 226894
rect 261822 226658 261854 226894
rect 261234 226574 261854 226658
rect 261234 226338 261266 226574
rect 261502 226338 261586 226574
rect 261822 226338 261854 226574
rect 261234 190894 261854 226338
rect 261234 190658 261266 190894
rect 261502 190658 261586 190894
rect 261822 190658 261854 190894
rect 261234 190574 261854 190658
rect 261234 190338 261266 190574
rect 261502 190338 261586 190574
rect 261822 190338 261854 190574
rect 261234 154894 261854 190338
rect 261234 154658 261266 154894
rect 261502 154658 261586 154894
rect 261822 154658 261854 154894
rect 261234 154574 261854 154658
rect 261234 154338 261266 154574
rect 261502 154338 261586 154574
rect 261822 154338 261854 154574
rect 258579 130660 258645 130661
rect 258579 130596 258580 130660
rect 258644 130596 258645 130660
rect 258579 130595 258645 130596
rect 257514 114938 257546 115174
rect 257782 114938 257866 115174
rect 258102 114938 258134 115174
rect 257514 114854 258134 114938
rect 257514 114618 257546 114854
rect 257782 114618 257866 114854
rect 258102 114618 258134 114854
rect 257514 79174 258134 114618
rect 257514 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 258134 79174
rect 257514 78854 258134 78938
rect 257514 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 258134 78854
rect 257514 43174 258134 78618
rect 258582 71093 258642 130595
rect 260051 126444 260117 126445
rect 260051 126380 260052 126444
rect 260116 126380 260117 126444
rect 260051 126379 260117 126380
rect 258579 71092 258645 71093
rect 258579 71028 258580 71092
rect 258644 71028 258645 71092
rect 258579 71027 258645 71028
rect 260054 55861 260114 126379
rect 261234 118894 261854 154338
rect 264954 374614 265574 375600
rect 264954 374378 264986 374614
rect 265222 374378 265306 374614
rect 265542 374378 265574 374614
rect 264954 374294 265574 374378
rect 264954 374058 264986 374294
rect 265222 374058 265306 374294
rect 265542 374058 265574 374294
rect 264954 338614 265574 374058
rect 267595 364444 267661 364445
rect 267595 364380 267596 364444
rect 267660 364380 267661 364444
rect 267595 364379 267661 364380
rect 264954 338378 264986 338614
rect 265222 338378 265306 338614
rect 265542 338378 265574 338614
rect 264954 338294 265574 338378
rect 264954 338058 264986 338294
rect 265222 338058 265306 338294
rect 265542 338058 265574 338294
rect 264954 302614 265574 338058
rect 264954 302378 264986 302614
rect 265222 302378 265306 302614
rect 265542 302378 265574 302614
rect 264954 302294 265574 302378
rect 264954 302058 264986 302294
rect 265222 302058 265306 302294
rect 265542 302058 265574 302294
rect 264954 266614 265574 302058
rect 264954 266378 264986 266614
rect 265222 266378 265306 266614
rect 265542 266378 265574 266614
rect 264954 266294 265574 266378
rect 264954 266058 264986 266294
rect 265222 266058 265306 266294
rect 265542 266058 265574 266294
rect 264954 230614 265574 266058
rect 264954 230378 264986 230614
rect 265222 230378 265306 230614
rect 265542 230378 265574 230614
rect 264954 230294 265574 230378
rect 264954 230058 264986 230294
rect 265222 230058 265306 230294
rect 265542 230058 265574 230294
rect 264954 194614 265574 230058
rect 264954 194378 264986 194614
rect 265222 194378 265306 194614
rect 265542 194378 265574 194614
rect 264954 194294 265574 194378
rect 264954 194058 264986 194294
rect 265222 194058 265306 194294
rect 265542 194058 265574 194294
rect 264954 158614 265574 194058
rect 264954 158378 264986 158614
rect 265222 158378 265306 158614
rect 265542 158378 265574 158614
rect 264954 158294 265574 158378
rect 264954 158058 264986 158294
rect 265222 158058 265306 158294
rect 265542 158058 265574 158294
rect 262811 134876 262877 134877
rect 262811 134812 262812 134876
rect 262876 134812 262877 134876
rect 262811 134811 262877 134812
rect 261234 118658 261266 118894
rect 261502 118658 261586 118894
rect 261822 118658 261854 118894
rect 261234 118574 261854 118658
rect 261234 118338 261266 118574
rect 261502 118338 261586 118574
rect 261822 118338 261854 118574
rect 261234 82894 261854 118338
rect 261234 82658 261266 82894
rect 261502 82658 261586 82894
rect 261822 82658 261854 82894
rect 261234 82574 261854 82658
rect 261234 82338 261266 82574
rect 261502 82338 261586 82574
rect 261822 82338 261854 82574
rect 260051 55860 260117 55861
rect 260051 55796 260052 55860
rect 260116 55796 260117 55860
rect 260051 55795 260117 55796
rect 257514 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 258134 43174
rect 257514 42854 258134 42938
rect 257514 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 258134 42854
rect 257514 7174 258134 42618
rect 257514 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 258134 7174
rect 257514 6854 258134 6938
rect 257514 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 258134 6854
rect 256555 3364 256621 3365
rect 256555 3300 256556 3364
rect 256620 3300 256621 3364
rect 256555 3299 256621 3300
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -1894 254414 -902
rect 257514 -2266 258134 6618
rect 257514 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 258134 -2266
rect 257514 -2586 258134 -2502
rect 257514 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 258134 -2586
rect 257514 -3814 258134 -2822
rect 261234 46894 261854 82338
rect 262814 59941 262874 134811
rect 264099 130116 264165 130117
rect 264099 130052 264100 130116
rect 264164 130052 264165 130116
rect 264099 130051 264165 130052
rect 264102 105637 264162 130051
rect 264954 122614 265574 158058
rect 266859 140452 266925 140453
rect 266859 140388 266860 140452
rect 266924 140388 266925 140452
rect 266859 140387 266925 140388
rect 264954 122378 264986 122614
rect 265222 122378 265306 122614
rect 265542 122378 265574 122614
rect 264954 122294 265574 122378
rect 264954 122058 264986 122294
rect 265222 122058 265306 122294
rect 265542 122058 265574 122294
rect 264099 105636 264165 105637
rect 264099 105572 264100 105636
rect 264164 105572 264165 105636
rect 264099 105571 264165 105572
rect 262995 102236 263061 102237
rect 262995 102172 262996 102236
rect 263060 102172 263061 102236
rect 262995 102171 263061 102172
rect 262998 100061 263058 102171
rect 262995 100060 263061 100061
rect 262995 99996 262996 100060
rect 263060 99996 263061 100060
rect 262995 99995 263061 99996
rect 264099 97476 264165 97477
rect 264099 97412 264100 97476
rect 264164 97412 264165 97476
rect 264099 97411 264165 97412
rect 264102 80749 264162 97411
rect 264954 86614 265574 122058
rect 264954 86378 264986 86614
rect 265222 86378 265306 86614
rect 265542 86378 265574 86614
rect 264954 86294 265574 86378
rect 264954 86058 264986 86294
rect 265222 86058 265306 86294
rect 265542 86058 265574 86294
rect 264099 80748 264165 80749
rect 264099 80684 264100 80748
rect 264164 80684 264165 80748
rect 264099 80683 264165 80684
rect 262811 59940 262877 59941
rect 262811 59876 262812 59940
rect 262876 59876 262877 59940
rect 262811 59875 262877 59876
rect 261234 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 261854 46894
rect 261234 46574 261854 46658
rect 261234 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 261854 46574
rect 261234 10894 261854 46338
rect 261234 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 261854 10894
rect 261234 10574 261854 10658
rect 261234 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 261854 10574
rect 261234 -4186 261854 10338
rect 261234 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 261854 -4186
rect 261234 -4506 261854 -4422
rect 261234 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 261854 -4506
rect 261234 -5734 261854 -4742
rect 264954 50614 265574 86058
rect 264954 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 265574 50614
rect 264954 50294 265574 50378
rect 264954 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 265574 50294
rect 264954 14614 265574 50058
rect 266862 17237 266922 140387
rect 267598 94621 267658 364379
rect 271794 345454 272414 375600
rect 271794 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 272414 345454
rect 271794 345134 272414 345218
rect 271794 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 272414 345134
rect 271794 309454 272414 344898
rect 271794 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 272414 309454
rect 271794 309134 272414 309218
rect 271794 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 272414 309134
rect 267779 295356 267845 295357
rect 267779 295292 267780 295356
rect 267844 295292 267845 295356
rect 267779 295291 267845 295292
rect 267782 108901 267842 295291
rect 271794 273454 272414 308898
rect 271794 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 272414 273454
rect 271794 273134 272414 273218
rect 271794 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 272414 273134
rect 271794 237454 272414 272898
rect 271794 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 272414 237454
rect 271794 237134 272414 237218
rect 271794 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 272414 237134
rect 271794 201454 272414 236898
rect 271794 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 272414 201454
rect 271794 201134 272414 201218
rect 271794 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 272414 201134
rect 271794 178000 272414 200898
rect 275514 349174 276134 375600
rect 275514 348938 275546 349174
rect 275782 348938 275866 349174
rect 276102 348938 276134 349174
rect 275514 348854 276134 348938
rect 275514 348618 275546 348854
rect 275782 348618 275866 348854
rect 276102 348618 276134 348854
rect 275514 313174 276134 348618
rect 275514 312938 275546 313174
rect 275782 312938 275866 313174
rect 276102 312938 276134 313174
rect 275514 312854 276134 312938
rect 275514 312618 275546 312854
rect 275782 312618 275866 312854
rect 276102 312618 276134 312854
rect 275514 277174 276134 312618
rect 275514 276938 275546 277174
rect 275782 276938 275866 277174
rect 276102 276938 276134 277174
rect 275514 276854 276134 276938
rect 275514 276618 275546 276854
rect 275782 276618 275866 276854
rect 276102 276618 276134 276854
rect 275514 241174 276134 276618
rect 275514 240938 275546 241174
rect 275782 240938 275866 241174
rect 276102 240938 276134 241174
rect 275514 240854 276134 240938
rect 275514 240618 275546 240854
rect 275782 240618 275866 240854
rect 276102 240618 276134 240854
rect 275514 205174 276134 240618
rect 275514 204938 275546 205174
rect 275782 204938 275866 205174
rect 276102 204938 276134 205174
rect 275514 204854 276134 204938
rect 275514 204618 275546 204854
rect 275782 204618 275866 204854
rect 276102 204618 276134 204854
rect 275514 178000 276134 204618
rect 279234 352894 279854 375600
rect 279234 352658 279266 352894
rect 279502 352658 279586 352894
rect 279822 352658 279854 352894
rect 279234 352574 279854 352658
rect 279234 352338 279266 352574
rect 279502 352338 279586 352574
rect 279822 352338 279854 352574
rect 279234 316894 279854 352338
rect 279234 316658 279266 316894
rect 279502 316658 279586 316894
rect 279822 316658 279854 316894
rect 279234 316574 279854 316658
rect 279234 316338 279266 316574
rect 279502 316338 279586 316574
rect 279822 316338 279854 316574
rect 279234 280894 279854 316338
rect 279234 280658 279266 280894
rect 279502 280658 279586 280894
rect 279822 280658 279854 280894
rect 279234 280574 279854 280658
rect 279234 280338 279266 280574
rect 279502 280338 279586 280574
rect 279822 280338 279854 280574
rect 279234 244894 279854 280338
rect 282954 356614 283574 375600
rect 287651 367572 287717 367573
rect 287651 367508 287652 367572
rect 287716 367508 287717 367572
rect 287651 367507 287717 367508
rect 282954 356378 282986 356614
rect 283222 356378 283306 356614
rect 283542 356378 283574 356614
rect 282954 356294 283574 356378
rect 282954 356058 282986 356294
rect 283222 356058 283306 356294
rect 283542 356058 283574 356294
rect 282954 320614 283574 356058
rect 282954 320378 282986 320614
rect 283222 320378 283306 320614
rect 283542 320378 283574 320614
rect 282954 320294 283574 320378
rect 282954 320058 282986 320294
rect 283222 320058 283306 320294
rect 283542 320058 283574 320294
rect 282954 284614 283574 320058
rect 286179 285700 286245 285701
rect 286179 285636 286180 285700
rect 286244 285636 286245 285700
rect 286179 285635 286245 285636
rect 282954 284378 282986 284614
rect 283222 284378 283306 284614
rect 283542 284378 283574 284614
rect 282954 284294 283574 284378
rect 282954 284058 282986 284294
rect 283222 284058 283306 284294
rect 283542 284058 283574 284294
rect 280291 280260 280357 280261
rect 280291 280196 280292 280260
rect 280356 280196 280357 280260
rect 280291 280195 280357 280196
rect 279234 244658 279266 244894
rect 279502 244658 279586 244894
rect 279822 244658 279854 244894
rect 279234 244574 279854 244658
rect 279234 244338 279266 244574
rect 279502 244338 279586 244574
rect 279822 244338 279854 244574
rect 279234 208894 279854 244338
rect 279234 208658 279266 208894
rect 279502 208658 279586 208894
rect 279822 208658 279854 208894
rect 279234 208574 279854 208658
rect 279234 208338 279266 208574
rect 279502 208338 279586 208574
rect 279822 208338 279854 208574
rect 277899 189956 277965 189957
rect 277899 189892 277900 189956
rect 277964 189892 277965 189956
rect 277899 189891 277965 189892
rect 277902 175813 277962 189891
rect 278819 181524 278885 181525
rect 278819 181460 278820 181524
rect 278884 181460 278885 181524
rect 278819 181459 278885 181460
rect 277899 175812 277965 175813
rect 277899 175748 277900 175812
rect 277964 175748 277965 175812
rect 277899 175747 277965 175748
rect 272207 165454 272527 165486
rect 272207 165218 272249 165454
rect 272485 165218 272527 165454
rect 272207 165134 272527 165218
rect 272207 164898 272249 165134
rect 272485 164898 272527 165134
rect 272207 164866 272527 164898
rect 275471 165454 275791 165486
rect 275471 165218 275513 165454
rect 275749 165218 275791 165454
rect 275471 165134 275791 165218
rect 275471 164898 275513 165134
rect 275749 164898 275791 165134
rect 275471 164866 275791 164898
rect 270575 147454 270895 147486
rect 270575 147218 270617 147454
rect 270853 147218 270895 147454
rect 270575 147134 270895 147218
rect 270575 146898 270617 147134
rect 270853 146898 270895 147134
rect 270575 146866 270895 146898
rect 273839 147454 274159 147486
rect 273839 147218 273881 147454
rect 274117 147218 274159 147454
rect 273839 147134 274159 147218
rect 273839 146898 273881 147134
rect 274117 146898 274159 147134
rect 273839 146866 274159 146898
rect 277103 147454 277423 147486
rect 277103 147218 277145 147454
rect 277381 147218 277423 147454
rect 277103 147134 277423 147218
rect 277103 146898 277145 147134
rect 277381 146898 277423 147134
rect 277103 146866 277423 146898
rect 272207 129454 272527 129486
rect 272207 129218 272249 129454
rect 272485 129218 272527 129454
rect 272207 129134 272527 129218
rect 272207 128898 272249 129134
rect 272485 128898 272527 129134
rect 272207 128866 272527 128898
rect 275471 129454 275791 129486
rect 275471 129218 275513 129454
rect 275749 129218 275791 129454
rect 275471 129134 275791 129218
rect 275471 128898 275513 129134
rect 275749 128898 275791 129134
rect 275471 128866 275791 128898
rect 278822 113190 278882 181459
rect 279234 178000 279854 208338
rect 280294 180810 280354 280195
rect 282131 270604 282197 270605
rect 282131 270540 282132 270604
rect 282196 270540 282197 270604
rect 282131 270539 282197 270540
rect 280475 182884 280541 182885
rect 280475 182820 280476 182884
rect 280540 182820 280541 182884
rect 280475 182819 280541 182820
rect 280110 180750 280354 180810
rect 279371 177172 279437 177173
rect 279371 177108 279372 177172
rect 279436 177108 279437 177172
rect 279371 177107 279437 177108
rect 279374 170645 279434 177107
rect 279371 170644 279437 170645
rect 279371 170580 279372 170644
rect 279436 170580 279437 170644
rect 279371 170579 279437 170580
rect 280110 139773 280170 180750
rect 280478 161490 280538 182819
rect 281579 180028 281645 180029
rect 281579 179964 281580 180028
rect 281644 179964 281645 180028
rect 281579 179963 281645 179964
rect 280294 161430 280538 161490
rect 280107 139772 280173 139773
rect 280107 139708 280108 139772
rect 280172 139708 280173 139772
rect 280107 139707 280173 139708
rect 278822 113130 279434 113190
rect 270575 111454 270895 111486
rect 270575 111218 270617 111454
rect 270853 111218 270895 111454
rect 270575 111134 270895 111218
rect 270575 110898 270617 111134
rect 270853 110898 270895 111134
rect 270575 110866 270895 110898
rect 273839 111454 274159 111486
rect 273839 111218 273881 111454
rect 274117 111218 274159 111454
rect 273839 111134 274159 111218
rect 273839 110898 273881 111134
rect 274117 110898 274159 111134
rect 273839 110866 274159 110898
rect 277103 111454 277423 111486
rect 277103 111218 277145 111454
rect 277381 111218 277423 111454
rect 277103 111134 277423 111218
rect 277103 110898 277145 111134
rect 277381 110898 277423 111134
rect 277103 110866 277423 110898
rect 267779 108900 267845 108901
rect 267779 108836 267780 108900
rect 267844 108836 267845 108900
rect 267779 108835 267845 108836
rect 267963 107132 268029 107133
rect 267963 107068 267964 107132
rect 268028 107068 268029 107132
rect 267963 107067 268029 107068
rect 267779 99244 267845 99245
rect 267779 99180 267780 99244
rect 267844 99180 267845 99244
rect 267779 99179 267845 99180
rect 267595 94620 267661 94621
rect 267595 94556 267596 94620
rect 267660 94556 267661 94620
rect 267595 94555 267661 94556
rect 267782 36549 267842 99179
rect 267966 62797 268026 107067
rect 279374 100605 279434 113130
rect 280294 105501 280354 161430
rect 281582 155005 281642 179963
rect 282134 179485 282194 270539
rect 282954 248614 283574 284058
rect 282954 248378 282986 248614
rect 283222 248378 283306 248614
rect 283542 248378 283574 248614
rect 282954 248294 283574 248378
rect 282954 248058 282986 248294
rect 283222 248058 283306 248294
rect 283542 248058 283574 248294
rect 282954 212614 283574 248058
rect 283787 225588 283853 225589
rect 283787 225524 283788 225588
rect 283852 225524 283853 225588
rect 283787 225523 283853 225524
rect 282954 212378 282986 212614
rect 283222 212378 283306 212614
rect 283542 212378 283574 212614
rect 282954 212294 283574 212378
rect 282954 212058 282986 212294
rect 283222 212058 283306 212294
rect 283542 212058 283574 212294
rect 282131 179484 282197 179485
rect 282131 179420 282132 179484
rect 282196 179420 282197 179484
rect 282131 179419 282197 179420
rect 282954 176614 283574 212058
rect 282954 176378 282986 176614
rect 283222 176378 283306 176614
rect 283542 176378 283574 176614
rect 282954 176294 283574 176378
rect 282954 176058 282986 176294
rect 283222 176058 283306 176294
rect 283542 176058 283574 176294
rect 281579 155004 281645 155005
rect 281579 154940 281580 155004
rect 281644 154940 281645 155004
rect 281579 154939 281645 154940
rect 282131 153780 282197 153781
rect 282131 153716 282132 153780
rect 282196 153716 282197 153780
rect 282131 153715 282197 153716
rect 282134 132157 282194 153715
rect 282954 140614 283574 176058
rect 283790 157317 283850 225523
rect 284523 207636 284589 207637
rect 284523 207572 284524 207636
rect 284588 207572 284589 207636
rect 284523 207571 284589 207572
rect 284339 176764 284405 176765
rect 284339 176700 284340 176764
rect 284404 176700 284405 176764
rect 284339 176699 284405 176700
rect 283787 157316 283853 157317
rect 283787 157252 283788 157316
rect 283852 157252 283853 157316
rect 283787 157251 283853 157252
rect 282954 140378 282986 140614
rect 283222 140378 283306 140614
rect 283542 140378 283574 140614
rect 282954 140294 283574 140378
rect 282954 140058 282986 140294
rect 283222 140058 283306 140294
rect 283542 140058 283574 140294
rect 282131 132156 282197 132157
rect 282131 132092 282132 132156
rect 282196 132092 282197 132156
rect 282131 132091 282197 132092
rect 280291 105500 280357 105501
rect 280291 105436 280292 105500
rect 280356 105436 280357 105500
rect 280291 105435 280357 105436
rect 282954 104614 283574 140058
rect 282954 104378 282986 104614
rect 283222 104378 283306 104614
rect 283542 104378 283574 104614
rect 282954 104294 283574 104378
rect 282954 104058 282986 104294
rect 283222 104058 283306 104294
rect 283542 104058 283574 104294
rect 279371 100604 279437 100605
rect 279371 100540 279372 100604
rect 279436 100540 279437 100604
rect 279371 100539 279437 100540
rect 271794 93454 272414 94000
rect 271794 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 272414 93454
rect 271794 93134 272414 93218
rect 271794 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 272414 93134
rect 267963 62796 268029 62797
rect 267963 62732 267964 62796
rect 268028 62732 268029 62796
rect 267963 62731 268029 62732
rect 271794 57454 272414 92898
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 267779 36548 267845 36549
rect 267779 36484 267780 36548
rect 267844 36484 267845 36548
rect 267779 36483 267845 36484
rect 271794 21454 272414 56898
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 266859 17236 266925 17237
rect 266859 17172 266860 17236
rect 266924 17172 266925 17236
rect 266859 17171 266925 17172
rect 264954 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 265574 14614
rect 264954 14294 265574 14378
rect 264954 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 265574 14294
rect 246954 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 247574 -7066
rect 246954 -7386 247574 -7302
rect 246954 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 247574 -7386
rect 246954 -7654 247574 -7622
rect 264954 -6106 265574 14058
rect 271794 -1306 272414 20898
rect 271794 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 272414 -1306
rect 271794 -1626 272414 -1542
rect 271794 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 272414 -1626
rect 271794 -1894 272414 -1862
rect 275514 61174 276134 94000
rect 275514 60938 275546 61174
rect 275782 60938 275866 61174
rect 276102 60938 276134 61174
rect 275514 60854 276134 60938
rect 275514 60618 275546 60854
rect 275782 60618 275866 60854
rect 276102 60618 276134 60854
rect 275514 25174 276134 60618
rect 275514 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 276134 25174
rect 275514 24854 276134 24938
rect 275514 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 276134 24854
rect 275514 -3226 276134 24618
rect 275514 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 276134 -3226
rect 275514 -3546 276134 -3462
rect 275514 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 276134 -3546
rect 275514 -3814 276134 -3782
rect 279234 64894 279854 94000
rect 279234 64658 279266 64894
rect 279502 64658 279586 64894
rect 279822 64658 279854 64894
rect 279234 64574 279854 64658
rect 279234 64338 279266 64574
rect 279502 64338 279586 64574
rect 279822 64338 279854 64574
rect 279234 28894 279854 64338
rect 279234 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 279854 28894
rect 279234 28574 279854 28658
rect 279234 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 279854 28574
rect 279234 -5146 279854 28338
rect 279234 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 279854 -5146
rect 279234 -5466 279854 -5382
rect 279234 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 279854 -5466
rect 279234 -5734 279854 -5702
rect 282954 68614 283574 104058
rect 284342 101693 284402 176699
rect 284526 133653 284586 207571
rect 285627 183020 285693 183021
rect 285627 182956 285628 183020
rect 285692 182956 285693 183020
rect 285627 182955 285693 182956
rect 284523 133652 284589 133653
rect 284523 133588 284524 133652
rect 284588 133588 284589 133652
rect 284523 133587 284589 133588
rect 285630 111621 285690 182955
rect 286182 160717 286242 285635
rect 287099 193900 287165 193901
rect 287099 193836 287100 193900
rect 287164 193836 287165 193900
rect 287099 193835 287165 193836
rect 286179 160716 286245 160717
rect 286179 160652 286180 160716
rect 286244 160652 286245 160716
rect 286179 160651 286245 160652
rect 285627 111620 285693 111621
rect 285627 111556 285628 111620
rect 285692 111556 285693 111620
rect 285627 111555 285693 111556
rect 287102 109445 287162 193835
rect 287099 109444 287165 109445
rect 287099 109380 287100 109444
rect 287164 109380 287165 109444
rect 287099 109379 287165 109380
rect 284339 101692 284405 101693
rect 284339 101628 284340 101692
rect 284404 101628 284405 101692
rect 284339 101627 284405 101628
rect 282954 68378 282986 68614
rect 283222 68378 283306 68614
rect 283542 68378 283574 68614
rect 282954 68294 283574 68378
rect 282954 68058 282986 68294
rect 283222 68058 283306 68294
rect 283542 68058 283574 68294
rect 282954 32614 283574 68058
rect 287654 64157 287714 367507
rect 289794 363454 290414 375600
rect 289794 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 290414 363454
rect 289794 363134 290414 363218
rect 289794 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 290414 363134
rect 289794 327454 290414 362898
rect 289794 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 290414 327454
rect 289794 327134 290414 327218
rect 289794 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 290414 327134
rect 289794 291454 290414 326898
rect 289794 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 290414 291454
rect 289794 291134 290414 291218
rect 289794 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 290414 291134
rect 289794 255454 290414 290898
rect 289794 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 290414 255454
rect 289794 255134 290414 255218
rect 289794 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 290414 255134
rect 289794 219454 290414 254898
rect 289794 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 290414 219454
rect 289794 219134 290414 219218
rect 289794 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 290414 219134
rect 288571 201516 288637 201517
rect 288571 201452 288572 201516
rect 288636 201452 288637 201516
rect 288571 201451 288637 201452
rect 288387 194444 288453 194445
rect 288387 194380 288388 194444
rect 288452 194380 288453 194444
rect 288387 194379 288453 194380
rect 287651 64156 287717 64157
rect 287651 64092 287652 64156
rect 287716 64092 287717 64156
rect 287651 64091 287717 64092
rect 288390 60485 288450 194379
rect 288574 62797 288634 201451
rect 289794 183454 290414 218898
rect 293514 367174 294134 375600
rect 293514 366938 293546 367174
rect 293782 366938 293866 367174
rect 294102 366938 294134 367174
rect 293514 366854 294134 366938
rect 293514 366618 293546 366854
rect 293782 366618 293866 366854
rect 294102 366618 294134 366854
rect 293514 331174 294134 366618
rect 297234 370894 297854 375600
rect 297234 370658 297266 370894
rect 297502 370658 297586 370894
rect 297822 370658 297854 370894
rect 297234 370574 297854 370658
rect 297234 370338 297266 370574
rect 297502 370338 297586 370574
rect 297822 370338 297854 370574
rect 295931 350572 295997 350573
rect 295931 350508 295932 350572
rect 295996 350508 295997 350572
rect 295931 350507 295997 350508
rect 293514 330938 293546 331174
rect 293782 330938 293866 331174
rect 294102 330938 294134 331174
rect 293514 330854 294134 330938
rect 293514 330618 293546 330854
rect 293782 330618 293866 330854
rect 294102 330618 294134 330854
rect 293514 295174 294134 330618
rect 293514 294938 293546 295174
rect 293782 294938 293866 295174
rect 294102 294938 294134 295174
rect 293514 294854 294134 294938
rect 293514 294618 293546 294854
rect 293782 294618 293866 294854
rect 294102 294618 294134 294854
rect 293514 259174 294134 294618
rect 293514 258938 293546 259174
rect 293782 258938 293866 259174
rect 294102 258938 294134 259174
rect 293514 258854 294134 258938
rect 293514 258618 293546 258854
rect 293782 258618 293866 258854
rect 294102 258618 294134 258854
rect 293514 223174 294134 258618
rect 293514 222938 293546 223174
rect 293782 222938 293866 223174
rect 294102 222938 294134 223174
rect 293514 222854 294134 222938
rect 293514 222618 293546 222854
rect 293782 222618 293866 222854
rect 294102 222618 294134 222854
rect 290595 207636 290661 207637
rect 290595 207572 290596 207636
rect 290660 207572 290661 207636
rect 290595 207571 290661 207572
rect 289794 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 290414 183454
rect 289794 183134 290414 183218
rect 289794 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 290414 183134
rect 289794 147454 290414 182898
rect 289794 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 290414 147454
rect 289794 147134 290414 147218
rect 289794 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 290414 147134
rect 289794 111454 290414 146898
rect 289794 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 290414 111454
rect 289794 111134 290414 111218
rect 289794 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 290414 111134
rect 289794 75454 290414 110898
rect 289794 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 290414 75454
rect 289794 75134 290414 75218
rect 289794 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 290414 75134
rect 288571 62796 288637 62797
rect 288571 62732 288572 62796
rect 288636 62732 288637 62796
rect 288571 62731 288637 62732
rect 288387 60484 288453 60485
rect 288387 60420 288388 60484
rect 288452 60420 288453 60484
rect 288387 60419 288453 60420
rect 282954 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 283574 32614
rect 282954 32294 283574 32378
rect 282954 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 283574 32294
rect 264954 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 265574 -6106
rect 264954 -6426 265574 -6342
rect 264954 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 265574 -6426
rect 264954 -7654 265574 -6662
rect 282954 -7066 283574 32058
rect 289794 39454 290414 74898
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 290598 3501 290658 207571
rect 291699 199476 291765 199477
rect 291699 199412 291700 199476
rect 291764 199412 291765 199476
rect 291699 199411 291765 199412
rect 291702 87005 291762 199411
rect 293514 187174 294134 222618
rect 293514 186938 293546 187174
rect 293782 186938 293866 187174
rect 294102 186938 294134 187174
rect 293514 186854 294134 186938
rect 293514 186618 293546 186854
rect 293782 186618 293866 186854
rect 294102 186618 294134 186854
rect 293514 151174 294134 186618
rect 293514 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 294134 151174
rect 293514 150854 294134 150938
rect 293514 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 294134 150854
rect 293514 115174 294134 150618
rect 293514 114938 293546 115174
rect 293782 114938 293866 115174
rect 294102 114938 294134 115174
rect 293514 114854 294134 114938
rect 293514 114618 293546 114854
rect 293782 114618 293866 114854
rect 294102 114618 294134 114854
rect 291699 87004 291765 87005
rect 291699 86940 291700 87004
rect 291764 86940 291765 87004
rect 291699 86939 291765 86940
rect 291702 3501 291762 86939
rect 293514 79174 294134 114618
rect 293514 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 294134 79174
rect 293514 78854 294134 78938
rect 293514 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 294134 78854
rect 293514 43174 294134 78618
rect 293514 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 294134 43174
rect 293514 42854 294134 42938
rect 293514 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 294134 42854
rect 293514 7174 294134 42618
rect 295934 13701 295994 350507
rect 297234 334894 297854 370338
rect 297234 334658 297266 334894
rect 297502 334658 297586 334894
rect 297822 334658 297854 334894
rect 297234 334574 297854 334658
rect 297234 334338 297266 334574
rect 297502 334338 297586 334574
rect 297822 334338 297854 334574
rect 297234 298894 297854 334338
rect 297234 298658 297266 298894
rect 297502 298658 297586 298894
rect 297822 298658 297854 298894
rect 297234 298574 297854 298658
rect 297234 298338 297266 298574
rect 297502 298338 297586 298574
rect 297822 298338 297854 298574
rect 297234 262894 297854 298338
rect 297234 262658 297266 262894
rect 297502 262658 297586 262894
rect 297822 262658 297854 262894
rect 297234 262574 297854 262658
rect 297234 262338 297266 262574
rect 297502 262338 297586 262574
rect 297822 262338 297854 262574
rect 297234 226894 297854 262338
rect 297234 226658 297266 226894
rect 297502 226658 297586 226894
rect 297822 226658 297854 226894
rect 297234 226574 297854 226658
rect 297234 226338 297266 226574
rect 297502 226338 297586 226574
rect 297822 226338 297854 226574
rect 297234 190894 297854 226338
rect 300954 374614 301574 375600
rect 300954 374378 300986 374614
rect 301222 374378 301306 374614
rect 301542 374378 301574 374614
rect 300954 374294 301574 374378
rect 300954 374058 300986 374294
rect 301222 374058 301306 374294
rect 301542 374058 301574 374294
rect 300954 338614 301574 374058
rect 300954 338378 300986 338614
rect 301222 338378 301306 338614
rect 301542 338378 301574 338614
rect 300954 338294 301574 338378
rect 300954 338058 300986 338294
rect 301222 338058 301306 338294
rect 301542 338058 301574 338294
rect 300954 302614 301574 338058
rect 300954 302378 300986 302614
rect 301222 302378 301306 302614
rect 301542 302378 301574 302614
rect 300954 302294 301574 302378
rect 300954 302058 300986 302294
rect 301222 302058 301306 302294
rect 301542 302058 301574 302294
rect 300954 266614 301574 302058
rect 300954 266378 300986 266614
rect 301222 266378 301306 266614
rect 301542 266378 301574 266614
rect 300954 266294 301574 266378
rect 300954 266058 300986 266294
rect 301222 266058 301306 266294
rect 301542 266058 301574 266294
rect 300954 230614 301574 266058
rect 300954 230378 300986 230614
rect 301222 230378 301306 230614
rect 301542 230378 301574 230614
rect 300954 230294 301574 230378
rect 300954 230058 300986 230294
rect 301222 230058 301306 230294
rect 301542 230058 301574 230294
rect 298139 217292 298205 217293
rect 298139 217228 298140 217292
rect 298204 217228 298205 217292
rect 298139 217227 298205 217228
rect 297234 190658 297266 190894
rect 297502 190658 297586 190894
rect 297822 190658 297854 190894
rect 297234 190574 297854 190658
rect 297234 190338 297266 190574
rect 297502 190338 297586 190574
rect 297822 190338 297854 190574
rect 297234 154894 297854 190338
rect 297234 154658 297266 154894
rect 297502 154658 297586 154894
rect 297822 154658 297854 154894
rect 297234 154574 297854 154658
rect 297234 154338 297266 154574
rect 297502 154338 297586 154574
rect 297822 154338 297854 154574
rect 297234 118894 297854 154338
rect 298142 147797 298202 217227
rect 300954 194614 301574 230058
rect 300954 194378 300986 194614
rect 301222 194378 301306 194614
rect 301542 194378 301574 194614
rect 300954 194294 301574 194378
rect 300954 194058 300986 194294
rect 301222 194058 301306 194294
rect 301542 194058 301574 194294
rect 299611 188460 299677 188461
rect 299611 188396 299612 188460
rect 299676 188396 299677 188460
rect 299611 188395 299677 188396
rect 298139 147796 298205 147797
rect 298139 147732 298140 147796
rect 298204 147732 298205 147796
rect 298139 147731 298205 147732
rect 297234 118658 297266 118894
rect 297502 118658 297586 118894
rect 297822 118658 297854 118894
rect 297234 118574 297854 118658
rect 297234 118338 297266 118574
rect 297502 118338 297586 118574
rect 297822 118338 297854 118574
rect 297234 82894 297854 118338
rect 297234 82658 297266 82894
rect 297502 82658 297586 82894
rect 297822 82658 297854 82894
rect 297234 82574 297854 82658
rect 297234 82338 297266 82574
rect 297502 82338 297586 82574
rect 297822 82338 297854 82574
rect 297234 46894 297854 82338
rect 297234 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 297854 46894
rect 297234 46574 297854 46658
rect 297234 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 297854 46574
rect 295931 13700 295997 13701
rect 295931 13636 295932 13700
rect 295996 13636 295997 13700
rect 295931 13635 295997 13636
rect 293514 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 294134 7174
rect 293514 6854 294134 6938
rect 293514 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 294134 6854
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 290595 3500 290661 3501
rect 290595 3436 290596 3500
rect 290660 3436 290661 3500
rect 290595 3435 290661 3436
rect 291699 3500 291765 3501
rect 291699 3436 291700 3500
rect 291764 3436 291765 3500
rect 291699 3435 291765 3436
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -1894 290414 -902
rect 293514 -2266 294134 6618
rect 293514 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 294134 -2266
rect 293514 -2586 294134 -2502
rect 293514 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 294134 -2586
rect 293514 -3814 294134 -2822
rect 297234 10894 297854 46338
rect 299614 13157 299674 188395
rect 300954 158614 301574 194058
rect 307794 345454 308414 375600
rect 307794 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 308414 345454
rect 307794 345134 308414 345218
rect 307794 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 308414 345134
rect 307794 309454 308414 344898
rect 307794 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 308414 309454
rect 307794 309134 308414 309218
rect 307794 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 308414 309134
rect 307794 273454 308414 308898
rect 307794 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 308414 273454
rect 307794 273134 308414 273218
rect 307794 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 308414 273134
rect 307794 237454 308414 272898
rect 307794 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 308414 237454
rect 307794 237134 308414 237218
rect 307794 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 308414 237134
rect 307794 201454 308414 236898
rect 307794 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 308414 201454
rect 307794 201134 308414 201218
rect 307794 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 308414 201134
rect 303659 187100 303725 187101
rect 303659 187036 303660 187100
rect 303724 187036 303725 187100
rect 303659 187035 303725 187036
rect 300954 158378 300986 158614
rect 301222 158378 301306 158614
rect 301542 158378 301574 158614
rect 300954 158294 301574 158378
rect 300954 158058 300986 158294
rect 301222 158058 301306 158294
rect 301542 158058 301574 158294
rect 300954 122614 301574 158058
rect 303662 140861 303722 187035
rect 307794 165454 308414 200898
rect 307794 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 308414 165454
rect 307794 165134 308414 165218
rect 307794 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 308414 165134
rect 303659 140860 303725 140861
rect 303659 140796 303660 140860
rect 303724 140796 303725 140860
rect 303659 140795 303725 140796
rect 300954 122378 300986 122614
rect 301222 122378 301306 122614
rect 301542 122378 301574 122614
rect 300954 122294 301574 122378
rect 300954 122058 300986 122294
rect 301222 122058 301306 122294
rect 301542 122058 301574 122294
rect 300954 86614 301574 122058
rect 300954 86378 300986 86614
rect 301222 86378 301306 86614
rect 301542 86378 301574 86614
rect 300954 86294 301574 86378
rect 300954 86058 300986 86294
rect 301222 86058 301306 86294
rect 301542 86058 301574 86294
rect 300954 50614 301574 86058
rect 300954 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 301574 50614
rect 300954 50294 301574 50378
rect 300954 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 301574 50294
rect 300954 14614 301574 50058
rect 300954 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 301574 14614
rect 300954 14294 301574 14378
rect 300954 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 301574 14294
rect 299611 13156 299677 13157
rect 299611 13092 299612 13156
rect 299676 13092 299677 13156
rect 299611 13091 299677 13092
rect 297234 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 297854 10894
rect 297234 10574 297854 10658
rect 297234 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 297854 10574
rect 297234 -4186 297854 10338
rect 299614 3501 299674 13091
rect 299611 3500 299677 3501
rect 299611 3436 299612 3500
rect 299676 3436 299677 3500
rect 299611 3435 299677 3436
rect 297234 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 297854 -4186
rect 297234 -4506 297854 -4422
rect 297234 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 297854 -4506
rect 297234 -5734 297854 -4742
rect 282954 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 283574 -7066
rect 282954 -7386 283574 -7302
rect 282954 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 283574 -7386
rect 282954 -7654 283574 -7622
rect 300954 -6106 301574 14058
rect 307794 129454 308414 164898
rect 307794 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 308414 129454
rect 307794 129134 308414 129218
rect 307794 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 308414 129134
rect 307794 93454 308414 128898
rect 307794 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 308414 93454
rect 307794 93134 308414 93218
rect 307794 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 308414 93134
rect 307794 57454 308414 92898
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -1306 308414 20898
rect 307794 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 308414 -1306
rect 307794 -1626 308414 -1542
rect 307794 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 308414 -1626
rect 307794 -1894 308414 -1862
rect 311514 349174 312134 375600
rect 311514 348938 311546 349174
rect 311782 348938 311866 349174
rect 312102 348938 312134 349174
rect 311514 348854 312134 348938
rect 311514 348618 311546 348854
rect 311782 348618 311866 348854
rect 312102 348618 312134 348854
rect 311514 313174 312134 348618
rect 311514 312938 311546 313174
rect 311782 312938 311866 313174
rect 312102 312938 312134 313174
rect 311514 312854 312134 312938
rect 311514 312618 311546 312854
rect 311782 312618 311866 312854
rect 312102 312618 312134 312854
rect 311514 277174 312134 312618
rect 311514 276938 311546 277174
rect 311782 276938 311866 277174
rect 312102 276938 312134 277174
rect 311514 276854 312134 276938
rect 311514 276618 311546 276854
rect 311782 276618 311866 276854
rect 312102 276618 312134 276854
rect 311514 241174 312134 276618
rect 311514 240938 311546 241174
rect 311782 240938 311866 241174
rect 312102 240938 312134 241174
rect 311514 240854 312134 240938
rect 311514 240618 311546 240854
rect 311782 240618 311866 240854
rect 312102 240618 312134 240854
rect 311514 205174 312134 240618
rect 311514 204938 311546 205174
rect 311782 204938 311866 205174
rect 312102 204938 312134 205174
rect 311514 204854 312134 204938
rect 311514 204618 311546 204854
rect 311782 204618 311866 204854
rect 312102 204618 312134 204854
rect 311514 169174 312134 204618
rect 311514 168938 311546 169174
rect 311782 168938 311866 169174
rect 312102 168938 312134 169174
rect 311514 168854 312134 168938
rect 311514 168618 311546 168854
rect 311782 168618 311866 168854
rect 312102 168618 312134 168854
rect 311514 133174 312134 168618
rect 311514 132938 311546 133174
rect 311782 132938 311866 133174
rect 312102 132938 312134 133174
rect 311514 132854 312134 132938
rect 311514 132618 311546 132854
rect 311782 132618 311866 132854
rect 312102 132618 312134 132854
rect 311514 97174 312134 132618
rect 311514 96938 311546 97174
rect 311782 96938 311866 97174
rect 312102 96938 312134 97174
rect 311514 96854 312134 96938
rect 311514 96618 311546 96854
rect 311782 96618 311866 96854
rect 312102 96618 312134 96854
rect 311514 61174 312134 96618
rect 311514 60938 311546 61174
rect 311782 60938 311866 61174
rect 312102 60938 312134 61174
rect 311514 60854 312134 60938
rect 311514 60618 311546 60854
rect 311782 60618 311866 60854
rect 312102 60618 312134 60854
rect 311514 25174 312134 60618
rect 311514 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 312134 25174
rect 311514 24854 312134 24938
rect 311514 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 312134 24854
rect 311514 -3226 312134 24618
rect 311514 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 312134 -3226
rect 311514 -3546 312134 -3462
rect 311514 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 312134 -3546
rect 311514 -3814 312134 -3782
rect 315234 352894 315854 375600
rect 315234 352658 315266 352894
rect 315502 352658 315586 352894
rect 315822 352658 315854 352894
rect 315234 352574 315854 352658
rect 315234 352338 315266 352574
rect 315502 352338 315586 352574
rect 315822 352338 315854 352574
rect 315234 316894 315854 352338
rect 315234 316658 315266 316894
rect 315502 316658 315586 316894
rect 315822 316658 315854 316894
rect 315234 316574 315854 316658
rect 315234 316338 315266 316574
rect 315502 316338 315586 316574
rect 315822 316338 315854 316574
rect 315234 280894 315854 316338
rect 315234 280658 315266 280894
rect 315502 280658 315586 280894
rect 315822 280658 315854 280894
rect 315234 280574 315854 280658
rect 315234 280338 315266 280574
rect 315502 280338 315586 280574
rect 315822 280338 315854 280574
rect 315234 244894 315854 280338
rect 315234 244658 315266 244894
rect 315502 244658 315586 244894
rect 315822 244658 315854 244894
rect 315234 244574 315854 244658
rect 315234 244338 315266 244574
rect 315502 244338 315586 244574
rect 315822 244338 315854 244574
rect 315234 208894 315854 244338
rect 315234 208658 315266 208894
rect 315502 208658 315586 208894
rect 315822 208658 315854 208894
rect 315234 208574 315854 208658
rect 315234 208338 315266 208574
rect 315502 208338 315586 208574
rect 315822 208338 315854 208574
rect 315234 172894 315854 208338
rect 315234 172658 315266 172894
rect 315502 172658 315586 172894
rect 315822 172658 315854 172894
rect 315234 172574 315854 172658
rect 315234 172338 315266 172574
rect 315502 172338 315586 172574
rect 315822 172338 315854 172574
rect 315234 136894 315854 172338
rect 315234 136658 315266 136894
rect 315502 136658 315586 136894
rect 315822 136658 315854 136894
rect 315234 136574 315854 136658
rect 315234 136338 315266 136574
rect 315502 136338 315586 136574
rect 315822 136338 315854 136574
rect 315234 100894 315854 136338
rect 315234 100658 315266 100894
rect 315502 100658 315586 100894
rect 315822 100658 315854 100894
rect 315234 100574 315854 100658
rect 315234 100338 315266 100574
rect 315502 100338 315586 100574
rect 315822 100338 315854 100574
rect 315234 64894 315854 100338
rect 315234 64658 315266 64894
rect 315502 64658 315586 64894
rect 315822 64658 315854 64894
rect 315234 64574 315854 64658
rect 315234 64338 315266 64574
rect 315502 64338 315586 64574
rect 315822 64338 315854 64574
rect 315234 28894 315854 64338
rect 315234 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 315854 28894
rect 315234 28574 315854 28658
rect 315234 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 315854 28574
rect 315234 -5146 315854 28338
rect 315234 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 315854 -5146
rect 315234 -5466 315854 -5382
rect 315234 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 315854 -5466
rect 315234 -5734 315854 -5702
rect 318954 356614 319574 375600
rect 318954 356378 318986 356614
rect 319222 356378 319306 356614
rect 319542 356378 319574 356614
rect 318954 356294 319574 356378
rect 318954 356058 318986 356294
rect 319222 356058 319306 356294
rect 319542 356058 319574 356294
rect 318954 320614 319574 356058
rect 318954 320378 318986 320614
rect 319222 320378 319306 320614
rect 319542 320378 319574 320614
rect 318954 320294 319574 320378
rect 318954 320058 318986 320294
rect 319222 320058 319306 320294
rect 319542 320058 319574 320294
rect 318954 284614 319574 320058
rect 318954 284378 318986 284614
rect 319222 284378 319306 284614
rect 319542 284378 319574 284614
rect 318954 284294 319574 284378
rect 318954 284058 318986 284294
rect 319222 284058 319306 284294
rect 319542 284058 319574 284294
rect 318954 248614 319574 284058
rect 318954 248378 318986 248614
rect 319222 248378 319306 248614
rect 319542 248378 319574 248614
rect 318954 248294 319574 248378
rect 318954 248058 318986 248294
rect 319222 248058 319306 248294
rect 319542 248058 319574 248294
rect 318954 212614 319574 248058
rect 318954 212378 318986 212614
rect 319222 212378 319306 212614
rect 319542 212378 319574 212614
rect 318954 212294 319574 212378
rect 318954 212058 318986 212294
rect 319222 212058 319306 212294
rect 319542 212058 319574 212294
rect 318954 176614 319574 212058
rect 318954 176378 318986 176614
rect 319222 176378 319306 176614
rect 319542 176378 319574 176614
rect 318954 176294 319574 176378
rect 318954 176058 318986 176294
rect 319222 176058 319306 176294
rect 319542 176058 319574 176294
rect 318954 140614 319574 176058
rect 318954 140378 318986 140614
rect 319222 140378 319306 140614
rect 319542 140378 319574 140614
rect 318954 140294 319574 140378
rect 318954 140058 318986 140294
rect 319222 140058 319306 140294
rect 319542 140058 319574 140294
rect 318954 104614 319574 140058
rect 318954 104378 318986 104614
rect 319222 104378 319306 104614
rect 319542 104378 319574 104614
rect 318954 104294 319574 104378
rect 318954 104058 318986 104294
rect 319222 104058 319306 104294
rect 319542 104058 319574 104294
rect 318954 68614 319574 104058
rect 318954 68378 318986 68614
rect 319222 68378 319306 68614
rect 319542 68378 319574 68614
rect 318954 68294 319574 68378
rect 318954 68058 318986 68294
rect 319222 68058 319306 68294
rect 319542 68058 319574 68294
rect 318954 32614 319574 68058
rect 318954 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 319574 32614
rect 318954 32294 319574 32378
rect 318954 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 319574 32294
rect 300954 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 301574 -6106
rect 300954 -6426 301574 -6342
rect 300954 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 301574 -6426
rect 300954 -7654 301574 -6662
rect 318954 -7066 319574 32058
rect 325794 363454 326414 375600
rect 325794 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 326414 363454
rect 325794 363134 326414 363218
rect 325794 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 326414 363134
rect 325794 327454 326414 362898
rect 325794 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 326414 327454
rect 325794 327134 326414 327218
rect 325794 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 326414 327134
rect 325794 291454 326414 326898
rect 325794 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 326414 291454
rect 325794 291134 326414 291218
rect 325794 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 326414 291134
rect 325794 255454 326414 290898
rect 325794 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 326414 255454
rect 325794 255134 326414 255218
rect 325794 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 326414 255134
rect 325794 219454 326414 254898
rect 325794 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 326414 219454
rect 325794 219134 326414 219218
rect 325794 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 326414 219134
rect 325794 183454 326414 218898
rect 325794 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 326414 183454
rect 325794 183134 326414 183218
rect 325794 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 326414 183134
rect 325794 147454 326414 182898
rect 325794 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 326414 147454
rect 325794 147134 326414 147218
rect 325794 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 326414 147134
rect 325794 111454 326414 146898
rect 325794 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 326414 111454
rect 325794 111134 326414 111218
rect 325794 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 326414 111134
rect 325794 75454 326414 110898
rect 325794 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 326414 75454
rect 325794 75134 326414 75218
rect 325794 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 326414 75134
rect 325794 39454 326414 74898
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -1894 326414 -902
rect 329514 367174 330134 375600
rect 329514 366938 329546 367174
rect 329782 366938 329866 367174
rect 330102 366938 330134 367174
rect 329514 366854 330134 366938
rect 329514 366618 329546 366854
rect 329782 366618 329866 366854
rect 330102 366618 330134 366854
rect 329514 331174 330134 366618
rect 329514 330938 329546 331174
rect 329782 330938 329866 331174
rect 330102 330938 330134 331174
rect 329514 330854 330134 330938
rect 329514 330618 329546 330854
rect 329782 330618 329866 330854
rect 330102 330618 330134 330854
rect 329514 295174 330134 330618
rect 329514 294938 329546 295174
rect 329782 294938 329866 295174
rect 330102 294938 330134 295174
rect 329514 294854 330134 294938
rect 329514 294618 329546 294854
rect 329782 294618 329866 294854
rect 330102 294618 330134 294854
rect 329514 259174 330134 294618
rect 329514 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 330134 259174
rect 329514 258854 330134 258938
rect 329514 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 330134 258854
rect 329514 223174 330134 258618
rect 329514 222938 329546 223174
rect 329782 222938 329866 223174
rect 330102 222938 330134 223174
rect 329514 222854 330134 222938
rect 329514 222618 329546 222854
rect 329782 222618 329866 222854
rect 330102 222618 330134 222854
rect 329514 187174 330134 222618
rect 329514 186938 329546 187174
rect 329782 186938 329866 187174
rect 330102 186938 330134 187174
rect 329514 186854 330134 186938
rect 329514 186618 329546 186854
rect 329782 186618 329866 186854
rect 330102 186618 330134 186854
rect 329514 151174 330134 186618
rect 329514 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 330134 151174
rect 329514 150854 330134 150938
rect 329514 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 330134 150854
rect 329514 115174 330134 150618
rect 329514 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 330134 115174
rect 329514 114854 330134 114938
rect 329514 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 330134 114854
rect 329514 79174 330134 114618
rect 329514 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 330134 79174
rect 329514 78854 330134 78938
rect 329514 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 330134 78854
rect 329514 43174 330134 78618
rect 329514 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 330134 43174
rect 329514 42854 330134 42938
rect 329514 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 330134 42854
rect 329514 7174 330134 42618
rect 329514 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 330134 7174
rect 329514 6854 330134 6938
rect 329514 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 330134 6854
rect 329514 -2266 330134 6618
rect 329514 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 330134 -2266
rect 329514 -2586 330134 -2502
rect 329514 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 330134 -2586
rect 329514 -3814 330134 -2822
rect 333234 370894 333854 375600
rect 333234 370658 333266 370894
rect 333502 370658 333586 370894
rect 333822 370658 333854 370894
rect 333234 370574 333854 370658
rect 333234 370338 333266 370574
rect 333502 370338 333586 370574
rect 333822 370338 333854 370574
rect 333234 334894 333854 370338
rect 333234 334658 333266 334894
rect 333502 334658 333586 334894
rect 333822 334658 333854 334894
rect 333234 334574 333854 334658
rect 333234 334338 333266 334574
rect 333502 334338 333586 334574
rect 333822 334338 333854 334574
rect 333234 298894 333854 334338
rect 333234 298658 333266 298894
rect 333502 298658 333586 298894
rect 333822 298658 333854 298894
rect 333234 298574 333854 298658
rect 333234 298338 333266 298574
rect 333502 298338 333586 298574
rect 333822 298338 333854 298574
rect 333234 262894 333854 298338
rect 333234 262658 333266 262894
rect 333502 262658 333586 262894
rect 333822 262658 333854 262894
rect 333234 262574 333854 262658
rect 333234 262338 333266 262574
rect 333502 262338 333586 262574
rect 333822 262338 333854 262574
rect 333234 226894 333854 262338
rect 333234 226658 333266 226894
rect 333502 226658 333586 226894
rect 333822 226658 333854 226894
rect 333234 226574 333854 226658
rect 333234 226338 333266 226574
rect 333502 226338 333586 226574
rect 333822 226338 333854 226574
rect 333234 190894 333854 226338
rect 333234 190658 333266 190894
rect 333502 190658 333586 190894
rect 333822 190658 333854 190894
rect 333234 190574 333854 190658
rect 333234 190338 333266 190574
rect 333502 190338 333586 190574
rect 333822 190338 333854 190574
rect 333234 154894 333854 190338
rect 333234 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 333854 154894
rect 333234 154574 333854 154658
rect 333234 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 333854 154574
rect 333234 118894 333854 154338
rect 333234 118658 333266 118894
rect 333502 118658 333586 118894
rect 333822 118658 333854 118894
rect 333234 118574 333854 118658
rect 333234 118338 333266 118574
rect 333502 118338 333586 118574
rect 333822 118338 333854 118574
rect 333234 82894 333854 118338
rect 333234 82658 333266 82894
rect 333502 82658 333586 82894
rect 333822 82658 333854 82894
rect 333234 82574 333854 82658
rect 333234 82338 333266 82574
rect 333502 82338 333586 82574
rect 333822 82338 333854 82574
rect 333234 46894 333854 82338
rect 333234 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 333854 46894
rect 333234 46574 333854 46658
rect 333234 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 333854 46574
rect 333234 10894 333854 46338
rect 333234 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 333854 10894
rect 333234 10574 333854 10658
rect 333234 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 333854 10574
rect 333234 -4186 333854 10338
rect 333234 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 333854 -4186
rect 333234 -4506 333854 -4422
rect 333234 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 333854 -4506
rect 333234 -5734 333854 -4742
rect 336954 374614 337574 375600
rect 336954 374378 336986 374614
rect 337222 374378 337306 374614
rect 337542 374378 337574 374614
rect 336954 374294 337574 374378
rect 336954 374058 336986 374294
rect 337222 374058 337306 374294
rect 337542 374058 337574 374294
rect 336954 338614 337574 374058
rect 336954 338378 336986 338614
rect 337222 338378 337306 338614
rect 337542 338378 337574 338614
rect 336954 338294 337574 338378
rect 336954 338058 336986 338294
rect 337222 338058 337306 338294
rect 337542 338058 337574 338294
rect 336954 302614 337574 338058
rect 336954 302378 336986 302614
rect 337222 302378 337306 302614
rect 337542 302378 337574 302614
rect 336954 302294 337574 302378
rect 336954 302058 336986 302294
rect 337222 302058 337306 302294
rect 337542 302058 337574 302294
rect 336954 266614 337574 302058
rect 336954 266378 336986 266614
rect 337222 266378 337306 266614
rect 337542 266378 337574 266614
rect 336954 266294 337574 266378
rect 336954 266058 336986 266294
rect 337222 266058 337306 266294
rect 337542 266058 337574 266294
rect 336954 230614 337574 266058
rect 336954 230378 336986 230614
rect 337222 230378 337306 230614
rect 337542 230378 337574 230614
rect 336954 230294 337574 230378
rect 336954 230058 336986 230294
rect 337222 230058 337306 230294
rect 337542 230058 337574 230294
rect 336954 194614 337574 230058
rect 336954 194378 336986 194614
rect 337222 194378 337306 194614
rect 337542 194378 337574 194614
rect 336954 194294 337574 194378
rect 336954 194058 336986 194294
rect 337222 194058 337306 194294
rect 337542 194058 337574 194294
rect 336954 158614 337574 194058
rect 336954 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 337574 158614
rect 336954 158294 337574 158378
rect 336954 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 337574 158294
rect 336954 122614 337574 158058
rect 336954 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 337574 122614
rect 336954 122294 337574 122378
rect 336954 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 337574 122294
rect 336954 86614 337574 122058
rect 336954 86378 336986 86614
rect 337222 86378 337306 86614
rect 337542 86378 337574 86614
rect 336954 86294 337574 86378
rect 336954 86058 336986 86294
rect 337222 86058 337306 86294
rect 337542 86058 337574 86294
rect 336954 50614 337574 86058
rect 336954 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 337574 50614
rect 336954 50294 337574 50378
rect 336954 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 337574 50294
rect 336954 14614 337574 50058
rect 336954 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 337574 14614
rect 336954 14294 337574 14378
rect 336954 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 337574 14294
rect 318954 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 319574 -7066
rect 318954 -7386 319574 -7302
rect 318954 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 319574 -7386
rect 318954 -7654 319574 -7622
rect 336954 -6106 337574 14058
rect 343794 345454 344414 375600
rect 343794 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 344414 345454
rect 343794 345134 344414 345218
rect 343794 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 344414 345134
rect 343794 309454 344414 344898
rect 343794 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 344414 309454
rect 343794 309134 344414 309218
rect 343794 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 344414 309134
rect 343794 273454 344414 308898
rect 343794 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 344414 273454
rect 343794 273134 344414 273218
rect 343794 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 344414 273134
rect 343794 237454 344414 272898
rect 343794 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 344414 237454
rect 343794 237134 344414 237218
rect 343794 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 344414 237134
rect 343794 201454 344414 236898
rect 343794 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 344414 201454
rect 343794 201134 344414 201218
rect 343794 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 344414 201134
rect 343794 165454 344414 200898
rect 343794 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 344414 165454
rect 343794 165134 344414 165218
rect 343794 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 344414 165134
rect 343794 129454 344414 164898
rect 343794 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 344414 129454
rect 343794 129134 344414 129218
rect 343794 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 344414 129134
rect 343794 93454 344414 128898
rect 343794 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 344414 93454
rect 343794 93134 344414 93218
rect 343794 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 344414 93134
rect 343794 57454 344414 92898
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -1306 344414 20898
rect 343794 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 344414 -1306
rect 343794 -1626 344414 -1542
rect 343794 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 344414 -1626
rect 343794 -1894 344414 -1862
rect 347514 349174 348134 375600
rect 347514 348938 347546 349174
rect 347782 348938 347866 349174
rect 348102 348938 348134 349174
rect 347514 348854 348134 348938
rect 347514 348618 347546 348854
rect 347782 348618 347866 348854
rect 348102 348618 348134 348854
rect 347514 313174 348134 348618
rect 347514 312938 347546 313174
rect 347782 312938 347866 313174
rect 348102 312938 348134 313174
rect 347514 312854 348134 312938
rect 347514 312618 347546 312854
rect 347782 312618 347866 312854
rect 348102 312618 348134 312854
rect 347514 277174 348134 312618
rect 347514 276938 347546 277174
rect 347782 276938 347866 277174
rect 348102 276938 348134 277174
rect 347514 276854 348134 276938
rect 347514 276618 347546 276854
rect 347782 276618 347866 276854
rect 348102 276618 348134 276854
rect 347514 241174 348134 276618
rect 347514 240938 347546 241174
rect 347782 240938 347866 241174
rect 348102 240938 348134 241174
rect 347514 240854 348134 240938
rect 347514 240618 347546 240854
rect 347782 240618 347866 240854
rect 348102 240618 348134 240854
rect 347514 205174 348134 240618
rect 347514 204938 347546 205174
rect 347782 204938 347866 205174
rect 348102 204938 348134 205174
rect 347514 204854 348134 204938
rect 347514 204618 347546 204854
rect 347782 204618 347866 204854
rect 348102 204618 348134 204854
rect 347514 169174 348134 204618
rect 347514 168938 347546 169174
rect 347782 168938 347866 169174
rect 348102 168938 348134 169174
rect 347514 168854 348134 168938
rect 347514 168618 347546 168854
rect 347782 168618 347866 168854
rect 348102 168618 348134 168854
rect 347514 133174 348134 168618
rect 347514 132938 347546 133174
rect 347782 132938 347866 133174
rect 348102 132938 348134 133174
rect 347514 132854 348134 132938
rect 347514 132618 347546 132854
rect 347782 132618 347866 132854
rect 348102 132618 348134 132854
rect 347514 97174 348134 132618
rect 347514 96938 347546 97174
rect 347782 96938 347866 97174
rect 348102 96938 348134 97174
rect 347514 96854 348134 96938
rect 347514 96618 347546 96854
rect 347782 96618 347866 96854
rect 348102 96618 348134 96854
rect 347514 61174 348134 96618
rect 347514 60938 347546 61174
rect 347782 60938 347866 61174
rect 348102 60938 348134 61174
rect 347514 60854 348134 60938
rect 347514 60618 347546 60854
rect 347782 60618 347866 60854
rect 348102 60618 348134 60854
rect 347514 25174 348134 60618
rect 347514 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 348134 25174
rect 347514 24854 348134 24938
rect 347514 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 348134 24854
rect 347514 -3226 348134 24618
rect 347514 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 348134 -3226
rect 347514 -3546 348134 -3462
rect 347514 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 348134 -3546
rect 347514 -3814 348134 -3782
rect 351234 352894 351854 375600
rect 353342 358053 353402 541315
rect 354954 537993 355574 572058
rect 361794 704838 362414 705830
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 358859 546548 358925 546549
rect 358859 546484 358860 546548
rect 358924 546484 358925 546548
rect 358859 546483 358925 546484
rect 356099 499900 356165 499901
rect 356099 499836 356100 499900
rect 356164 499836 356165 499900
rect 356099 499835 356165 499836
rect 356102 476130 356162 499835
rect 356102 476070 356530 476130
rect 356283 467940 356349 467941
rect 356283 467876 356284 467940
rect 356348 467876 356349 467940
rect 356283 467875 356349 467876
rect 356286 467530 356346 467875
rect 354814 467470 356346 467530
rect 354814 463710 354874 467470
rect 356470 466470 356530 476070
rect 356651 475556 356717 475557
rect 356651 475492 356652 475556
rect 356716 475492 356717 475556
rect 356651 475491 356717 475492
rect 354446 463650 354874 463710
rect 356102 466410 356530 466470
rect 354446 361045 354506 463650
rect 354443 361044 354509 361045
rect 354443 360980 354444 361044
rect 354508 360980 354509 361044
rect 354443 360979 354509 360980
rect 353339 358052 353405 358053
rect 353339 357988 353340 358052
rect 353404 357988 353405 358052
rect 353339 357987 353405 357988
rect 351234 352658 351266 352894
rect 351502 352658 351586 352894
rect 351822 352658 351854 352894
rect 351234 352574 351854 352658
rect 351234 352338 351266 352574
rect 351502 352338 351586 352574
rect 351822 352338 351854 352574
rect 351234 316894 351854 352338
rect 351234 316658 351266 316894
rect 351502 316658 351586 316894
rect 351822 316658 351854 316894
rect 351234 316574 351854 316658
rect 351234 316338 351266 316574
rect 351502 316338 351586 316574
rect 351822 316338 351854 316574
rect 351234 280894 351854 316338
rect 351234 280658 351266 280894
rect 351502 280658 351586 280894
rect 351822 280658 351854 280894
rect 351234 280574 351854 280658
rect 351234 280338 351266 280574
rect 351502 280338 351586 280574
rect 351822 280338 351854 280574
rect 351234 244894 351854 280338
rect 351234 244658 351266 244894
rect 351502 244658 351586 244894
rect 351822 244658 351854 244894
rect 351234 244574 351854 244658
rect 351234 244338 351266 244574
rect 351502 244338 351586 244574
rect 351822 244338 351854 244574
rect 351234 208894 351854 244338
rect 351234 208658 351266 208894
rect 351502 208658 351586 208894
rect 351822 208658 351854 208894
rect 351234 208574 351854 208658
rect 351234 208338 351266 208574
rect 351502 208338 351586 208574
rect 351822 208338 351854 208574
rect 351234 172894 351854 208338
rect 351234 172658 351266 172894
rect 351502 172658 351586 172894
rect 351822 172658 351854 172894
rect 351234 172574 351854 172658
rect 351234 172338 351266 172574
rect 351502 172338 351586 172574
rect 351822 172338 351854 172574
rect 351234 136894 351854 172338
rect 351234 136658 351266 136894
rect 351502 136658 351586 136894
rect 351822 136658 351854 136894
rect 351234 136574 351854 136658
rect 351234 136338 351266 136574
rect 351502 136338 351586 136574
rect 351822 136338 351854 136574
rect 351234 100894 351854 136338
rect 351234 100658 351266 100894
rect 351502 100658 351586 100894
rect 351822 100658 351854 100894
rect 351234 100574 351854 100658
rect 351234 100338 351266 100574
rect 351502 100338 351586 100574
rect 351822 100338 351854 100574
rect 351234 64894 351854 100338
rect 351234 64658 351266 64894
rect 351502 64658 351586 64894
rect 351822 64658 351854 64894
rect 351234 64574 351854 64658
rect 351234 64338 351266 64574
rect 351502 64338 351586 64574
rect 351822 64338 351854 64574
rect 351234 28894 351854 64338
rect 351234 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 351854 28894
rect 351234 28574 351854 28658
rect 351234 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 351854 28574
rect 351234 -5146 351854 28338
rect 351234 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 351854 -5146
rect 351234 -5466 351854 -5382
rect 351234 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 351854 -5466
rect 351234 -5734 351854 -5702
rect 354954 356614 355574 375600
rect 356102 359413 356162 466410
rect 356654 451290 356714 475491
rect 356286 451230 356714 451290
rect 356286 360909 356346 451230
rect 358862 375189 358922 546483
rect 361794 543454 362414 578898
rect 361794 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 362414 543454
rect 361794 543134 362414 543218
rect 361794 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 362414 543134
rect 361794 507454 362414 542898
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 361619 487252 361685 487253
rect 361619 487188 361620 487252
rect 361684 487188 361685 487252
rect 361619 487187 361685 487188
rect 358859 375188 358925 375189
rect 358859 375124 358860 375188
rect 358924 375124 358925 375188
rect 358859 375123 358925 375124
rect 356283 360908 356349 360909
rect 356283 360844 356284 360908
rect 356348 360844 356349 360908
rect 356283 360843 356349 360844
rect 356099 359412 356165 359413
rect 356099 359348 356100 359412
rect 356164 359348 356165 359412
rect 356099 359347 356165 359348
rect 354954 356378 354986 356614
rect 355222 356378 355306 356614
rect 355542 356378 355574 356614
rect 354954 356294 355574 356378
rect 354954 356058 354986 356294
rect 355222 356058 355306 356294
rect 355542 356058 355574 356294
rect 354954 320614 355574 356058
rect 354954 320378 354986 320614
rect 355222 320378 355306 320614
rect 355542 320378 355574 320614
rect 354954 320294 355574 320378
rect 354954 320058 354986 320294
rect 355222 320058 355306 320294
rect 355542 320058 355574 320294
rect 354954 284614 355574 320058
rect 354954 284378 354986 284614
rect 355222 284378 355306 284614
rect 355542 284378 355574 284614
rect 354954 284294 355574 284378
rect 354954 284058 354986 284294
rect 355222 284058 355306 284294
rect 355542 284058 355574 284294
rect 354954 248614 355574 284058
rect 354954 248378 354986 248614
rect 355222 248378 355306 248614
rect 355542 248378 355574 248614
rect 354954 248294 355574 248378
rect 354954 248058 354986 248294
rect 355222 248058 355306 248294
rect 355542 248058 355574 248294
rect 354954 212614 355574 248058
rect 354954 212378 354986 212614
rect 355222 212378 355306 212614
rect 355542 212378 355574 212614
rect 354954 212294 355574 212378
rect 354954 212058 354986 212294
rect 355222 212058 355306 212294
rect 355542 212058 355574 212294
rect 354954 176614 355574 212058
rect 354954 176378 354986 176614
rect 355222 176378 355306 176614
rect 355542 176378 355574 176614
rect 354954 176294 355574 176378
rect 354954 176058 354986 176294
rect 355222 176058 355306 176294
rect 355542 176058 355574 176294
rect 354954 140614 355574 176058
rect 354954 140378 354986 140614
rect 355222 140378 355306 140614
rect 355542 140378 355574 140614
rect 354954 140294 355574 140378
rect 354954 140058 354986 140294
rect 355222 140058 355306 140294
rect 355542 140058 355574 140294
rect 354954 104614 355574 140058
rect 361622 117197 361682 487187
rect 361794 471454 362414 506898
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 361794 435454 362414 470898
rect 361794 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 362414 435454
rect 361794 435134 362414 435218
rect 361794 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 362414 435134
rect 361794 399454 362414 434898
rect 361794 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 362414 399454
rect 361794 399134 362414 399218
rect 361794 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 362414 399134
rect 361794 363454 362414 398898
rect 361794 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 362414 363454
rect 361794 363134 362414 363218
rect 361794 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 362414 363134
rect 361794 327454 362414 362898
rect 361794 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 362414 327454
rect 361794 327134 362414 327218
rect 361794 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 362414 327134
rect 361794 291454 362414 326898
rect 361794 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 362414 291454
rect 361794 291134 362414 291218
rect 361794 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 362414 291134
rect 361794 255454 362414 290898
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 361794 219454 362414 254898
rect 361794 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 362414 219454
rect 361794 219134 362414 219218
rect 361794 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 362414 219134
rect 361794 183454 362414 218898
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 361794 147454 362414 182898
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 361619 117196 361685 117197
rect 361619 117132 361620 117196
rect 361684 117132 361685 117196
rect 361619 117131 361685 117132
rect 354954 104378 354986 104614
rect 355222 104378 355306 104614
rect 355542 104378 355574 104614
rect 354954 104294 355574 104378
rect 354954 104058 354986 104294
rect 355222 104058 355306 104294
rect 355542 104058 355574 104294
rect 354954 68614 355574 104058
rect 354954 68378 354986 68614
rect 355222 68378 355306 68614
rect 355542 68378 355574 68614
rect 354954 68294 355574 68378
rect 354954 68058 354986 68294
rect 355222 68058 355306 68294
rect 355542 68058 355574 68294
rect 354954 32614 355574 68058
rect 354954 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 355574 32614
rect 354954 32294 355574 32378
rect 354954 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 355574 32294
rect 336954 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 337574 -6106
rect 336954 -6426 337574 -6342
rect 336954 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 337574 -6426
rect 336954 -7654 337574 -6662
rect 354954 -7066 355574 32058
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -1894 362414 -902
rect 365514 691174 366134 706202
rect 365514 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 366134 691174
rect 365514 690854 366134 690938
rect 365514 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 366134 690854
rect 365514 655174 366134 690618
rect 365514 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 366134 655174
rect 365514 654854 366134 654938
rect 365514 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 366134 654854
rect 365514 619174 366134 654618
rect 365514 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 366134 619174
rect 365514 618854 366134 618938
rect 365514 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 366134 618854
rect 365514 583174 366134 618618
rect 365514 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 366134 583174
rect 365514 582854 366134 582938
rect 365514 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 366134 582854
rect 365514 547174 366134 582618
rect 365514 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 366134 547174
rect 365514 546854 366134 546938
rect 365514 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 366134 546854
rect 365514 511174 366134 546618
rect 365514 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 366134 511174
rect 365514 510854 366134 510938
rect 365514 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 366134 510854
rect 365514 475174 366134 510618
rect 365514 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 366134 475174
rect 365514 474854 366134 474938
rect 365514 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 366134 474854
rect 365514 439174 366134 474618
rect 365514 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 366134 439174
rect 365514 438854 366134 438938
rect 365514 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 366134 438854
rect 365514 403174 366134 438618
rect 365514 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 366134 403174
rect 365514 402854 366134 402938
rect 365514 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 366134 402854
rect 365514 367174 366134 402618
rect 365514 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 366134 367174
rect 365514 366854 366134 366938
rect 365514 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 366134 366854
rect 365514 331174 366134 366618
rect 365514 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 366134 331174
rect 365514 330854 366134 330938
rect 365514 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 366134 330854
rect 365514 295174 366134 330618
rect 365514 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 366134 295174
rect 365514 294854 366134 294938
rect 365514 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 366134 294854
rect 365514 259174 366134 294618
rect 365514 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 366134 259174
rect 365514 258854 366134 258938
rect 365514 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 366134 258854
rect 365514 223174 366134 258618
rect 365514 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 366134 223174
rect 365514 222854 366134 222938
rect 365514 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 366134 222854
rect 365514 187174 366134 222618
rect 365514 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 366134 187174
rect 365514 186854 366134 186938
rect 365514 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 366134 186854
rect 365514 151174 366134 186618
rect 365514 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 366134 151174
rect 365514 150854 366134 150938
rect 365514 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 366134 150854
rect 365514 115174 366134 150618
rect 365514 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 366134 115174
rect 365514 114854 366134 114938
rect 365514 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 366134 114854
rect 365514 79174 366134 114618
rect 365514 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 366134 79174
rect 365514 78854 366134 78938
rect 365514 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 366134 78854
rect 365514 43174 366134 78618
rect 365514 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 366134 43174
rect 365514 42854 366134 42938
rect 365514 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 366134 42854
rect 365514 7174 366134 42618
rect 365514 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 366134 7174
rect 365514 6854 366134 6938
rect 365514 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 366134 6854
rect 365514 -2266 366134 6618
rect 365514 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 366134 -2266
rect 365514 -2586 366134 -2502
rect 365514 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 366134 -2586
rect 365514 -3814 366134 -2822
rect 369234 694894 369854 708122
rect 369234 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 369854 694894
rect 369234 694574 369854 694658
rect 369234 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 369854 694574
rect 369234 658894 369854 694338
rect 369234 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 369854 658894
rect 369234 658574 369854 658658
rect 369234 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 369854 658574
rect 369234 622894 369854 658338
rect 369234 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 369854 622894
rect 369234 622574 369854 622658
rect 369234 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 369854 622574
rect 369234 586894 369854 622338
rect 369234 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 369854 586894
rect 369234 586574 369854 586658
rect 369234 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 369854 586574
rect 369234 550894 369854 586338
rect 369234 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 369854 550894
rect 369234 550574 369854 550658
rect 369234 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 369854 550574
rect 369234 514894 369854 550338
rect 369234 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 369854 514894
rect 369234 514574 369854 514658
rect 369234 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 369854 514574
rect 369234 478894 369854 514338
rect 369234 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 369854 478894
rect 369234 478574 369854 478658
rect 369234 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 369854 478574
rect 369234 442894 369854 478338
rect 369234 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 369854 442894
rect 369234 442574 369854 442658
rect 369234 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 369854 442574
rect 369234 406894 369854 442338
rect 369234 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 369854 406894
rect 369234 406574 369854 406658
rect 369234 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 369854 406574
rect 369234 370894 369854 406338
rect 369234 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 369854 370894
rect 369234 370574 369854 370658
rect 369234 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 369854 370574
rect 369234 334894 369854 370338
rect 369234 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 369854 334894
rect 369234 334574 369854 334658
rect 369234 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 369854 334574
rect 369234 298894 369854 334338
rect 369234 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 369854 298894
rect 369234 298574 369854 298658
rect 369234 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 369854 298574
rect 369234 262894 369854 298338
rect 369234 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 369854 262894
rect 369234 262574 369854 262658
rect 369234 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 369854 262574
rect 369234 226894 369854 262338
rect 369234 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 369854 226894
rect 369234 226574 369854 226658
rect 369234 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 369854 226574
rect 369234 190894 369854 226338
rect 369234 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 369854 190894
rect 369234 190574 369854 190658
rect 369234 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 369854 190574
rect 369234 154894 369854 190338
rect 369234 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 369854 154894
rect 369234 154574 369854 154658
rect 369234 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 369854 154574
rect 369234 118894 369854 154338
rect 369234 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 369854 118894
rect 369234 118574 369854 118658
rect 369234 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 369854 118574
rect 369234 82894 369854 118338
rect 369234 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 369854 82894
rect 369234 82574 369854 82658
rect 369234 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 369854 82574
rect 369234 46894 369854 82338
rect 369234 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 369854 46894
rect 369234 46574 369854 46658
rect 369234 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 369854 46574
rect 369234 10894 369854 46338
rect 369234 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 369854 10894
rect 369234 10574 369854 10658
rect 369234 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 369854 10574
rect 369234 -4186 369854 10338
rect 369234 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 369854 -4186
rect 369234 -4506 369854 -4422
rect 369234 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 369854 -4506
rect 369234 -5734 369854 -4742
rect 372954 698614 373574 710042
rect 390954 711558 391574 711590
rect 390954 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 391574 711558
rect 390954 711238 391574 711322
rect 390954 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 391574 711238
rect 387234 709638 387854 709670
rect 387234 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 387854 709638
rect 387234 709318 387854 709402
rect 387234 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 387854 709318
rect 383514 707718 384134 707750
rect 383514 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 384134 707718
rect 383514 707398 384134 707482
rect 383514 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 384134 707398
rect 372954 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 373574 698614
rect 372954 698294 373574 698378
rect 372954 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 373574 698294
rect 372954 662614 373574 698058
rect 372954 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 373574 662614
rect 372954 662294 373574 662378
rect 372954 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 373574 662294
rect 372954 626614 373574 662058
rect 372954 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 373574 626614
rect 372954 626294 373574 626378
rect 372954 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 373574 626294
rect 372954 590614 373574 626058
rect 372954 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 373574 590614
rect 372954 590294 373574 590378
rect 372954 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 373574 590294
rect 372954 554614 373574 590058
rect 372954 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 373574 554614
rect 372954 554294 373574 554378
rect 372954 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 373574 554294
rect 372954 518614 373574 554058
rect 372954 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 373574 518614
rect 372954 518294 373574 518378
rect 372954 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 373574 518294
rect 372954 482614 373574 518058
rect 372954 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 373574 482614
rect 372954 482294 373574 482378
rect 372954 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 373574 482294
rect 372954 446614 373574 482058
rect 372954 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 373574 446614
rect 372954 446294 373574 446378
rect 372954 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 373574 446294
rect 372954 410614 373574 446058
rect 372954 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 373574 410614
rect 372954 410294 373574 410378
rect 372954 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 373574 410294
rect 372954 374614 373574 410058
rect 372954 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 373574 374614
rect 372954 374294 373574 374378
rect 372954 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 373574 374294
rect 372954 338614 373574 374058
rect 372954 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 373574 338614
rect 372954 338294 373574 338378
rect 372954 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 373574 338294
rect 372954 302614 373574 338058
rect 372954 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 373574 302614
rect 372954 302294 373574 302378
rect 372954 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 373574 302294
rect 372954 266614 373574 302058
rect 372954 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 373574 266614
rect 372954 266294 373574 266378
rect 372954 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 373574 266294
rect 372954 230614 373574 266058
rect 372954 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 373574 230614
rect 372954 230294 373574 230378
rect 372954 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 373574 230294
rect 372954 194614 373574 230058
rect 372954 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 373574 194614
rect 372954 194294 373574 194378
rect 372954 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 373574 194294
rect 372954 158614 373574 194058
rect 372954 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 373574 158614
rect 372954 158294 373574 158378
rect 372954 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 373574 158294
rect 372954 122614 373574 158058
rect 372954 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 373574 122614
rect 372954 122294 373574 122378
rect 372954 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 373574 122294
rect 372954 86614 373574 122058
rect 372954 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 373574 86614
rect 372954 86294 373574 86378
rect 372954 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 373574 86294
rect 372954 50614 373574 86058
rect 372954 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 373574 50614
rect 372954 50294 373574 50378
rect 372954 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 373574 50294
rect 372954 14614 373574 50058
rect 372954 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 373574 14614
rect 372954 14294 373574 14378
rect 372954 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 373574 14294
rect 354954 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 355574 -7066
rect 354954 -7386 355574 -7302
rect 354954 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 355574 -7386
rect 354954 -7654 355574 -7622
rect 372954 -6106 373574 14058
rect 379794 705798 380414 705830
rect 379794 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 380414 705798
rect 379794 705478 380414 705562
rect 379794 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 380414 705478
rect 379794 669454 380414 705242
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 633454 380414 668898
rect 379794 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 380414 633454
rect 379794 633134 380414 633218
rect 379794 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 380414 633134
rect 379794 597454 380414 632898
rect 379794 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 380414 597454
rect 379794 597134 380414 597218
rect 379794 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 380414 597134
rect 379794 561454 380414 596898
rect 379794 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 380414 561454
rect 379794 561134 380414 561218
rect 379794 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 380414 561134
rect 379794 525454 380414 560898
rect 379794 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 380414 525454
rect 379794 525134 380414 525218
rect 379794 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 380414 525134
rect 379794 489454 380414 524898
rect 379794 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 380414 489454
rect 379794 489134 380414 489218
rect 379794 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 380414 489134
rect 379794 453454 380414 488898
rect 379794 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 380414 453454
rect 379794 453134 380414 453218
rect 379794 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 380414 453134
rect 379794 417454 380414 452898
rect 379794 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 380414 417454
rect 379794 417134 380414 417218
rect 379794 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 380414 417134
rect 379794 381454 380414 416898
rect 379794 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 380414 381454
rect 379794 381134 380414 381218
rect 379794 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 380414 381134
rect 379794 345454 380414 380898
rect 379794 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 380414 345454
rect 379794 345134 380414 345218
rect 379794 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 380414 345134
rect 379794 309454 380414 344898
rect 379794 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 380414 309454
rect 379794 309134 380414 309218
rect 379794 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 380414 309134
rect 379794 273454 380414 308898
rect 379794 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 380414 273454
rect 379794 273134 380414 273218
rect 379794 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 380414 273134
rect 379794 237454 380414 272898
rect 379794 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 380414 237454
rect 379794 237134 380414 237218
rect 379794 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 380414 237134
rect 379794 201454 380414 236898
rect 379794 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 380414 201454
rect 379794 201134 380414 201218
rect 379794 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 380414 201134
rect 379794 165454 380414 200898
rect 379794 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 380414 165454
rect 379794 165134 380414 165218
rect 379794 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 380414 165134
rect 379794 129454 380414 164898
rect 379794 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 380414 129454
rect 379794 129134 380414 129218
rect 379794 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 380414 129134
rect 379794 93454 380414 128898
rect 379794 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 380414 93454
rect 379794 93134 380414 93218
rect 379794 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 380414 93134
rect 379794 57454 380414 92898
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -1306 380414 20898
rect 379794 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 380414 -1306
rect 379794 -1626 380414 -1542
rect 379794 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 380414 -1626
rect 379794 -1894 380414 -1862
rect 383514 673174 384134 707162
rect 383514 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 384134 673174
rect 383514 672854 384134 672938
rect 383514 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 384134 672854
rect 383514 637174 384134 672618
rect 383514 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 384134 637174
rect 383514 636854 384134 636938
rect 383514 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 384134 636854
rect 383514 601174 384134 636618
rect 383514 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 384134 601174
rect 383514 600854 384134 600938
rect 383514 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 384134 600854
rect 383514 565174 384134 600618
rect 383514 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 384134 565174
rect 383514 564854 384134 564938
rect 383514 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 384134 564854
rect 383514 529174 384134 564618
rect 383514 528938 383546 529174
rect 383782 528938 383866 529174
rect 384102 528938 384134 529174
rect 383514 528854 384134 528938
rect 383514 528618 383546 528854
rect 383782 528618 383866 528854
rect 384102 528618 384134 528854
rect 383514 493174 384134 528618
rect 383514 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 384134 493174
rect 383514 492854 384134 492938
rect 383514 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 384134 492854
rect 383514 457174 384134 492618
rect 383514 456938 383546 457174
rect 383782 456938 383866 457174
rect 384102 456938 384134 457174
rect 383514 456854 384134 456938
rect 383514 456618 383546 456854
rect 383782 456618 383866 456854
rect 384102 456618 384134 456854
rect 383514 421174 384134 456618
rect 383514 420938 383546 421174
rect 383782 420938 383866 421174
rect 384102 420938 384134 421174
rect 383514 420854 384134 420938
rect 383514 420618 383546 420854
rect 383782 420618 383866 420854
rect 384102 420618 384134 420854
rect 383514 385174 384134 420618
rect 383514 384938 383546 385174
rect 383782 384938 383866 385174
rect 384102 384938 384134 385174
rect 383514 384854 384134 384938
rect 383514 384618 383546 384854
rect 383782 384618 383866 384854
rect 384102 384618 384134 384854
rect 383514 349174 384134 384618
rect 383514 348938 383546 349174
rect 383782 348938 383866 349174
rect 384102 348938 384134 349174
rect 383514 348854 384134 348938
rect 383514 348618 383546 348854
rect 383782 348618 383866 348854
rect 384102 348618 384134 348854
rect 383514 313174 384134 348618
rect 383514 312938 383546 313174
rect 383782 312938 383866 313174
rect 384102 312938 384134 313174
rect 383514 312854 384134 312938
rect 383514 312618 383546 312854
rect 383782 312618 383866 312854
rect 384102 312618 384134 312854
rect 383514 277174 384134 312618
rect 383514 276938 383546 277174
rect 383782 276938 383866 277174
rect 384102 276938 384134 277174
rect 383514 276854 384134 276938
rect 383514 276618 383546 276854
rect 383782 276618 383866 276854
rect 384102 276618 384134 276854
rect 383514 241174 384134 276618
rect 383514 240938 383546 241174
rect 383782 240938 383866 241174
rect 384102 240938 384134 241174
rect 383514 240854 384134 240938
rect 383514 240618 383546 240854
rect 383782 240618 383866 240854
rect 384102 240618 384134 240854
rect 383514 205174 384134 240618
rect 383514 204938 383546 205174
rect 383782 204938 383866 205174
rect 384102 204938 384134 205174
rect 383514 204854 384134 204938
rect 383514 204618 383546 204854
rect 383782 204618 383866 204854
rect 384102 204618 384134 204854
rect 383514 169174 384134 204618
rect 383514 168938 383546 169174
rect 383782 168938 383866 169174
rect 384102 168938 384134 169174
rect 383514 168854 384134 168938
rect 383514 168618 383546 168854
rect 383782 168618 383866 168854
rect 384102 168618 384134 168854
rect 383514 133174 384134 168618
rect 383514 132938 383546 133174
rect 383782 132938 383866 133174
rect 384102 132938 384134 133174
rect 383514 132854 384134 132938
rect 383514 132618 383546 132854
rect 383782 132618 383866 132854
rect 384102 132618 384134 132854
rect 383514 97174 384134 132618
rect 383514 96938 383546 97174
rect 383782 96938 383866 97174
rect 384102 96938 384134 97174
rect 383514 96854 384134 96938
rect 383514 96618 383546 96854
rect 383782 96618 383866 96854
rect 384102 96618 384134 96854
rect 383514 61174 384134 96618
rect 383514 60938 383546 61174
rect 383782 60938 383866 61174
rect 384102 60938 384134 61174
rect 383514 60854 384134 60938
rect 383514 60618 383546 60854
rect 383782 60618 383866 60854
rect 384102 60618 384134 60854
rect 383514 25174 384134 60618
rect 383514 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 384134 25174
rect 383514 24854 384134 24938
rect 383514 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 384134 24854
rect 383514 -3226 384134 24618
rect 383514 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 384134 -3226
rect 383514 -3546 384134 -3462
rect 383514 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 384134 -3546
rect 383514 -3814 384134 -3782
rect 387234 676894 387854 709082
rect 387234 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 387854 676894
rect 387234 676574 387854 676658
rect 387234 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 387854 676574
rect 387234 640894 387854 676338
rect 387234 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 387854 640894
rect 387234 640574 387854 640658
rect 387234 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 387854 640574
rect 387234 604894 387854 640338
rect 387234 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 387854 604894
rect 387234 604574 387854 604658
rect 387234 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 387854 604574
rect 387234 568894 387854 604338
rect 387234 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 387854 568894
rect 387234 568574 387854 568658
rect 387234 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 387854 568574
rect 387234 532894 387854 568338
rect 387234 532658 387266 532894
rect 387502 532658 387586 532894
rect 387822 532658 387854 532894
rect 387234 532574 387854 532658
rect 387234 532338 387266 532574
rect 387502 532338 387586 532574
rect 387822 532338 387854 532574
rect 387234 496894 387854 532338
rect 387234 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 387854 496894
rect 387234 496574 387854 496658
rect 387234 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 387854 496574
rect 387234 460894 387854 496338
rect 387234 460658 387266 460894
rect 387502 460658 387586 460894
rect 387822 460658 387854 460894
rect 387234 460574 387854 460658
rect 387234 460338 387266 460574
rect 387502 460338 387586 460574
rect 387822 460338 387854 460574
rect 387234 424894 387854 460338
rect 387234 424658 387266 424894
rect 387502 424658 387586 424894
rect 387822 424658 387854 424894
rect 387234 424574 387854 424658
rect 387234 424338 387266 424574
rect 387502 424338 387586 424574
rect 387822 424338 387854 424574
rect 387234 388894 387854 424338
rect 387234 388658 387266 388894
rect 387502 388658 387586 388894
rect 387822 388658 387854 388894
rect 387234 388574 387854 388658
rect 387234 388338 387266 388574
rect 387502 388338 387586 388574
rect 387822 388338 387854 388574
rect 387234 352894 387854 388338
rect 387234 352658 387266 352894
rect 387502 352658 387586 352894
rect 387822 352658 387854 352894
rect 387234 352574 387854 352658
rect 387234 352338 387266 352574
rect 387502 352338 387586 352574
rect 387822 352338 387854 352574
rect 387234 316894 387854 352338
rect 387234 316658 387266 316894
rect 387502 316658 387586 316894
rect 387822 316658 387854 316894
rect 387234 316574 387854 316658
rect 387234 316338 387266 316574
rect 387502 316338 387586 316574
rect 387822 316338 387854 316574
rect 387234 280894 387854 316338
rect 387234 280658 387266 280894
rect 387502 280658 387586 280894
rect 387822 280658 387854 280894
rect 387234 280574 387854 280658
rect 387234 280338 387266 280574
rect 387502 280338 387586 280574
rect 387822 280338 387854 280574
rect 387234 244894 387854 280338
rect 387234 244658 387266 244894
rect 387502 244658 387586 244894
rect 387822 244658 387854 244894
rect 387234 244574 387854 244658
rect 387234 244338 387266 244574
rect 387502 244338 387586 244574
rect 387822 244338 387854 244574
rect 387234 208894 387854 244338
rect 387234 208658 387266 208894
rect 387502 208658 387586 208894
rect 387822 208658 387854 208894
rect 387234 208574 387854 208658
rect 387234 208338 387266 208574
rect 387502 208338 387586 208574
rect 387822 208338 387854 208574
rect 387234 172894 387854 208338
rect 387234 172658 387266 172894
rect 387502 172658 387586 172894
rect 387822 172658 387854 172894
rect 387234 172574 387854 172658
rect 387234 172338 387266 172574
rect 387502 172338 387586 172574
rect 387822 172338 387854 172574
rect 387234 136894 387854 172338
rect 387234 136658 387266 136894
rect 387502 136658 387586 136894
rect 387822 136658 387854 136894
rect 387234 136574 387854 136658
rect 387234 136338 387266 136574
rect 387502 136338 387586 136574
rect 387822 136338 387854 136574
rect 387234 100894 387854 136338
rect 387234 100658 387266 100894
rect 387502 100658 387586 100894
rect 387822 100658 387854 100894
rect 387234 100574 387854 100658
rect 387234 100338 387266 100574
rect 387502 100338 387586 100574
rect 387822 100338 387854 100574
rect 387234 64894 387854 100338
rect 387234 64658 387266 64894
rect 387502 64658 387586 64894
rect 387822 64658 387854 64894
rect 387234 64574 387854 64658
rect 387234 64338 387266 64574
rect 387502 64338 387586 64574
rect 387822 64338 387854 64574
rect 387234 28894 387854 64338
rect 387234 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 387854 28894
rect 387234 28574 387854 28658
rect 387234 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 387854 28574
rect 387234 -5146 387854 28338
rect 387234 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 387854 -5146
rect 387234 -5466 387854 -5382
rect 387234 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 387854 -5466
rect 387234 -5734 387854 -5702
rect 390954 680614 391574 711002
rect 408954 710598 409574 711590
rect 408954 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 409574 710598
rect 408954 710278 409574 710362
rect 408954 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 409574 710278
rect 405234 708678 405854 709670
rect 405234 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 405854 708678
rect 405234 708358 405854 708442
rect 405234 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 405854 708358
rect 401514 706758 402134 707750
rect 401514 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 402134 706758
rect 401514 706438 402134 706522
rect 401514 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 402134 706438
rect 390954 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 391574 680614
rect 390954 680294 391574 680378
rect 390954 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 391574 680294
rect 390954 644614 391574 680058
rect 390954 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 391574 644614
rect 390954 644294 391574 644378
rect 390954 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 391574 644294
rect 390954 608614 391574 644058
rect 390954 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 391574 608614
rect 390954 608294 391574 608378
rect 390954 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 391574 608294
rect 390954 572614 391574 608058
rect 390954 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 391574 572614
rect 390954 572294 391574 572378
rect 390954 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 391574 572294
rect 390954 536614 391574 572058
rect 390954 536378 390986 536614
rect 391222 536378 391306 536614
rect 391542 536378 391574 536614
rect 390954 536294 391574 536378
rect 390954 536058 390986 536294
rect 391222 536058 391306 536294
rect 391542 536058 391574 536294
rect 390954 500614 391574 536058
rect 390954 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 391574 500614
rect 390954 500294 391574 500378
rect 390954 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 391574 500294
rect 390954 464614 391574 500058
rect 390954 464378 390986 464614
rect 391222 464378 391306 464614
rect 391542 464378 391574 464614
rect 390954 464294 391574 464378
rect 390954 464058 390986 464294
rect 391222 464058 391306 464294
rect 391542 464058 391574 464294
rect 390954 428614 391574 464058
rect 390954 428378 390986 428614
rect 391222 428378 391306 428614
rect 391542 428378 391574 428614
rect 390954 428294 391574 428378
rect 390954 428058 390986 428294
rect 391222 428058 391306 428294
rect 391542 428058 391574 428294
rect 390954 392614 391574 428058
rect 390954 392378 390986 392614
rect 391222 392378 391306 392614
rect 391542 392378 391574 392614
rect 390954 392294 391574 392378
rect 390954 392058 390986 392294
rect 391222 392058 391306 392294
rect 391542 392058 391574 392294
rect 390954 356614 391574 392058
rect 390954 356378 390986 356614
rect 391222 356378 391306 356614
rect 391542 356378 391574 356614
rect 390954 356294 391574 356378
rect 390954 356058 390986 356294
rect 391222 356058 391306 356294
rect 391542 356058 391574 356294
rect 390954 320614 391574 356058
rect 390954 320378 390986 320614
rect 391222 320378 391306 320614
rect 391542 320378 391574 320614
rect 390954 320294 391574 320378
rect 390954 320058 390986 320294
rect 391222 320058 391306 320294
rect 391542 320058 391574 320294
rect 390954 284614 391574 320058
rect 390954 284378 390986 284614
rect 391222 284378 391306 284614
rect 391542 284378 391574 284614
rect 390954 284294 391574 284378
rect 390954 284058 390986 284294
rect 391222 284058 391306 284294
rect 391542 284058 391574 284294
rect 390954 248614 391574 284058
rect 390954 248378 390986 248614
rect 391222 248378 391306 248614
rect 391542 248378 391574 248614
rect 390954 248294 391574 248378
rect 390954 248058 390986 248294
rect 391222 248058 391306 248294
rect 391542 248058 391574 248294
rect 390954 212614 391574 248058
rect 390954 212378 390986 212614
rect 391222 212378 391306 212614
rect 391542 212378 391574 212614
rect 390954 212294 391574 212378
rect 390954 212058 390986 212294
rect 391222 212058 391306 212294
rect 391542 212058 391574 212294
rect 390954 176614 391574 212058
rect 390954 176378 390986 176614
rect 391222 176378 391306 176614
rect 391542 176378 391574 176614
rect 390954 176294 391574 176378
rect 390954 176058 390986 176294
rect 391222 176058 391306 176294
rect 391542 176058 391574 176294
rect 390954 140614 391574 176058
rect 397794 704838 398414 705830
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 543454 398414 578898
rect 397794 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 398414 543454
rect 397794 543134 398414 543218
rect 397794 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 398414 543134
rect 397794 507454 398414 542898
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 435454 398414 470898
rect 397794 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 398414 435454
rect 397794 435134 398414 435218
rect 397794 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 398414 435134
rect 397794 399454 398414 434898
rect 397794 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 398414 399454
rect 397794 399134 398414 399218
rect 397794 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 398414 399134
rect 397794 363454 398414 398898
rect 401514 691174 402134 706202
rect 401514 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 402134 691174
rect 401514 690854 402134 690938
rect 401514 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 402134 690854
rect 401514 655174 402134 690618
rect 401514 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 402134 655174
rect 401514 654854 402134 654938
rect 401514 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 402134 654854
rect 401514 619174 402134 654618
rect 401514 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 402134 619174
rect 401514 618854 402134 618938
rect 401514 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 402134 618854
rect 401514 583174 402134 618618
rect 401514 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 402134 583174
rect 401514 582854 402134 582938
rect 401514 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 402134 582854
rect 401514 547174 402134 582618
rect 401514 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 402134 547174
rect 401514 546854 402134 546938
rect 401514 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 402134 546854
rect 401514 511174 402134 546618
rect 401514 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 402134 511174
rect 401514 510854 402134 510938
rect 401514 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 402134 510854
rect 401514 475174 402134 510618
rect 401514 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 402134 475174
rect 401514 474854 402134 474938
rect 401514 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 402134 474854
rect 401514 439174 402134 474618
rect 401514 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 402134 439174
rect 401514 438854 402134 438938
rect 401514 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 402134 438854
rect 401514 403174 402134 438618
rect 401514 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 402134 403174
rect 401514 402854 402134 402938
rect 401514 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 402134 402854
rect 400259 393412 400325 393413
rect 400259 393348 400260 393412
rect 400324 393348 400325 393412
rect 400259 393347 400325 393348
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 397794 327454 398414 362898
rect 397794 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 398414 327454
rect 397794 327134 398414 327218
rect 397794 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 398414 327134
rect 397794 291454 398414 326898
rect 397794 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 398414 291454
rect 397794 291134 398414 291218
rect 397794 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 398414 291134
rect 397794 255454 398414 290898
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 219454 398414 254898
rect 397794 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 398414 219454
rect 397794 219134 398414 219218
rect 397794 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 398414 219134
rect 397794 183454 398414 218898
rect 397794 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 398414 183454
rect 397794 183134 398414 183218
rect 397794 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 398414 183134
rect 397794 147454 398414 182898
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 142000 398414 146898
rect 390954 140378 390986 140614
rect 391222 140378 391306 140614
rect 391542 140378 391574 140614
rect 390954 140294 391574 140378
rect 390954 140058 390986 140294
rect 391222 140058 391306 140294
rect 391542 140058 391574 140294
rect 390954 104614 391574 140058
rect 400262 135149 400322 393347
rect 401514 367174 402134 402618
rect 401514 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 402134 367174
rect 401514 366854 402134 366938
rect 401514 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 402134 366854
rect 401514 331174 402134 366618
rect 401514 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 402134 331174
rect 401514 330854 402134 330938
rect 401514 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 402134 330854
rect 401514 295174 402134 330618
rect 401514 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 402134 295174
rect 401514 294854 402134 294938
rect 401514 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 402134 294854
rect 401514 259174 402134 294618
rect 401514 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 402134 259174
rect 401514 258854 402134 258938
rect 401514 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 402134 258854
rect 401514 223174 402134 258618
rect 401514 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 402134 223174
rect 401514 222854 402134 222938
rect 401514 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 402134 222854
rect 401514 187174 402134 222618
rect 401514 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 402134 187174
rect 401514 186854 402134 186938
rect 401514 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 402134 186854
rect 401514 151174 402134 186618
rect 401514 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 402134 151174
rect 401514 150854 402134 150938
rect 401514 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 402134 150854
rect 401514 142000 402134 150618
rect 405234 694894 405854 708122
rect 405234 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 405854 694894
rect 405234 694574 405854 694658
rect 405234 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 405854 694574
rect 405234 658894 405854 694338
rect 405234 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 405854 658894
rect 405234 658574 405854 658658
rect 405234 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 405854 658574
rect 405234 622894 405854 658338
rect 405234 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 405854 622894
rect 405234 622574 405854 622658
rect 405234 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 405854 622574
rect 405234 586894 405854 622338
rect 405234 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 405854 586894
rect 405234 586574 405854 586658
rect 405234 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 405854 586574
rect 405234 550894 405854 586338
rect 405234 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 405854 550894
rect 405234 550574 405854 550658
rect 405234 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 405854 550574
rect 405234 514894 405854 550338
rect 405234 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 405854 514894
rect 405234 514574 405854 514658
rect 405234 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 405854 514574
rect 405234 478894 405854 514338
rect 405234 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 405854 478894
rect 405234 478574 405854 478658
rect 405234 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 405854 478574
rect 405234 442894 405854 478338
rect 405234 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 405854 442894
rect 405234 442574 405854 442658
rect 405234 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 405854 442574
rect 405234 406894 405854 442338
rect 405234 406658 405266 406894
rect 405502 406658 405586 406894
rect 405822 406658 405854 406894
rect 405234 406574 405854 406658
rect 405234 406338 405266 406574
rect 405502 406338 405586 406574
rect 405822 406338 405854 406574
rect 405234 370894 405854 406338
rect 405234 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 405854 370894
rect 405234 370574 405854 370658
rect 405234 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 405854 370574
rect 405234 334894 405854 370338
rect 405234 334658 405266 334894
rect 405502 334658 405586 334894
rect 405822 334658 405854 334894
rect 405234 334574 405854 334658
rect 405234 334338 405266 334574
rect 405502 334338 405586 334574
rect 405822 334338 405854 334574
rect 405234 298894 405854 334338
rect 405234 298658 405266 298894
rect 405502 298658 405586 298894
rect 405822 298658 405854 298894
rect 405234 298574 405854 298658
rect 405234 298338 405266 298574
rect 405502 298338 405586 298574
rect 405822 298338 405854 298574
rect 405234 262894 405854 298338
rect 405234 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 405854 262894
rect 405234 262574 405854 262658
rect 405234 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 405854 262574
rect 405234 226894 405854 262338
rect 405234 226658 405266 226894
rect 405502 226658 405586 226894
rect 405822 226658 405854 226894
rect 405234 226574 405854 226658
rect 405234 226338 405266 226574
rect 405502 226338 405586 226574
rect 405822 226338 405854 226574
rect 405234 190894 405854 226338
rect 405234 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 405854 190894
rect 405234 190574 405854 190658
rect 405234 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 405854 190574
rect 405234 154894 405854 190338
rect 405234 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 405854 154894
rect 405234 154574 405854 154658
rect 405234 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 405854 154574
rect 405234 142000 405854 154338
rect 408954 698614 409574 710042
rect 426954 711558 427574 711590
rect 426954 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 427574 711558
rect 426954 711238 427574 711322
rect 426954 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 427574 711238
rect 423234 709638 423854 709670
rect 423234 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 423854 709638
rect 423234 709318 423854 709402
rect 423234 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 423854 709318
rect 419514 707718 420134 707750
rect 419514 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 420134 707718
rect 419514 707398 420134 707482
rect 419514 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 420134 707398
rect 408954 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 409574 698614
rect 408954 698294 409574 698378
rect 408954 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 409574 698294
rect 408954 662614 409574 698058
rect 408954 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 409574 662614
rect 408954 662294 409574 662378
rect 408954 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 409574 662294
rect 408954 626614 409574 662058
rect 408954 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 409574 626614
rect 408954 626294 409574 626378
rect 408954 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 409574 626294
rect 408954 590614 409574 626058
rect 408954 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 409574 590614
rect 408954 590294 409574 590378
rect 408954 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 409574 590294
rect 408954 554614 409574 590058
rect 408954 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 409574 554614
rect 408954 554294 409574 554378
rect 408954 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 409574 554294
rect 408954 518614 409574 554058
rect 408954 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 409574 518614
rect 408954 518294 409574 518378
rect 408954 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 409574 518294
rect 408954 482614 409574 518058
rect 408954 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 409574 482614
rect 408954 482294 409574 482378
rect 408954 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 409574 482294
rect 408954 446614 409574 482058
rect 408954 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 409574 446614
rect 408954 446294 409574 446378
rect 408954 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 409574 446294
rect 408954 410614 409574 446058
rect 408954 410378 408986 410614
rect 409222 410378 409306 410614
rect 409542 410378 409574 410614
rect 408954 410294 409574 410378
rect 408954 410058 408986 410294
rect 409222 410058 409306 410294
rect 409542 410058 409574 410294
rect 408954 374614 409574 410058
rect 408954 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 409574 374614
rect 408954 374294 409574 374378
rect 408954 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 409574 374294
rect 408954 338614 409574 374058
rect 408954 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 409574 338614
rect 408954 338294 409574 338378
rect 408954 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 409574 338294
rect 408954 302614 409574 338058
rect 408954 302378 408986 302614
rect 409222 302378 409306 302614
rect 409542 302378 409574 302614
rect 408954 302294 409574 302378
rect 408954 302058 408986 302294
rect 409222 302058 409306 302294
rect 409542 302058 409574 302294
rect 408954 266614 409574 302058
rect 408954 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 409574 266614
rect 408954 266294 409574 266378
rect 408954 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 409574 266294
rect 408954 230614 409574 266058
rect 408954 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 409574 230614
rect 408954 230294 409574 230378
rect 408954 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 409574 230294
rect 408954 194614 409574 230058
rect 408954 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 409574 194614
rect 408954 194294 409574 194378
rect 408954 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 409574 194294
rect 408954 158614 409574 194058
rect 408954 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 409574 158614
rect 408954 158294 409574 158378
rect 408954 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 409574 158294
rect 408954 142000 409574 158058
rect 415794 705798 416414 705830
rect 415794 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 416414 705798
rect 415794 705478 416414 705562
rect 415794 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 416414 705478
rect 415794 669454 416414 705242
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 633454 416414 668898
rect 415794 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 416414 633454
rect 415794 633134 416414 633218
rect 415794 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 416414 633134
rect 415794 597454 416414 632898
rect 415794 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 416414 597454
rect 415794 597134 416414 597218
rect 415794 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 416414 597134
rect 415794 561454 416414 596898
rect 415794 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 416414 561454
rect 415794 561134 416414 561218
rect 415794 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 416414 561134
rect 415794 525454 416414 560898
rect 415794 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 416414 525454
rect 415794 525134 416414 525218
rect 415794 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 416414 525134
rect 415794 489454 416414 524898
rect 415794 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 416414 489454
rect 415794 489134 416414 489218
rect 415794 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 416414 489134
rect 415794 453454 416414 488898
rect 415794 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 416414 453454
rect 415794 453134 416414 453218
rect 415794 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 416414 453134
rect 415794 417454 416414 452898
rect 415794 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 416414 417454
rect 415794 417134 416414 417218
rect 415794 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 416414 417134
rect 415794 381454 416414 416898
rect 415794 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 416414 381454
rect 415794 381134 416414 381218
rect 415794 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 416414 381134
rect 415794 345454 416414 380898
rect 415794 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 416414 345454
rect 415794 345134 416414 345218
rect 415794 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 416414 345134
rect 415794 309454 416414 344898
rect 415794 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 416414 309454
rect 415794 309134 416414 309218
rect 415794 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 416414 309134
rect 415794 273454 416414 308898
rect 415794 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 416414 273454
rect 415794 273134 416414 273218
rect 415794 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 416414 273134
rect 415794 237454 416414 272898
rect 415794 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 416414 237454
rect 415794 237134 416414 237218
rect 415794 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 416414 237134
rect 415794 201454 416414 236898
rect 415794 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 416414 201454
rect 415794 201134 416414 201218
rect 415794 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 416414 201134
rect 415794 165454 416414 200898
rect 415794 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 416414 165454
rect 415794 165134 416414 165218
rect 415794 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 416414 165134
rect 409827 143444 409893 143445
rect 409827 143380 409828 143444
rect 409892 143380 409893 143444
rect 409827 143379 409893 143380
rect 400259 135148 400325 135149
rect 400259 135084 400260 135148
rect 400324 135084 400325 135148
rect 400259 135083 400325 135084
rect 402544 129454 402864 129486
rect 402544 129218 402586 129454
rect 402822 129218 402864 129454
rect 402544 129134 402864 129218
rect 402544 128898 402586 129134
rect 402822 128898 402864 129134
rect 402544 128866 402864 128898
rect 405744 129454 406064 129486
rect 405744 129218 405786 129454
rect 406022 129218 406064 129454
rect 405744 129134 406064 129218
rect 405744 128898 405786 129134
rect 406022 128898 406064 129134
rect 405744 128866 406064 128898
rect 408944 129454 409264 129486
rect 408944 129218 408986 129454
rect 409222 129218 409264 129454
rect 408944 129134 409264 129218
rect 408944 128898 408986 129134
rect 409222 128898 409264 129134
rect 408944 128866 409264 128898
rect 404144 111454 404464 111486
rect 404144 111218 404186 111454
rect 404422 111218 404464 111454
rect 404144 111134 404464 111218
rect 404144 110898 404186 111134
rect 404422 110898 404464 111134
rect 404144 110866 404464 110898
rect 407344 111454 407664 111486
rect 407344 111218 407386 111454
rect 407622 111218 407664 111454
rect 407344 111134 407664 111218
rect 407344 110898 407386 111134
rect 407622 110898 407664 111134
rect 407344 110866 407664 110898
rect 390954 104378 390986 104614
rect 391222 104378 391306 104614
rect 391542 104378 391574 104614
rect 390954 104294 391574 104378
rect 390954 104058 390986 104294
rect 391222 104058 391306 104294
rect 391542 104058 391574 104294
rect 390954 68614 391574 104058
rect 398787 102780 398853 102781
rect 398787 102716 398788 102780
rect 398852 102716 398853 102780
rect 398787 102715 398853 102716
rect 398790 99381 398850 102715
rect 398787 99380 398853 99381
rect 398787 99316 398788 99380
rect 398852 99316 398853 99380
rect 398787 99315 398853 99316
rect 390954 68378 390986 68614
rect 391222 68378 391306 68614
rect 391542 68378 391574 68614
rect 390954 68294 391574 68378
rect 390954 68058 390986 68294
rect 391222 68058 391306 68294
rect 391542 68058 391574 68294
rect 390954 32614 391574 68058
rect 390954 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 391574 32614
rect 390954 32294 391574 32378
rect 390954 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 391574 32294
rect 372954 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 373574 -6106
rect 372954 -6426 373574 -6342
rect 372954 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 373574 -6426
rect 372954 -7654 373574 -6662
rect 390954 -7066 391574 32058
rect 397794 75454 398414 98000
rect 397794 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 398414 75454
rect 397794 75134 398414 75218
rect 397794 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 398414 75134
rect 397794 39454 398414 74898
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -1894 398414 -902
rect 401514 79174 402134 98000
rect 401514 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 402134 79174
rect 401514 78854 402134 78938
rect 401514 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 402134 78854
rect 401514 43174 402134 78618
rect 401514 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 402134 43174
rect 401514 42854 402134 42938
rect 401514 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 402134 42854
rect 401514 7174 402134 42618
rect 401514 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 402134 7174
rect 401514 6854 402134 6938
rect 401514 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 402134 6854
rect 401514 -2266 402134 6618
rect 401514 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 402134 -2266
rect 401514 -2586 402134 -2502
rect 401514 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 402134 -2586
rect 401514 -3814 402134 -2822
rect 405234 82894 405854 98000
rect 405234 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 405854 82894
rect 405234 82574 405854 82658
rect 405234 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 405854 82574
rect 405234 46894 405854 82338
rect 405234 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 405854 46894
rect 405234 46574 405854 46658
rect 405234 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 405854 46574
rect 405234 10894 405854 46338
rect 405234 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 405854 10894
rect 405234 10574 405854 10658
rect 405234 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 405854 10574
rect 405234 -4186 405854 10338
rect 405234 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 405854 -4186
rect 405234 -4506 405854 -4422
rect 405234 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 405854 -4506
rect 405234 -5734 405854 -4742
rect 408954 86614 409574 98000
rect 408954 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 409574 86614
rect 408954 86294 409574 86378
rect 408954 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 409574 86294
rect 408954 50614 409574 86058
rect 409830 57221 409890 143379
rect 415794 142000 416414 164898
rect 419514 673174 420134 707162
rect 419514 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 420134 673174
rect 419514 672854 420134 672938
rect 419514 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 420134 672854
rect 419514 637174 420134 672618
rect 419514 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 420134 637174
rect 419514 636854 420134 636938
rect 419514 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 420134 636854
rect 419514 601174 420134 636618
rect 419514 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 420134 601174
rect 419514 600854 420134 600938
rect 419514 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 420134 600854
rect 419514 565174 420134 600618
rect 419514 564938 419546 565174
rect 419782 564938 419866 565174
rect 420102 564938 420134 565174
rect 419514 564854 420134 564938
rect 419514 564618 419546 564854
rect 419782 564618 419866 564854
rect 420102 564618 420134 564854
rect 419514 529174 420134 564618
rect 419514 528938 419546 529174
rect 419782 528938 419866 529174
rect 420102 528938 420134 529174
rect 419514 528854 420134 528938
rect 419514 528618 419546 528854
rect 419782 528618 419866 528854
rect 420102 528618 420134 528854
rect 419514 493174 420134 528618
rect 419514 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 420134 493174
rect 419514 492854 420134 492938
rect 419514 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 420134 492854
rect 419514 457174 420134 492618
rect 419514 456938 419546 457174
rect 419782 456938 419866 457174
rect 420102 456938 420134 457174
rect 419514 456854 420134 456938
rect 419514 456618 419546 456854
rect 419782 456618 419866 456854
rect 420102 456618 420134 456854
rect 419514 421174 420134 456618
rect 419514 420938 419546 421174
rect 419782 420938 419866 421174
rect 420102 420938 420134 421174
rect 419514 420854 420134 420938
rect 419514 420618 419546 420854
rect 419782 420618 419866 420854
rect 420102 420618 420134 420854
rect 419514 385174 420134 420618
rect 419514 384938 419546 385174
rect 419782 384938 419866 385174
rect 420102 384938 420134 385174
rect 419514 384854 420134 384938
rect 419514 384618 419546 384854
rect 419782 384618 419866 384854
rect 420102 384618 420134 384854
rect 419514 349174 420134 384618
rect 419514 348938 419546 349174
rect 419782 348938 419866 349174
rect 420102 348938 420134 349174
rect 419514 348854 420134 348938
rect 419514 348618 419546 348854
rect 419782 348618 419866 348854
rect 420102 348618 420134 348854
rect 419514 313174 420134 348618
rect 419514 312938 419546 313174
rect 419782 312938 419866 313174
rect 420102 312938 420134 313174
rect 419514 312854 420134 312938
rect 419514 312618 419546 312854
rect 419782 312618 419866 312854
rect 420102 312618 420134 312854
rect 419514 277174 420134 312618
rect 419514 276938 419546 277174
rect 419782 276938 419866 277174
rect 420102 276938 420134 277174
rect 419514 276854 420134 276938
rect 419514 276618 419546 276854
rect 419782 276618 419866 276854
rect 420102 276618 420134 276854
rect 419514 241174 420134 276618
rect 419514 240938 419546 241174
rect 419782 240938 419866 241174
rect 420102 240938 420134 241174
rect 419514 240854 420134 240938
rect 419514 240618 419546 240854
rect 419782 240618 419866 240854
rect 420102 240618 420134 240854
rect 419514 205174 420134 240618
rect 419514 204938 419546 205174
rect 419782 204938 419866 205174
rect 420102 204938 420134 205174
rect 419514 204854 420134 204938
rect 419514 204618 419546 204854
rect 419782 204618 419866 204854
rect 420102 204618 420134 204854
rect 419514 169174 420134 204618
rect 419514 168938 419546 169174
rect 419782 168938 419866 169174
rect 420102 168938 420134 169174
rect 419514 168854 420134 168938
rect 419514 168618 419546 168854
rect 419782 168618 419866 168854
rect 420102 168618 420134 168854
rect 417371 143444 417437 143445
rect 417371 143380 417372 143444
rect 417436 143380 417437 143444
rect 417371 143379 417437 143380
rect 412144 129454 412464 129486
rect 412144 129218 412186 129454
rect 412422 129218 412464 129454
rect 412144 129134 412464 129218
rect 412144 128898 412186 129134
rect 412422 128898 412464 129134
rect 412144 128866 412464 128898
rect 415344 129454 415664 129486
rect 415344 129218 415386 129454
rect 415622 129218 415664 129454
rect 415344 129134 415664 129218
rect 415344 128898 415386 129134
rect 415622 128898 415664 129134
rect 415344 128866 415664 128898
rect 410544 111454 410864 111486
rect 410544 111218 410586 111454
rect 410822 111218 410864 111454
rect 410544 111134 410864 111218
rect 410544 110898 410586 111134
rect 410822 110898 410864 111134
rect 410544 110866 410864 110898
rect 413744 111454 414064 111486
rect 413744 111218 413786 111454
rect 414022 111218 414064 111454
rect 413744 111134 414064 111218
rect 413744 110898 413786 111134
rect 414022 110898 414064 111134
rect 413744 110866 414064 110898
rect 416944 111454 417264 111486
rect 416944 111218 416986 111454
rect 417222 111218 417264 111454
rect 416944 111134 417264 111218
rect 416944 110898 416986 111134
rect 417222 110898 417264 111134
rect 416944 110866 417264 110898
rect 415794 93454 416414 98000
rect 415794 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 416414 93454
rect 415794 93134 416414 93218
rect 415794 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 416414 93134
rect 415794 57454 416414 92898
rect 409827 57220 409893 57221
rect 409827 57156 409828 57220
rect 409892 57156 409893 57220
rect 409827 57155 409893 57156
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 408954 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 409574 50614
rect 408954 50294 409574 50378
rect 408954 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 409574 50294
rect 408954 14614 409574 50058
rect 408954 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 409574 14614
rect 408954 14294 409574 14378
rect 408954 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 409574 14294
rect 390954 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 391574 -7066
rect 390954 -7386 391574 -7302
rect 390954 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 391574 -7386
rect 390954 -7654 391574 -7622
rect 408954 -6106 409574 14058
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 415794 21454 416414 56898
rect 417374 33829 417434 143379
rect 419514 142000 420134 168618
rect 423234 676894 423854 709082
rect 423234 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 423854 676894
rect 423234 676574 423854 676658
rect 423234 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 423854 676574
rect 423234 640894 423854 676338
rect 423234 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 423854 640894
rect 423234 640574 423854 640658
rect 423234 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 423854 640574
rect 423234 604894 423854 640338
rect 423234 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 423854 604894
rect 423234 604574 423854 604658
rect 423234 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 423854 604574
rect 423234 568894 423854 604338
rect 423234 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 423854 568894
rect 423234 568574 423854 568658
rect 423234 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 423854 568574
rect 423234 532894 423854 568338
rect 423234 532658 423266 532894
rect 423502 532658 423586 532894
rect 423822 532658 423854 532894
rect 423234 532574 423854 532658
rect 423234 532338 423266 532574
rect 423502 532338 423586 532574
rect 423822 532338 423854 532574
rect 423234 496894 423854 532338
rect 423234 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 423854 496894
rect 423234 496574 423854 496658
rect 423234 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 423854 496574
rect 423234 460894 423854 496338
rect 423234 460658 423266 460894
rect 423502 460658 423586 460894
rect 423822 460658 423854 460894
rect 423234 460574 423854 460658
rect 423234 460338 423266 460574
rect 423502 460338 423586 460574
rect 423822 460338 423854 460574
rect 423234 424894 423854 460338
rect 423234 424658 423266 424894
rect 423502 424658 423586 424894
rect 423822 424658 423854 424894
rect 423234 424574 423854 424658
rect 423234 424338 423266 424574
rect 423502 424338 423586 424574
rect 423822 424338 423854 424574
rect 423234 388894 423854 424338
rect 423234 388658 423266 388894
rect 423502 388658 423586 388894
rect 423822 388658 423854 388894
rect 423234 388574 423854 388658
rect 423234 388338 423266 388574
rect 423502 388338 423586 388574
rect 423822 388338 423854 388574
rect 423234 352894 423854 388338
rect 423234 352658 423266 352894
rect 423502 352658 423586 352894
rect 423822 352658 423854 352894
rect 423234 352574 423854 352658
rect 423234 352338 423266 352574
rect 423502 352338 423586 352574
rect 423822 352338 423854 352574
rect 423234 316894 423854 352338
rect 423234 316658 423266 316894
rect 423502 316658 423586 316894
rect 423822 316658 423854 316894
rect 423234 316574 423854 316658
rect 423234 316338 423266 316574
rect 423502 316338 423586 316574
rect 423822 316338 423854 316574
rect 423234 280894 423854 316338
rect 426954 680614 427574 711002
rect 444954 710598 445574 711590
rect 444954 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 445574 710598
rect 444954 710278 445574 710362
rect 444954 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 445574 710278
rect 441234 708678 441854 709670
rect 441234 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 441854 708678
rect 441234 708358 441854 708442
rect 441234 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 441854 708358
rect 437514 706758 438134 707750
rect 437514 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 438134 706758
rect 437514 706438 438134 706522
rect 437514 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 438134 706438
rect 426954 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 427574 680614
rect 426954 680294 427574 680378
rect 426954 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 427574 680294
rect 426954 644614 427574 680058
rect 426954 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 427574 644614
rect 426954 644294 427574 644378
rect 426954 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 427574 644294
rect 426954 608614 427574 644058
rect 426954 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 427574 608614
rect 426954 608294 427574 608378
rect 426954 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 427574 608294
rect 426954 572614 427574 608058
rect 426954 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 427574 572614
rect 426954 572294 427574 572378
rect 426954 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 427574 572294
rect 426954 536614 427574 572058
rect 426954 536378 426986 536614
rect 427222 536378 427306 536614
rect 427542 536378 427574 536614
rect 426954 536294 427574 536378
rect 426954 536058 426986 536294
rect 427222 536058 427306 536294
rect 427542 536058 427574 536294
rect 426954 500614 427574 536058
rect 426954 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 427574 500614
rect 426954 500294 427574 500378
rect 426954 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 427574 500294
rect 426954 464614 427574 500058
rect 426954 464378 426986 464614
rect 427222 464378 427306 464614
rect 427542 464378 427574 464614
rect 426954 464294 427574 464378
rect 426954 464058 426986 464294
rect 427222 464058 427306 464294
rect 427542 464058 427574 464294
rect 426954 428614 427574 464058
rect 426954 428378 426986 428614
rect 427222 428378 427306 428614
rect 427542 428378 427574 428614
rect 426954 428294 427574 428378
rect 426954 428058 426986 428294
rect 427222 428058 427306 428294
rect 427542 428058 427574 428294
rect 426954 392614 427574 428058
rect 426954 392378 426986 392614
rect 427222 392378 427306 392614
rect 427542 392378 427574 392614
rect 426954 392294 427574 392378
rect 426954 392058 426986 392294
rect 427222 392058 427306 392294
rect 427542 392058 427574 392294
rect 426954 356614 427574 392058
rect 426954 356378 426986 356614
rect 427222 356378 427306 356614
rect 427542 356378 427574 356614
rect 426954 356294 427574 356378
rect 426954 356058 426986 356294
rect 427222 356058 427306 356294
rect 427542 356058 427574 356294
rect 426954 320614 427574 356058
rect 426954 320378 426986 320614
rect 427222 320378 427306 320614
rect 427542 320378 427574 320614
rect 426954 320294 427574 320378
rect 426954 320058 426986 320294
rect 427222 320058 427306 320294
rect 427542 320058 427574 320294
rect 425651 285020 425717 285021
rect 425651 284956 425652 285020
rect 425716 284956 425717 285020
rect 425651 284955 425717 284956
rect 423234 280658 423266 280894
rect 423502 280658 423586 280894
rect 423822 280658 423854 280894
rect 423234 280574 423854 280658
rect 423234 280338 423266 280574
rect 423502 280338 423586 280574
rect 423822 280338 423854 280574
rect 423234 244894 423854 280338
rect 423234 244658 423266 244894
rect 423502 244658 423586 244894
rect 423822 244658 423854 244894
rect 423234 244574 423854 244658
rect 423234 244338 423266 244574
rect 423502 244338 423586 244574
rect 423822 244338 423854 244574
rect 423234 208894 423854 244338
rect 423234 208658 423266 208894
rect 423502 208658 423586 208894
rect 423822 208658 423854 208894
rect 423234 208574 423854 208658
rect 423234 208338 423266 208574
rect 423502 208338 423586 208574
rect 423822 208338 423854 208574
rect 423234 172894 423854 208338
rect 423995 207636 424061 207637
rect 423995 207572 423996 207636
rect 424060 207572 424061 207636
rect 423995 207571 424061 207572
rect 423234 172658 423266 172894
rect 423502 172658 423586 172894
rect 423822 172658 423854 172894
rect 423234 172574 423854 172658
rect 423234 172338 423266 172574
rect 423502 172338 423586 172574
rect 423822 172338 423854 172574
rect 423234 142000 423854 172338
rect 419027 139772 419093 139773
rect 419027 139708 419028 139772
rect 419092 139708 419093 139772
rect 419027 139707 419093 139708
rect 418544 129454 418864 129486
rect 418544 129218 418586 129454
rect 418822 129218 418864 129454
rect 418544 129134 418864 129218
rect 418544 128898 418586 129134
rect 418822 128898 418864 129134
rect 418544 128866 418864 128898
rect 417371 33828 417437 33829
rect 417371 33764 417372 33828
rect 417436 33764 417437 33828
rect 417371 33763 417437 33764
rect 419030 23357 419090 139707
rect 420683 139636 420749 139637
rect 420683 139572 420684 139636
rect 420748 139572 420749 139636
rect 420683 139571 420749 139572
rect 420144 111454 420464 111486
rect 420144 111218 420186 111454
rect 420422 111218 420464 111454
rect 420144 111134 420464 111218
rect 420144 110898 420186 111134
rect 420422 110898 420464 111134
rect 420144 110866 420464 110898
rect 419514 97174 420134 98000
rect 419514 96938 419546 97174
rect 419782 96938 419866 97174
rect 420102 96938 420134 97174
rect 419514 96854 420134 96938
rect 419514 96618 419546 96854
rect 419782 96618 419866 96854
rect 420102 96618 420134 96854
rect 419514 61174 420134 96618
rect 420686 90405 420746 139571
rect 421051 139500 421117 139501
rect 421051 139436 421052 139500
rect 421116 139436 421117 139500
rect 421051 139435 421117 139436
rect 420683 90404 420749 90405
rect 420683 90340 420684 90404
rect 420748 90340 420749 90404
rect 420683 90339 420749 90340
rect 421054 73813 421114 139435
rect 421744 129454 422064 129486
rect 421744 129218 421786 129454
rect 422022 129218 422064 129454
rect 421744 129134 422064 129218
rect 421744 128898 421786 129134
rect 422022 128898 422064 129134
rect 421744 128866 422064 128898
rect 423344 111454 423664 111486
rect 423344 111218 423386 111454
rect 423622 111218 423664 111454
rect 423344 111134 423664 111218
rect 423344 110898 423386 111134
rect 423622 110898 423664 111134
rect 423344 110866 423664 110898
rect 423998 100741 424058 207571
rect 424944 129454 425264 129486
rect 424944 129218 424986 129454
rect 425222 129218 425264 129454
rect 424944 129134 425264 129218
rect 424944 128898 424986 129134
rect 425222 128898 425264 129134
rect 424944 128866 425264 128898
rect 425654 100741 425714 284955
rect 426954 284614 427574 320058
rect 426954 284378 426986 284614
rect 427222 284378 427306 284614
rect 427542 284378 427574 284614
rect 426954 284294 427574 284378
rect 426954 284058 426986 284294
rect 427222 284058 427306 284294
rect 427542 284058 427574 284294
rect 426954 248614 427574 284058
rect 426954 248378 426986 248614
rect 427222 248378 427306 248614
rect 427542 248378 427574 248614
rect 426954 248294 427574 248378
rect 426954 248058 426986 248294
rect 427222 248058 427306 248294
rect 427542 248058 427574 248294
rect 426954 212614 427574 248058
rect 426954 212378 426986 212614
rect 427222 212378 427306 212614
rect 427542 212378 427574 212614
rect 426954 212294 427574 212378
rect 426954 212058 426986 212294
rect 427222 212058 427306 212294
rect 427542 212058 427574 212294
rect 426954 176614 427574 212058
rect 426954 176378 426986 176614
rect 427222 176378 427306 176614
rect 427542 176378 427574 176614
rect 426954 176294 427574 176378
rect 426954 176058 426986 176294
rect 427222 176058 427306 176294
rect 427542 176058 427574 176294
rect 426954 142000 427574 176058
rect 433794 704838 434414 705830
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 433794 507454 434414 542898
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 471454 434414 506898
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 435454 434414 470898
rect 433794 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 434414 435454
rect 433794 435134 434414 435218
rect 433794 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 434414 435134
rect 433794 399454 434414 434898
rect 433794 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 434414 399454
rect 433794 399134 434414 399218
rect 433794 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 434414 399134
rect 433794 363454 434414 398898
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 433794 327454 434414 362898
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 433794 291454 434414 326898
rect 433794 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 434414 291454
rect 433794 291134 434414 291218
rect 433794 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 434414 291134
rect 433794 255454 434414 290898
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 219454 434414 254898
rect 433794 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 434414 219454
rect 433794 219134 434414 219218
rect 433794 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 434414 219134
rect 433794 183454 434414 218898
rect 433794 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 434414 183454
rect 433794 183134 434414 183218
rect 433794 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 434414 183134
rect 433794 147454 434414 182898
rect 433794 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 434414 147454
rect 433794 147134 434414 147218
rect 433794 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 434414 147134
rect 431907 142220 431973 142221
rect 431907 142156 431908 142220
rect 431972 142156 431973 142220
rect 431907 142155 431973 142156
rect 426387 139500 426453 139501
rect 426387 139436 426388 139500
rect 426452 139436 426453 139500
rect 426387 139435 426453 139436
rect 427859 139500 427925 139501
rect 427859 139436 427860 139500
rect 427924 139436 427925 139500
rect 427859 139435 427925 139436
rect 429147 139500 429213 139501
rect 429147 139436 429148 139500
rect 429212 139436 429213 139500
rect 429147 139435 429213 139436
rect 423995 100740 424061 100741
rect 423995 100676 423996 100740
rect 424060 100676 424061 100740
rect 423995 100675 424061 100676
rect 425651 100740 425717 100741
rect 425651 100676 425652 100740
rect 425716 100676 425717 100740
rect 425651 100675 425717 100676
rect 421051 73812 421117 73813
rect 421051 73748 421052 73812
rect 421116 73748 421117 73812
rect 421051 73747 421117 73748
rect 419514 60938 419546 61174
rect 419782 60938 419866 61174
rect 420102 60938 420134 61174
rect 419514 60854 420134 60938
rect 419514 60618 419546 60854
rect 419782 60618 419866 60854
rect 420102 60618 420134 60854
rect 419514 25174 420134 60618
rect 419514 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 420134 25174
rect 419514 24854 420134 24938
rect 419514 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 420134 24854
rect 419027 23356 419093 23357
rect 419027 23292 419028 23356
rect 419092 23292 419093 23356
rect 419027 23291 419093 23292
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -1306 416414 20898
rect 415794 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 416414 -1306
rect 415794 -1626 416414 -1542
rect 415794 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 416414 -1626
rect 415794 -1894 416414 -1862
rect 419514 -3226 420134 24618
rect 419514 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 420134 -3226
rect 419514 -3546 420134 -3462
rect 419514 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 420134 -3546
rect 419514 -3814 420134 -3782
rect 423234 64894 423854 98000
rect 423234 64658 423266 64894
rect 423502 64658 423586 64894
rect 423822 64658 423854 64894
rect 423234 64574 423854 64658
rect 423234 64338 423266 64574
rect 423502 64338 423586 64574
rect 423822 64338 423854 64574
rect 423234 28894 423854 64338
rect 426390 33149 426450 139435
rect 426544 111454 426864 111486
rect 426544 111218 426586 111454
rect 426822 111218 426864 111454
rect 426544 111134 426864 111218
rect 426544 110898 426586 111134
rect 426822 110898 426864 111134
rect 426544 110866 426864 110898
rect 426954 68614 427574 98000
rect 426954 68378 426986 68614
rect 427222 68378 427306 68614
rect 427542 68378 427574 68614
rect 426954 68294 427574 68378
rect 426954 68058 426986 68294
rect 427222 68058 427306 68294
rect 427542 68058 427574 68294
rect 426387 33148 426453 33149
rect 426387 33084 426388 33148
rect 426452 33084 426453 33148
rect 426387 33083 426453 33084
rect 423234 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 423854 28894
rect 423234 28574 423854 28658
rect 423234 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 423854 28574
rect 423234 -5146 423854 28338
rect 423234 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 423854 -5146
rect 423234 -5466 423854 -5382
rect 423234 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 423854 -5466
rect 423234 -5734 423854 -5702
rect 426954 32614 427574 68058
rect 426954 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 427574 32614
rect 426954 32294 427574 32378
rect 426954 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 427574 32294
rect 408954 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 409574 -6106
rect 408954 -6426 409574 -6342
rect 408954 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 409574 -6426
rect 408954 -7654 409574 -6662
rect 426954 -7066 427574 32058
rect 427862 17917 427922 139435
rect 428144 129454 428464 129486
rect 428144 129218 428186 129454
rect 428422 129218 428464 129454
rect 428144 129134 428464 129218
rect 428144 128898 428186 129134
rect 428422 128898 428464 129134
rect 428144 128866 428464 128898
rect 429150 53141 429210 139435
rect 431910 138030 431970 142155
rect 433794 142000 434414 146898
rect 437514 691174 438134 706202
rect 437514 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 438134 691174
rect 437514 690854 438134 690938
rect 437514 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 438134 690854
rect 437514 655174 438134 690618
rect 437514 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 438134 655174
rect 437514 654854 438134 654938
rect 437514 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 438134 654854
rect 437514 619174 438134 654618
rect 437514 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 438134 619174
rect 437514 618854 438134 618938
rect 437514 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 438134 618854
rect 437514 583174 438134 618618
rect 437514 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 438134 583174
rect 437514 582854 438134 582938
rect 437514 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 438134 582854
rect 437514 547174 438134 582618
rect 437514 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 438134 547174
rect 437514 546854 438134 546938
rect 437514 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 438134 546854
rect 437514 511174 438134 546618
rect 437514 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 438134 511174
rect 437514 510854 438134 510938
rect 437514 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 438134 510854
rect 437514 475174 438134 510618
rect 437514 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 438134 475174
rect 437514 474854 438134 474938
rect 437514 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 438134 474854
rect 437514 439174 438134 474618
rect 437514 438938 437546 439174
rect 437782 438938 437866 439174
rect 438102 438938 438134 439174
rect 437514 438854 438134 438938
rect 437514 438618 437546 438854
rect 437782 438618 437866 438854
rect 438102 438618 438134 438854
rect 437514 403174 438134 438618
rect 437514 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 438134 403174
rect 437514 402854 438134 402938
rect 437514 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 438134 402854
rect 437514 367174 438134 402618
rect 437514 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 438134 367174
rect 437514 366854 438134 366938
rect 437514 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 438134 366854
rect 437514 331174 438134 366618
rect 437514 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 438134 331174
rect 437514 330854 438134 330938
rect 437514 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 438134 330854
rect 437514 295174 438134 330618
rect 437514 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 438134 295174
rect 437514 294854 438134 294938
rect 437514 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 438134 294854
rect 437514 259174 438134 294618
rect 441234 694894 441854 708122
rect 441234 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 441854 694894
rect 441234 694574 441854 694658
rect 441234 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 441854 694574
rect 441234 658894 441854 694338
rect 441234 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 441854 658894
rect 441234 658574 441854 658658
rect 441234 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 441854 658574
rect 441234 622894 441854 658338
rect 441234 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 441854 622894
rect 441234 622574 441854 622658
rect 441234 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 441854 622574
rect 441234 586894 441854 622338
rect 441234 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 441854 586894
rect 441234 586574 441854 586658
rect 441234 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 441854 586574
rect 441234 550894 441854 586338
rect 441234 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 441854 550894
rect 441234 550574 441854 550658
rect 441234 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 441854 550574
rect 441234 514894 441854 550338
rect 441234 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 441854 514894
rect 441234 514574 441854 514658
rect 441234 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 441854 514574
rect 441234 478894 441854 514338
rect 441234 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 441854 478894
rect 441234 478574 441854 478658
rect 441234 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 441854 478574
rect 441234 442894 441854 478338
rect 441234 442658 441266 442894
rect 441502 442658 441586 442894
rect 441822 442658 441854 442894
rect 441234 442574 441854 442658
rect 441234 442338 441266 442574
rect 441502 442338 441586 442574
rect 441822 442338 441854 442574
rect 441234 406894 441854 442338
rect 441234 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 441854 406894
rect 441234 406574 441854 406658
rect 441234 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 441854 406574
rect 441234 370894 441854 406338
rect 441234 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 441854 370894
rect 441234 370574 441854 370658
rect 441234 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 441854 370574
rect 441234 334894 441854 370338
rect 441234 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 441854 334894
rect 441234 334574 441854 334658
rect 441234 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 441854 334574
rect 441234 298894 441854 334338
rect 441234 298658 441266 298894
rect 441502 298658 441586 298894
rect 441822 298658 441854 298894
rect 441234 298574 441854 298658
rect 441234 298338 441266 298574
rect 441502 298338 441586 298574
rect 441822 298338 441854 298574
rect 438899 286380 438965 286381
rect 438899 286316 438900 286380
rect 438964 286316 438965 286380
rect 438899 286315 438965 286316
rect 437514 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 438134 259174
rect 437514 258854 438134 258938
rect 437514 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 438134 258854
rect 437514 223174 438134 258618
rect 437514 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 438134 223174
rect 437514 222854 438134 222938
rect 437514 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 438134 222854
rect 437514 187174 438134 222618
rect 437514 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 438134 187174
rect 437514 186854 438134 186938
rect 437514 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 438134 186854
rect 437514 151174 438134 186618
rect 437514 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 438134 151174
rect 437514 150854 438134 150938
rect 437514 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 438134 150854
rect 437514 142000 438134 150618
rect 435035 139500 435101 139501
rect 435035 139436 435036 139500
rect 435100 139436 435101 139500
rect 435035 139435 435101 139436
rect 431726 137970 431970 138030
rect 431344 129454 431664 129486
rect 431344 129218 431386 129454
rect 431622 129218 431664 129454
rect 431344 129134 431664 129218
rect 431344 128898 431386 129134
rect 431622 128898 431664 129134
rect 431344 128866 431664 128898
rect 429744 111454 430064 111486
rect 429744 111218 429786 111454
rect 430022 111218 430064 111454
rect 429744 111134 430064 111218
rect 429744 110898 429786 111134
rect 430022 110898 430064 111134
rect 429744 110866 430064 110898
rect 431726 65517 431786 137970
rect 434544 129454 434864 129486
rect 434544 129218 434586 129454
rect 434822 129218 434864 129454
rect 434544 129134 434864 129218
rect 434544 128898 434586 129134
rect 434822 128898 434864 129134
rect 434544 128866 434864 128898
rect 432944 111454 433264 111486
rect 432944 111218 432986 111454
rect 433222 111218 433264 111454
rect 432944 111134 433264 111218
rect 432944 110898 432986 111134
rect 433222 110898 433264 111134
rect 432944 110866 433264 110898
rect 433794 75454 434414 98000
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 431723 65516 431789 65517
rect 431723 65452 431724 65516
rect 431788 65452 431789 65516
rect 431723 65451 431789 65452
rect 429147 53140 429213 53141
rect 429147 53076 429148 53140
rect 429212 53076 429213 53140
rect 429147 53075 429213 53076
rect 433794 39454 434414 74898
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 427859 17916 427925 17917
rect 427859 17852 427860 17916
rect 427924 17852 427925 17916
rect 427859 17851 427925 17852
rect 433794 3454 434414 38898
rect 435038 24173 435098 139435
rect 437744 129454 438064 129486
rect 437744 129218 437786 129454
rect 438022 129218 438064 129454
rect 437744 129134 438064 129218
rect 437744 128898 437786 129134
rect 438022 128898 438064 129134
rect 437744 128866 438064 128898
rect 438902 125490 438962 286315
rect 441234 262894 441854 298338
rect 441234 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 441854 262894
rect 441234 262574 441854 262658
rect 441234 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 441854 262574
rect 441234 226894 441854 262338
rect 441234 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 441854 226894
rect 441234 226574 441854 226658
rect 441234 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 441854 226574
rect 441234 190894 441854 226338
rect 444954 698614 445574 710042
rect 462954 711558 463574 711590
rect 462954 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 463574 711558
rect 462954 711238 463574 711322
rect 462954 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 463574 711238
rect 459234 709638 459854 709670
rect 459234 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 459854 709638
rect 459234 709318 459854 709402
rect 459234 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 459854 709318
rect 455514 707718 456134 707750
rect 455514 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 456134 707718
rect 455514 707398 456134 707482
rect 455514 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 456134 707398
rect 444954 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 445574 698614
rect 444954 698294 445574 698378
rect 444954 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 445574 698294
rect 444954 662614 445574 698058
rect 444954 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 445574 662614
rect 444954 662294 445574 662378
rect 444954 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 445574 662294
rect 444954 626614 445574 662058
rect 444954 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 445574 626614
rect 444954 626294 445574 626378
rect 444954 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 445574 626294
rect 444954 590614 445574 626058
rect 444954 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 445574 590614
rect 444954 590294 445574 590378
rect 444954 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 445574 590294
rect 444954 554614 445574 590058
rect 444954 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 445574 554614
rect 444954 554294 445574 554378
rect 444954 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 445574 554294
rect 444954 518614 445574 554058
rect 444954 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 445574 518614
rect 444954 518294 445574 518378
rect 444954 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 445574 518294
rect 444954 482614 445574 518058
rect 444954 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 445574 482614
rect 444954 482294 445574 482378
rect 444954 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 445574 482294
rect 444954 446614 445574 482058
rect 444954 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 445574 446614
rect 444954 446294 445574 446378
rect 444954 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 445574 446294
rect 444954 410614 445574 446058
rect 444954 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 445574 410614
rect 444954 410294 445574 410378
rect 444954 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 445574 410294
rect 444954 374614 445574 410058
rect 444954 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 445574 374614
rect 444954 374294 445574 374378
rect 444954 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 445574 374294
rect 444954 338614 445574 374058
rect 444954 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 445574 338614
rect 444954 338294 445574 338378
rect 444954 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 445574 338294
rect 444954 302614 445574 338058
rect 444954 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 445574 302614
rect 444954 302294 445574 302378
rect 444954 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 445574 302294
rect 444954 266614 445574 302058
rect 444954 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 445574 266614
rect 444954 266294 445574 266378
rect 444954 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 445574 266294
rect 444954 230614 445574 266058
rect 444954 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 445574 230614
rect 444954 230294 445574 230378
rect 444954 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 445574 230294
rect 442027 215932 442093 215933
rect 442027 215868 442028 215932
rect 442092 215868 442093 215932
rect 442027 215867 442093 215868
rect 441234 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 441854 190894
rect 441234 190574 441854 190658
rect 441234 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 441854 190574
rect 441234 154894 441854 190338
rect 441234 154658 441266 154894
rect 441502 154658 441586 154894
rect 441822 154658 441854 154894
rect 441234 154574 441854 154658
rect 441234 154338 441266 154574
rect 441502 154338 441586 154574
rect 441822 154338 441854 154574
rect 441234 142000 441854 154338
rect 441659 140860 441725 140861
rect 441659 140796 441660 140860
rect 441724 140796 441725 140860
rect 441659 140795 441725 140796
rect 439083 139500 439149 139501
rect 439083 139436 439084 139500
rect 439148 139436 439149 139500
rect 439083 139435 439149 139436
rect 439086 125610 439146 139435
rect 441662 138685 441722 140795
rect 441659 138684 441725 138685
rect 441659 138620 441660 138684
rect 441724 138620 441725 138684
rect 441659 138619 441725 138620
rect 439086 125550 439698 125610
rect 438902 125430 439146 125490
rect 439086 125082 439146 125430
rect 439086 125022 439514 125082
rect 439267 120596 439333 120597
rect 439267 120532 439268 120596
rect 439332 120532 439333 120596
rect 439267 120531 439333 120532
rect 439270 119370 439330 120531
rect 438902 119310 439330 119370
rect 438902 115950 438962 119310
rect 439454 115970 439514 125022
rect 439638 120597 439698 125550
rect 439635 120596 439701 120597
rect 439635 120532 439636 120596
rect 439700 120532 439701 120596
rect 439635 120531 439701 120532
rect 438902 115890 439146 115950
rect 436144 111454 436464 111486
rect 436144 111218 436186 111454
rect 436422 111218 436464 111454
rect 436144 111134 436464 111218
rect 436144 110898 436186 111134
rect 436422 110898 436464 111134
rect 436144 110866 436464 110898
rect 437514 79174 438134 98000
rect 437514 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 438134 79174
rect 437514 78854 438134 78938
rect 437514 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 438134 78854
rect 437514 43174 438134 78618
rect 437514 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 438134 43174
rect 437514 42854 438134 42938
rect 437514 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 438134 42854
rect 435035 24172 435101 24173
rect 435035 24108 435036 24172
rect 435100 24108 435101 24172
rect 435035 24107 435101 24108
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -1894 434414 -902
rect 437514 7174 438134 42618
rect 439086 9621 439146 115890
rect 439270 115910 439514 115970
rect 439270 113117 439330 115910
rect 439267 113116 439333 113117
rect 439267 113052 439268 113116
rect 439332 113052 439333 113116
rect 439267 113051 439333 113052
rect 442030 105365 442090 215867
rect 444954 194614 445574 230058
rect 444954 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 445574 194614
rect 444954 194294 445574 194378
rect 444954 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 445574 194294
rect 444954 158614 445574 194058
rect 444954 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 445574 158614
rect 444954 158294 445574 158378
rect 444954 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 445574 158294
rect 442211 125084 442277 125085
rect 442211 125020 442212 125084
rect 442276 125020 442277 125084
rect 442211 125019 442277 125020
rect 442027 105364 442093 105365
rect 442027 105300 442028 105364
rect 442092 105300 442093 105364
rect 442027 105299 442093 105300
rect 441234 82894 441854 98000
rect 442214 95845 442274 125019
rect 444954 122614 445574 158058
rect 444954 122378 444986 122614
rect 445222 122378 445306 122614
rect 445542 122378 445574 122614
rect 444954 122294 445574 122378
rect 444954 122058 444986 122294
rect 445222 122058 445306 122294
rect 445542 122058 445574 122294
rect 442211 95844 442277 95845
rect 442211 95780 442212 95844
rect 442276 95780 442277 95844
rect 442211 95779 442277 95780
rect 441234 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 441854 82894
rect 441234 82574 441854 82658
rect 441234 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 441854 82574
rect 441234 46894 441854 82338
rect 441234 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 441854 46894
rect 441234 46574 441854 46658
rect 441234 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 441854 46574
rect 441234 10894 441854 46338
rect 441234 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 441854 10894
rect 441234 10574 441854 10658
rect 441234 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 441854 10574
rect 439083 9620 439149 9621
rect 439083 9556 439084 9620
rect 439148 9556 439149 9620
rect 439083 9555 439149 9556
rect 437514 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 438134 7174
rect 437514 6854 438134 6938
rect 437514 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 438134 6854
rect 437514 -2266 438134 6618
rect 437514 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 438134 -2266
rect 437514 -2586 438134 -2502
rect 437514 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 438134 -2586
rect 437514 -3814 438134 -2822
rect 441234 -4186 441854 10338
rect 441234 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 441854 -4186
rect 441234 -4506 441854 -4422
rect 441234 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 441854 -4506
rect 441234 -5734 441854 -4742
rect 444954 86614 445574 122058
rect 444954 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 445574 86614
rect 444954 86294 445574 86378
rect 444954 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 445574 86294
rect 444954 50614 445574 86058
rect 444954 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 445574 50614
rect 444954 50294 445574 50378
rect 444954 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 445574 50294
rect 444954 14614 445574 50058
rect 444954 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 445574 14614
rect 444954 14294 445574 14378
rect 444954 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 445574 14294
rect 426954 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 427574 -7066
rect 426954 -7386 427574 -7302
rect 426954 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 427574 -7386
rect 426954 -7654 427574 -7622
rect 444954 -6106 445574 14058
rect 451794 705798 452414 705830
rect 451794 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 452414 705798
rect 451794 705478 452414 705562
rect 451794 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 452414 705478
rect 451794 669454 452414 705242
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597454 452414 632898
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 561454 452414 596898
rect 451794 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 452414 561454
rect 451794 561134 452414 561218
rect 451794 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 452414 561134
rect 451794 525454 452414 560898
rect 451794 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 452414 525454
rect 451794 525134 452414 525218
rect 451794 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 452414 525134
rect 451794 489454 452414 524898
rect 451794 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 452414 489454
rect 451794 489134 452414 489218
rect 451794 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 452414 489134
rect 451794 453454 452414 488898
rect 451794 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 452414 453454
rect 451794 453134 452414 453218
rect 451794 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 452414 453134
rect 451794 417454 452414 452898
rect 451794 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 452414 417454
rect 451794 417134 452414 417218
rect 451794 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 452414 417134
rect 451794 381454 452414 416898
rect 451794 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 452414 381454
rect 451794 381134 452414 381218
rect 451794 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 452414 381134
rect 451794 345454 452414 380898
rect 451794 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 452414 345454
rect 451794 345134 452414 345218
rect 451794 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 452414 345134
rect 451794 309454 452414 344898
rect 451794 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 452414 309454
rect 451794 309134 452414 309218
rect 451794 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 452414 309134
rect 451794 273454 452414 308898
rect 451794 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 452414 273454
rect 451794 273134 452414 273218
rect 451794 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 452414 273134
rect 451794 237454 452414 272898
rect 451794 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 452414 237454
rect 451794 237134 452414 237218
rect 451794 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 452414 237134
rect 451794 201454 452414 236898
rect 451794 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 452414 201454
rect 451794 201134 452414 201218
rect 451794 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 452414 201134
rect 451794 165454 452414 200898
rect 451794 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 452414 165454
rect 451794 165134 452414 165218
rect 451794 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 452414 165134
rect 451794 129454 452414 164898
rect 451794 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 452414 129454
rect 451794 129134 452414 129218
rect 451794 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 452414 129134
rect 451794 93454 452414 128898
rect 451794 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 452414 93454
rect 451794 93134 452414 93218
rect 451794 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 452414 93134
rect 451794 57454 452414 92898
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -1306 452414 20898
rect 451794 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 452414 -1306
rect 451794 -1626 452414 -1542
rect 451794 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 452414 -1626
rect 451794 -1894 452414 -1862
rect 455514 673174 456134 707162
rect 455514 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 456134 673174
rect 455514 672854 456134 672938
rect 455514 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 456134 672854
rect 455514 637174 456134 672618
rect 455514 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 456134 637174
rect 455514 636854 456134 636938
rect 455514 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 456134 636854
rect 455514 601174 456134 636618
rect 455514 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 456134 601174
rect 455514 600854 456134 600938
rect 455514 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 456134 600854
rect 455514 565174 456134 600618
rect 455514 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 456134 565174
rect 455514 564854 456134 564938
rect 455514 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 456134 564854
rect 455514 529174 456134 564618
rect 455514 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 456134 529174
rect 455514 528854 456134 528938
rect 455514 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 456134 528854
rect 455514 493174 456134 528618
rect 455514 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 456134 493174
rect 455514 492854 456134 492938
rect 455514 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 456134 492854
rect 455514 457174 456134 492618
rect 455514 456938 455546 457174
rect 455782 456938 455866 457174
rect 456102 456938 456134 457174
rect 455514 456854 456134 456938
rect 455514 456618 455546 456854
rect 455782 456618 455866 456854
rect 456102 456618 456134 456854
rect 455514 421174 456134 456618
rect 455514 420938 455546 421174
rect 455782 420938 455866 421174
rect 456102 420938 456134 421174
rect 455514 420854 456134 420938
rect 455514 420618 455546 420854
rect 455782 420618 455866 420854
rect 456102 420618 456134 420854
rect 455514 385174 456134 420618
rect 455514 384938 455546 385174
rect 455782 384938 455866 385174
rect 456102 384938 456134 385174
rect 455514 384854 456134 384938
rect 455514 384618 455546 384854
rect 455782 384618 455866 384854
rect 456102 384618 456134 384854
rect 455514 349174 456134 384618
rect 455514 348938 455546 349174
rect 455782 348938 455866 349174
rect 456102 348938 456134 349174
rect 455514 348854 456134 348938
rect 455514 348618 455546 348854
rect 455782 348618 455866 348854
rect 456102 348618 456134 348854
rect 455514 313174 456134 348618
rect 455514 312938 455546 313174
rect 455782 312938 455866 313174
rect 456102 312938 456134 313174
rect 455514 312854 456134 312938
rect 455514 312618 455546 312854
rect 455782 312618 455866 312854
rect 456102 312618 456134 312854
rect 455514 277174 456134 312618
rect 455514 276938 455546 277174
rect 455782 276938 455866 277174
rect 456102 276938 456134 277174
rect 455514 276854 456134 276938
rect 455514 276618 455546 276854
rect 455782 276618 455866 276854
rect 456102 276618 456134 276854
rect 455514 241174 456134 276618
rect 455514 240938 455546 241174
rect 455782 240938 455866 241174
rect 456102 240938 456134 241174
rect 455514 240854 456134 240938
rect 455514 240618 455546 240854
rect 455782 240618 455866 240854
rect 456102 240618 456134 240854
rect 455514 205174 456134 240618
rect 455514 204938 455546 205174
rect 455782 204938 455866 205174
rect 456102 204938 456134 205174
rect 455514 204854 456134 204938
rect 455514 204618 455546 204854
rect 455782 204618 455866 204854
rect 456102 204618 456134 204854
rect 455514 169174 456134 204618
rect 455514 168938 455546 169174
rect 455782 168938 455866 169174
rect 456102 168938 456134 169174
rect 455514 168854 456134 168938
rect 455514 168618 455546 168854
rect 455782 168618 455866 168854
rect 456102 168618 456134 168854
rect 455514 133174 456134 168618
rect 455514 132938 455546 133174
rect 455782 132938 455866 133174
rect 456102 132938 456134 133174
rect 455514 132854 456134 132938
rect 455514 132618 455546 132854
rect 455782 132618 455866 132854
rect 456102 132618 456134 132854
rect 455514 97174 456134 132618
rect 455514 96938 455546 97174
rect 455782 96938 455866 97174
rect 456102 96938 456134 97174
rect 455514 96854 456134 96938
rect 455514 96618 455546 96854
rect 455782 96618 455866 96854
rect 456102 96618 456134 96854
rect 455514 61174 456134 96618
rect 455514 60938 455546 61174
rect 455782 60938 455866 61174
rect 456102 60938 456134 61174
rect 455514 60854 456134 60938
rect 455514 60618 455546 60854
rect 455782 60618 455866 60854
rect 456102 60618 456134 60854
rect 455514 25174 456134 60618
rect 455514 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 456134 25174
rect 455514 24854 456134 24938
rect 455514 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 456134 24854
rect 455514 -3226 456134 24618
rect 455514 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 456134 -3226
rect 455514 -3546 456134 -3462
rect 455514 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 456134 -3546
rect 455514 -3814 456134 -3782
rect 459234 676894 459854 709082
rect 459234 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 459854 676894
rect 459234 676574 459854 676658
rect 459234 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 459854 676574
rect 459234 640894 459854 676338
rect 459234 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 459854 640894
rect 459234 640574 459854 640658
rect 459234 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 459854 640574
rect 459234 604894 459854 640338
rect 459234 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 459854 604894
rect 459234 604574 459854 604658
rect 459234 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 459854 604574
rect 459234 568894 459854 604338
rect 459234 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 459854 568894
rect 459234 568574 459854 568658
rect 459234 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 459854 568574
rect 459234 532894 459854 568338
rect 459234 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 459854 532894
rect 459234 532574 459854 532658
rect 459234 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 459854 532574
rect 459234 496894 459854 532338
rect 459234 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 459854 496894
rect 459234 496574 459854 496658
rect 459234 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 459854 496574
rect 459234 460894 459854 496338
rect 459234 460658 459266 460894
rect 459502 460658 459586 460894
rect 459822 460658 459854 460894
rect 459234 460574 459854 460658
rect 459234 460338 459266 460574
rect 459502 460338 459586 460574
rect 459822 460338 459854 460574
rect 459234 424894 459854 460338
rect 459234 424658 459266 424894
rect 459502 424658 459586 424894
rect 459822 424658 459854 424894
rect 459234 424574 459854 424658
rect 459234 424338 459266 424574
rect 459502 424338 459586 424574
rect 459822 424338 459854 424574
rect 459234 388894 459854 424338
rect 459234 388658 459266 388894
rect 459502 388658 459586 388894
rect 459822 388658 459854 388894
rect 459234 388574 459854 388658
rect 459234 388338 459266 388574
rect 459502 388338 459586 388574
rect 459822 388338 459854 388574
rect 459234 352894 459854 388338
rect 459234 352658 459266 352894
rect 459502 352658 459586 352894
rect 459822 352658 459854 352894
rect 459234 352574 459854 352658
rect 459234 352338 459266 352574
rect 459502 352338 459586 352574
rect 459822 352338 459854 352574
rect 459234 316894 459854 352338
rect 459234 316658 459266 316894
rect 459502 316658 459586 316894
rect 459822 316658 459854 316894
rect 459234 316574 459854 316658
rect 459234 316338 459266 316574
rect 459502 316338 459586 316574
rect 459822 316338 459854 316574
rect 459234 280894 459854 316338
rect 459234 280658 459266 280894
rect 459502 280658 459586 280894
rect 459822 280658 459854 280894
rect 459234 280574 459854 280658
rect 459234 280338 459266 280574
rect 459502 280338 459586 280574
rect 459822 280338 459854 280574
rect 459234 244894 459854 280338
rect 459234 244658 459266 244894
rect 459502 244658 459586 244894
rect 459822 244658 459854 244894
rect 459234 244574 459854 244658
rect 459234 244338 459266 244574
rect 459502 244338 459586 244574
rect 459822 244338 459854 244574
rect 459234 208894 459854 244338
rect 459234 208658 459266 208894
rect 459502 208658 459586 208894
rect 459822 208658 459854 208894
rect 459234 208574 459854 208658
rect 459234 208338 459266 208574
rect 459502 208338 459586 208574
rect 459822 208338 459854 208574
rect 459234 172894 459854 208338
rect 459234 172658 459266 172894
rect 459502 172658 459586 172894
rect 459822 172658 459854 172894
rect 459234 172574 459854 172658
rect 459234 172338 459266 172574
rect 459502 172338 459586 172574
rect 459822 172338 459854 172574
rect 459234 136894 459854 172338
rect 459234 136658 459266 136894
rect 459502 136658 459586 136894
rect 459822 136658 459854 136894
rect 459234 136574 459854 136658
rect 459234 136338 459266 136574
rect 459502 136338 459586 136574
rect 459822 136338 459854 136574
rect 459234 100894 459854 136338
rect 459234 100658 459266 100894
rect 459502 100658 459586 100894
rect 459822 100658 459854 100894
rect 459234 100574 459854 100658
rect 459234 100338 459266 100574
rect 459502 100338 459586 100574
rect 459822 100338 459854 100574
rect 459234 64894 459854 100338
rect 459234 64658 459266 64894
rect 459502 64658 459586 64894
rect 459822 64658 459854 64894
rect 459234 64574 459854 64658
rect 459234 64338 459266 64574
rect 459502 64338 459586 64574
rect 459822 64338 459854 64574
rect 459234 28894 459854 64338
rect 459234 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 459854 28894
rect 459234 28574 459854 28658
rect 459234 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 459854 28574
rect 459234 -5146 459854 28338
rect 459234 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 459854 -5146
rect 459234 -5466 459854 -5382
rect 459234 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 459854 -5466
rect 459234 -5734 459854 -5702
rect 462954 680614 463574 711002
rect 480954 710598 481574 711590
rect 480954 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 481574 710598
rect 480954 710278 481574 710362
rect 480954 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 481574 710278
rect 477234 708678 477854 709670
rect 477234 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 477854 708678
rect 477234 708358 477854 708442
rect 477234 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 477854 708358
rect 473514 706758 474134 707750
rect 473514 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 474134 706758
rect 473514 706438 474134 706522
rect 473514 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 474134 706438
rect 462954 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 463574 680614
rect 462954 680294 463574 680378
rect 462954 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 463574 680294
rect 462954 644614 463574 680058
rect 462954 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 463574 644614
rect 462954 644294 463574 644378
rect 462954 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 463574 644294
rect 462954 608614 463574 644058
rect 462954 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 463574 608614
rect 462954 608294 463574 608378
rect 462954 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 463574 608294
rect 462954 572614 463574 608058
rect 462954 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 463574 572614
rect 462954 572294 463574 572378
rect 462954 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 463574 572294
rect 462954 536614 463574 572058
rect 462954 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 463574 536614
rect 462954 536294 463574 536378
rect 462954 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 463574 536294
rect 462954 500614 463574 536058
rect 462954 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 463574 500614
rect 462954 500294 463574 500378
rect 462954 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 463574 500294
rect 462954 464614 463574 500058
rect 462954 464378 462986 464614
rect 463222 464378 463306 464614
rect 463542 464378 463574 464614
rect 462954 464294 463574 464378
rect 462954 464058 462986 464294
rect 463222 464058 463306 464294
rect 463542 464058 463574 464294
rect 462954 428614 463574 464058
rect 462954 428378 462986 428614
rect 463222 428378 463306 428614
rect 463542 428378 463574 428614
rect 462954 428294 463574 428378
rect 462954 428058 462986 428294
rect 463222 428058 463306 428294
rect 463542 428058 463574 428294
rect 462954 392614 463574 428058
rect 462954 392378 462986 392614
rect 463222 392378 463306 392614
rect 463542 392378 463574 392614
rect 462954 392294 463574 392378
rect 462954 392058 462986 392294
rect 463222 392058 463306 392294
rect 463542 392058 463574 392294
rect 462954 356614 463574 392058
rect 462954 356378 462986 356614
rect 463222 356378 463306 356614
rect 463542 356378 463574 356614
rect 462954 356294 463574 356378
rect 462954 356058 462986 356294
rect 463222 356058 463306 356294
rect 463542 356058 463574 356294
rect 462954 320614 463574 356058
rect 462954 320378 462986 320614
rect 463222 320378 463306 320614
rect 463542 320378 463574 320614
rect 462954 320294 463574 320378
rect 462954 320058 462986 320294
rect 463222 320058 463306 320294
rect 463542 320058 463574 320294
rect 462954 284614 463574 320058
rect 462954 284378 462986 284614
rect 463222 284378 463306 284614
rect 463542 284378 463574 284614
rect 462954 284294 463574 284378
rect 462954 284058 462986 284294
rect 463222 284058 463306 284294
rect 463542 284058 463574 284294
rect 462954 248614 463574 284058
rect 462954 248378 462986 248614
rect 463222 248378 463306 248614
rect 463542 248378 463574 248614
rect 462954 248294 463574 248378
rect 462954 248058 462986 248294
rect 463222 248058 463306 248294
rect 463542 248058 463574 248294
rect 462954 212614 463574 248058
rect 462954 212378 462986 212614
rect 463222 212378 463306 212614
rect 463542 212378 463574 212614
rect 462954 212294 463574 212378
rect 462954 212058 462986 212294
rect 463222 212058 463306 212294
rect 463542 212058 463574 212294
rect 462954 176614 463574 212058
rect 462954 176378 462986 176614
rect 463222 176378 463306 176614
rect 463542 176378 463574 176614
rect 462954 176294 463574 176378
rect 462954 176058 462986 176294
rect 463222 176058 463306 176294
rect 463542 176058 463574 176294
rect 462954 140614 463574 176058
rect 462954 140378 462986 140614
rect 463222 140378 463306 140614
rect 463542 140378 463574 140614
rect 462954 140294 463574 140378
rect 462954 140058 462986 140294
rect 463222 140058 463306 140294
rect 463542 140058 463574 140294
rect 462954 104614 463574 140058
rect 462954 104378 462986 104614
rect 463222 104378 463306 104614
rect 463542 104378 463574 104614
rect 462954 104294 463574 104378
rect 462954 104058 462986 104294
rect 463222 104058 463306 104294
rect 463542 104058 463574 104294
rect 462954 68614 463574 104058
rect 462954 68378 462986 68614
rect 463222 68378 463306 68614
rect 463542 68378 463574 68614
rect 462954 68294 463574 68378
rect 462954 68058 462986 68294
rect 463222 68058 463306 68294
rect 463542 68058 463574 68294
rect 462954 32614 463574 68058
rect 462954 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 463574 32614
rect 462954 32294 463574 32378
rect 462954 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 463574 32294
rect 444954 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 445574 -6106
rect 444954 -6426 445574 -6342
rect 444954 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 445574 -6426
rect 444954 -7654 445574 -6662
rect 462954 -7066 463574 32058
rect 469794 704838 470414 705830
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 579454 470414 614898
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 399454 470414 434898
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 469794 363454 470414 398898
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 469794 327454 470414 362898
rect 469794 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 470414 327454
rect 469794 327134 470414 327218
rect 469794 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 470414 327134
rect 469794 291454 470414 326898
rect 469794 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 470414 291454
rect 469794 291134 470414 291218
rect 469794 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 470414 291134
rect 469794 255454 470414 290898
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 219454 470414 254898
rect 469794 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 470414 219454
rect 469794 219134 470414 219218
rect 469794 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 470414 219134
rect 469794 183454 470414 218898
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 147454 470414 182898
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 111454 470414 146898
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -1894 470414 -902
rect 473514 691174 474134 706202
rect 473514 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 474134 691174
rect 473514 690854 474134 690938
rect 473514 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 474134 690854
rect 473514 655174 474134 690618
rect 473514 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 474134 655174
rect 473514 654854 474134 654938
rect 473514 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 474134 654854
rect 473514 619174 474134 654618
rect 473514 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 474134 619174
rect 473514 618854 474134 618938
rect 473514 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 474134 618854
rect 473514 583174 474134 618618
rect 473514 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 474134 583174
rect 473514 582854 474134 582938
rect 473514 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 474134 582854
rect 473514 547174 474134 582618
rect 473514 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 474134 547174
rect 473514 546854 474134 546938
rect 473514 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 474134 546854
rect 473514 511174 474134 546618
rect 473514 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 474134 511174
rect 473514 510854 474134 510938
rect 473514 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 474134 510854
rect 473514 475174 474134 510618
rect 473514 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 474134 475174
rect 473514 474854 474134 474938
rect 473514 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 474134 474854
rect 473514 439174 474134 474618
rect 473514 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 474134 439174
rect 473514 438854 474134 438938
rect 473514 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 474134 438854
rect 473514 403174 474134 438618
rect 473514 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 474134 403174
rect 473514 402854 474134 402938
rect 473514 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 474134 402854
rect 473514 367174 474134 402618
rect 473514 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 474134 367174
rect 473514 366854 474134 366938
rect 473514 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 474134 366854
rect 473514 331174 474134 366618
rect 473514 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 474134 331174
rect 473514 330854 474134 330938
rect 473514 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 474134 330854
rect 473514 295174 474134 330618
rect 473514 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 474134 295174
rect 473514 294854 474134 294938
rect 473514 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 474134 294854
rect 473514 259174 474134 294618
rect 473514 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 474134 259174
rect 473514 258854 474134 258938
rect 473514 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 474134 258854
rect 473514 223174 474134 258618
rect 473514 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 474134 223174
rect 473514 222854 474134 222938
rect 473514 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 474134 222854
rect 473514 187174 474134 222618
rect 473514 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 474134 187174
rect 473514 186854 474134 186938
rect 473514 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 474134 186854
rect 473514 151174 474134 186618
rect 473514 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 474134 151174
rect 473514 150854 474134 150938
rect 473514 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 474134 150854
rect 473514 115174 474134 150618
rect 473514 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 474134 115174
rect 473514 114854 474134 114938
rect 473514 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 474134 114854
rect 473514 79174 474134 114618
rect 473514 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 474134 79174
rect 473514 78854 474134 78938
rect 473514 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 474134 78854
rect 473514 43174 474134 78618
rect 473514 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 474134 43174
rect 473514 42854 474134 42938
rect 473514 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 474134 42854
rect 473514 7174 474134 42618
rect 473514 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 474134 7174
rect 473514 6854 474134 6938
rect 473514 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 474134 6854
rect 473514 -2266 474134 6618
rect 473514 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 474134 -2266
rect 473514 -2586 474134 -2502
rect 473514 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 474134 -2586
rect 473514 -3814 474134 -2822
rect 477234 694894 477854 708122
rect 477234 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 477854 694894
rect 477234 694574 477854 694658
rect 477234 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 477854 694574
rect 477234 658894 477854 694338
rect 477234 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 477854 658894
rect 477234 658574 477854 658658
rect 477234 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 477854 658574
rect 477234 622894 477854 658338
rect 477234 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 477854 622894
rect 477234 622574 477854 622658
rect 477234 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 477854 622574
rect 477234 586894 477854 622338
rect 477234 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 477854 586894
rect 477234 586574 477854 586658
rect 477234 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 477854 586574
rect 477234 550894 477854 586338
rect 477234 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 477854 550894
rect 477234 550574 477854 550658
rect 477234 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 477854 550574
rect 477234 514894 477854 550338
rect 477234 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 477854 514894
rect 477234 514574 477854 514658
rect 477234 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 477854 514574
rect 477234 478894 477854 514338
rect 477234 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 477854 478894
rect 477234 478574 477854 478658
rect 477234 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 477854 478574
rect 477234 442894 477854 478338
rect 477234 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 477854 442894
rect 477234 442574 477854 442658
rect 477234 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 477854 442574
rect 477234 406894 477854 442338
rect 477234 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 477854 406894
rect 477234 406574 477854 406658
rect 477234 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 477854 406574
rect 477234 370894 477854 406338
rect 477234 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 477854 370894
rect 477234 370574 477854 370658
rect 477234 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 477854 370574
rect 477234 334894 477854 370338
rect 477234 334658 477266 334894
rect 477502 334658 477586 334894
rect 477822 334658 477854 334894
rect 477234 334574 477854 334658
rect 477234 334338 477266 334574
rect 477502 334338 477586 334574
rect 477822 334338 477854 334574
rect 477234 298894 477854 334338
rect 477234 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 477854 298894
rect 477234 298574 477854 298658
rect 477234 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 477854 298574
rect 477234 262894 477854 298338
rect 477234 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 477854 262894
rect 477234 262574 477854 262658
rect 477234 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 477854 262574
rect 477234 226894 477854 262338
rect 477234 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 477854 226894
rect 477234 226574 477854 226658
rect 477234 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 477854 226574
rect 477234 190894 477854 226338
rect 477234 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 477854 190894
rect 477234 190574 477854 190658
rect 477234 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 477854 190574
rect 477234 154894 477854 190338
rect 477234 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 477854 154894
rect 477234 154574 477854 154658
rect 477234 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 477854 154574
rect 477234 118894 477854 154338
rect 477234 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 477854 118894
rect 477234 118574 477854 118658
rect 477234 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 477854 118574
rect 477234 82894 477854 118338
rect 477234 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 477854 82894
rect 477234 82574 477854 82658
rect 477234 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 477854 82574
rect 477234 46894 477854 82338
rect 477234 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 477854 46894
rect 477234 46574 477854 46658
rect 477234 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 477854 46574
rect 477234 10894 477854 46338
rect 477234 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 477854 10894
rect 477234 10574 477854 10658
rect 477234 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 477854 10574
rect 477234 -4186 477854 10338
rect 477234 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 477854 -4186
rect 477234 -4506 477854 -4422
rect 477234 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 477854 -4506
rect 477234 -5734 477854 -4742
rect 480954 698614 481574 710042
rect 498954 711558 499574 711590
rect 498954 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 499574 711558
rect 498954 711238 499574 711322
rect 498954 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 499574 711238
rect 495234 709638 495854 709670
rect 495234 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 495854 709638
rect 495234 709318 495854 709402
rect 495234 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 495854 709318
rect 491514 707718 492134 707750
rect 491514 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 492134 707718
rect 491514 707398 492134 707482
rect 491514 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 492134 707398
rect 480954 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 481574 698614
rect 480954 698294 481574 698378
rect 480954 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 481574 698294
rect 480954 662614 481574 698058
rect 480954 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 481574 662614
rect 480954 662294 481574 662378
rect 480954 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 481574 662294
rect 480954 626614 481574 662058
rect 480954 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 481574 626614
rect 480954 626294 481574 626378
rect 480954 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 481574 626294
rect 480954 590614 481574 626058
rect 480954 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 481574 590614
rect 480954 590294 481574 590378
rect 480954 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 481574 590294
rect 480954 554614 481574 590058
rect 480954 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 481574 554614
rect 480954 554294 481574 554378
rect 480954 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 481574 554294
rect 480954 518614 481574 554058
rect 480954 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 481574 518614
rect 480954 518294 481574 518378
rect 480954 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 481574 518294
rect 480954 482614 481574 518058
rect 480954 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 481574 482614
rect 480954 482294 481574 482378
rect 480954 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 481574 482294
rect 480954 446614 481574 482058
rect 480954 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 481574 446614
rect 480954 446294 481574 446378
rect 480954 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 481574 446294
rect 480954 410614 481574 446058
rect 480954 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 481574 410614
rect 480954 410294 481574 410378
rect 480954 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 481574 410294
rect 480954 374614 481574 410058
rect 480954 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 481574 374614
rect 480954 374294 481574 374378
rect 480954 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 481574 374294
rect 480954 338614 481574 374058
rect 480954 338378 480986 338614
rect 481222 338378 481306 338614
rect 481542 338378 481574 338614
rect 480954 338294 481574 338378
rect 480954 338058 480986 338294
rect 481222 338058 481306 338294
rect 481542 338058 481574 338294
rect 480954 302614 481574 338058
rect 480954 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 481574 302614
rect 480954 302294 481574 302378
rect 480954 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 481574 302294
rect 480954 266614 481574 302058
rect 480954 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 481574 266614
rect 480954 266294 481574 266378
rect 480954 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 481574 266294
rect 480954 230614 481574 266058
rect 480954 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 481574 230614
rect 480954 230294 481574 230378
rect 480954 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 481574 230294
rect 480954 194614 481574 230058
rect 480954 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 481574 194614
rect 480954 194294 481574 194378
rect 480954 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 481574 194294
rect 480954 158614 481574 194058
rect 480954 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 481574 158614
rect 480954 158294 481574 158378
rect 480954 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 481574 158294
rect 480954 122614 481574 158058
rect 480954 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 481574 122614
rect 480954 122294 481574 122378
rect 480954 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 481574 122294
rect 480954 86614 481574 122058
rect 480954 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 481574 86614
rect 480954 86294 481574 86378
rect 480954 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 481574 86294
rect 480954 50614 481574 86058
rect 480954 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 481574 50614
rect 480954 50294 481574 50378
rect 480954 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 481574 50294
rect 480954 14614 481574 50058
rect 480954 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 481574 14614
rect 480954 14294 481574 14378
rect 480954 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 481574 14294
rect 462954 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 463574 -7066
rect 462954 -7386 463574 -7302
rect 462954 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 463574 -7386
rect 462954 -7654 463574 -7622
rect 480954 -6106 481574 14058
rect 487794 705798 488414 705830
rect 487794 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 488414 705798
rect 487794 705478 488414 705562
rect 487794 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 488414 705478
rect 487794 669454 488414 705242
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 633454 488414 668898
rect 487794 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 488414 633454
rect 487794 633134 488414 633218
rect 487794 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 488414 633134
rect 487794 597454 488414 632898
rect 487794 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 488414 597454
rect 487794 597134 488414 597218
rect 487794 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 488414 597134
rect 487794 561454 488414 596898
rect 487794 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 488414 561454
rect 487794 561134 488414 561218
rect 487794 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 488414 561134
rect 487794 525454 488414 560898
rect 487794 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 488414 525454
rect 487794 525134 488414 525218
rect 487794 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 488414 525134
rect 487794 489454 488414 524898
rect 487794 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 488414 489454
rect 487794 489134 488414 489218
rect 487794 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 488414 489134
rect 487794 453454 488414 488898
rect 487794 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 488414 453454
rect 487794 453134 488414 453218
rect 487794 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 488414 453134
rect 487794 417454 488414 452898
rect 487794 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 488414 417454
rect 487794 417134 488414 417218
rect 487794 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 488414 417134
rect 487794 381454 488414 416898
rect 487794 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 488414 381454
rect 487794 381134 488414 381218
rect 487794 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 488414 381134
rect 487794 345454 488414 380898
rect 487794 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 488414 345454
rect 487794 345134 488414 345218
rect 487794 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 488414 345134
rect 487794 309454 488414 344898
rect 487794 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 488414 309454
rect 487794 309134 488414 309218
rect 487794 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 488414 309134
rect 487794 273454 488414 308898
rect 487794 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 488414 273454
rect 487794 273134 488414 273218
rect 487794 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 488414 273134
rect 487794 237454 488414 272898
rect 487794 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 488414 237454
rect 487794 237134 488414 237218
rect 487794 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 488414 237134
rect 487794 201454 488414 236898
rect 487794 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 488414 201454
rect 487794 201134 488414 201218
rect 487794 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 488414 201134
rect 487794 165454 488414 200898
rect 487794 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 488414 165454
rect 487794 165134 488414 165218
rect 487794 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 488414 165134
rect 487794 129454 488414 164898
rect 487794 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 488414 129454
rect 487794 129134 488414 129218
rect 487794 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 488414 129134
rect 487794 93454 488414 128898
rect 487794 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 488414 93454
rect 487794 93134 488414 93218
rect 487794 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 488414 93134
rect 487794 57454 488414 92898
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -1306 488414 20898
rect 487794 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 488414 -1306
rect 487794 -1626 488414 -1542
rect 487794 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 488414 -1626
rect 487794 -1894 488414 -1862
rect 491514 673174 492134 707162
rect 491514 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 492134 673174
rect 491514 672854 492134 672938
rect 491514 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 492134 672854
rect 491514 637174 492134 672618
rect 491514 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 492134 637174
rect 491514 636854 492134 636938
rect 491514 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 492134 636854
rect 491514 601174 492134 636618
rect 491514 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 492134 601174
rect 491514 600854 492134 600938
rect 491514 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 492134 600854
rect 491514 565174 492134 600618
rect 491514 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 492134 565174
rect 491514 564854 492134 564938
rect 491514 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 492134 564854
rect 491514 529174 492134 564618
rect 491514 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 492134 529174
rect 491514 528854 492134 528938
rect 491514 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 492134 528854
rect 491514 493174 492134 528618
rect 491514 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 492134 493174
rect 491514 492854 492134 492938
rect 491514 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 492134 492854
rect 491514 457174 492134 492618
rect 491514 456938 491546 457174
rect 491782 456938 491866 457174
rect 492102 456938 492134 457174
rect 491514 456854 492134 456938
rect 491514 456618 491546 456854
rect 491782 456618 491866 456854
rect 492102 456618 492134 456854
rect 491514 421174 492134 456618
rect 491514 420938 491546 421174
rect 491782 420938 491866 421174
rect 492102 420938 492134 421174
rect 491514 420854 492134 420938
rect 491514 420618 491546 420854
rect 491782 420618 491866 420854
rect 492102 420618 492134 420854
rect 491514 385174 492134 420618
rect 491514 384938 491546 385174
rect 491782 384938 491866 385174
rect 492102 384938 492134 385174
rect 491514 384854 492134 384938
rect 491514 384618 491546 384854
rect 491782 384618 491866 384854
rect 492102 384618 492134 384854
rect 491514 349174 492134 384618
rect 491514 348938 491546 349174
rect 491782 348938 491866 349174
rect 492102 348938 492134 349174
rect 491514 348854 492134 348938
rect 491514 348618 491546 348854
rect 491782 348618 491866 348854
rect 492102 348618 492134 348854
rect 491514 313174 492134 348618
rect 491514 312938 491546 313174
rect 491782 312938 491866 313174
rect 492102 312938 492134 313174
rect 491514 312854 492134 312938
rect 491514 312618 491546 312854
rect 491782 312618 491866 312854
rect 492102 312618 492134 312854
rect 491514 277174 492134 312618
rect 491514 276938 491546 277174
rect 491782 276938 491866 277174
rect 492102 276938 492134 277174
rect 491514 276854 492134 276938
rect 491514 276618 491546 276854
rect 491782 276618 491866 276854
rect 492102 276618 492134 276854
rect 491514 241174 492134 276618
rect 491514 240938 491546 241174
rect 491782 240938 491866 241174
rect 492102 240938 492134 241174
rect 491514 240854 492134 240938
rect 491514 240618 491546 240854
rect 491782 240618 491866 240854
rect 492102 240618 492134 240854
rect 491514 205174 492134 240618
rect 491514 204938 491546 205174
rect 491782 204938 491866 205174
rect 492102 204938 492134 205174
rect 491514 204854 492134 204938
rect 491514 204618 491546 204854
rect 491782 204618 491866 204854
rect 492102 204618 492134 204854
rect 491514 169174 492134 204618
rect 491514 168938 491546 169174
rect 491782 168938 491866 169174
rect 492102 168938 492134 169174
rect 491514 168854 492134 168938
rect 491514 168618 491546 168854
rect 491782 168618 491866 168854
rect 492102 168618 492134 168854
rect 491514 133174 492134 168618
rect 491514 132938 491546 133174
rect 491782 132938 491866 133174
rect 492102 132938 492134 133174
rect 491514 132854 492134 132938
rect 491514 132618 491546 132854
rect 491782 132618 491866 132854
rect 492102 132618 492134 132854
rect 491514 97174 492134 132618
rect 491514 96938 491546 97174
rect 491782 96938 491866 97174
rect 492102 96938 492134 97174
rect 491514 96854 492134 96938
rect 491514 96618 491546 96854
rect 491782 96618 491866 96854
rect 492102 96618 492134 96854
rect 491514 61174 492134 96618
rect 491514 60938 491546 61174
rect 491782 60938 491866 61174
rect 492102 60938 492134 61174
rect 491514 60854 492134 60938
rect 491514 60618 491546 60854
rect 491782 60618 491866 60854
rect 492102 60618 492134 60854
rect 491514 25174 492134 60618
rect 491514 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 492134 25174
rect 491514 24854 492134 24938
rect 491514 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 492134 24854
rect 491514 -3226 492134 24618
rect 491514 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 492134 -3226
rect 491514 -3546 492134 -3462
rect 491514 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 492134 -3546
rect 491514 -3814 492134 -3782
rect 495234 676894 495854 709082
rect 495234 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 495854 676894
rect 495234 676574 495854 676658
rect 495234 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 495854 676574
rect 495234 640894 495854 676338
rect 495234 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 495854 640894
rect 495234 640574 495854 640658
rect 495234 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 495854 640574
rect 495234 604894 495854 640338
rect 495234 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 495854 604894
rect 495234 604574 495854 604658
rect 495234 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 495854 604574
rect 495234 568894 495854 604338
rect 495234 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 495854 568894
rect 495234 568574 495854 568658
rect 495234 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 495854 568574
rect 495234 532894 495854 568338
rect 495234 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 495854 532894
rect 495234 532574 495854 532658
rect 495234 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 495854 532574
rect 495234 496894 495854 532338
rect 495234 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 495854 496894
rect 495234 496574 495854 496658
rect 495234 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 495854 496574
rect 495234 460894 495854 496338
rect 495234 460658 495266 460894
rect 495502 460658 495586 460894
rect 495822 460658 495854 460894
rect 495234 460574 495854 460658
rect 495234 460338 495266 460574
rect 495502 460338 495586 460574
rect 495822 460338 495854 460574
rect 495234 424894 495854 460338
rect 495234 424658 495266 424894
rect 495502 424658 495586 424894
rect 495822 424658 495854 424894
rect 495234 424574 495854 424658
rect 495234 424338 495266 424574
rect 495502 424338 495586 424574
rect 495822 424338 495854 424574
rect 495234 388894 495854 424338
rect 495234 388658 495266 388894
rect 495502 388658 495586 388894
rect 495822 388658 495854 388894
rect 495234 388574 495854 388658
rect 495234 388338 495266 388574
rect 495502 388338 495586 388574
rect 495822 388338 495854 388574
rect 495234 352894 495854 388338
rect 495234 352658 495266 352894
rect 495502 352658 495586 352894
rect 495822 352658 495854 352894
rect 495234 352574 495854 352658
rect 495234 352338 495266 352574
rect 495502 352338 495586 352574
rect 495822 352338 495854 352574
rect 495234 316894 495854 352338
rect 495234 316658 495266 316894
rect 495502 316658 495586 316894
rect 495822 316658 495854 316894
rect 495234 316574 495854 316658
rect 495234 316338 495266 316574
rect 495502 316338 495586 316574
rect 495822 316338 495854 316574
rect 495234 280894 495854 316338
rect 495234 280658 495266 280894
rect 495502 280658 495586 280894
rect 495822 280658 495854 280894
rect 495234 280574 495854 280658
rect 495234 280338 495266 280574
rect 495502 280338 495586 280574
rect 495822 280338 495854 280574
rect 495234 244894 495854 280338
rect 495234 244658 495266 244894
rect 495502 244658 495586 244894
rect 495822 244658 495854 244894
rect 495234 244574 495854 244658
rect 495234 244338 495266 244574
rect 495502 244338 495586 244574
rect 495822 244338 495854 244574
rect 495234 208894 495854 244338
rect 495234 208658 495266 208894
rect 495502 208658 495586 208894
rect 495822 208658 495854 208894
rect 495234 208574 495854 208658
rect 495234 208338 495266 208574
rect 495502 208338 495586 208574
rect 495822 208338 495854 208574
rect 495234 172894 495854 208338
rect 495234 172658 495266 172894
rect 495502 172658 495586 172894
rect 495822 172658 495854 172894
rect 495234 172574 495854 172658
rect 495234 172338 495266 172574
rect 495502 172338 495586 172574
rect 495822 172338 495854 172574
rect 495234 136894 495854 172338
rect 495234 136658 495266 136894
rect 495502 136658 495586 136894
rect 495822 136658 495854 136894
rect 495234 136574 495854 136658
rect 495234 136338 495266 136574
rect 495502 136338 495586 136574
rect 495822 136338 495854 136574
rect 495234 100894 495854 136338
rect 495234 100658 495266 100894
rect 495502 100658 495586 100894
rect 495822 100658 495854 100894
rect 495234 100574 495854 100658
rect 495234 100338 495266 100574
rect 495502 100338 495586 100574
rect 495822 100338 495854 100574
rect 495234 64894 495854 100338
rect 495234 64658 495266 64894
rect 495502 64658 495586 64894
rect 495822 64658 495854 64894
rect 495234 64574 495854 64658
rect 495234 64338 495266 64574
rect 495502 64338 495586 64574
rect 495822 64338 495854 64574
rect 495234 28894 495854 64338
rect 495234 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 495854 28894
rect 495234 28574 495854 28658
rect 495234 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 495854 28574
rect 495234 -5146 495854 28338
rect 495234 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 495854 -5146
rect 495234 -5466 495854 -5382
rect 495234 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 495854 -5466
rect 495234 -5734 495854 -5702
rect 498954 680614 499574 711002
rect 516954 710598 517574 711590
rect 516954 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 517574 710598
rect 516954 710278 517574 710362
rect 516954 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 517574 710278
rect 513234 708678 513854 709670
rect 513234 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 513854 708678
rect 513234 708358 513854 708442
rect 513234 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 513854 708358
rect 509514 706758 510134 707750
rect 509514 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 510134 706758
rect 509514 706438 510134 706522
rect 509514 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 510134 706438
rect 498954 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 499574 680614
rect 498954 680294 499574 680378
rect 498954 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 499574 680294
rect 498954 644614 499574 680058
rect 498954 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 499574 644614
rect 498954 644294 499574 644378
rect 498954 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 499574 644294
rect 498954 608614 499574 644058
rect 498954 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 499574 608614
rect 498954 608294 499574 608378
rect 498954 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 499574 608294
rect 498954 572614 499574 608058
rect 498954 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 499574 572614
rect 498954 572294 499574 572378
rect 498954 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 499574 572294
rect 498954 536614 499574 572058
rect 498954 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 499574 536614
rect 498954 536294 499574 536378
rect 498954 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 499574 536294
rect 498954 500614 499574 536058
rect 498954 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 499574 500614
rect 498954 500294 499574 500378
rect 498954 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 499574 500294
rect 498954 464614 499574 500058
rect 498954 464378 498986 464614
rect 499222 464378 499306 464614
rect 499542 464378 499574 464614
rect 498954 464294 499574 464378
rect 498954 464058 498986 464294
rect 499222 464058 499306 464294
rect 499542 464058 499574 464294
rect 498954 428614 499574 464058
rect 498954 428378 498986 428614
rect 499222 428378 499306 428614
rect 499542 428378 499574 428614
rect 498954 428294 499574 428378
rect 498954 428058 498986 428294
rect 499222 428058 499306 428294
rect 499542 428058 499574 428294
rect 498954 392614 499574 428058
rect 498954 392378 498986 392614
rect 499222 392378 499306 392614
rect 499542 392378 499574 392614
rect 498954 392294 499574 392378
rect 498954 392058 498986 392294
rect 499222 392058 499306 392294
rect 499542 392058 499574 392294
rect 498954 356614 499574 392058
rect 498954 356378 498986 356614
rect 499222 356378 499306 356614
rect 499542 356378 499574 356614
rect 498954 356294 499574 356378
rect 498954 356058 498986 356294
rect 499222 356058 499306 356294
rect 499542 356058 499574 356294
rect 498954 320614 499574 356058
rect 498954 320378 498986 320614
rect 499222 320378 499306 320614
rect 499542 320378 499574 320614
rect 498954 320294 499574 320378
rect 498954 320058 498986 320294
rect 499222 320058 499306 320294
rect 499542 320058 499574 320294
rect 498954 284614 499574 320058
rect 498954 284378 498986 284614
rect 499222 284378 499306 284614
rect 499542 284378 499574 284614
rect 498954 284294 499574 284378
rect 498954 284058 498986 284294
rect 499222 284058 499306 284294
rect 499542 284058 499574 284294
rect 498954 248614 499574 284058
rect 498954 248378 498986 248614
rect 499222 248378 499306 248614
rect 499542 248378 499574 248614
rect 498954 248294 499574 248378
rect 498954 248058 498986 248294
rect 499222 248058 499306 248294
rect 499542 248058 499574 248294
rect 498954 212614 499574 248058
rect 498954 212378 498986 212614
rect 499222 212378 499306 212614
rect 499542 212378 499574 212614
rect 498954 212294 499574 212378
rect 498954 212058 498986 212294
rect 499222 212058 499306 212294
rect 499542 212058 499574 212294
rect 498954 176614 499574 212058
rect 498954 176378 498986 176614
rect 499222 176378 499306 176614
rect 499542 176378 499574 176614
rect 498954 176294 499574 176378
rect 498954 176058 498986 176294
rect 499222 176058 499306 176294
rect 499542 176058 499574 176294
rect 498954 140614 499574 176058
rect 498954 140378 498986 140614
rect 499222 140378 499306 140614
rect 499542 140378 499574 140614
rect 498954 140294 499574 140378
rect 498954 140058 498986 140294
rect 499222 140058 499306 140294
rect 499542 140058 499574 140294
rect 498954 104614 499574 140058
rect 498954 104378 498986 104614
rect 499222 104378 499306 104614
rect 499542 104378 499574 104614
rect 498954 104294 499574 104378
rect 498954 104058 498986 104294
rect 499222 104058 499306 104294
rect 499542 104058 499574 104294
rect 498954 68614 499574 104058
rect 498954 68378 498986 68614
rect 499222 68378 499306 68614
rect 499542 68378 499574 68614
rect 498954 68294 499574 68378
rect 498954 68058 498986 68294
rect 499222 68058 499306 68294
rect 499542 68058 499574 68294
rect 498954 32614 499574 68058
rect 498954 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 499574 32614
rect 498954 32294 499574 32378
rect 498954 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 499574 32294
rect 480954 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 481574 -6106
rect 480954 -6426 481574 -6342
rect 480954 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 481574 -6426
rect 480954 -7654 481574 -6662
rect 498954 -7066 499574 32058
rect 505794 704838 506414 705830
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 505794 579454 506414 614898
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 291454 506414 326898
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 255454 506414 290898
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 219454 506414 254898
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 111454 506414 146898
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -1894 506414 -902
rect 509514 691174 510134 706202
rect 509514 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 510134 691174
rect 509514 690854 510134 690938
rect 509514 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 510134 690854
rect 509514 655174 510134 690618
rect 509514 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 510134 655174
rect 509514 654854 510134 654938
rect 509514 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 510134 654854
rect 509514 619174 510134 654618
rect 509514 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 510134 619174
rect 509514 618854 510134 618938
rect 509514 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 510134 618854
rect 509514 583174 510134 618618
rect 509514 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 510134 583174
rect 509514 582854 510134 582938
rect 509514 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 510134 582854
rect 509514 547174 510134 582618
rect 509514 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 510134 547174
rect 509514 546854 510134 546938
rect 509514 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 510134 546854
rect 509514 511174 510134 546618
rect 509514 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 510134 511174
rect 509514 510854 510134 510938
rect 509514 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 510134 510854
rect 509514 475174 510134 510618
rect 509514 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 510134 475174
rect 509514 474854 510134 474938
rect 509514 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 510134 474854
rect 509514 439174 510134 474618
rect 509514 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 510134 439174
rect 509514 438854 510134 438938
rect 509514 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 510134 438854
rect 509514 403174 510134 438618
rect 509514 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 510134 403174
rect 509514 402854 510134 402938
rect 509514 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 510134 402854
rect 509514 367174 510134 402618
rect 509514 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 510134 367174
rect 509514 366854 510134 366938
rect 509514 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 510134 366854
rect 509514 331174 510134 366618
rect 509514 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 510134 331174
rect 509514 330854 510134 330938
rect 509514 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 510134 330854
rect 509514 295174 510134 330618
rect 509514 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 510134 295174
rect 509514 294854 510134 294938
rect 509514 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 510134 294854
rect 509514 259174 510134 294618
rect 509514 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 510134 259174
rect 509514 258854 510134 258938
rect 509514 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 510134 258854
rect 509514 223174 510134 258618
rect 509514 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 510134 223174
rect 509514 222854 510134 222938
rect 509514 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 510134 222854
rect 509514 187174 510134 222618
rect 509514 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 510134 187174
rect 509514 186854 510134 186938
rect 509514 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 510134 186854
rect 509514 151174 510134 186618
rect 509514 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 510134 151174
rect 509514 150854 510134 150938
rect 509514 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 510134 150854
rect 509514 115174 510134 150618
rect 509514 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 510134 115174
rect 509514 114854 510134 114938
rect 509514 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 510134 114854
rect 509514 79174 510134 114618
rect 509514 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 510134 79174
rect 509514 78854 510134 78938
rect 509514 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 510134 78854
rect 509514 43174 510134 78618
rect 509514 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 510134 43174
rect 509514 42854 510134 42938
rect 509514 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 510134 42854
rect 509514 7174 510134 42618
rect 509514 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 510134 7174
rect 509514 6854 510134 6938
rect 509514 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 510134 6854
rect 509514 -2266 510134 6618
rect 509514 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 510134 -2266
rect 509514 -2586 510134 -2502
rect 509514 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 510134 -2586
rect 509514 -3814 510134 -2822
rect 513234 694894 513854 708122
rect 513234 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 513854 694894
rect 513234 694574 513854 694658
rect 513234 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 513854 694574
rect 513234 658894 513854 694338
rect 513234 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 513854 658894
rect 513234 658574 513854 658658
rect 513234 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 513854 658574
rect 513234 622894 513854 658338
rect 513234 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 513854 622894
rect 513234 622574 513854 622658
rect 513234 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 513854 622574
rect 513234 586894 513854 622338
rect 513234 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 513854 586894
rect 513234 586574 513854 586658
rect 513234 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 513854 586574
rect 513234 550894 513854 586338
rect 513234 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 513854 550894
rect 513234 550574 513854 550658
rect 513234 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 513854 550574
rect 513234 514894 513854 550338
rect 513234 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 513854 514894
rect 513234 514574 513854 514658
rect 513234 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 513854 514574
rect 513234 478894 513854 514338
rect 513234 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 513854 478894
rect 513234 478574 513854 478658
rect 513234 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 513854 478574
rect 513234 442894 513854 478338
rect 513234 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 513854 442894
rect 513234 442574 513854 442658
rect 513234 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 513854 442574
rect 513234 406894 513854 442338
rect 513234 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 513854 406894
rect 513234 406574 513854 406658
rect 513234 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 513854 406574
rect 513234 370894 513854 406338
rect 513234 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 513854 370894
rect 513234 370574 513854 370658
rect 513234 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 513854 370574
rect 513234 334894 513854 370338
rect 513234 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 513854 334894
rect 513234 334574 513854 334658
rect 513234 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 513854 334574
rect 513234 298894 513854 334338
rect 513234 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 513854 298894
rect 513234 298574 513854 298658
rect 513234 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 513854 298574
rect 513234 262894 513854 298338
rect 513234 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 513854 262894
rect 513234 262574 513854 262658
rect 513234 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 513854 262574
rect 513234 226894 513854 262338
rect 513234 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 513854 226894
rect 513234 226574 513854 226658
rect 513234 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 513854 226574
rect 513234 190894 513854 226338
rect 513234 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 513854 190894
rect 513234 190574 513854 190658
rect 513234 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 513854 190574
rect 513234 154894 513854 190338
rect 513234 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 513854 154894
rect 513234 154574 513854 154658
rect 513234 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 513854 154574
rect 513234 118894 513854 154338
rect 513234 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 513854 118894
rect 513234 118574 513854 118658
rect 513234 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 513854 118574
rect 513234 82894 513854 118338
rect 513234 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 513854 82894
rect 513234 82574 513854 82658
rect 513234 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 513854 82574
rect 513234 46894 513854 82338
rect 513234 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 513854 46894
rect 513234 46574 513854 46658
rect 513234 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 513854 46574
rect 513234 10894 513854 46338
rect 513234 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 513854 10894
rect 513234 10574 513854 10658
rect 513234 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 513854 10574
rect 513234 -4186 513854 10338
rect 513234 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 513854 -4186
rect 513234 -4506 513854 -4422
rect 513234 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 513854 -4506
rect 513234 -5734 513854 -4742
rect 516954 698614 517574 710042
rect 534954 711558 535574 711590
rect 534954 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 535574 711558
rect 534954 711238 535574 711322
rect 534954 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 535574 711238
rect 531234 709638 531854 709670
rect 531234 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 531854 709638
rect 531234 709318 531854 709402
rect 531234 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 531854 709318
rect 527514 707718 528134 707750
rect 527514 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 528134 707718
rect 527514 707398 528134 707482
rect 527514 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 528134 707398
rect 516954 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 517574 698614
rect 516954 698294 517574 698378
rect 516954 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 517574 698294
rect 516954 662614 517574 698058
rect 516954 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 517574 662614
rect 516954 662294 517574 662378
rect 516954 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 517574 662294
rect 516954 626614 517574 662058
rect 516954 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 517574 626614
rect 516954 626294 517574 626378
rect 516954 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 517574 626294
rect 516954 590614 517574 626058
rect 516954 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 517574 590614
rect 516954 590294 517574 590378
rect 516954 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 517574 590294
rect 516954 554614 517574 590058
rect 516954 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 517574 554614
rect 516954 554294 517574 554378
rect 516954 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 517574 554294
rect 516954 518614 517574 554058
rect 516954 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 517574 518614
rect 516954 518294 517574 518378
rect 516954 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 517574 518294
rect 516954 482614 517574 518058
rect 516954 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 517574 482614
rect 516954 482294 517574 482378
rect 516954 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 517574 482294
rect 516954 446614 517574 482058
rect 516954 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 517574 446614
rect 516954 446294 517574 446378
rect 516954 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 517574 446294
rect 516954 410614 517574 446058
rect 516954 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 517574 410614
rect 516954 410294 517574 410378
rect 516954 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 517574 410294
rect 516954 374614 517574 410058
rect 516954 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 517574 374614
rect 516954 374294 517574 374378
rect 516954 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 517574 374294
rect 516954 338614 517574 374058
rect 516954 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 517574 338614
rect 516954 338294 517574 338378
rect 516954 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 517574 338294
rect 516954 302614 517574 338058
rect 516954 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 517574 302614
rect 516954 302294 517574 302378
rect 516954 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 517574 302294
rect 516954 266614 517574 302058
rect 516954 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 517574 266614
rect 516954 266294 517574 266378
rect 516954 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 517574 266294
rect 516954 230614 517574 266058
rect 516954 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 517574 230614
rect 516954 230294 517574 230378
rect 516954 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 517574 230294
rect 516954 194614 517574 230058
rect 516954 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 517574 194614
rect 516954 194294 517574 194378
rect 516954 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 517574 194294
rect 516954 158614 517574 194058
rect 516954 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 517574 158614
rect 516954 158294 517574 158378
rect 516954 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 517574 158294
rect 516954 122614 517574 158058
rect 516954 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 517574 122614
rect 516954 122294 517574 122378
rect 516954 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 517574 122294
rect 516954 86614 517574 122058
rect 516954 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 517574 86614
rect 516954 86294 517574 86378
rect 516954 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 517574 86294
rect 516954 50614 517574 86058
rect 516954 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 517574 50614
rect 516954 50294 517574 50378
rect 516954 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 517574 50294
rect 516954 14614 517574 50058
rect 516954 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 517574 14614
rect 516954 14294 517574 14378
rect 516954 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 517574 14294
rect 498954 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 499574 -7066
rect 498954 -7386 499574 -7302
rect 498954 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 499574 -7386
rect 498954 -7654 499574 -7622
rect 516954 -6106 517574 14058
rect 523794 705798 524414 705830
rect 523794 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 524414 705798
rect 523794 705478 524414 705562
rect 523794 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 524414 705478
rect 523794 669454 524414 705242
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 523794 309454 524414 344898
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 523794 273454 524414 308898
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -1306 524414 20898
rect 523794 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 524414 -1306
rect 523794 -1626 524414 -1542
rect 523794 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 524414 -1626
rect 523794 -1894 524414 -1862
rect 527514 673174 528134 707162
rect 527514 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 528134 673174
rect 527514 672854 528134 672938
rect 527514 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 528134 672854
rect 527514 637174 528134 672618
rect 527514 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 528134 637174
rect 527514 636854 528134 636938
rect 527514 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 528134 636854
rect 527514 601174 528134 636618
rect 527514 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 528134 601174
rect 527514 600854 528134 600938
rect 527514 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 528134 600854
rect 527514 565174 528134 600618
rect 527514 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 528134 565174
rect 527514 564854 528134 564938
rect 527514 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 528134 564854
rect 527514 529174 528134 564618
rect 527514 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 528134 529174
rect 527514 528854 528134 528938
rect 527514 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 528134 528854
rect 527514 493174 528134 528618
rect 527514 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 528134 493174
rect 527514 492854 528134 492938
rect 527514 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 528134 492854
rect 527514 457174 528134 492618
rect 527514 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 528134 457174
rect 527514 456854 528134 456938
rect 527514 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 528134 456854
rect 527514 421174 528134 456618
rect 527514 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 528134 421174
rect 527514 420854 528134 420938
rect 527514 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 528134 420854
rect 527514 385174 528134 420618
rect 527514 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 528134 385174
rect 527514 384854 528134 384938
rect 527514 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 528134 384854
rect 527514 349174 528134 384618
rect 527514 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 528134 349174
rect 527514 348854 528134 348938
rect 527514 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 528134 348854
rect 527514 313174 528134 348618
rect 527514 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 528134 313174
rect 527514 312854 528134 312938
rect 527514 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 528134 312854
rect 527514 277174 528134 312618
rect 527514 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 528134 277174
rect 527514 276854 528134 276938
rect 527514 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 528134 276854
rect 527514 241174 528134 276618
rect 527514 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 528134 241174
rect 527514 240854 528134 240938
rect 527514 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 528134 240854
rect 527514 205174 528134 240618
rect 527514 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 528134 205174
rect 527514 204854 528134 204938
rect 527514 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 528134 204854
rect 527514 169174 528134 204618
rect 527514 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 528134 169174
rect 527514 168854 528134 168938
rect 527514 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 528134 168854
rect 527514 133174 528134 168618
rect 527514 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 528134 133174
rect 527514 132854 528134 132938
rect 527514 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 528134 132854
rect 527514 97174 528134 132618
rect 527514 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 528134 97174
rect 527514 96854 528134 96938
rect 527514 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 528134 96854
rect 527514 61174 528134 96618
rect 527514 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 528134 61174
rect 527514 60854 528134 60938
rect 527514 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 528134 60854
rect 527514 25174 528134 60618
rect 527514 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 528134 25174
rect 527514 24854 528134 24938
rect 527514 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 528134 24854
rect 527514 -3226 528134 24618
rect 527514 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 528134 -3226
rect 527514 -3546 528134 -3462
rect 527514 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 528134 -3546
rect 527514 -3814 528134 -3782
rect 531234 676894 531854 709082
rect 531234 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 531854 676894
rect 531234 676574 531854 676658
rect 531234 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 531854 676574
rect 531234 640894 531854 676338
rect 531234 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 531854 640894
rect 531234 640574 531854 640658
rect 531234 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 531854 640574
rect 531234 604894 531854 640338
rect 531234 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 531854 604894
rect 531234 604574 531854 604658
rect 531234 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 531854 604574
rect 531234 568894 531854 604338
rect 531234 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 531854 568894
rect 531234 568574 531854 568658
rect 531234 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 531854 568574
rect 531234 532894 531854 568338
rect 531234 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 531854 532894
rect 531234 532574 531854 532658
rect 531234 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 531854 532574
rect 531234 496894 531854 532338
rect 531234 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 531854 496894
rect 531234 496574 531854 496658
rect 531234 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 531854 496574
rect 531234 460894 531854 496338
rect 531234 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 531854 460894
rect 531234 460574 531854 460658
rect 531234 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 531854 460574
rect 531234 424894 531854 460338
rect 531234 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 531854 424894
rect 531234 424574 531854 424658
rect 531234 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 531854 424574
rect 531234 388894 531854 424338
rect 531234 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 531854 388894
rect 531234 388574 531854 388658
rect 531234 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 531854 388574
rect 531234 352894 531854 388338
rect 531234 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 531854 352894
rect 531234 352574 531854 352658
rect 531234 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 531854 352574
rect 531234 316894 531854 352338
rect 531234 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 531854 316894
rect 531234 316574 531854 316658
rect 531234 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 531854 316574
rect 531234 280894 531854 316338
rect 531234 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 531854 280894
rect 531234 280574 531854 280658
rect 531234 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 531854 280574
rect 531234 244894 531854 280338
rect 531234 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 531854 244894
rect 531234 244574 531854 244658
rect 531234 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 531854 244574
rect 531234 208894 531854 244338
rect 531234 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 531854 208894
rect 531234 208574 531854 208658
rect 531234 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 531854 208574
rect 531234 172894 531854 208338
rect 531234 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 531854 172894
rect 531234 172574 531854 172658
rect 531234 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 531854 172574
rect 531234 136894 531854 172338
rect 531234 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 531854 136894
rect 531234 136574 531854 136658
rect 531234 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 531854 136574
rect 531234 100894 531854 136338
rect 531234 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 531854 100894
rect 531234 100574 531854 100658
rect 531234 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 531854 100574
rect 531234 64894 531854 100338
rect 531234 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 531854 64894
rect 531234 64574 531854 64658
rect 531234 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 531854 64574
rect 531234 28894 531854 64338
rect 531234 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 531854 28894
rect 531234 28574 531854 28658
rect 531234 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 531854 28574
rect 531234 -5146 531854 28338
rect 531234 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 531854 -5146
rect 531234 -5466 531854 -5382
rect 531234 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 531854 -5466
rect 531234 -5734 531854 -5702
rect 534954 680614 535574 711002
rect 552954 710598 553574 711590
rect 552954 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 553574 710598
rect 552954 710278 553574 710362
rect 552954 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 553574 710278
rect 549234 708678 549854 709670
rect 549234 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 549854 708678
rect 549234 708358 549854 708442
rect 549234 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 549854 708358
rect 545514 706758 546134 707750
rect 545514 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 546134 706758
rect 545514 706438 546134 706522
rect 545514 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 546134 706438
rect 534954 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 535574 680614
rect 534954 680294 535574 680378
rect 534954 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 535574 680294
rect 534954 644614 535574 680058
rect 534954 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 535574 644614
rect 534954 644294 535574 644378
rect 534954 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 535574 644294
rect 534954 608614 535574 644058
rect 534954 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 535574 608614
rect 534954 608294 535574 608378
rect 534954 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 535574 608294
rect 534954 572614 535574 608058
rect 534954 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 535574 572614
rect 534954 572294 535574 572378
rect 534954 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 535574 572294
rect 534954 536614 535574 572058
rect 534954 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 535574 536614
rect 534954 536294 535574 536378
rect 534954 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 535574 536294
rect 534954 500614 535574 536058
rect 534954 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 535574 500614
rect 534954 500294 535574 500378
rect 534954 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 535574 500294
rect 534954 464614 535574 500058
rect 534954 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 535574 464614
rect 534954 464294 535574 464378
rect 534954 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 535574 464294
rect 534954 428614 535574 464058
rect 534954 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 535574 428614
rect 534954 428294 535574 428378
rect 534954 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 535574 428294
rect 534954 392614 535574 428058
rect 534954 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 535574 392614
rect 534954 392294 535574 392378
rect 534954 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 535574 392294
rect 534954 356614 535574 392058
rect 534954 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 535574 356614
rect 534954 356294 535574 356378
rect 534954 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 535574 356294
rect 534954 320614 535574 356058
rect 534954 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 535574 320614
rect 534954 320294 535574 320378
rect 534954 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 535574 320294
rect 534954 284614 535574 320058
rect 534954 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 535574 284614
rect 534954 284294 535574 284378
rect 534954 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 535574 284294
rect 534954 248614 535574 284058
rect 534954 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 535574 248614
rect 534954 248294 535574 248378
rect 534954 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 535574 248294
rect 534954 212614 535574 248058
rect 534954 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 535574 212614
rect 534954 212294 535574 212378
rect 534954 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 535574 212294
rect 534954 176614 535574 212058
rect 534954 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 535574 176614
rect 534954 176294 535574 176378
rect 534954 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 535574 176294
rect 534954 140614 535574 176058
rect 534954 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 535574 140614
rect 534954 140294 535574 140378
rect 534954 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 535574 140294
rect 534954 104614 535574 140058
rect 534954 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 535574 104614
rect 534954 104294 535574 104378
rect 534954 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 535574 104294
rect 534954 68614 535574 104058
rect 534954 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 535574 68614
rect 534954 68294 535574 68378
rect 534954 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 535574 68294
rect 534954 32614 535574 68058
rect 534954 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 535574 32614
rect 534954 32294 535574 32378
rect 534954 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 535574 32294
rect 516954 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 517574 -6106
rect 516954 -6426 517574 -6342
rect 516954 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 517574 -6426
rect 516954 -7654 517574 -6662
rect 534954 -7066 535574 32058
rect 541794 704838 542414 705830
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -1894 542414 -902
rect 545514 691174 546134 706202
rect 545514 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 546134 691174
rect 545514 690854 546134 690938
rect 545514 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 546134 690854
rect 545514 655174 546134 690618
rect 545514 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 546134 655174
rect 545514 654854 546134 654938
rect 545514 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 546134 654854
rect 545514 619174 546134 654618
rect 545514 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 546134 619174
rect 545514 618854 546134 618938
rect 545514 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 546134 618854
rect 545514 583174 546134 618618
rect 545514 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 546134 583174
rect 545514 582854 546134 582938
rect 545514 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 546134 582854
rect 545514 547174 546134 582618
rect 545514 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 546134 547174
rect 545514 546854 546134 546938
rect 545514 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 546134 546854
rect 545514 511174 546134 546618
rect 545514 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 546134 511174
rect 545514 510854 546134 510938
rect 545514 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 546134 510854
rect 545514 475174 546134 510618
rect 545514 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 546134 475174
rect 545514 474854 546134 474938
rect 545514 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 546134 474854
rect 545514 439174 546134 474618
rect 545514 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 546134 439174
rect 545514 438854 546134 438938
rect 545514 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 546134 438854
rect 545514 403174 546134 438618
rect 545514 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 546134 403174
rect 545514 402854 546134 402938
rect 545514 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 546134 402854
rect 545514 367174 546134 402618
rect 545514 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 546134 367174
rect 545514 366854 546134 366938
rect 545514 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 546134 366854
rect 545514 331174 546134 366618
rect 545514 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 546134 331174
rect 545514 330854 546134 330938
rect 545514 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 546134 330854
rect 545514 295174 546134 330618
rect 545514 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 546134 295174
rect 545514 294854 546134 294938
rect 545514 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 546134 294854
rect 545514 259174 546134 294618
rect 545514 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 546134 259174
rect 545514 258854 546134 258938
rect 545514 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 546134 258854
rect 545514 223174 546134 258618
rect 545514 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 546134 223174
rect 545514 222854 546134 222938
rect 545514 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 546134 222854
rect 545514 187174 546134 222618
rect 545514 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 546134 187174
rect 545514 186854 546134 186938
rect 545514 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 546134 186854
rect 545514 151174 546134 186618
rect 545514 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 546134 151174
rect 545514 150854 546134 150938
rect 545514 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 546134 150854
rect 545514 115174 546134 150618
rect 545514 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 546134 115174
rect 545514 114854 546134 114938
rect 545514 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 546134 114854
rect 545514 79174 546134 114618
rect 545514 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 546134 79174
rect 545514 78854 546134 78938
rect 545514 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 546134 78854
rect 545514 43174 546134 78618
rect 545514 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 546134 43174
rect 545514 42854 546134 42938
rect 545514 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 546134 42854
rect 545514 7174 546134 42618
rect 545514 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 546134 7174
rect 545514 6854 546134 6938
rect 545514 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 546134 6854
rect 545514 -2266 546134 6618
rect 545514 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 546134 -2266
rect 545514 -2586 546134 -2502
rect 545514 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 546134 -2586
rect 545514 -3814 546134 -2822
rect 549234 694894 549854 708122
rect 549234 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 549854 694894
rect 549234 694574 549854 694658
rect 549234 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 549854 694574
rect 549234 658894 549854 694338
rect 549234 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 549854 658894
rect 549234 658574 549854 658658
rect 549234 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 549854 658574
rect 549234 622894 549854 658338
rect 549234 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 549854 622894
rect 549234 622574 549854 622658
rect 549234 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 549854 622574
rect 549234 586894 549854 622338
rect 549234 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 549854 586894
rect 549234 586574 549854 586658
rect 549234 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 549854 586574
rect 549234 550894 549854 586338
rect 549234 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 549854 550894
rect 549234 550574 549854 550658
rect 549234 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 549854 550574
rect 549234 514894 549854 550338
rect 549234 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 549854 514894
rect 549234 514574 549854 514658
rect 549234 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 549854 514574
rect 549234 478894 549854 514338
rect 549234 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 549854 478894
rect 549234 478574 549854 478658
rect 549234 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 549854 478574
rect 549234 442894 549854 478338
rect 549234 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 549854 442894
rect 549234 442574 549854 442658
rect 549234 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 549854 442574
rect 549234 406894 549854 442338
rect 549234 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 549854 406894
rect 549234 406574 549854 406658
rect 549234 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 549854 406574
rect 549234 370894 549854 406338
rect 549234 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 549854 370894
rect 549234 370574 549854 370658
rect 549234 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 549854 370574
rect 549234 334894 549854 370338
rect 549234 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 549854 334894
rect 549234 334574 549854 334658
rect 549234 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 549854 334574
rect 549234 298894 549854 334338
rect 549234 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 549854 298894
rect 549234 298574 549854 298658
rect 549234 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 549854 298574
rect 549234 262894 549854 298338
rect 549234 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 549854 262894
rect 549234 262574 549854 262658
rect 549234 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 549854 262574
rect 549234 226894 549854 262338
rect 549234 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 549854 226894
rect 549234 226574 549854 226658
rect 549234 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 549854 226574
rect 549234 190894 549854 226338
rect 549234 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 549854 190894
rect 549234 190574 549854 190658
rect 549234 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 549854 190574
rect 549234 154894 549854 190338
rect 549234 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 549854 154894
rect 549234 154574 549854 154658
rect 549234 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 549854 154574
rect 549234 118894 549854 154338
rect 549234 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 549854 118894
rect 549234 118574 549854 118658
rect 549234 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 549854 118574
rect 549234 82894 549854 118338
rect 549234 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 549854 82894
rect 549234 82574 549854 82658
rect 549234 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 549854 82574
rect 549234 46894 549854 82338
rect 549234 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 549854 46894
rect 549234 46574 549854 46658
rect 549234 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 549854 46574
rect 549234 10894 549854 46338
rect 549234 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 549854 10894
rect 549234 10574 549854 10658
rect 549234 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 549854 10574
rect 549234 -4186 549854 10338
rect 549234 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 549854 -4186
rect 549234 -4506 549854 -4422
rect 549234 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 549854 -4506
rect 549234 -5734 549854 -4742
rect 552954 698614 553574 710042
rect 570954 711558 571574 711590
rect 570954 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 571574 711558
rect 570954 711238 571574 711322
rect 570954 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 571574 711238
rect 567234 709638 567854 709670
rect 567234 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 567854 709638
rect 567234 709318 567854 709402
rect 567234 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 567854 709318
rect 563514 707718 564134 707750
rect 563514 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 564134 707718
rect 563514 707398 564134 707482
rect 563514 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 564134 707398
rect 552954 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 553574 698614
rect 552954 698294 553574 698378
rect 552954 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 553574 698294
rect 552954 662614 553574 698058
rect 552954 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 553574 662614
rect 552954 662294 553574 662378
rect 552954 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 553574 662294
rect 552954 626614 553574 662058
rect 552954 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 553574 626614
rect 552954 626294 553574 626378
rect 552954 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 553574 626294
rect 552954 590614 553574 626058
rect 552954 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 553574 590614
rect 552954 590294 553574 590378
rect 552954 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 553574 590294
rect 552954 554614 553574 590058
rect 552954 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 553574 554614
rect 552954 554294 553574 554378
rect 552954 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 553574 554294
rect 552954 518614 553574 554058
rect 552954 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 553574 518614
rect 552954 518294 553574 518378
rect 552954 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 553574 518294
rect 552954 482614 553574 518058
rect 552954 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 553574 482614
rect 552954 482294 553574 482378
rect 552954 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 553574 482294
rect 552954 446614 553574 482058
rect 552954 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 553574 446614
rect 552954 446294 553574 446378
rect 552954 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 553574 446294
rect 552954 410614 553574 446058
rect 552954 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 553574 410614
rect 552954 410294 553574 410378
rect 552954 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 553574 410294
rect 552954 374614 553574 410058
rect 552954 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 553574 374614
rect 552954 374294 553574 374378
rect 552954 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 553574 374294
rect 552954 338614 553574 374058
rect 552954 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 553574 338614
rect 552954 338294 553574 338378
rect 552954 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 553574 338294
rect 552954 302614 553574 338058
rect 552954 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 553574 302614
rect 552954 302294 553574 302378
rect 552954 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 553574 302294
rect 552954 266614 553574 302058
rect 552954 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 553574 266614
rect 552954 266294 553574 266378
rect 552954 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 553574 266294
rect 552954 230614 553574 266058
rect 552954 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 553574 230614
rect 552954 230294 553574 230378
rect 552954 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 553574 230294
rect 552954 194614 553574 230058
rect 552954 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 553574 194614
rect 552954 194294 553574 194378
rect 552954 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 553574 194294
rect 552954 158614 553574 194058
rect 552954 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 553574 158614
rect 552954 158294 553574 158378
rect 552954 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 553574 158294
rect 552954 122614 553574 158058
rect 552954 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 553574 122614
rect 552954 122294 553574 122378
rect 552954 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 553574 122294
rect 552954 86614 553574 122058
rect 552954 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 553574 86614
rect 552954 86294 553574 86378
rect 552954 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 553574 86294
rect 552954 50614 553574 86058
rect 552954 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 553574 50614
rect 552954 50294 553574 50378
rect 552954 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 553574 50294
rect 552954 14614 553574 50058
rect 552954 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 553574 14614
rect 552954 14294 553574 14378
rect 552954 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 553574 14294
rect 534954 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 535574 -7066
rect 534954 -7386 535574 -7302
rect 534954 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 535574 -7386
rect 534954 -7654 535574 -7622
rect 552954 -6106 553574 14058
rect 559794 705798 560414 705830
rect 559794 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 560414 705798
rect 559794 705478 560414 705562
rect 559794 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 560414 705478
rect 559794 669454 560414 705242
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -1306 560414 20898
rect 559794 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 560414 -1306
rect 559794 -1626 560414 -1542
rect 559794 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 560414 -1626
rect 559794 -1894 560414 -1862
rect 563514 673174 564134 707162
rect 563514 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 564134 673174
rect 563514 672854 564134 672938
rect 563514 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 564134 672854
rect 563514 637174 564134 672618
rect 563514 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 564134 637174
rect 563514 636854 564134 636938
rect 563514 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 564134 636854
rect 563514 601174 564134 636618
rect 563514 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 564134 601174
rect 563514 600854 564134 600938
rect 563514 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 564134 600854
rect 563514 565174 564134 600618
rect 563514 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 564134 565174
rect 563514 564854 564134 564938
rect 563514 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 564134 564854
rect 563514 529174 564134 564618
rect 563514 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 564134 529174
rect 563514 528854 564134 528938
rect 563514 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 564134 528854
rect 563514 493174 564134 528618
rect 563514 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 564134 493174
rect 563514 492854 564134 492938
rect 563514 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 564134 492854
rect 563514 457174 564134 492618
rect 563514 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 564134 457174
rect 563514 456854 564134 456938
rect 563514 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 564134 456854
rect 563514 421174 564134 456618
rect 563514 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 564134 421174
rect 563514 420854 564134 420938
rect 563514 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 564134 420854
rect 563514 385174 564134 420618
rect 563514 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 564134 385174
rect 563514 384854 564134 384938
rect 563514 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 564134 384854
rect 563514 349174 564134 384618
rect 563514 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 564134 349174
rect 563514 348854 564134 348938
rect 563514 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 564134 348854
rect 563514 313174 564134 348618
rect 563514 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 564134 313174
rect 563514 312854 564134 312938
rect 563514 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 564134 312854
rect 563514 277174 564134 312618
rect 563514 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 564134 277174
rect 563514 276854 564134 276938
rect 563514 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 564134 276854
rect 563514 241174 564134 276618
rect 563514 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 564134 241174
rect 563514 240854 564134 240938
rect 563514 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 564134 240854
rect 563514 205174 564134 240618
rect 563514 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 564134 205174
rect 563514 204854 564134 204938
rect 563514 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 564134 204854
rect 563514 169174 564134 204618
rect 563514 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 564134 169174
rect 563514 168854 564134 168938
rect 563514 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 564134 168854
rect 563514 133174 564134 168618
rect 563514 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 564134 133174
rect 563514 132854 564134 132938
rect 563514 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 564134 132854
rect 563514 97174 564134 132618
rect 563514 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 564134 97174
rect 563514 96854 564134 96938
rect 563514 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 564134 96854
rect 563514 61174 564134 96618
rect 563514 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 564134 61174
rect 563514 60854 564134 60938
rect 563514 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 564134 60854
rect 563514 25174 564134 60618
rect 563514 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 564134 25174
rect 563514 24854 564134 24938
rect 563514 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 564134 24854
rect 563514 -3226 564134 24618
rect 563514 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 564134 -3226
rect 563514 -3546 564134 -3462
rect 563514 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 564134 -3546
rect 563514 -3814 564134 -3782
rect 567234 676894 567854 709082
rect 567234 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 567854 676894
rect 567234 676574 567854 676658
rect 567234 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 567854 676574
rect 567234 640894 567854 676338
rect 567234 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 567854 640894
rect 567234 640574 567854 640658
rect 567234 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 567854 640574
rect 567234 604894 567854 640338
rect 567234 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 567854 604894
rect 567234 604574 567854 604658
rect 567234 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 567854 604574
rect 567234 568894 567854 604338
rect 567234 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 567854 568894
rect 567234 568574 567854 568658
rect 567234 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 567854 568574
rect 567234 532894 567854 568338
rect 567234 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 567854 532894
rect 567234 532574 567854 532658
rect 567234 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 567854 532574
rect 567234 496894 567854 532338
rect 567234 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 567854 496894
rect 567234 496574 567854 496658
rect 567234 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 567854 496574
rect 567234 460894 567854 496338
rect 567234 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 567854 460894
rect 567234 460574 567854 460658
rect 567234 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 567854 460574
rect 567234 424894 567854 460338
rect 567234 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 567854 424894
rect 567234 424574 567854 424658
rect 567234 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 567854 424574
rect 567234 388894 567854 424338
rect 567234 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 567854 388894
rect 567234 388574 567854 388658
rect 567234 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 567854 388574
rect 567234 352894 567854 388338
rect 567234 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 567854 352894
rect 567234 352574 567854 352658
rect 567234 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 567854 352574
rect 567234 316894 567854 352338
rect 567234 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 567854 316894
rect 567234 316574 567854 316658
rect 567234 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 567854 316574
rect 567234 280894 567854 316338
rect 567234 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 567854 280894
rect 567234 280574 567854 280658
rect 567234 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 567854 280574
rect 567234 244894 567854 280338
rect 567234 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 567854 244894
rect 567234 244574 567854 244658
rect 567234 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 567854 244574
rect 567234 208894 567854 244338
rect 567234 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 567854 208894
rect 567234 208574 567854 208658
rect 567234 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 567854 208574
rect 567234 172894 567854 208338
rect 567234 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 567854 172894
rect 567234 172574 567854 172658
rect 567234 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 567854 172574
rect 567234 136894 567854 172338
rect 567234 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 567854 136894
rect 567234 136574 567854 136658
rect 567234 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 567854 136574
rect 567234 100894 567854 136338
rect 567234 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 567854 100894
rect 567234 100574 567854 100658
rect 567234 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 567854 100574
rect 567234 64894 567854 100338
rect 567234 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 567854 64894
rect 567234 64574 567854 64658
rect 567234 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 567854 64574
rect 567234 28894 567854 64338
rect 567234 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 567854 28894
rect 567234 28574 567854 28658
rect 567234 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 567854 28574
rect 567234 -5146 567854 28338
rect 567234 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 567854 -5146
rect 567234 -5466 567854 -5382
rect 567234 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 567854 -5466
rect 567234 -5734 567854 -5702
rect 570954 680614 571574 711002
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 581514 706758 582134 707750
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 581514 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 582134 706758
rect 581514 706438 582134 706522
rect 581514 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 582134 706438
rect 570954 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 571574 680614
rect 570954 680294 571574 680378
rect 570954 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 571574 680294
rect 570954 644614 571574 680058
rect 570954 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 571574 644614
rect 570954 644294 571574 644378
rect 570954 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 571574 644294
rect 570954 608614 571574 644058
rect 570954 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 571574 608614
rect 570954 608294 571574 608378
rect 570954 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 571574 608294
rect 570954 572614 571574 608058
rect 570954 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 571574 572614
rect 570954 572294 571574 572378
rect 570954 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 571574 572294
rect 570954 536614 571574 572058
rect 570954 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 571574 536614
rect 570954 536294 571574 536378
rect 570954 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 571574 536294
rect 570954 500614 571574 536058
rect 570954 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 571574 500614
rect 570954 500294 571574 500378
rect 570954 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 571574 500294
rect 570954 464614 571574 500058
rect 570954 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 571574 464614
rect 570954 464294 571574 464378
rect 570954 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 571574 464294
rect 570954 428614 571574 464058
rect 570954 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 571574 428614
rect 570954 428294 571574 428378
rect 570954 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 571574 428294
rect 570954 392614 571574 428058
rect 570954 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 571574 392614
rect 570954 392294 571574 392378
rect 570954 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 571574 392294
rect 570954 356614 571574 392058
rect 570954 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 571574 356614
rect 570954 356294 571574 356378
rect 570954 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 571574 356294
rect 570954 320614 571574 356058
rect 570954 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 571574 320614
rect 570954 320294 571574 320378
rect 570954 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 571574 320294
rect 570954 284614 571574 320058
rect 570954 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 571574 284614
rect 570954 284294 571574 284378
rect 570954 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 571574 284294
rect 570954 248614 571574 284058
rect 570954 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 571574 248614
rect 570954 248294 571574 248378
rect 570954 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 571574 248294
rect 570954 212614 571574 248058
rect 570954 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 571574 212614
rect 570954 212294 571574 212378
rect 570954 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 571574 212294
rect 570954 176614 571574 212058
rect 570954 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 571574 176614
rect 570954 176294 571574 176378
rect 570954 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 571574 176294
rect 570954 140614 571574 176058
rect 570954 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 571574 140614
rect 570954 140294 571574 140378
rect 570954 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 571574 140294
rect 570954 104614 571574 140058
rect 570954 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 571574 104614
rect 570954 104294 571574 104378
rect 570954 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 571574 104294
rect 570954 68614 571574 104058
rect 570954 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 571574 68614
rect 570954 68294 571574 68378
rect 570954 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 571574 68294
rect 570954 32614 571574 68058
rect 570954 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 571574 32614
rect 570954 32294 571574 32378
rect 570954 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 571574 32294
rect 552954 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 553574 -6106
rect 552954 -6426 553574 -6342
rect 552954 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 553574 -6426
rect 552954 -7654 553574 -6662
rect 570954 -7066 571574 32058
rect 577794 704838 578414 705830
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -1894 578414 -902
rect 581514 691174 582134 706202
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581514 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 582134 691174
rect 581514 690854 582134 690938
rect 581514 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 582134 690854
rect 581514 655174 582134 690618
rect 581514 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 582134 655174
rect 581514 654854 582134 654938
rect 581514 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 582134 654854
rect 581514 619174 582134 654618
rect 581514 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 582134 619174
rect 581514 618854 582134 618938
rect 581514 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 582134 618854
rect 581514 583174 582134 618618
rect 581514 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 582134 583174
rect 581514 582854 582134 582938
rect 581514 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 582134 582854
rect 581514 547174 582134 582618
rect 581514 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 582134 547174
rect 581514 546854 582134 546938
rect 581514 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 582134 546854
rect 581514 511174 582134 546618
rect 581514 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 582134 511174
rect 581514 510854 582134 510938
rect 581514 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 582134 510854
rect 581514 475174 582134 510618
rect 581514 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 582134 475174
rect 581514 474854 582134 474938
rect 581514 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 582134 474854
rect 581514 439174 582134 474618
rect 581514 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 582134 439174
rect 581514 438854 582134 438938
rect 581514 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 582134 438854
rect 581514 403174 582134 438618
rect 581514 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 582134 403174
rect 581514 402854 582134 402938
rect 581514 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 582134 402854
rect 581514 367174 582134 402618
rect 581514 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 582134 367174
rect 581514 366854 582134 366938
rect 581514 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 582134 366854
rect 581514 331174 582134 366618
rect 581514 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 582134 331174
rect 581514 330854 582134 330938
rect 581514 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 582134 330854
rect 581514 295174 582134 330618
rect 581514 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 582134 295174
rect 581514 294854 582134 294938
rect 581514 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 582134 294854
rect 581514 259174 582134 294618
rect 581514 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 582134 259174
rect 581514 258854 582134 258938
rect 581514 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 582134 258854
rect 581514 223174 582134 258618
rect 581514 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 582134 223174
rect 581514 222854 582134 222938
rect 581514 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 582134 222854
rect 581514 187174 582134 222618
rect 581514 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 582134 187174
rect 581514 186854 582134 186938
rect 581514 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 582134 186854
rect 581514 151174 582134 186618
rect 581514 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 582134 151174
rect 581514 150854 582134 150938
rect 581514 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 582134 150854
rect 581514 115174 582134 150618
rect 581514 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 582134 115174
rect 581514 114854 582134 114938
rect 581514 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 582134 114854
rect 581514 79174 582134 114618
rect 581514 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 582134 79174
rect 581514 78854 582134 78938
rect 581514 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 582134 78854
rect 581514 43174 582134 78618
rect 581514 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 582134 43174
rect 581514 42854 582134 42938
rect 581514 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 582134 42854
rect 581514 7174 582134 42618
rect 581514 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 582134 7174
rect 581514 6854 582134 6938
rect 581514 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 582134 6854
rect 581514 -2266 582134 6618
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 669454 586890 705242
rect 586270 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect 586270 669134 586890 669218
rect 586270 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect 586270 633454 586890 668898
rect 586270 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect 586270 633134 586890 633218
rect 586270 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect 586270 597454 586890 632898
rect 586270 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect 586270 597134 586890 597218
rect 586270 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect 586270 561454 586890 596898
rect 586270 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect 586270 561134 586890 561218
rect 586270 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect 586270 525454 586890 560898
rect 586270 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect 586270 525134 586890 525218
rect 586270 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect 586270 489454 586890 524898
rect 586270 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect 586270 489134 586890 489218
rect 586270 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect 586270 453454 586890 488898
rect 586270 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect 586270 453134 586890 453218
rect 586270 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect 586270 417454 586890 452898
rect 586270 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect 586270 417134 586890 417218
rect 586270 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect 586270 381454 586890 416898
rect 586270 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect 586270 381134 586890 381218
rect 586270 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect 586270 345454 586890 380898
rect 586270 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect 586270 345134 586890 345218
rect 586270 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect 586270 309454 586890 344898
rect 586270 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect 586270 309134 586890 309218
rect 586270 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect 586270 273454 586890 308898
rect 586270 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect 586270 273134 586890 273218
rect 586270 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect 586270 237454 586890 272898
rect 586270 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect 586270 237134 586890 237218
rect 586270 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect 586270 201454 586890 236898
rect 586270 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect 586270 201134 586890 201218
rect 586270 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect 586270 165454 586890 200898
rect 586270 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect 586270 165134 586890 165218
rect 586270 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect 586270 129454 586890 164898
rect 586270 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect 586270 129134 586890 129218
rect 586270 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect 586270 93454 586890 128898
rect 586270 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect 586270 93134 586890 93218
rect 586270 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect 586270 57454 586890 92898
rect 586270 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect 586270 57134 586890 57218
rect 586270 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect 586270 21454 586890 56898
rect 586270 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect 586270 21134 586890 21218
rect 586270 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect 586270 -1306 586890 20898
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 691174 587850 706202
rect 587230 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 587850 691174
rect 587230 690854 587850 690938
rect 587230 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 587850 690854
rect 587230 655174 587850 690618
rect 587230 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 587850 655174
rect 587230 654854 587850 654938
rect 587230 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 587850 654854
rect 587230 619174 587850 654618
rect 587230 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 587850 619174
rect 587230 618854 587850 618938
rect 587230 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 587850 618854
rect 587230 583174 587850 618618
rect 587230 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 587850 583174
rect 587230 582854 587850 582938
rect 587230 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 587850 582854
rect 587230 547174 587850 582618
rect 587230 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 587850 547174
rect 587230 546854 587850 546938
rect 587230 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 587850 546854
rect 587230 511174 587850 546618
rect 587230 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 587850 511174
rect 587230 510854 587850 510938
rect 587230 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 587850 510854
rect 587230 475174 587850 510618
rect 587230 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 587850 475174
rect 587230 474854 587850 474938
rect 587230 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 587850 474854
rect 587230 439174 587850 474618
rect 587230 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 587850 439174
rect 587230 438854 587850 438938
rect 587230 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 587850 438854
rect 587230 403174 587850 438618
rect 587230 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 587850 403174
rect 587230 402854 587850 402938
rect 587230 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 587850 402854
rect 587230 367174 587850 402618
rect 587230 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 587850 367174
rect 587230 366854 587850 366938
rect 587230 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 587850 366854
rect 587230 331174 587850 366618
rect 587230 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 587850 331174
rect 587230 330854 587850 330938
rect 587230 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 587850 330854
rect 587230 295174 587850 330618
rect 587230 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 587850 295174
rect 587230 294854 587850 294938
rect 587230 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 587850 294854
rect 587230 259174 587850 294618
rect 587230 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 587850 259174
rect 587230 258854 587850 258938
rect 587230 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 587850 258854
rect 587230 223174 587850 258618
rect 587230 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 587850 223174
rect 587230 222854 587850 222938
rect 587230 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 587850 222854
rect 587230 187174 587850 222618
rect 587230 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 587850 187174
rect 587230 186854 587850 186938
rect 587230 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 587850 186854
rect 587230 151174 587850 186618
rect 587230 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 587850 151174
rect 587230 150854 587850 150938
rect 587230 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 587850 150854
rect 587230 115174 587850 150618
rect 587230 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 587850 115174
rect 587230 114854 587850 114938
rect 587230 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 587850 114854
rect 587230 79174 587850 114618
rect 587230 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 587850 79174
rect 587230 78854 587850 78938
rect 587230 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 587850 78854
rect 587230 43174 587850 78618
rect 587230 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 587850 43174
rect 587230 42854 587850 42938
rect 587230 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 587850 42854
rect 587230 7174 587850 42618
rect 587230 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 587850 7174
rect 587230 6854 587850 6938
rect 587230 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 587850 6854
rect 581514 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 582134 -2266
rect 581514 -2586 582134 -2502
rect 581514 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 582134 -2586
rect 581514 -3814 582134 -2822
rect 587230 -2266 587850 6618
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 673174 588810 707162
rect 588190 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect 588190 672854 588810 672938
rect 588190 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect 588190 637174 588810 672618
rect 588190 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect 588190 636854 588810 636938
rect 588190 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect 588190 601174 588810 636618
rect 588190 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect 588190 600854 588810 600938
rect 588190 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect 588190 565174 588810 600618
rect 588190 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect 588190 564854 588810 564938
rect 588190 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect 588190 529174 588810 564618
rect 588190 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect 588190 528854 588810 528938
rect 588190 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect 588190 493174 588810 528618
rect 588190 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect 588190 492854 588810 492938
rect 588190 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect 588190 457174 588810 492618
rect 588190 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect 588190 456854 588810 456938
rect 588190 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect 588190 421174 588810 456618
rect 588190 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect 588190 420854 588810 420938
rect 588190 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect 588190 385174 588810 420618
rect 588190 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect 588190 384854 588810 384938
rect 588190 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect 588190 349174 588810 384618
rect 588190 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect 588190 348854 588810 348938
rect 588190 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect 588190 313174 588810 348618
rect 588190 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect 588190 312854 588810 312938
rect 588190 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect 588190 277174 588810 312618
rect 588190 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect 588190 276854 588810 276938
rect 588190 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect 588190 241174 588810 276618
rect 588190 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect 588190 240854 588810 240938
rect 588190 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect 588190 205174 588810 240618
rect 588190 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect 588190 204854 588810 204938
rect 588190 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect 588190 169174 588810 204618
rect 588190 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect 588190 168854 588810 168938
rect 588190 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect 588190 133174 588810 168618
rect 588190 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect 588190 132854 588810 132938
rect 588190 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect 588190 97174 588810 132618
rect 588190 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect 588190 96854 588810 96938
rect 588190 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect 588190 61174 588810 96618
rect 588190 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect 588190 60854 588810 60938
rect 588190 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect 588190 25174 588810 60618
rect 588190 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect 588190 24854 588810 24938
rect 588190 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect 588190 -3226 588810 24618
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 694894 589770 708122
rect 589150 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 589770 694894
rect 589150 694574 589770 694658
rect 589150 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 589770 694574
rect 589150 658894 589770 694338
rect 589150 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 589770 658894
rect 589150 658574 589770 658658
rect 589150 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 589770 658574
rect 589150 622894 589770 658338
rect 589150 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 589770 622894
rect 589150 622574 589770 622658
rect 589150 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 589770 622574
rect 589150 586894 589770 622338
rect 589150 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 589770 586894
rect 589150 586574 589770 586658
rect 589150 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 589770 586574
rect 589150 550894 589770 586338
rect 589150 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 589770 550894
rect 589150 550574 589770 550658
rect 589150 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 589770 550574
rect 589150 514894 589770 550338
rect 589150 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 589770 514894
rect 589150 514574 589770 514658
rect 589150 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 589770 514574
rect 589150 478894 589770 514338
rect 589150 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 589770 478894
rect 589150 478574 589770 478658
rect 589150 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 589770 478574
rect 589150 442894 589770 478338
rect 589150 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 589770 442894
rect 589150 442574 589770 442658
rect 589150 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 589770 442574
rect 589150 406894 589770 442338
rect 589150 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 589770 406894
rect 589150 406574 589770 406658
rect 589150 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 589770 406574
rect 589150 370894 589770 406338
rect 589150 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 589770 370894
rect 589150 370574 589770 370658
rect 589150 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 589770 370574
rect 589150 334894 589770 370338
rect 589150 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 589770 334894
rect 589150 334574 589770 334658
rect 589150 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 589770 334574
rect 589150 298894 589770 334338
rect 589150 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 589770 298894
rect 589150 298574 589770 298658
rect 589150 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 589770 298574
rect 589150 262894 589770 298338
rect 589150 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 589770 262894
rect 589150 262574 589770 262658
rect 589150 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 589770 262574
rect 589150 226894 589770 262338
rect 589150 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 589770 226894
rect 589150 226574 589770 226658
rect 589150 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 589770 226574
rect 589150 190894 589770 226338
rect 589150 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 589770 190894
rect 589150 190574 589770 190658
rect 589150 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 589770 190574
rect 589150 154894 589770 190338
rect 589150 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 589770 154894
rect 589150 154574 589770 154658
rect 589150 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 589770 154574
rect 589150 118894 589770 154338
rect 589150 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 589770 118894
rect 589150 118574 589770 118658
rect 589150 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 589770 118574
rect 589150 82894 589770 118338
rect 589150 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 589770 82894
rect 589150 82574 589770 82658
rect 589150 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 589770 82574
rect 589150 46894 589770 82338
rect 589150 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 589770 46894
rect 589150 46574 589770 46658
rect 589150 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 589770 46574
rect 589150 10894 589770 46338
rect 589150 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 589770 10894
rect 589150 10574 589770 10658
rect 589150 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 589770 10574
rect 589150 -4186 589770 10338
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 676894 590730 709082
rect 590110 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect 590110 676574 590730 676658
rect 590110 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect 590110 640894 590730 676338
rect 590110 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect 590110 640574 590730 640658
rect 590110 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect 590110 604894 590730 640338
rect 590110 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect 590110 604574 590730 604658
rect 590110 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect 590110 568894 590730 604338
rect 590110 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect 590110 568574 590730 568658
rect 590110 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect 590110 532894 590730 568338
rect 590110 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect 590110 532574 590730 532658
rect 590110 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect 590110 496894 590730 532338
rect 590110 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect 590110 496574 590730 496658
rect 590110 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect 590110 460894 590730 496338
rect 590110 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect 590110 460574 590730 460658
rect 590110 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect 590110 424894 590730 460338
rect 590110 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect 590110 424574 590730 424658
rect 590110 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect 590110 388894 590730 424338
rect 590110 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect 590110 388574 590730 388658
rect 590110 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect 590110 352894 590730 388338
rect 590110 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect 590110 352574 590730 352658
rect 590110 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect 590110 316894 590730 352338
rect 590110 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect 590110 316574 590730 316658
rect 590110 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect 590110 280894 590730 316338
rect 590110 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect 590110 280574 590730 280658
rect 590110 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect 590110 244894 590730 280338
rect 590110 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect 590110 244574 590730 244658
rect 590110 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect 590110 208894 590730 244338
rect 590110 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect 590110 208574 590730 208658
rect 590110 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect 590110 172894 590730 208338
rect 590110 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect 590110 172574 590730 172658
rect 590110 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect 590110 136894 590730 172338
rect 590110 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect 590110 136574 590730 136658
rect 590110 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect 590110 100894 590730 136338
rect 590110 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect 590110 100574 590730 100658
rect 590110 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect 590110 64894 590730 100338
rect 590110 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect 590110 64574 590730 64658
rect 590110 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect 590110 28894 590730 64338
rect 590110 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect 590110 28574 590730 28658
rect 590110 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect 590110 -5146 590730 28338
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 698614 591690 710042
rect 591070 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 591690 698614
rect 591070 698294 591690 698378
rect 591070 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 591690 698294
rect 591070 662614 591690 698058
rect 591070 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 591690 662614
rect 591070 662294 591690 662378
rect 591070 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 591690 662294
rect 591070 626614 591690 662058
rect 591070 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 591690 626614
rect 591070 626294 591690 626378
rect 591070 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 591690 626294
rect 591070 590614 591690 626058
rect 591070 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 591690 590614
rect 591070 590294 591690 590378
rect 591070 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 591690 590294
rect 591070 554614 591690 590058
rect 591070 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 591690 554614
rect 591070 554294 591690 554378
rect 591070 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 591690 554294
rect 591070 518614 591690 554058
rect 591070 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 591690 518614
rect 591070 518294 591690 518378
rect 591070 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 591690 518294
rect 591070 482614 591690 518058
rect 591070 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 591690 482614
rect 591070 482294 591690 482378
rect 591070 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 591690 482294
rect 591070 446614 591690 482058
rect 591070 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 591690 446614
rect 591070 446294 591690 446378
rect 591070 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 591690 446294
rect 591070 410614 591690 446058
rect 591070 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 591690 410614
rect 591070 410294 591690 410378
rect 591070 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 591690 410294
rect 591070 374614 591690 410058
rect 591070 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 591690 374614
rect 591070 374294 591690 374378
rect 591070 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 591690 374294
rect 591070 338614 591690 374058
rect 591070 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 591690 338614
rect 591070 338294 591690 338378
rect 591070 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 591690 338294
rect 591070 302614 591690 338058
rect 591070 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 591690 302614
rect 591070 302294 591690 302378
rect 591070 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 591690 302294
rect 591070 266614 591690 302058
rect 591070 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 591690 266614
rect 591070 266294 591690 266378
rect 591070 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 591690 266294
rect 591070 230614 591690 266058
rect 591070 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 591690 230614
rect 591070 230294 591690 230378
rect 591070 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 591690 230294
rect 591070 194614 591690 230058
rect 591070 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 591690 194614
rect 591070 194294 591690 194378
rect 591070 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 591690 194294
rect 591070 158614 591690 194058
rect 591070 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 591690 158614
rect 591070 158294 591690 158378
rect 591070 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 591690 158294
rect 591070 122614 591690 158058
rect 591070 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 591690 122614
rect 591070 122294 591690 122378
rect 591070 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 591690 122294
rect 591070 86614 591690 122058
rect 591070 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 591690 86614
rect 591070 86294 591690 86378
rect 591070 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 591690 86294
rect 591070 50614 591690 86058
rect 591070 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 591690 50614
rect 591070 50294 591690 50378
rect 591070 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 591690 50294
rect 591070 14614 591690 50058
rect 591070 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 591690 14614
rect 591070 14294 591690 14378
rect 591070 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 591690 14294
rect 591070 -6106 591690 14058
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 680614 592650 711002
rect 592030 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect 592030 680294 592650 680378
rect 592030 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect 592030 644614 592650 680058
rect 592030 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect 592030 644294 592650 644378
rect 592030 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect 592030 608614 592650 644058
rect 592030 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect 592030 608294 592650 608378
rect 592030 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect 592030 572614 592650 608058
rect 592030 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect 592030 572294 592650 572378
rect 592030 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect 592030 536614 592650 572058
rect 592030 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect 592030 536294 592650 536378
rect 592030 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect 592030 500614 592650 536058
rect 592030 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect 592030 500294 592650 500378
rect 592030 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect 592030 464614 592650 500058
rect 592030 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect 592030 464294 592650 464378
rect 592030 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect 592030 428614 592650 464058
rect 592030 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect 592030 428294 592650 428378
rect 592030 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect 592030 392614 592650 428058
rect 592030 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect 592030 392294 592650 392378
rect 592030 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect 592030 356614 592650 392058
rect 592030 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect 592030 356294 592650 356378
rect 592030 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect 592030 320614 592650 356058
rect 592030 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect 592030 320294 592650 320378
rect 592030 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect 592030 284614 592650 320058
rect 592030 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect 592030 284294 592650 284378
rect 592030 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect 592030 248614 592650 284058
rect 592030 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect 592030 248294 592650 248378
rect 592030 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect 592030 212614 592650 248058
rect 592030 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect 592030 212294 592650 212378
rect 592030 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect 592030 176614 592650 212058
rect 592030 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect 592030 176294 592650 176378
rect 592030 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect 592030 140614 592650 176058
rect 592030 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect 592030 140294 592650 140378
rect 592030 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect 592030 104614 592650 140058
rect 592030 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect 592030 104294 592650 104378
rect 592030 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect 592030 68614 592650 104058
rect 592030 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect 592030 68294 592650 68378
rect 592030 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect 592030 32614 592650 68058
rect 592030 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect 592030 32294 592650 32378
rect 592030 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect 570954 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 571574 -7066
rect 570954 -7386 571574 -7302
rect 570954 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 571574 -7386
rect 570954 -7654 571574 -7622
rect 592030 -7066 592650 32058
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 680378 -8458 680614
rect -8374 680378 -8138 680614
rect -8694 680058 -8458 680294
rect -8374 680058 -8138 680294
rect -8694 644378 -8458 644614
rect -8374 644378 -8138 644614
rect -8694 644058 -8458 644294
rect -8374 644058 -8138 644294
rect -8694 608378 -8458 608614
rect -8374 608378 -8138 608614
rect -8694 608058 -8458 608294
rect -8374 608058 -8138 608294
rect -8694 572378 -8458 572614
rect -8374 572378 -8138 572614
rect -8694 572058 -8458 572294
rect -8374 572058 -8138 572294
rect -8694 536378 -8458 536614
rect -8374 536378 -8138 536614
rect -8694 536058 -8458 536294
rect -8374 536058 -8138 536294
rect -8694 500378 -8458 500614
rect -8374 500378 -8138 500614
rect -8694 500058 -8458 500294
rect -8374 500058 -8138 500294
rect -8694 464378 -8458 464614
rect -8374 464378 -8138 464614
rect -8694 464058 -8458 464294
rect -8374 464058 -8138 464294
rect -8694 428378 -8458 428614
rect -8374 428378 -8138 428614
rect -8694 428058 -8458 428294
rect -8374 428058 -8138 428294
rect -8694 392378 -8458 392614
rect -8374 392378 -8138 392614
rect -8694 392058 -8458 392294
rect -8374 392058 -8138 392294
rect -8694 356378 -8458 356614
rect -8374 356378 -8138 356614
rect -8694 356058 -8458 356294
rect -8374 356058 -8138 356294
rect -8694 320378 -8458 320614
rect -8374 320378 -8138 320614
rect -8694 320058 -8458 320294
rect -8374 320058 -8138 320294
rect -8694 284378 -8458 284614
rect -8374 284378 -8138 284614
rect -8694 284058 -8458 284294
rect -8374 284058 -8138 284294
rect -8694 248378 -8458 248614
rect -8374 248378 -8138 248614
rect -8694 248058 -8458 248294
rect -8374 248058 -8138 248294
rect -8694 212378 -8458 212614
rect -8374 212378 -8138 212614
rect -8694 212058 -8458 212294
rect -8374 212058 -8138 212294
rect -8694 176378 -8458 176614
rect -8374 176378 -8138 176614
rect -8694 176058 -8458 176294
rect -8374 176058 -8138 176294
rect -8694 140378 -8458 140614
rect -8374 140378 -8138 140614
rect -8694 140058 -8458 140294
rect -8374 140058 -8138 140294
rect -8694 104378 -8458 104614
rect -8374 104378 -8138 104614
rect -8694 104058 -8458 104294
rect -8374 104058 -8138 104294
rect -8694 68378 -8458 68614
rect -8374 68378 -8138 68614
rect -8694 68058 -8458 68294
rect -8374 68058 -8138 68294
rect -8694 32378 -8458 32614
rect -8374 32378 -8138 32614
rect -8694 32058 -8458 32294
rect -8374 32058 -8138 32294
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect 12986 710362 13222 710598
rect 13306 710362 13542 710598
rect 12986 710042 13222 710278
rect 13306 710042 13542 710278
rect -7734 698378 -7498 698614
rect -7414 698378 -7178 698614
rect -7734 698058 -7498 698294
rect -7414 698058 -7178 698294
rect -7734 662378 -7498 662614
rect -7414 662378 -7178 662614
rect -7734 662058 -7498 662294
rect -7414 662058 -7178 662294
rect -7734 626378 -7498 626614
rect -7414 626378 -7178 626614
rect -7734 626058 -7498 626294
rect -7414 626058 -7178 626294
rect -7734 590378 -7498 590614
rect -7414 590378 -7178 590614
rect -7734 590058 -7498 590294
rect -7414 590058 -7178 590294
rect -7734 554378 -7498 554614
rect -7414 554378 -7178 554614
rect -7734 554058 -7498 554294
rect -7414 554058 -7178 554294
rect -7734 518378 -7498 518614
rect -7414 518378 -7178 518614
rect -7734 518058 -7498 518294
rect -7414 518058 -7178 518294
rect -7734 482378 -7498 482614
rect -7414 482378 -7178 482614
rect -7734 482058 -7498 482294
rect -7414 482058 -7178 482294
rect -7734 446378 -7498 446614
rect -7414 446378 -7178 446614
rect -7734 446058 -7498 446294
rect -7414 446058 -7178 446294
rect -7734 410378 -7498 410614
rect -7414 410378 -7178 410614
rect -7734 410058 -7498 410294
rect -7414 410058 -7178 410294
rect -7734 374378 -7498 374614
rect -7414 374378 -7178 374614
rect -7734 374058 -7498 374294
rect -7414 374058 -7178 374294
rect -7734 338378 -7498 338614
rect -7414 338378 -7178 338614
rect -7734 338058 -7498 338294
rect -7414 338058 -7178 338294
rect -7734 302378 -7498 302614
rect -7414 302378 -7178 302614
rect -7734 302058 -7498 302294
rect -7414 302058 -7178 302294
rect -7734 266378 -7498 266614
rect -7414 266378 -7178 266614
rect -7734 266058 -7498 266294
rect -7414 266058 -7178 266294
rect -7734 230378 -7498 230614
rect -7414 230378 -7178 230614
rect -7734 230058 -7498 230294
rect -7414 230058 -7178 230294
rect -7734 194378 -7498 194614
rect -7414 194378 -7178 194614
rect -7734 194058 -7498 194294
rect -7414 194058 -7178 194294
rect -7734 158378 -7498 158614
rect -7414 158378 -7178 158614
rect -7734 158058 -7498 158294
rect -7414 158058 -7178 158294
rect -7734 122378 -7498 122614
rect -7414 122378 -7178 122614
rect -7734 122058 -7498 122294
rect -7414 122058 -7178 122294
rect -7734 86378 -7498 86614
rect -7414 86378 -7178 86614
rect -7734 86058 -7498 86294
rect -7414 86058 -7178 86294
rect -7734 50378 -7498 50614
rect -7414 50378 -7178 50614
rect -7734 50058 -7498 50294
rect -7414 50058 -7178 50294
rect -7734 14378 -7498 14614
rect -7414 14378 -7178 14614
rect -7734 14058 -7498 14294
rect -7414 14058 -7178 14294
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 676658 -6538 676894
rect -6454 676658 -6218 676894
rect -6774 676338 -6538 676574
rect -6454 676338 -6218 676574
rect -6774 640658 -6538 640894
rect -6454 640658 -6218 640894
rect -6774 640338 -6538 640574
rect -6454 640338 -6218 640574
rect -6774 604658 -6538 604894
rect -6454 604658 -6218 604894
rect -6774 604338 -6538 604574
rect -6454 604338 -6218 604574
rect -6774 568658 -6538 568894
rect -6454 568658 -6218 568894
rect -6774 568338 -6538 568574
rect -6454 568338 -6218 568574
rect -6774 532658 -6538 532894
rect -6454 532658 -6218 532894
rect -6774 532338 -6538 532574
rect -6454 532338 -6218 532574
rect -6774 496658 -6538 496894
rect -6454 496658 -6218 496894
rect -6774 496338 -6538 496574
rect -6454 496338 -6218 496574
rect -6774 460658 -6538 460894
rect -6454 460658 -6218 460894
rect -6774 460338 -6538 460574
rect -6454 460338 -6218 460574
rect -6774 424658 -6538 424894
rect -6454 424658 -6218 424894
rect -6774 424338 -6538 424574
rect -6454 424338 -6218 424574
rect -6774 388658 -6538 388894
rect -6454 388658 -6218 388894
rect -6774 388338 -6538 388574
rect -6454 388338 -6218 388574
rect -6774 352658 -6538 352894
rect -6454 352658 -6218 352894
rect -6774 352338 -6538 352574
rect -6454 352338 -6218 352574
rect -6774 316658 -6538 316894
rect -6454 316658 -6218 316894
rect -6774 316338 -6538 316574
rect -6454 316338 -6218 316574
rect -6774 280658 -6538 280894
rect -6454 280658 -6218 280894
rect -6774 280338 -6538 280574
rect -6454 280338 -6218 280574
rect -6774 244658 -6538 244894
rect -6454 244658 -6218 244894
rect -6774 244338 -6538 244574
rect -6454 244338 -6218 244574
rect -6774 208658 -6538 208894
rect -6454 208658 -6218 208894
rect -6774 208338 -6538 208574
rect -6454 208338 -6218 208574
rect -6774 172658 -6538 172894
rect -6454 172658 -6218 172894
rect -6774 172338 -6538 172574
rect -6454 172338 -6218 172574
rect -6774 136658 -6538 136894
rect -6454 136658 -6218 136894
rect -6774 136338 -6538 136574
rect -6454 136338 -6218 136574
rect -6774 100658 -6538 100894
rect -6454 100658 -6218 100894
rect -6774 100338 -6538 100574
rect -6454 100338 -6218 100574
rect -6774 64658 -6538 64894
rect -6454 64658 -6218 64894
rect -6774 64338 -6538 64574
rect -6454 64338 -6218 64574
rect -6774 28658 -6538 28894
rect -6454 28658 -6218 28894
rect -6774 28338 -6538 28574
rect -6454 28338 -6218 28574
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect 9266 708442 9502 708678
rect 9586 708442 9822 708678
rect 9266 708122 9502 708358
rect 9586 708122 9822 708358
rect -5814 694658 -5578 694894
rect -5494 694658 -5258 694894
rect -5814 694338 -5578 694574
rect -5494 694338 -5258 694574
rect -5814 658658 -5578 658894
rect -5494 658658 -5258 658894
rect -5814 658338 -5578 658574
rect -5494 658338 -5258 658574
rect -5814 622658 -5578 622894
rect -5494 622658 -5258 622894
rect -5814 622338 -5578 622574
rect -5494 622338 -5258 622574
rect -5814 586658 -5578 586894
rect -5494 586658 -5258 586894
rect -5814 586338 -5578 586574
rect -5494 586338 -5258 586574
rect -5814 550658 -5578 550894
rect -5494 550658 -5258 550894
rect -5814 550338 -5578 550574
rect -5494 550338 -5258 550574
rect -5814 514658 -5578 514894
rect -5494 514658 -5258 514894
rect -5814 514338 -5578 514574
rect -5494 514338 -5258 514574
rect -5814 478658 -5578 478894
rect -5494 478658 -5258 478894
rect -5814 478338 -5578 478574
rect -5494 478338 -5258 478574
rect -5814 442658 -5578 442894
rect -5494 442658 -5258 442894
rect -5814 442338 -5578 442574
rect -5494 442338 -5258 442574
rect -5814 406658 -5578 406894
rect -5494 406658 -5258 406894
rect -5814 406338 -5578 406574
rect -5494 406338 -5258 406574
rect -5814 370658 -5578 370894
rect -5494 370658 -5258 370894
rect -5814 370338 -5578 370574
rect -5494 370338 -5258 370574
rect -5814 334658 -5578 334894
rect -5494 334658 -5258 334894
rect -5814 334338 -5578 334574
rect -5494 334338 -5258 334574
rect -5814 298658 -5578 298894
rect -5494 298658 -5258 298894
rect -5814 298338 -5578 298574
rect -5494 298338 -5258 298574
rect -5814 262658 -5578 262894
rect -5494 262658 -5258 262894
rect -5814 262338 -5578 262574
rect -5494 262338 -5258 262574
rect -5814 226658 -5578 226894
rect -5494 226658 -5258 226894
rect -5814 226338 -5578 226574
rect -5494 226338 -5258 226574
rect -5814 190658 -5578 190894
rect -5494 190658 -5258 190894
rect -5814 190338 -5578 190574
rect -5494 190338 -5258 190574
rect -5814 154658 -5578 154894
rect -5494 154658 -5258 154894
rect -5814 154338 -5578 154574
rect -5494 154338 -5258 154574
rect -5814 118658 -5578 118894
rect -5494 118658 -5258 118894
rect -5814 118338 -5578 118574
rect -5494 118338 -5258 118574
rect -5814 82658 -5578 82894
rect -5494 82658 -5258 82894
rect -5814 82338 -5578 82574
rect -5494 82338 -5258 82574
rect -5814 46658 -5578 46894
rect -5494 46658 -5258 46894
rect -5814 46338 -5578 46574
rect -5494 46338 -5258 46574
rect -5814 10658 -5578 10894
rect -5494 10658 -5258 10894
rect -5814 10338 -5578 10574
rect -5494 10338 -5258 10574
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 672938 -4618 673174
rect -4534 672938 -4298 673174
rect -4854 672618 -4618 672854
rect -4534 672618 -4298 672854
rect -4854 636938 -4618 637174
rect -4534 636938 -4298 637174
rect -4854 636618 -4618 636854
rect -4534 636618 -4298 636854
rect -4854 600938 -4618 601174
rect -4534 600938 -4298 601174
rect -4854 600618 -4618 600854
rect -4534 600618 -4298 600854
rect -4854 564938 -4618 565174
rect -4534 564938 -4298 565174
rect -4854 564618 -4618 564854
rect -4534 564618 -4298 564854
rect -4854 528938 -4618 529174
rect -4534 528938 -4298 529174
rect -4854 528618 -4618 528854
rect -4534 528618 -4298 528854
rect -4854 492938 -4618 493174
rect -4534 492938 -4298 493174
rect -4854 492618 -4618 492854
rect -4534 492618 -4298 492854
rect -4854 456938 -4618 457174
rect -4534 456938 -4298 457174
rect -4854 456618 -4618 456854
rect -4534 456618 -4298 456854
rect -4854 420938 -4618 421174
rect -4534 420938 -4298 421174
rect -4854 420618 -4618 420854
rect -4534 420618 -4298 420854
rect -4854 384938 -4618 385174
rect -4534 384938 -4298 385174
rect -4854 384618 -4618 384854
rect -4534 384618 -4298 384854
rect -4854 348938 -4618 349174
rect -4534 348938 -4298 349174
rect -4854 348618 -4618 348854
rect -4534 348618 -4298 348854
rect -4854 312938 -4618 313174
rect -4534 312938 -4298 313174
rect -4854 312618 -4618 312854
rect -4534 312618 -4298 312854
rect -4854 276938 -4618 277174
rect -4534 276938 -4298 277174
rect -4854 276618 -4618 276854
rect -4534 276618 -4298 276854
rect -4854 240938 -4618 241174
rect -4534 240938 -4298 241174
rect -4854 240618 -4618 240854
rect -4534 240618 -4298 240854
rect -4854 204938 -4618 205174
rect -4534 204938 -4298 205174
rect -4854 204618 -4618 204854
rect -4534 204618 -4298 204854
rect -4854 168938 -4618 169174
rect -4534 168938 -4298 169174
rect -4854 168618 -4618 168854
rect -4534 168618 -4298 168854
rect -4854 132938 -4618 133174
rect -4534 132938 -4298 133174
rect -4854 132618 -4618 132854
rect -4534 132618 -4298 132854
rect -4854 96938 -4618 97174
rect -4534 96938 -4298 97174
rect -4854 96618 -4618 96854
rect -4534 96618 -4298 96854
rect -4854 60938 -4618 61174
rect -4534 60938 -4298 61174
rect -4854 60618 -4618 60854
rect -4534 60618 -4298 60854
rect -4854 24938 -4618 25174
rect -4534 24938 -4298 25174
rect -4854 24618 -4618 24854
rect -4534 24618 -4298 24854
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect 5546 706522 5782 706758
rect 5866 706522 6102 706758
rect 5546 706202 5782 706438
rect 5866 706202 6102 706438
rect -3894 690938 -3658 691174
rect -3574 690938 -3338 691174
rect -3894 690618 -3658 690854
rect -3574 690618 -3338 690854
rect -3894 654938 -3658 655174
rect -3574 654938 -3338 655174
rect -3894 654618 -3658 654854
rect -3574 654618 -3338 654854
rect -3894 618938 -3658 619174
rect -3574 618938 -3338 619174
rect -3894 618618 -3658 618854
rect -3574 618618 -3338 618854
rect -3894 582938 -3658 583174
rect -3574 582938 -3338 583174
rect -3894 582618 -3658 582854
rect -3574 582618 -3338 582854
rect -3894 546938 -3658 547174
rect -3574 546938 -3338 547174
rect -3894 546618 -3658 546854
rect -3574 546618 -3338 546854
rect -3894 510938 -3658 511174
rect -3574 510938 -3338 511174
rect -3894 510618 -3658 510854
rect -3574 510618 -3338 510854
rect -3894 474938 -3658 475174
rect -3574 474938 -3338 475174
rect -3894 474618 -3658 474854
rect -3574 474618 -3338 474854
rect -3894 438938 -3658 439174
rect -3574 438938 -3338 439174
rect -3894 438618 -3658 438854
rect -3574 438618 -3338 438854
rect -3894 402938 -3658 403174
rect -3574 402938 -3338 403174
rect -3894 402618 -3658 402854
rect -3574 402618 -3338 402854
rect -3894 366938 -3658 367174
rect -3574 366938 -3338 367174
rect -3894 366618 -3658 366854
rect -3574 366618 -3338 366854
rect -3894 330938 -3658 331174
rect -3574 330938 -3338 331174
rect -3894 330618 -3658 330854
rect -3574 330618 -3338 330854
rect -3894 294938 -3658 295174
rect -3574 294938 -3338 295174
rect -3894 294618 -3658 294854
rect -3574 294618 -3338 294854
rect -3894 258938 -3658 259174
rect -3574 258938 -3338 259174
rect -3894 258618 -3658 258854
rect -3574 258618 -3338 258854
rect -3894 222938 -3658 223174
rect -3574 222938 -3338 223174
rect -3894 222618 -3658 222854
rect -3574 222618 -3338 222854
rect -3894 186938 -3658 187174
rect -3574 186938 -3338 187174
rect -3894 186618 -3658 186854
rect -3574 186618 -3338 186854
rect -3894 150938 -3658 151174
rect -3574 150938 -3338 151174
rect -3894 150618 -3658 150854
rect -3574 150618 -3338 150854
rect -3894 114938 -3658 115174
rect -3574 114938 -3338 115174
rect -3894 114618 -3658 114854
rect -3574 114618 -3338 114854
rect -3894 78938 -3658 79174
rect -3574 78938 -3338 79174
rect -3894 78618 -3658 78854
rect -3574 78618 -3338 78854
rect -3894 42938 -3658 43174
rect -3574 42938 -3338 43174
rect -3894 42618 -3658 42854
rect -3574 42618 -3338 42854
rect -3894 6938 -3658 7174
rect -3574 6938 -3338 7174
rect -3894 6618 -3658 6854
rect -3574 6618 -3338 6854
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 669218 -2698 669454
rect -2614 669218 -2378 669454
rect -2934 668898 -2698 669134
rect -2614 668898 -2378 669134
rect -2934 633218 -2698 633454
rect -2614 633218 -2378 633454
rect -2934 632898 -2698 633134
rect -2614 632898 -2378 633134
rect -2934 597218 -2698 597454
rect -2614 597218 -2378 597454
rect -2934 596898 -2698 597134
rect -2614 596898 -2378 597134
rect -2934 561218 -2698 561454
rect -2614 561218 -2378 561454
rect -2934 560898 -2698 561134
rect -2614 560898 -2378 561134
rect -2934 525218 -2698 525454
rect -2614 525218 -2378 525454
rect -2934 524898 -2698 525134
rect -2614 524898 -2378 525134
rect -2934 489218 -2698 489454
rect -2614 489218 -2378 489454
rect -2934 488898 -2698 489134
rect -2614 488898 -2378 489134
rect -2934 453218 -2698 453454
rect -2614 453218 -2378 453454
rect -2934 452898 -2698 453134
rect -2614 452898 -2378 453134
rect -2934 417218 -2698 417454
rect -2614 417218 -2378 417454
rect -2934 416898 -2698 417134
rect -2614 416898 -2378 417134
rect -2934 381218 -2698 381454
rect -2614 381218 -2378 381454
rect -2934 380898 -2698 381134
rect -2614 380898 -2378 381134
rect -2934 345218 -2698 345454
rect -2614 345218 -2378 345454
rect -2934 344898 -2698 345134
rect -2614 344898 -2378 345134
rect -2934 309218 -2698 309454
rect -2614 309218 -2378 309454
rect -2934 308898 -2698 309134
rect -2614 308898 -2378 309134
rect -2934 273218 -2698 273454
rect -2614 273218 -2378 273454
rect -2934 272898 -2698 273134
rect -2614 272898 -2378 273134
rect -2934 237218 -2698 237454
rect -2614 237218 -2378 237454
rect -2934 236898 -2698 237134
rect -2614 236898 -2378 237134
rect -2934 201218 -2698 201454
rect -2614 201218 -2378 201454
rect -2934 200898 -2698 201134
rect -2614 200898 -2378 201134
rect -2934 165218 -2698 165454
rect -2614 165218 -2378 165454
rect -2934 164898 -2698 165134
rect -2614 164898 -2378 165134
rect -2934 129218 -2698 129454
rect -2614 129218 -2378 129454
rect -2934 128898 -2698 129134
rect -2614 128898 -2378 129134
rect -2934 93218 -2698 93454
rect -2614 93218 -2378 93454
rect -2934 92898 -2698 93134
rect -2614 92898 -2378 93134
rect -2934 57218 -2698 57454
rect -2614 57218 -2378 57454
rect -2934 56898 -2698 57134
rect -2614 56898 -2378 57134
rect -2934 21218 -2698 21454
rect -2614 21218 -2378 21454
rect -2934 20898 -2698 21134
rect -2614 20898 -2378 21134
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect 5546 690938 5782 691174
rect 5866 690938 6102 691174
rect 5546 690618 5782 690854
rect 5866 690618 6102 690854
rect 5546 654938 5782 655174
rect 5866 654938 6102 655174
rect 5546 654618 5782 654854
rect 5866 654618 6102 654854
rect 5546 618938 5782 619174
rect 5866 618938 6102 619174
rect 5546 618618 5782 618854
rect 5866 618618 6102 618854
rect 5546 582938 5782 583174
rect 5866 582938 6102 583174
rect 5546 582618 5782 582854
rect 5866 582618 6102 582854
rect 5546 546938 5782 547174
rect 5866 546938 6102 547174
rect 5546 546618 5782 546854
rect 5866 546618 6102 546854
rect 5546 510938 5782 511174
rect 5866 510938 6102 511174
rect 5546 510618 5782 510854
rect 5866 510618 6102 510854
rect 5546 474938 5782 475174
rect 5866 474938 6102 475174
rect 5546 474618 5782 474854
rect 5866 474618 6102 474854
rect 5546 438938 5782 439174
rect 5866 438938 6102 439174
rect 5546 438618 5782 438854
rect 5866 438618 6102 438854
rect 5546 402938 5782 403174
rect 5866 402938 6102 403174
rect 5546 402618 5782 402854
rect 5866 402618 6102 402854
rect 5546 366938 5782 367174
rect 5866 366938 6102 367174
rect 5546 366618 5782 366854
rect 5866 366618 6102 366854
rect 5546 330938 5782 331174
rect 5866 330938 6102 331174
rect 5546 330618 5782 330854
rect 5866 330618 6102 330854
rect 5546 294938 5782 295174
rect 5866 294938 6102 295174
rect 5546 294618 5782 294854
rect 5866 294618 6102 294854
rect 5546 258938 5782 259174
rect 5866 258938 6102 259174
rect 5546 258618 5782 258854
rect 5866 258618 6102 258854
rect 5546 222938 5782 223174
rect 5866 222938 6102 223174
rect 5546 222618 5782 222854
rect 5866 222618 6102 222854
rect 5546 186938 5782 187174
rect 5866 186938 6102 187174
rect 5546 186618 5782 186854
rect 5866 186618 6102 186854
rect 5546 150938 5782 151174
rect 5866 150938 6102 151174
rect 5546 150618 5782 150854
rect 5866 150618 6102 150854
rect 5546 114938 5782 115174
rect 5866 114938 6102 115174
rect 5546 114618 5782 114854
rect 5866 114618 6102 114854
rect 5546 78938 5782 79174
rect 5866 78938 6102 79174
rect 5546 78618 5782 78854
rect 5866 78618 6102 78854
rect 5546 42938 5782 43174
rect 5866 42938 6102 43174
rect 5546 42618 5782 42854
rect 5866 42618 6102 42854
rect 5546 6938 5782 7174
rect 5866 6938 6102 7174
rect 5546 6618 5782 6854
rect 5866 6618 6102 6854
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect 5546 -2502 5782 -2266
rect 5866 -2502 6102 -2266
rect 5546 -2822 5782 -2586
rect 5866 -2822 6102 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect 9266 694658 9502 694894
rect 9586 694658 9822 694894
rect 9266 694338 9502 694574
rect 9586 694338 9822 694574
rect 9266 658658 9502 658894
rect 9586 658658 9822 658894
rect 9266 658338 9502 658574
rect 9586 658338 9822 658574
rect 9266 622658 9502 622894
rect 9586 622658 9822 622894
rect 9266 622338 9502 622574
rect 9586 622338 9822 622574
rect 9266 586658 9502 586894
rect 9586 586658 9822 586894
rect 9266 586338 9502 586574
rect 9586 586338 9822 586574
rect 9266 550658 9502 550894
rect 9586 550658 9822 550894
rect 9266 550338 9502 550574
rect 9586 550338 9822 550574
rect 9266 514658 9502 514894
rect 9586 514658 9822 514894
rect 9266 514338 9502 514574
rect 9586 514338 9822 514574
rect 9266 478658 9502 478894
rect 9586 478658 9822 478894
rect 9266 478338 9502 478574
rect 9586 478338 9822 478574
rect 9266 442658 9502 442894
rect 9586 442658 9822 442894
rect 9266 442338 9502 442574
rect 9586 442338 9822 442574
rect 9266 406658 9502 406894
rect 9586 406658 9822 406894
rect 9266 406338 9502 406574
rect 9586 406338 9822 406574
rect 9266 370658 9502 370894
rect 9586 370658 9822 370894
rect 9266 370338 9502 370574
rect 9586 370338 9822 370574
rect 9266 334658 9502 334894
rect 9586 334658 9822 334894
rect 9266 334338 9502 334574
rect 9586 334338 9822 334574
rect 9266 298658 9502 298894
rect 9586 298658 9822 298894
rect 9266 298338 9502 298574
rect 9586 298338 9822 298574
rect 9266 262658 9502 262894
rect 9586 262658 9822 262894
rect 9266 262338 9502 262574
rect 9586 262338 9822 262574
rect 9266 226658 9502 226894
rect 9586 226658 9822 226894
rect 9266 226338 9502 226574
rect 9586 226338 9822 226574
rect 9266 190658 9502 190894
rect 9586 190658 9822 190894
rect 9266 190338 9502 190574
rect 9586 190338 9822 190574
rect 9266 154658 9502 154894
rect 9586 154658 9822 154894
rect 9266 154338 9502 154574
rect 9586 154338 9822 154574
rect 9266 118658 9502 118894
rect 9586 118658 9822 118894
rect 9266 118338 9502 118574
rect 9586 118338 9822 118574
rect 9266 82658 9502 82894
rect 9586 82658 9822 82894
rect 9266 82338 9502 82574
rect 9586 82338 9822 82574
rect 9266 46658 9502 46894
rect 9586 46658 9822 46894
rect 9266 46338 9502 46574
rect 9586 46338 9822 46574
rect 9266 10658 9502 10894
rect 9586 10658 9822 10894
rect 9266 10338 9502 10574
rect 9586 10338 9822 10574
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect 9266 -4422 9502 -4186
rect 9586 -4422 9822 -4186
rect 9266 -4742 9502 -4506
rect 9586 -4742 9822 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect 30986 711322 31222 711558
rect 31306 711322 31542 711558
rect 30986 711002 31222 711238
rect 31306 711002 31542 711238
rect 27266 709402 27502 709638
rect 27586 709402 27822 709638
rect 27266 709082 27502 709318
rect 27586 709082 27822 709318
rect 23546 707482 23782 707718
rect 23866 707482 24102 707718
rect 23546 707162 23782 707398
rect 23866 707162 24102 707398
rect 12986 698378 13222 698614
rect 13306 698378 13542 698614
rect 12986 698058 13222 698294
rect 13306 698058 13542 698294
rect 12986 662378 13222 662614
rect 13306 662378 13542 662614
rect 12986 662058 13222 662294
rect 13306 662058 13542 662294
rect 12986 626378 13222 626614
rect 13306 626378 13542 626614
rect 12986 626058 13222 626294
rect 13306 626058 13542 626294
rect 12986 590378 13222 590614
rect 13306 590378 13542 590614
rect 12986 590058 13222 590294
rect 13306 590058 13542 590294
rect 12986 554378 13222 554614
rect 13306 554378 13542 554614
rect 12986 554058 13222 554294
rect 13306 554058 13542 554294
rect 12986 518378 13222 518614
rect 13306 518378 13542 518614
rect 12986 518058 13222 518294
rect 13306 518058 13542 518294
rect 12986 482378 13222 482614
rect 13306 482378 13542 482614
rect 12986 482058 13222 482294
rect 13306 482058 13542 482294
rect 12986 446378 13222 446614
rect 13306 446378 13542 446614
rect 12986 446058 13222 446294
rect 13306 446058 13542 446294
rect 12986 410378 13222 410614
rect 13306 410378 13542 410614
rect 12986 410058 13222 410294
rect 13306 410058 13542 410294
rect 12986 374378 13222 374614
rect 13306 374378 13542 374614
rect 12986 374058 13222 374294
rect 13306 374058 13542 374294
rect 12986 338378 13222 338614
rect 13306 338378 13542 338614
rect 12986 338058 13222 338294
rect 13306 338058 13542 338294
rect 12986 302378 13222 302614
rect 13306 302378 13542 302614
rect 12986 302058 13222 302294
rect 13306 302058 13542 302294
rect 12986 266378 13222 266614
rect 13306 266378 13542 266614
rect 12986 266058 13222 266294
rect 13306 266058 13542 266294
rect 12986 230378 13222 230614
rect 13306 230378 13542 230614
rect 12986 230058 13222 230294
rect 13306 230058 13542 230294
rect 12986 194378 13222 194614
rect 13306 194378 13542 194614
rect 12986 194058 13222 194294
rect 13306 194058 13542 194294
rect 12986 158378 13222 158614
rect 13306 158378 13542 158614
rect 12986 158058 13222 158294
rect 13306 158058 13542 158294
rect 12986 122378 13222 122614
rect 13306 122378 13542 122614
rect 12986 122058 13222 122294
rect 13306 122058 13542 122294
rect 12986 86378 13222 86614
rect 13306 86378 13542 86614
rect 12986 86058 13222 86294
rect 13306 86058 13542 86294
rect 12986 50378 13222 50614
rect 13306 50378 13542 50614
rect 12986 50058 13222 50294
rect 13306 50058 13542 50294
rect 12986 14378 13222 14614
rect 13306 14378 13542 14614
rect 12986 14058 13222 14294
rect 13306 14058 13542 14294
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect 19826 705562 20062 705798
rect 20146 705562 20382 705798
rect 19826 705242 20062 705478
rect 20146 705242 20382 705478
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -1542 20062 -1306
rect 20146 -1542 20382 -1306
rect 19826 -1862 20062 -1626
rect 20146 -1862 20382 -1626
rect 23546 672938 23782 673174
rect 23866 672938 24102 673174
rect 23546 672618 23782 672854
rect 23866 672618 24102 672854
rect 23546 636938 23782 637174
rect 23866 636938 24102 637174
rect 23546 636618 23782 636854
rect 23866 636618 24102 636854
rect 23546 600938 23782 601174
rect 23866 600938 24102 601174
rect 23546 600618 23782 600854
rect 23866 600618 24102 600854
rect 23546 564938 23782 565174
rect 23866 564938 24102 565174
rect 23546 564618 23782 564854
rect 23866 564618 24102 564854
rect 23546 528938 23782 529174
rect 23866 528938 24102 529174
rect 23546 528618 23782 528854
rect 23866 528618 24102 528854
rect 23546 492938 23782 493174
rect 23866 492938 24102 493174
rect 23546 492618 23782 492854
rect 23866 492618 24102 492854
rect 23546 456938 23782 457174
rect 23866 456938 24102 457174
rect 23546 456618 23782 456854
rect 23866 456618 24102 456854
rect 23546 420938 23782 421174
rect 23866 420938 24102 421174
rect 23546 420618 23782 420854
rect 23866 420618 24102 420854
rect 23546 384938 23782 385174
rect 23866 384938 24102 385174
rect 23546 384618 23782 384854
rect 23866 384618 24102 384854
rect 23546 348938 23782 349174
rect 23866 348938 24102 349174
rect 23546 348618 23782 348854
rect 23866 348618 24102 348854
rect 23546 312938 23782 313174
rect 23866 312938 24102 313174
rect 23546 312618 23782 312854
rect 23866 312618 24102 312854
rect 23546 276938 23782 277174
rect 23866 276938 24102 277174
rect 23546 276618 23782 276854
rect 23866 276618 24102 276854
rect 23546 240938 23782 241174
rect 23866 240938 24102 241174
rect 23546 240618 23782 240854
rect 23866 240618 24102 240854
rect 23546 204938 23782 205174
rect 23866 204938 24102 205174
rect 23546 204618 23782 204854
rect 23866 204618 24102 204854
rect 23546 168938 23782 169174
rect 23866 168938 24102 169174
rect 23546 168618 23782 168854
rect 23866 168618 24102 168854
rect 23546 132938 23782 133174
rect 23866 132938 24102 133174
rect 23546 132618 23782 132854
rect 23866 132618 24102 132854
rect 23546 96938 23782 97174
rect 23866 96938 24102 97174
rect 23546 96618 23782 96854
rect 23866 96618 24102 96854
rect 23546 60938 23782 61174
rect 23866 60938 24102 61174
rect 23546 60618 23782 60854
rect 23866 60618 24102 60854
rect 23546 24938 23782 25174
rect 23866 24938 24102 25174
rect 23546 24618 23782 24854
rect 23866 24618 24102 24854
rect 23546 -3462 23782 -3226
rect 23866 -3462 24102 -3226
rect 23546 -3782 23782 -3546
rect 23866 -3782 24102 -3546
rect 27266 676658 27502 676894
rect 27586 676658 27822 676894
rect 27266 676338 27502 676574
rect 27586 676338 27822 676574
rect 27266 640658 27502 640894
rect 27586 640658 27822 640894
rect 27266 640338 27502 640574
rect 27586 640338 27822 640574
rect 27266 604658 27502 604894
rect 27586 604658 27822 604894
rect 27266 604338 27502 604574
rect 27586 604338 27822 604574
rect 27266 568658 27502 568894
rect 27586 568658 27822 568894
rect 27266 568338 27502 568574
rect 27586 568338 27822 568574
rect 27266 532658 27502 532894
rect 27586 532658 27822 532894
rect 27266 532338 27502 532574
rect 27586 532338 27822 532574
rect 27266 496658 27502 496894
rect 27586 496658 27822 496894
rect 27266 496338 27502 496574
rect 27586 496338 27822 496574
rect 27266 460658 27502 460894
rect 27586 460658 27822 460894
rect 27266 460338 27502 460574
rect 27586 460338 27822 460574
rect 27266 424658 27502 424894
rect 27586 424658 27822 424894
rect 27266 424338 27502 424574
rect 27586 424338 27822 424574
rect 27266 388658 27502 388894
rect 27586 388658 27822 388894
rect 27266 388338 27502 388574
rect 27586 388338 27822 388574
rect 27266 352658 27502 352894
rect 27586 352658 27822 352894
rect 27266 352338 27502 352574
rect 27586 352338 27822 352574
rect 27266 316658 27502 316894
rect 27586 316658 27822 316894
rect 27266 316338 27502 316574
rect 27586 316338 27822 316574
rect 27266 280658 27502 280894
rect 27586 280658 27822 280894
rect 27266 280338 27502 280574
rect 27586 280338 27822 280574
rect 27266 244658 27502 244894
rect 27586 244658 27822 244894
rect 27266 244338 27502 244574
rect 27586 244338 27822 244574
rect 27266 208658 27502 208894
rect 27586 208658 27822 208894
rect 27266 208338 27502 208574
rect 27586 208338 27822 208574
rect 27266 172658 27502 172894
rect 27586 172658 27822 172894
rect 27266 172338 27502 172574
rect 27586 172338 27822 172574
rect 27266 136658 27502 136894
rect 27586 136658 27822 136894
rect 27266 136338 27502 136574
rect 27586 136338 27822 136574
rect 27266 100658 27502 100894
rect 27586 100658 27822 100894
rect 27266 100338 27502 100574
rect 27586 100338 27822 100574
rect 27266 64658 27502 64894
rect 27586 64658 27822 64894
rect 27266 64338 27502 64574
rect 27586 64338 27822 64574
rect 27266 28658 27502 28894
rect 27586 28658 27822 28894
rect 27266 28338 27502 28574
rect 27586 28338 27822 28574
rect 27266 -5382 27502 -5146
rect 27586 -5382 27822 -5146
rect 27266 -5702 27502 -5466
rect 27586 -5702 27822 -5466
rect 48986 710362 49222 710598
rect 49306 710362 49542 710598
rect 48986 710042 49222 710278
rect 49306 710042 49542 710278
rect 45266 708442 45502 708678
rect 45586 708442 45822 708678
rect 45266 708122 45502 708358
rect 45586 708122 45822 708358
rect 41546 706522 41782 706758
rect 41866 706522 42102 706758
rect 41546 706202 41782 706438
rect 41866 706202 42102 706438
rect 30986 680378 31222 680614
rect 31306 680378 31542 680614
rect 30986 680058 31222 680294
rect 31306 680058 31542 680294
rect 30986 644378 31222 644614
rect 31306 644378 31542 644614
rect 30986 644058 31222 644294
rect 31306 644058 31542 644294
rect 30986 608378 31222 608614
rect 31306 608378 31542 608614
rect 30986 608058 31222 608294
rect 31306 608058 31542 608294
rect 30986 572378 31222 572614
rect 31306 572378 31542 572614
rect 30986 572058 31222 572294
rect 31306 572058 31542 572294
rect 30986 536378 31222 536614
rect 31306 536378 31542 536614
rect 30986 536058 31222 536294
rect 31306 536058 31542 536294
rect 30986 500378 31222 500614
rect 31306 500378 31542 500614
rect 30986 500058 31222 500294
rect 31306 500058 31542 500294
rect 30986 464378 31222 464614
rect 31306 464378 31542 464614
rect 30986 464058 31222 464294
rect 31306 464058 31542 464294
rect 30986 428378 31222 428614
rect 31306 428378 31542 428614
rect 30986 428058 31222 428294
rect 31306 428058 31542 428294
rect 30986 392378 31222 392614
rect 31306 392378 31542 392614
rect 30986 392058 31222 392294
rect 31306 392058 31542 392294
rect 30986 356378 31222 356614
rect 31306 356378 31542 356614
rect 30986 356058 31222 356294
rect 31306 356058 31542 356294
rect 30986 320378 31222 320614
rect 31306 320378 31542 320614
rect 30986 320058 31222 320294
rect 31306 320058 31542 320294
rect 30986 284378 31222 284614
rect 31306 284378 31542 284614
rect 30986 284058 31222 284294
rect 31306 284058 31542 284294
rect 30986 248378 31222 248614
rect 31306 248378 31542 248614
rect 30986 248058 31222 248294
rect 31306 248058 31542 248294
rect 30986 212378 31222 212614
rect 31306 212378 31542 212614
rect 30986 212058 31222 212294
rect 31306 212058 31542 212294
rect 30986 176378 31222 176614
rect 31306 176378 31542 176614
rect 30986 176058 31222 176294
rect 31306 176058 31542 176294
rect 30986 140378 31222 140614
rect 31306 140378 31542 140614
rect 30986 140058 31222 140294
rect 31306 140058 31542 140294
rect 30986 104378 31222 104614
rect 31306 104378 31542 104614
rect 30986 104058 31222 104294
rect 31306 104058 31542 104294
rect 30986 68378 31222 68614
rect 31306 68378 31542 68614
rect 30986 68058 31222 68294
rect 31306 68058 31542 68294
rect 30986 32378 31222 32614
rect 31306 32378 31542 32614
rect 30986 32058 31222 32294
rect 31306 32058 31542 32294
rect 12986 -6342 13222 -6106
rect 13306 -6342 13542 -6106
rect 12986 -6662 13222 -6426
rect 13306 -6662 13542 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 41546 690938 41782 691174
rect 41866 690938 42102 691174
rect 41546 690618 41782 690854
rect 41866 690618 42102 690854
rect 41546 654938 41782 655174
rect 41866 654938 42102 655174
rect 41546 654618 41782 654854
rect 41866 654618 42102 654854
rect 41546 618938 41782 619174
rect 41866 618938 42102 619174
rect 41546 618618 41782 618854
rect 41866 618618 42102 618854
rect 41546 582938 41782 583174
rect 41866 582938 42102 583174
rect 41546 582618 41782 582854
rect 41866 582618 42102 582854
rect 41546 546938 41782 547174
rect 41866 546938 42102 547174
rect 41546 546618 41782 546854
rect 41866 546618 42102 546854
rect 41546 510938 41782 511174
rect 41866 510938 42102 511174
rect 41546 510618 41782 510854
rect 41866 510618 42102 510854
rect 41546 474938 41782 475174
rect 41866 474938 42102 475174
rect 41546 474618 41782 474854
rect 41866 474618 42102 474854
rect 41546 438938 41782 439174
rect 41866 438938 42102 439174
rect 41546 438618 41782 438854
rect 41866 438618 42102 438854
rect 41546 402938 41782 403174
rect 41866 402938 42102 403174
rect 41546 402618 41782 402854
rect 41866 402618 42102 402854
rect 41546 366938 41782 367174
rect 41866 366938 42102 367174
rect 41546 366618 41782 366854
rect 41866 366618 42102 366854
rect 41546 330938 41782 331174
rect 41866 330938 42102 331174
rect 41546 330618 41782 330854
rect 41866 330618 42102 330854
rect 41546 294938 41782 295174
rect 41866 294938 42102 295174
rect 41546 294618 41782 294854
rect 41866 294618 42102 294854
rect 41546 258938 41782 259174
rect 41866 258938 42102 259174
rect 41546 258618 41782 258854
rect 41866 258618 42102 258854
rect 41546 222938 41782 223174
rect 41866 222938 42102 223174
rect 41546 222618 41782 222854
rect 41866 222618 42102 222854
rect 41546 186938 41782 187174
rect 41866 186938 42102 187174
rect 41546 186618 41782 186854
rect 41866 186618 42102 186854
rect 41546 150938 41782 151174
rect 41866 150938 42102 151174
rect 41546 150618 41782 150854
rect 41866 150618 42102 150854
rect 41546 114938 41782 115174
rect 41866 114938 42102 115174
rect 41546 114618 41782 114854
rect 41866 114618 42102 114854
rect 41546 78938 41782 79174
rect 41866 78938 42102 79174
rect 41546 78618 41782 78854
rect 41866 78618 42102 78854
rect 41546 42938 41782 43174
rect 41866 42938 42102 43174
rect 41546 42618 41782 42854
rect 41866 42618 42102 42854
rect 41546 6938 41782 7174
rect 41866 6938 42102 7174
rect 41546 6618 41782 6854
rect 41866 6618 42102 6854
rect 41546 -2502 41782 -2266
rect 41866 -2502 42102 -2266
rect 41546 -2822 41782 -2586
rect 41866 -2822 42102 -2586
rect 45266 694658 45502 694894
rect 45586 694658 45822 694894
rect 45266 694338 45502 694574
rect 45586 694338 45822 694574
rect 45266 658658 45502 658894
rect 45586 658658 45822 658894
rect 45266 658338 45502 658574
rect 45586 658338 45822 658574
rect 45266 622658 45502 622894
rect 45586 622658 45822 622894
rect 45266 622338 45502 622574
rect 45586 622338 45822 622574
rect 45266 586658 45502 586894
rect 45586 586658 45822 586894
rect 45266 586338 45502 586574
rect 45586 586338 45822 586574
rect 45266 550658 45502 550894
rect 45586 550658 45822 550894
rect 45266 550338 45502 550574
rect 45586 550338 45822 550574
rect 45266 514658 45502 514894
rect 45586 514658 45822 514894
rect 45266 514338 45502 514574
rect 45586 514338 45822 514574
rect 45266 478658 45502 478894
rect 45586 478658 45822 478894
rect 45266 478338 45502 478574
rect 45586 478338 45822 478574
rect 45266 442658 45502 442894
rect 45586 442658 45822 442894
rect 45266 442338 45502 442574
rect 45586 442338 45822 442574
rect 45266 406658 45502 406894
rect 45586 406658 45822 406894
rect 45266 406338 45502 406574
rect 45586 406338 45822 406574
rect 45266 370658 45502 370894
rect 45586 370658 45822 370894
rect 45266 370338 45502 370574
rect 45586 370338 45822 370574
rect 45266 334658 45502 334894
rect 45586 334658 45822 334894
rect 45266 334338 45502 334574
rect 45586 334338 45822 334574
rect 45266 298658 45502 298894
rect 45586 298658 45822 298894
rect 45266 298338 45502 298574
rect 45586 298338 45822 298574
rect 45266 262658 45502 262894
rect 45586 262658 45822 262894
rect 45266 262338 45502 262574
rect 45586 262338 45822 262574
rect 45266 226658 45502 226894
rect 45586 226658 45822 226894
rect 45266 226338 45502 226574
rect 45586 226338 45822 226574
rect 45266 190658 45502 190894
rect 45586 190658 45822 190894
rect 45266 190338 45502 190574
rect 45586 190338 45822 190574
rect 45266 154658 45502 154894
rect 45586 154658 45822 154894
rect 45266 154338 45502 154574
rect 45586 154338 45822 154574
rect 45266 118658 45502 118894
rect 45586 118658 45822 118894
rect 45266 118338 45502 118574
rect 45586 118338 45822 118574
rect 45266 82658 45502 82894
rect 45586 82658 45822 82894
rect 45266 82338 45502 82574
rect 45586 82338 45822 82574
rect 45266 46658 45502 46894
rect 45586 46658 45822 46894
rect 45266 46338 45502 46574
rect 45586 46338 45822 46574
rect 45266 10658 45502 10894
rect 45586 10658 45822 10894
rect 45266 10338 45502 10574
rect 45586 10338 45822 10574
rect 45266 -4422 45502 -4186
rect 45586 -4422 45822 -4186
rect 45266 -4742 45502 -4506
rect 45586 -4742 45822 -4506
rect 66986 711322 67222 711558
rect 67306 711322 67542 711558
rect 66986 711002 67222 711238
rect 67306 711002 67542 711238
rect 63266 709402 63502 709638
rect 63586 709402 63822 709638
rect 63266 709082 63502 709318
rect 63586 709082 63822 709318
rect 59546 707482 59782 707718
rect 59866 707482 60102 707718
rect 59546 707162 59782 707398
rect 59866 707162 60102 707398
rect 48986 698378 49222 698614
rect 49306 698378 49542 698614
rect 48986 698058 49222 698294
rect 49306 698058 49542 698294
rect 48986 662378 49222 662614
rect 49306 662378 49542 662614
rect 48986 662058 49222 662294
rect 49306 662058 49542 662294
rect 48986 626378 49222 626614
rect 49306 626378 49542 626614
rect 48986 626058 49222 626294
rect 49306 626058 49542 626294
rect 48986 590378 49222 590614
rect 49306 590378 49542 590614
rect 48986 590058 49222 590294
rect 49306 590058 49542 590294
rect 48986 554378 49222 554614
rect 49306 554378 49542 554614
rect 48986 554058 49222 554294
rect 49306 554058 49542 554294
rect 48986 518378 49222 518614
rect 49306 518378 49542 518614
rect 48986 518058 49222 518294
rect 49306 518058 49542 518294
rect 48986 482378 49222 482614
rect 49306 482378 49542 482614
rect 48986 482058 49222 482294
rect 49306 482058 49542 482294
rect 48986 446378 49222 446614
rect 49306 446378 49542 446614
rect 48986 446058 49222 446294
rect 49306 446058 49542 446294
rect 48986 410378 49222 410614
rect 49306 410378 49542 410614
rect 48986 410058 49222 410294
rect 49306 410058 49542 410294
rect 48986 374378 49222 374614
rect 49306 374378 49542 374614
rect 48986 374058 49222 374294
rect 49306 374058 49542 374294
rect 48986 338378 49222 338614
rect 49306 338378 49542 338614
rect 48986 338058 49222 338294
rect 49306 338058 49542 338294
rect 48986 302378 49222 302614
rect 49306 302378 49542 302614
rect 48986 302058 49222 302294
rect 49306 302058 49542 302294
rect 48986 266378 49222 266614
rect 49306 266378 49542 266614
rect 48986 266058 49222 266294
rect 49306 266058 49542 266294
rect 48986 230378 49222 230614
rect 49306 230378 49542 230614
rect 48986 230058 49222 230294
rect 49306 230058 49542 230294
rect 48986 194378 49222 194614
rect 49306 194378 49542 194614
rect 48986 194058 49222 194294
rect 49306 194058 49542 194294
rect 48986 158378 49222 158614
rect 49306 158378 49542 158614
rect 48986 158058 49222 158294
rect 49306 158058 49542 158294
rect 48986 122378 49222 122614
rect 49306 122378 49542 122614
rect 48986 122058 49222 122294
rect 49306 122058 49542 122294
rect 48986 86378 49222 86614
rect 49306 86378 49542 86614
rect 48986 86058 49222 86294
rect 49306 86058 49542 86294
rect 48986 50378 49222 50614
rect 49306 50378 49542 50614
rect 48986 50058 49222 50294
rect 49306 50058 49542 50294
rect 48986 14378 49222 14614
rect 49306 14378 49542 14614
rect 48986 14058 49222 14294
rect 49306 14058 49542 14294
rect 30986 -7302 31222 -7066
rect 31306 -7302 31542 -7066
rect 30986 -7622 31222 -7386
rect 31306 -7622 31542 -7386
rect 55826 705562 56062 705798
rect 56146 705562 56382 705798
rect 55826 705242 56062 705478
rect 56146 705242 56382 705478
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 55826 381218 56062 381454
rect 56146 381218 56382 381454
rect 55826 380898 56062 381134
rect 56146 380898 56382 381134
rect 55826 345218 56062 345454
rect 56146 345218 56382 345454
rect 55826 344898 56062 345134
rect 56146 344898 56382 345134
rect 55826 309218 56062 309454
rect 56146 309218 56382 309454
rect 55826 308898 56062 309134
rect 56146 308898 56382 309134
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 59546 672938 59782 673174
rect 59866 672938 60102 673174
rect 59546 672618 59782 672854
rect 59866 672618 60102 672854
rect 59546 636938 59782 637174
rect 59866 636938 60102 637174
rect 59546 636618 59782 636854
rect 59866 636618 60102 636854
rect 59546 600938 59782 601174
rect 59866 600938 60102 601174
rect 59546 600618 59782 600854
rect 59866 600618 60102 600854
rect 59546 564938 59782 565174
rect 59866 564938 60102 565174
rect 59546 564618 59782 564854
rect 59866 564618 60102 564854
rect 59546 528938 59782 529174
rect 59866 528938 60102 529174
rect 59546 528618 59782 528854
rect 59866 528618 60102 528854
rect 59546 492938 59782 493174
rect 59866 492938 60102 493174
rect 59546 492618 59782 492854
rect 59866 492618 60102 492854
rect 59546 456938 59782 457174
rect 59866 456938 60102 457174
rect 59546 456618 59782 456854
rect 59866 456618 60102 456854
rect 59546 420938 59782 421174
rect 59866 420938 60102 421174
rect 59546 420618 59782 420854
rect 59866 420618 60102 420854
rect 59546 384938 59782 385174
rect 59866 384938 60102 385174
rect 59546 384618 59782 384854
rect 59866 384618 60102 384854
rect 59546 348938 59782 349174
rect 59866 348938 60102 349174
rect 59546 348618 59782 348854
rect 59866 348618 60102 348854
rect 59546 312938 59782 313174
rect 59866 312938 60102 313174
rect 59546 312618 59782 312854
rect 59866 312618 60102 312854
rect 63266 676658 63502 676894
rect 63586 676658 63822 676894
rect 63266 676338 63502 676574
rect 63586 676338 63822 676574
rect 63266 640658 63502 640894
rect 63586 640658 63822 640894
rect 63266 640338 63502 640574
rect 63586 640338 63822 640574
rect 63266 604658 63502 604894
rect 63586 604658 63822 604894
rect 63266 604338 63502 604574
rect 63586 604338 63822 604574
rect 84986 710362 85222 710598
rect 85306 710362 85542 710598
rect 84986 710042 85222 710278
rect 85306 710042 85542 710278
rect 81266 708442 81502 708678
rect 81586 708442 81822 708678
rect 81266 708122 81502 708358
rect 81586 708122 81822 708358
rect 77546 706522 77782 706758
rect 77866 706522 78102 706758
rect 77546 706202 77782 706438
rect 77866 706202 78102 706438
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 66986 680378 67222 680614
rect 67306 680378 67542 680614
rect 66986 680058 67222 680294
rect 67306 680058 67542 680294
rect 66986 644378 67222 644614
rect 67306 644378 67542 644614
rect 66986 644058 67222 644294
rect 67306 644058 67542 644294
rect 66986 608378 67222 608614
rect 67306 608378 67542 608614
rect 66986 608058 67222 608294
rect 67306 608058 67542 608294
rect 63266 568658 63502 568894
rect 63586 568658 63822 568894
rect 63266 568338 63502 568574
rect 63586 568338 63822 568574
rect 63266 532658 63502 532894
rect 63586 532658 63822 532894
rect 63266 532338 63502 532574
rect 63586 532338 63822 532574
rect 63266 496658 63502 496894
rect 63586 496658 63822 496894
rect 63266 496338 63502 496574
rect 63586 496338 63822 496574
rect 63266 460658 63502 460894
rect 63586 460658 63822 460894
rect 63266 460338 63502 460574
rect 63586 460338 63822 460574
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 77546 690938 77782 691174
rect 77866 690938 78102 691174
rect 77546 690618 77782 690854
rect 77866 690618 78102 690854
rect 77546 654938 77782 655174
rect 77866 654938 78102 655174
rect 77546 654618 77782 654854
rect 77866 654618 78102 654854
rect 77546 618938 77782 619174
rect 77866 618938 78102 619174
rect 77546 618618 77782 618854
rect 77866 618618 78102 618854
rect 81266 694658 81502 694894
rect 81586 694658 81822 694894
rect 81266 694338 81502 694574
rect 81586 694338 81822 694574
rect 81266 658658 81502 658894
rect 81586 658658 81822 658894
rect 81266 658338 81502 658574
rect 81586 658338 81822 658574
rect 81266 622658 81502 622894
rect 81586 622658 81822 622894
rect 81266 622338 81502 622574
rect 81586 622338 81822 622574
rect 102986 711322 103222 711558
rect 103306 711322 103542 711558
rect 102986 711002 103222 711238
rect 103306 711002 103542 711238
rect 99266 709402 99502 709638
rect 99586 709402 99822 709638
rect 99266 709082 99502 709318
rect 99586 709082 99822 709318
rect 95546 707482 95782 707718
rect 95866 707482 96102 707718
rect 95546 707162 95782 707398
rect 95866 707162 96102 707398
rect 84986 698378 85222 698614
rect 85306 698378 85542 698614
rect 84986 698058 85222 698294
rect 85306 698058 85542 698294
rect 84986 662378 85222 662614
rect 85306 662378 85542 662614
rect 84986 662058 85222 662294
rect 85306 662058 85542 662294
rect 84986 626378 85222 626614
rect 85306 626378 85542 626614
rect 84986 626058 85222 626294
rect 85306 626058 85542 626294
rect 91826 705562 92062 705798
rect 92146 705562 92382 705798
rect 91826 705242 92062 705478
rect 92146 705242 92382 705478
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 91826 633218 92062 633454
rect 92146 633218 92382 633454
rect 91826 632898 92062 633134
rect 92146 632898 92382 633134
rect 91826 597218 92062 597454
rect 92146 597218 92382 597454
rect 91826 596898 92062 597134
rect 92146 596898 92382 597134
rect 72721 579218 72957 579454
rect 72721 578898 72957 579134
rect 78651 579218 78887 579454
rect 78651 578898 78887 579134
rect 84582 579218 84818 579454
rect 84582 578898 84818 579134
rect 75686 561218 75922 561454
rect 75686 560898 75922 561134
rect 81617 561218 81853 561454
rect 81617 560898 81853 561134
rect 72721 543218 72957 543454
rect 72721 542898 72957 543134
rect 78651 543218 78887 543454
rect 78651 542898 78887 543134
rect 84582 543218 84818 543454
rect 84582 542898 84818 543134
rect 91826 561218 92062 561454
rect 92146 561218 92382 561454
rect 91826 560898 92062 561134
rect 92146 560898 92382 561134
rect 66986 536378 67222 536614
rect 67306 536378 67542 536614
rect 66986 536058 67222 536294
rect 67306 536058 67542 536294
rect 63266 424658 63502 424894
rect 63586 424658 63822 424894
rect 63266 424338 63502 424574
rect 63586 424338 63822 424574
rect 66986 500378 67222 500614
rect 67306 500378 67542 500614
rect 66986 500058 67222 500294
rect 67306 500058 67542 500294
rect 66986 464378 67222 464614
rect 67306 464378 67542 464614
rect 66986 464058 67222 464294
rect 67306 464058 67542 464294
rect 63266 388658 63502 388894
rect 63586 388658 63822 388894
rect 63266 388338 63502 388574
rect 63586 388338 63822 388574
rect 63266 352658 63502 352894
rect 63586 352658 63822 352894
rect 63266 352338 63502 352574
rect 63586 352338 63822 352574
rect 66986 356378 67222 356614
rect 67306 356378 67542 356614
rect 66986 356058 67222 356294
rect 67306 356058 67542 356294
rect 63266 316658 63502 316894
rect 63586 316658 63822 316894
rect 63266 316338 63502 316574
rect 63586 316338 63822 316574
rect 59546 276938 59782 277174
rect 59866 276938 60102 277174
rect 59546 276618 59782 276854
rect 59866 276618 60102 276854
rect 55826 237218 56062 237454
rect 56146 237218 56382 237454
rect 55826 236898 56062 237134
rect 56146 236898 56382 237134
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 59546 240938 59782 241174
rect 59866 240938 60102 241174
rect 59546 240618 59782 240854
rect 59866 240618 60102 240854
rect 59546 204938 59782 205174
rect 59866 204938 60102 205174
rect 59546 204618 59782 204854
rect 59866 204618 60102 204854
rect 59546 168938 59782 169174
rect 59866 168938 60102 169174
rect 59546 168618 59782 168854
rect 59866 168618 60102 168854
rect 59546 132938 59782 133174
rect 59866 132938 60102 133174
rect 59546 132618 59782 132854
rect 59866 132618 60102 132854
rect 59546 96938 59782 97174
rect 59866 96938 60102 97174
rect 59546 96618 59782 96854
rect 59866 96618 60102 96854
rect 59546 60938 59782 61174
rect 59866 60938 60102 61174
rect 59546 60618 59782 60854
rect 59866 60618 60102 60854
rect 73826 507218 74062 507454
rect 74146 507218 74382 507454
rect 73826 506898 74062 507134
rect 74146 506898 74382 507134
rect 73826 471218 74062 471454
rect 74146 471218 74382 471454
rect 73826 470898 74062 471134
rect 74146 470898 74382 471134
rect 63266 280658 63502 280894
rect 63586 280658 63822 280894
rect 63266 280338 63502 280574
rect 63586 280338 63822 280574
rect 63266 244658 63502 244894
rect 63586 244658 63822 244894
rect 63266 244338 63502 244574
rect 63586 244338 63822 244574
rect 63266 208658 63502 208894
rect 63586 208658 63822 208894
rect 63266 208338 63502 208574
rect 63586 208338 63822 208574
rect 63266 172658 63502 172894
rect 63586 172658 63822 172894
rect 63266 172338 63502 172574
rect 63586 172338 63822 172574
rect 63266 136658 63502 136894
rect 63586 136658 63822 136894
rect 63266 136338 63502 136574
rect 63586 136338 63822 136574
rect 63266 100658 63502 100894
rect 63586 100658 63822 100894
rect 63266 100338 63502 100574
rect 63586 100338 63822 100574
rect 63266 64658 63502 64894
rect 63586 64658 63822 64894
rect 63266 64338 63502 64574
rect 63586 64338 63822 64574
rect 59546 24938 59782 25174
rect 59866 24938 60102 25174
rect 59546 24618 59782 24854
rect 59866 24618 60102 24854
rect 55826 -1542 56062 -1306
rect 56146 -1542 56382 -1306
rect 55826 -1862 56062 -1626
rect 56146 -1862 56382 -1626
rect 59546 -3462 59782 -3226
rect 59866 -3462 60102 -3226
rect 59546 -3782 59782 -3546
rect 59866 -3782 60102 -3546
rect 66986 212378 67222 212614
rect 67306 212378 67542 212614
rect 66986 212058 67222 212294
rect 67306 212058 67542 212294
rect 66986 68378 67222 68614
rect 67306 68378 67542 68614
rect 66986 68058 67222 68294
rect 67306 68058 67542 68294
rect 63266 28658 63502 28894
rect 63586 28658 63822 28894
rect 63266 28338 63502 28574
rect 63586 28338 63822 28574
rect 63266 -5382 63502 -5146
rect 63586 -5382 63822 -5146
rect 63266 -5702 63502 -5466
rect 63586 -5702 63822 -5466
rect 66986 32378 67222 32614
rect 67306 32378 67542 32614
rect 66986 32058 67222 32294
rect 67306 32058 67542 32294
rect 48986 -6342 49222 -6106
rect 49306 -6342 49542 -6106
rect 48986 -6662 49222 -6426
rect 49306 -6662 49542 -6426
rect 77546 510938 77782 511174
rect 77866 510938 78102 511174
rect 77546 510618 77782 510854
rect 77866 510618 78102 510854
rect 77546 474938 77782 475174
rect 77866 474938 78102 475174
rect 77546 474618 77782 474854
rect 77866 474618 78102 474854
rect 81266 514658 81502 514894
rect 81586 514658 81822 514894
rect 81266 514338 81502 514574
rect 81586 514338 81822 514574
rect 81266 478658 81502 478894
rect 81586 478658 81822 478894
rect 81266 478338 81502 478574
rect 81586 478338 81822 478574
rect 84986 518378 85222 518614
rect 85306 518378 85542 518614
rect 84986 518058 85222 518294
rect 85306 518058 85542 518294
rect 84986 482378 85222 482614
rect 85306 482378 85542 482614
rect 84986 482058 85222 482294
rect 85306 482058 85542 482294
rect 91826 525218 92062 525454
rect 92146 525218 92382 525454
rect 91826 524898 92062 525134
rect 92146 524898 92382 525134
rect 91826 489218 92062 489454
rect 92146 489218 92382 489454
rect 91826 488898 92062 489134
rect 92146 488898 92382 489134
rect 73020 435218 73256 435454
rect 73020 434898 73256 435134
rect 88380 417218 88616 417454
rect 88380 416898 88616 417134
rect 73020 399218 73256 399454
rect 73020 398898 73256 399134
rect 95546 672938 95782 673174
rect 95866 672938 96102 673174
rect 95546 672618 95782 672854
rect 95866 672618 96102 672854
rect 95546 636938 95782 637174
rect 95866 636938 96102 637174
rect 95546 636618 95782 636854
rect 95866 636618 96102 636854
rect 95546 600938 95782 601174
rect 95866 600938 96102 601174
rect 95546 600618 95782 600854
rect 95866 600618 96102 600854
rect 95546 564938 95782 565174
rect 95866 564938 96102 565174
rect 95546 564618 95782 564854
rect 95866 564618 96102 564854
rect 99266 676658 99502 676894
rect 99586 676658 99822 676894
rect 99266 676338 99502 676574
rect 99586 676338 99822 676574
rect 99266 640658 99502 640894
rect 99586 640658 99822 640894
rect 99266 640338 99502 640574
rect 99586 640338 99822 640574
rect 99266 604658 99502 604894
rect 99586 604658 99822 604894
rect 99266 604338 99502 604574
rect 99586 604338 99822 604574
rect 99266 568658 99502 568894
rect 99586 568658 99822 568894
rect 99266 568338 99502 568574
rect 99586 568338 99822 568574
rect 99266 532658 99502 532894
rect 99586 532658 99822 532894
rect 99266 532338 99502 532574
rect 99586 532338 99822 532574
rect 95546 528938 95782 529174
rect 95866 528938 96102 529174
rect 95546 528618 95782 528854
rect 95866 528618 96102 528854
rect 95546 492938 95782 493174
rect 95866 492938 96102 493174
rect 95546 492618 95782 492854
rect 95866 492618 96102 492854
rect 91826 453218 92062 453454
rect 92146 453218 92382 453454
rect 91826 452898 92062 453134
rect 92146 452898 92382 453134
rect 95546 456938 95782 457174
rect 95866 456938 96102 457174
rect 95546 456618 95782 456854
rect 95866 456618 96102 456854
rect 73826 363218 74062 363454
rect 74146 363218 74382 363454
rect 73826 362898 74062 363134
rect 74146 362898 74382 363134
rect 77546 366938 77782 367174
rect 77866 366938 78102 367174
rect 77546 366618 77782 366854
rect 77866 366618 78102 366854
rect 81266 370658 81502 370894
rect 81586 370658 81822 370894
rect 81266 370338 81502 370574
rect 81586 370338 81822 370574
rect 73020 291218 73256 291454
rect 73020 290898 73256 291134
rect 73020 255218 73256 255454
rect 73020 254898 73256 255134
rect 73826 219218 74062 219454
rect 74146 219218 74382 219454
rect 73826 218898 74062 219134
rect 74146 218898 74382 219134
rect 81266 334658 81502 334894
rect 81586 334658 81822 334894
rect 81266 334338 81502 334574
rect 81586 334338 81822 334574
rect 77546 222938 77782 223174
rect 77866 222938 78102 223174
rect 77546 222618 77782 222854
rect 77866 222618 78102 222854
rect 73826 183218 74062 183454
rect 74146 183218 74382 183454
rect 73826 182898 74062 183134
rect 74146 182898 74382 183134
rect 77546 186938 77782 187174
rect 77866 186938 78102 187174
rect 77546 186618 77782 186854
rect 77866 186618 78102 186854
rect 84986 374378 85222 374614
rect 85306 374378 85542 374614
rect 84986 374058 85222 374294
rect 85306 374058 85542 374294
rect 84986 338378 85222 338614
rect 85306 338378 85542 338614
rect 84986 338058 85222 338294
rect 85306 338058 85542 338294
rect 91826 381218 92062 381454
rect 92146 381218 92382 381454
rect 91826 380898 92062 381134
rect 92146 380898 92382 381134
rect 99266 496658 99502 496894
rect 99586 496658 99822 496894
rect 99266 496338 99502 496574
rect 99586 496338 99822 496574
rect 99266 460658 99502 460894
rect 99586 460658 99822 460894
rect 99266 460338 99502 460574
rect 99586 460338 99822 460574
rect 120986 710362 121222 710598
rect 121306 710362 121542 710598
rect 120986 710042 121222 710278
rect 121306 710042 121542 710278
rect 117266 708442 117502 708678
rect 117586 708442 117822 708678
rect 117266 708122 117502 708358
rect 117586 708122 117822 708358
rect 113546 706522 113782 706758
rect 113866 706522 114102 706758
rect 113546 706202 113782 706438
rect 113866 706202 114102 706438
rect 102986 680378 103222 680614
rect 103306 680378 103542 680614
rect 102986 680058 103222 680294
rect 103306 680058 103542 680294
rect 102986 644378 103222 644614
rect 103306 644378 103542 644614
rect 102986 644058 103222 644294
rect 103306 644058 103542 644294
rect 102986 608378 103222 608614
rect 103306 608378 103542 608614
rect 102986 608058 103222 608294
rect 103306 608058 103542 608294
rect 102986 572378 103222 572614
rect 103306 572378 103542 572614
rect 102986 572058 103222 572294
rect 103306 572058 103542 572294
rect 102986 536378 103222 536614
rect 103306 536378 103542 536614
rect 102986 536058 103222 536294
rect 103306 536058 103542 536294
rect 102986 500378 103222 500614
rect 103306 500378 103542 500614
rect 102986 500058 103222 500294
rect 103306 500058 103542 500294
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 109826 615218 110062 615454
rect 110146 615218 110382 615454
rect 109826 614898 110062 615134
rect 110146 614898 110382 615134
rect 109826 579218 110062 579454
rect 110146 579218 110382 579454
rect 109826 578898 110062 579134
rect 110146 578898 110382 579134
rect 109826 543218 110062 543454
rect 110146 543218 110382 543454
rect 109826 542898 110062 543134
rect 110146 542898 110382 543134
rect 109826 507218 110062 507454
rect 110146 507218 110382 507454
rect 109826 506898 110062 507134
rect 110146 506898 110382 507134
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 102986 464378 103222 464614
rect 103306 464378 103542 464614
rect 102986 464058 103222 464294
rect 103306 464058 103542 464294
rect 95546 384938 95782 385174
rect 95866 384938 96102 385174
rect 95546 384618 95782 384854
rect 95866 384618 96102 384854
rect 95546 348938 95782 349174
rect 95866 348938 96102 349174
rect 95546 348618 95782 348854
rect 95866 348618 96102 348854
rect 91826 345218 92062 345454
rect 92146 345218 92382 345454
rect 91826 344898 92062 345134
rect 92146 344898 92382 345134
rect 103740 435218 103976 435454
rect 103740 434898 103976 435134
rect 103740 399218 103976 399454
rect 103740 398898 103976 399134
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 113546 690938 113782 691174
rect 113866 690938 114102 691174
rect 113546 690618 113782 690854
rect 113866 690618 114102 690854
rect 113546 654938 113782 655174
rect 113866 654938 114102 655174
rect 113546 654618 113782 654854
rect 113866 654618 114102 654854
rect 113546 618938 113782 619174
rect 113866 618938 114102 619174
rect 113546 618618 113782 618854
rect 113866 618618 114102 618854
rect 113546 582938 113782 583174
rect 113866 582938 114102 583174
rect 113546 582618 113782 582854
rect 113866 582618 114102 582854
rect 113546 546938 113782 547174
rect 113866 546938 114102 547174
rect 113546 546618 113782 546854
rect 113866 546618 114102 546854
rect 113546 510938 113782 511174
rect 113866 510938 114102 511174
rect 113546 510618 113782 510854
rect 113866 510618 114102 510854
rect 113546 474938 113782 475174
rect 113866 474938 114102 475174
rect 113546 474618 113782 474854
rect 113866 474618 114102 474854
rect 109826 363218 110062 363454
rect 110146 363218 110382 363454
rect 109826 362898 110062 363134
rect 110146 362898 110382 363134
rect 102986 356378 103222 356614
rect 103306 356378 103542 356614
rect 102986 356058 103222 356294
rect 103306 356058 103542 356294
rect 99266 352658 99502 352894
rect 99586 352658 99822 352894
rect 99266 352338 99502 352574
rect 99586 352338 99822 352574
rect 117266 694658 117502 694894
rect 117586 694658 117822 694894
rect 117266 694338 117502 694574
rect 117586 694338 117822 694574
rect 117266 658658 117502 658894
rect 117586 658658 117822 658894
rect 117266 658338 117502 658574
rect 117586 658338 117822 658574
rect 117266 622658 117502 622894
rect 117586 622658 117822 622894
rect 117266 622338 117502 622574
rect 117586 622338 117822 622574
rect 117266 586658 117502 586894
rect 117586 586658 117822 586894
rect 117266 586338 117502 586574
rect 117586 586338 117822 586574
rect 117266 550658 117502 550894
rect 117586 550658 117822 550894
rect 117266 550338 117502 550574
rect 117586 550338 117822 550574
rect 117266 514658 117502 514894
rect 117586 514658 117822 514894
rect 117266 514338 117502 514574
rect 117586 514338 117822 514574
rect 117266 478658 117502 478894
rect 117586 478658 117822 478894
rect 117266 478338 117502 478574
rect 117586 478338 117822 478574
rect 113546 366938 113782 367174
rect 113866 366938 114102 367174
rect 113546 366618 113782 366854
rect 113866 366618 114102 366854
rect 138986 711322 139222 711558
rect 139306 711322 139542 711558
rect 138986 711002 139222 711238
rect 139306 711002 139542 711238
rect 135266 709402 135502 709638
rect 135586 709402 135822 709638
rect 135266 709082 135502 709318
rect 135586 709082 135822 709318
rect 131546 707482 131782 707718
rect 131866 707482 132102 707718
rect 131546 707162 131782 707398
rect 131866 707162 132102 707398
rect 120986 698378 121222 698614
rect 121306 698378 121542 698614
rect 120986 698058 121222 698294
rect 121306 698058 121542 698294
rect 120986 662378 121222 662614
rect 121306 662378 121542 662614
rect 120986 662058 121222 662294
rect 121306 662058 121542 662294
rect 120986 626378 121222 626614
rect 121306 626378 121542 626614
rect 120986 626058 121222 626294
rect 121306 626058 121542 626294
rect 120986 590378 121222 590614
rect 121306 590378 121542 590614
rect 120986 590058 121222 590294
rect 121306 590058 121542 590294
rect 120986 554378 121222 554614
rect 121306 554378 121542 554614
rect 120986 554058 121222 554294
rect 121306 554058 121542 554294
rect 120986 518378 121222 518614
rect 121306 518378 121542 518614
rect 120986 518058 121222 518294
rect 121306 518058 121542 518294
rect 120986 482378 121222 482614
rect 121306 482378 121542 482614
rect 120986 482058 121222 482294
rect 121306 482058 121542 482294
rect 117266 370658 117502 370894
rect 117586 370658 117822 370894
rect 117266 370338 117502 370574
rect 117586 370338 117822 370574
rect 119100 417218 119336 417454
rect 119100 416898 119336 417134
rect 127826 705562 128062 705798
rect 128146 705562 128382 705798
rect 127826 705242 128062 705478
rect 128146 705242 128382 705478
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 127826 597218 128062 597454
rect 128146 597218 128382 597454
rect 127826 596898 128062 597134
rect 128146 596898 128382 597134
rect 127826 561218 128062 561454
rect 128146 561218 128382 561454
rect 127826 560898 128062 561134
rect 128146 560898 128382 561134
rect 127826 525218 128062 525454
rect 128146 525218 128382 525454
rect 127826 524898 128062 525134
rect 128146 524898 128382 525134
rect 127826 489218 128062 489454
rect 128146 489218 128382 489454
rect 127826 488898 128062 489134
rect 128146 488898 128382 489134
rect 120986 374378 121222 374614
rect 121306 374378 121542 374614
rect 120986 374058 121222 374294
rect 121306 374058 121542 374294
rect 117266 334658 117502 334894
rect 117586 334658 117822 334894
rect 117266 334338 117502 334574
rect 117586 334338 117822 334574
rect 127826 453218 128062 453454
rect 128146 453218 128382 453454
rect 127826 452898 128062 453134
rect 128146 452898 128382 453134
rect 127826 417218 128062 417454
rect 128146 417218 128382 417454
rect 127826 416898 128062 417134
rect 128146 416898 128382 417134
rect 127826 381218 128062 381454
rect 128146 381218 128382 381454
rect 127826 380898 128062 381134
rect 128146 380898 128382 381134
rect 120986 338378 121222 338614
rect 121306 338378 121542 338614
rect 120986 338058 121222 338294
rect 121306 338058 121542 338294
rect 127826 345218 128062 345454
rect 128146 345218 128382 345454
rect 127826 344898 128062 345134
rect 128146 344898 128382 345134
rect 131546 672938 131782 673174
rect 131866 672938 132102 673174
rect 131546 672618 131782 672854
rect 131866 672618 132102 672854
rect 131546 636938 131782 637174
rect 131866 636938 132102 637174
rect 131546 636618 131782 636854
rect 131866 636618 132102 636854
rect 131546 600938 131782 601174
rect 131866 600938 132102 601174
rect 131546 600618 131782 600854
rect 131866 600618 132102 600854
rect 131546 564938 131782 565174
rect 131866 564938 132102 565174
rect 131546 564618 131782 564854
rect 131866 564618 132102 564854
rect 131546 528938 131782 529174
rect 131866 528938 132102 529174
rect 131546 528618 131782 528854
rect 131866 528618 132102 528854
rect 131546 492938 131782 493174
rect 131866 492938 132102 493174
rect 131546 492618 131782 492854
rect 131866 492618 132102 492854
rect 131546 456938 131782 457174
rect 131866 456938 132102 457174
rect 131546 456618 131782 456854
rect 131866 456618 132102 456854
rect 131546 420938 131782 421174
rect 131866 420938 132102 421174
rect 131546 420618 131782 420854
rect 131866 420618 132102 420854
rect 131546 384938 131782 385174
rect 131866 384938 132102 385174
rect 131546 384618 131782 384854
rect 131866 384618 132102 384854
rect 131546 348938 131782 349174
rect 131866 348938 132102 349174
rect 131546 348618 131782 348854
rect 131866 348618 132102 348854
rect 135266 676658 135502 676894
rect 135586 676658 135822 676894
rect 135266 676338 135502 676574
rect 135586 676338 135822 676574
rect 135266 640658 135502 640894
rect 135586 640658 135822 640894
rect 135266 640338 135502 640574
rect 135586 640338 135822 640574
rect 135266 604658 135502 604894
rect 135586 604658 135822 604894
rect 135266 604338 135502 604574
rect 135586 604338 135822 604574
rect 135266 568658 135502 568894
rect 135586 568658 135822 568894
rect 135266 568338 135502 568574
rect 135586 568338 135822 568574
rect 135266 532658 135502 532894
rect 135586 532658 135822 532894
rect 135266 532338 135502 532574
rect 135586 532338 135822 532574
rect 135266 496658 135502 496894
rect 135586 496658 135822 496894
rect 135266 496338 135502 496574
rect 135586 496338 135822 496574
rect 135266 460658 135502 460894
rect 135586 460658 135822 460894
rect 135266 460338 135502 460574
rect 135586 460338 135822 460574
rect 135266 424658 135502 424894
rect 135586 424658 135822 424894
rect 135266 424338 135502 424574
rect 135586 424338 135822 424574
rect 135266 388658 135502 388894
rect 135586 388658 135822 388894
rect 135266 388338 135502 388574
rect 135586 388338 135822 388574
rect 135266 352658 135502 352894
rect 135586 352658 135822 352894
rect 135266 352338 135502 352574
rect 135586 352338 135822 352574
rect 156986 710362 157222 710598
rect 157306 710362 157542 710598
rect 156986 710042 157222 710278
rect 157306 710042 157542 710278
rect 153266 708442 153502 708678
rect 153586 708442 153822 708678
rect 153266 708122 153502 708358
rect 153586 708122 153822 708358
rect 149546 706522 149782 706758
rect 149866 706522 150102 706758
rect 149546 706202 149782 706438
rect 149866 706202 150102 706438
rect 138986 680378 139222 680614
rect 139306 680378 139542 680614
rect 138986 680058 139222 680294
rect 139306 680058 139542 680294
rect 138986 644378 139222 644614
rect 139306 644378 139542 644614
rect 138986 644058 139222 644294
rect 139306 644058 139542 644294
rect 138986 608378 139222 608614
rect 139306 608378 139542 608614
rect 138986 608058 139222 608294
rect 139306 608058 139542 608294
rect 138986 572378 139222 572614
rect 139306 572378 139542 572614
rect 138986 572058 139222 572294
rect 139306 572058 139542 572294
rect 138986 536378 139222 536614
rect 139306 536378 139542 536614
rect 138986 536058 139222 536294
rect 139306 536058 139542 536294
rect 138986 500378 139222 500614
rect 139306 500378 139542 500614
rect 138986 500058 139222 500294
rect 139306 500058 139542 500294
rect 138986 464378 139222 464614
rect 139306 464378 139542 464614
rect 138986 464058 139222 464294
rect 139306 464058 139542 464294
rect 138986 428378 139222 428614
rect 139306 428378 139542 428614
rect 138986 428058 139222 428294
rect 139306 428058 139542 428294
rect 138986 392378 139222 392614
rect 139306 392378 139542 392614
rect 138986 392058 139222 392294
rect 139306 392058 139542 392294
rect 138986 356378 139222 356614
rect 139306 356378 139542 356614
rect 138986 356058 139222 356294
rect 139306 356058 139542 356294
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 145826 543218 146062 543454
rect 146146 543218 146382 543454
rect 145826 542898 146062 543134
rect 146146 542898 146382 543134
rect 145826 507218 146062 507454
rect 146146 507218 146382 507454
rect 145826 506898 146062 507134
rect 146146 506898 146382 507134
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 145826 435218 146062 435454
rect 146146 435218 146382 435454
rect 145826 434898 146062 435134
rect 146146 434898 146382 435134
rect 145826 399218 146062 399454
rect 146146 399218 146382 399454
rect 145826 398898 146062 399134
rect 146146 398898 146382 399134
rect 145826 363218 146062 363454
rect 146146 363218 146382 363454
rect 145826 362898 146062 363134
rect 146146 362898 146382 363134
rect 149546 690938 149782 691174
rect 149866 690938 150102 691174
rect 149546 690618 149782 690854
rect 149866 690618 150102 690854
rect 149546 654938 149782 655174
rect 149866 654938 150102 655174
rect 149546 654618 149782 654854
rect 149866 654618 150102 654854
rect 149546 618938 149782 619174
rect 149866 618938 150102 619174
rect 149546 618618 149782 618854
rect 149866 618618 150102 618854
rect 149546 582938 149782 583174
rect 149866 582938 150102 583174
rect 149546 582618 149782 582854
rect 149866 582618 150102 582854
rect 149546 546938 149782 547174
rect 149866 546938 150102 547174
rect 149546 546618 149782 546854
rect 149866 546618 150102 546854
rect 149546 510938 149782 511174
rect 149866 510938 150102 511174
rect 149546 510618 149782 510854
rect 149866 510618 150102 510854
rect 149546 474938 149782 475174
rect 149866 474938 150102 475174
rect 149546 474618 149782 474854
rect 149866 474618 150102 474854
rect 149546 438938 149782 439174
rect 149866 438938 150102 439174
rect 149546 438618 149782 438854
rect 149866 438618 150102 438854
rect 149546 402938 149782 403174
rect 149866 402938 150102 403174
rect 149546 402618 149782 402854
rect 149866 402618 150102 402854
rect 149546 366938 149782 367174
rect 149866 366938 150102 367174
rect 149546 366618 149782 366854
rect 149866 366618 150102 366854
rect 153266 694658 153502 694894
rect 153586 694658 153822 694894
rect 153266 694338 153502 694574
rect 153586 694338 153822 694574
rect 153266 658658 153502 658894
rect 153586 658658 153822 658894
rect 153266 658338 153502 658574
rect 153586 658338 153822 658574
rect 153266 622658 153502 622894
rect 153586 622658 153822 622894
rect 153266 622338 153502 622574
rect 153586 622338 153822 622574
rect 153266 586658 153502 586894
rect 153586 586658 153822 586894
rect 153266 586338 153502 586574
rect 153586 586338 153822 586574
rect 153266 550658 153502 550894
rect 153586 550658 153822 550894
rect 153266 550338 153502 550574
rect 153586 550338 153822 550574
rect 153266 514658 153502 514894
rect 153586 514658 153822 514894
rect 153266 514338 153502 514574
rect 153586 514338 153822 514574
rect 153266 478658 153502 478894
rect 153586 478658 153822 478894
rect 153266 478338 153502 478574
rect 153586 478338 153822 478574
rect 153266 442658 153502 442894
rect 153586 442658 153822 442894
rect 153266 442338 153502 442574
rect 153586 442338 153822 442574
rect 174986 711322 175222 711558
rect 175306 711322 175542 711558
rect 174986 711002 175222 711238
rect 175306 711002 175542 711238
rect 171266 709402 171502 709638
rect 171586 709402 171822 709638
rect 171266 709082 171502 709318
rect 171586 709082 171822 709318
rect 167546 707482 167782 707718
rect 167866 707482 168102 707718
rect 167546 707162 167782 707398
rect 167866 707162 168102 707398
rect 156986 698378 157222 698614
rect 157306 698378 157542 698614
rect 156986 698058 157222 698294
rect 157306 698058 157542 698294
rect 156986 662378 157222 662614
rect 157306 662378 157542 662614
rect 156986 662058 157222 662294
rect 157306 662058 157542 662294
rect 156986 626378 157222 626614
rect 157306 626378 157542 626614
rect 156986 626058 157222 626294
rect 157306 626058 157542 626294
rect 156986 590378 157222 590614
rect 157306 590378 157542 590614
rect 156986 590058 157222 590294
rect 157306 590058 157542 590294
rect 156986 554378 157222 554614
rect 157306 554378 157542 554614
rect 156986 554058 157222 554294
rect 157306 554058 157542 554294
rect 163826 705562 164062 705798
rect 164146 705562 164382 705798
rect 163826 705242 164062 705478
rect 164146 705242 164382 705478
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 163826 633218 164062 633454
rect 164146 633218 164382 633454
rect 163826 632898 164062 633134
rect 164146 632898 164382 633134
rect 163826 597218 164062 597454
rect 164146 597218 164382 597454
rect 163826 596898 164062 597134
rect 164146 596898 164382 597134
rect 163826 561218 164062 561454
rect 164146 561218 164382 561454
rect 163826 560898 164062 561134
rect 164146 560898 164382 561134
rect 163826 525218 164062 525454
rect 164146 525218 164382 525454
rect 163826 524898 164062 525134
rect 164146 524898 164382 525134
rect 156986 518378 157222 518614
rect 157306 518378 157542 518614
rect 156986 518058 157222 518294
rect 157306 518058 157542 518294
rect 156986 482378 157222 482614
rect 157306 482378 157542 482614
rect 156986 482058 157222 482294
rect 157306 482058 157542 482294
rect 156986 446378 157222 446614
rect 157306 446378 157542 446614
rect 156986 446058 157222 446294
rect 157306 446058 157542 446294
rect 153266 406658 153502 406894
rect 153586 406658 153822 406894
rect 153266 406338 153502 406574
rect 153586 406338 153822 406574
rect 153266 370658 153502 370894
rect 153586 370658 153822 370894
rect 153266 370338 153502 370574
rect 153586 370338 153822 370574
rect 153266 334658 153502 334894
rect 153586 334658 153822 334894
rect 153266 334338 153502 334574
rect 153586 334338 153822 334574
rect 88380 309218 88616 309454
rect 88380 308898 88616 309134
rect 119100 309218 119336 309454
rect 119100 308898 119336 309134
rect 149820 309218 150056 309454
rect 149820 308898 150056 309134
rect 103740 291218 103976 291454
rect 103740 290898 103976 291134
rect 134460 291218 134696 291454
rect 134460 290898 134696 291134
rect 88380 273218 88616 273454
rect 88380 272898 88616 273134
rect 119100 273218 119336 273454
rect 119100 272898 119336 273134
rect 149820 273218 150056 273454
rect 149820 272898 150056 273134
rect 103740 255218 103976 255454
rect 103740 254898 103976 255134
rect 134460 255218 134696 255454
rect 134460 254898 134696 255134
rect 81266 226658 81502 226894
rect 81586 226658 81822 226894
rect 81266 226338 81502 226574
rect 81586 226338 81822 226574
rect 81266 190658 81502 190894
rect 81586 190658 81822 190894
rect 81266 190338 81502 190574
rect 81586 190338 81822 190574
rect 84986 230378 85222 230614
rect 85306 230378 85542 230614
rect 84986 230058 85222 230294
rect 85306 230058 85542 230294
rect 84986 194378 85222 194614
rect 85306 194378 85542 194614
rect 84986 194058 85222 194294
rect 85306 194058 85542 194294
rect 91826 237218 92062 237454
rect 92146 237218 92382 237454
rect 91826 236898 92062 237134
rect 92146 236898 92382 237134
rect 91826 201218 92062 201454
rect 92146 201218 92382 201454
rect 91826 200898 92062 201134
rect 92146 200898 92382 201134
rect 95546 204938 95782 205174
rect 95866 204938 96102 205174
rect 95546 204618 95782 204854
rect 95866 204618 96102 204854
rect 99266 208658 99502 208894
rect 99586 208658 99822 208894
rect 99266 208338 99502 208574
rect 99586 208338 99822 208574
rect 102986 212378 103222 212614
rect 103306 212378 103542 212614
rect 102986 212058 103222 212294
rect 103306 212058 103542 212294
rect 109826 219218 110062 219454
rect 110146 219218 110382 219454
rect 109826 218898 110062 219134
rect 110146 218898 110382 219134
rect 109826 183218 110062 183454
rect 110146 183218 110382 183454
rect 109826 182898 110062 183134
rect 110146 182898 110382 183134
rect 113546 222938 113782 223174
rect 113866 222938 114102 223174
rect 113546 222618 113782 222854
rect 113866 222618 114102 222854
rect 113546 186938 113782 187174
rect 113866 186938 114102 187174
rect 113546 186618 113782 186854
rect 113866 186618 114102 186854
rect 117266 226658 117502 226894
rect 117586 226658 117822 226894
rect 117266 226338 117502 226574
rect 117586 226338 117822 226574
rect 117266 190658 117502 190894
rect 117586 190658 117822 190894
rect 117266 190338 117502 190574
rect 117586 190338 117822 190574
rect 120986 230378 121222 230614
rect 121306 230378 121542 230614
rect 120986 230058 121222 230294
rect 121306 230058 121542 230294
rect 120986 194378 121222 194614
rect 121306 194378 121542 194614
rect 120986 194058 121222 194294
rect 121306 194058 121542 194294
rect 127826 237218 128062 237454
rect 128146 237218 128382 237454
rect 127826 236898 128062 237134
rect 128146 236898 128382 237134
rect 127826 201218 128062 201454
rect 128146 201218 128382 201454
rect 127826 200898 128062 201134
rect 128146 200898 128382 201134
rect 131546 204938 131782 205174
rect 131866 204938 132102 205174
rect 131546 204618 131782 204854
rect 131866 204618 132102 204854
rect 135266 208658 135502 208894
rect 135586 208658 135822 208894
rect 135266 208338 135502 208574
rect 135586 208338 135822 208574
rect 138986 212378 139222 212614
rect 139306 212378 139542 212614
rect 138986 212058 139222 212294
rect 139306 212058 139542 212294
rect 145826 219218 146062 219454
rect 146146 219218 146382 219454
rect 145826 218898 146062 219134
rect 146146 218898 146382 219134
rect 145826 183218 146062 183454
rect 146146 183218 146382 183454
rect 145826 182898 146062 183134
rect 146146 182898 146382 183134
rect 149546 222938 149782 223174
rect 149866 222938 150102 223174
rect 149546 222618 149782 222854
rect 149866 222618 150102 222854
rect 149546 186938 149782 187174
rect 149866 186938 150102 187174
rect 149546 186618 149782 186854
rect 149866 186618 150102 186854
rect 156986 410378 157222 410614
rect 157306 410378 157542 410614
rect 156986 410058 157222 410294
rect 157306 410058 157542 410294
rect 156986 374378 157222 374614
rect 157306 374378 157542 374614
rect 156986 374058 157222 374294
rect 157306 374058 157542 374294
rect 156986 338378 157222 338614
rect 157306 338378 157542 338614
rect 156986 338058 157222 338294
rect 157306 338058 157542 338294
rect 153266 226658 153502 226894
rect 153586 226658 153822 226894
rect 153266 226338 153502 226574
rect 153586 226338 153822 226574
rect 153266 190658 153502 190894
rect 153586 190658 153822 190894
rect 153266 190338 153502 190574
rect 153586 190338 153822 190574
rect 156986 230378 157222 230614
rect 157306 230378 157542 230614
rect 156986 230058 157222 230294
rect 157306 230058 157542 230294
rect 163826 489218 164062 489454
rect 164146 489218 164382 489454
rect 163826 488898 164062 489134
rect 164146 488898 164382 489134
rect 163826 453218 164062 453454
rect 164146 453218 164382 453454
rect 163826 452898 164062 453134
rect 164146 452898 164382 453134
rect 163826 417218 164062 417454
rect 164146 417218 164382 417454
rect 163826 416898 164062 417134
rect 164146 416898 164382 417134
rect 163826 381218 164062 381454
rect 164146 381218 164382 381454
rect 163826 380898 164062 381134
rect 164146 380898 164382 381134
rect 167546 672938 167782 673174
rect 167866 672938 168102 673174
rect 167546 672618 167782 672854
rect 167866 672618 168102 672854
rect 167546 636938 167782 637174
rect 167866 636938 168102 637174
rect 167546 636618 167782 636854
rect 167866 636618 168102 636854
rect 167546 600938 167782 601174
rect 167866 600938 168102 601174
rect 167546 600618 167782 600854
rect 167866 600618 168102 600854
rect 167546 564938 167782 565174
rect 167866 564938 168102 565174
rect 167546 564618 167782 564854
rect 167866 564618 168102 564854
rect 171266 676658 171502 676894
rect 171586 676658 171822 676894
rect 171266 676338 171502 676574
rect 171586 676338 171822 676574
rect 171266 640658 171502 640894
rect 171586 640658 171822 640894
rect 171266 640338 171502 640574
rect 171586 640338 171822 640574
rect 171266 604658 171502 604894
rect 171586 604658 171822 604894
rect 171266 604338 171502 604574
rect 171586 604338 171822 604574
rect 171266 568658 171502 568894
rect 171586 568658 171822 568894
rect 171266 568338 171502 568574
rect 171586 568338 171822 568574
rect 167546 528938 167782 529174
rect 167866 528938 168102 529174
rect 167546 528618 167782 528854
rect 167866 528618 168102 528854
rect 167546 492938 167782 493174
rect 167866 492938 168102 493174
rect 167546 492618 167782 492854
rect 167866 492618 168102 492854
rect 167546 456938 167782 457174
rect 167866 456938 168102 457174
rect 167546 456618 167782 456854
rect 167866 456618 168102 456854
rect 167546 420938 167782 421174
rect 167866 420938 168102 421174
rect 167546 420618 167782 420854
rect 167866 420618 168102 420854
rect 167546 384938 167782 385174
rect 167866 384938 168102 385174
rect 167546 384618 167782 384854
rect 167866 384618 168102 384854
rect 163826 345218 164062 345454
rect 164146 345218 164382 345454
rect 163826 344898 164062 345134
rect 164146 344898 164382 345134
rect 167546 348938 167782 349174
rect 167866 348938 168102 349174
rect 167546 348618 167782 348854
rect 167866 348618 168102 348854
rect 163826 309218 164062 309454
rect 164146 309218 164382 309454
rect 163826 308898 164062 309134
rect 164146 308898 164382 309134
rect 163826 273218 164062 273454
rect 164146 273218 164382 273454
rect 163826 272898 164062 273134
rect 164146 272898 164382 273134
rect 156986 194378 157222 194614
rect 157306 194378 157542 194614
rect 156986 194058 157222 194294
rect 157306 194058 157542 194294
rect 163826 237218 164062 237454
rect 164146 237218 164382 237454
rect 163826 236898 164062 237134
rect 164146 236898 164382 237134
rect 163826 201218 164062 201454
rect 164146 201218 164382 201454
rect 163826 200898 164062 201134
rect 164146 200898 164382 201134
rect 69128 165218 69364 165454
rect 69128 164898 69364 165134
rect 164192 165218 164428 165454
rect 164192 164898 164428 165134
rect 69808 147218 70044 147454
rect 69808 146898 70044 147134
rect 163512 147218 163748 147454
rect 163512 146898 163748 147134
rect 69128 129218 69364 129454
rect 69128 128898 69364 129134
rect 164192 129218 164428 129454
rect 164192 128898 164428 129134
rect 69808 111218 70044 111454
rect 69808 110898 70044 111134
rect 163512 111218 163748 111454
rect 163512 110898 163748 111134
rect 73826 75218 74062 75454
rect 74146 75218 74382 75454
rect 73826 74898 74062 75134
rect 74146 74898 74382 75134
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 77546 78938 77782 79174
rect 77866 78938 78102 79174
rect 77546 78618 77782 78854
rect 77866 78618 78102 78854
rect 77546 42938 77782 43174
rect 77866 42938 78102 43174
rect 77546 42618 77782 42854
rect 77866 42618 78102 42854
rect 77546 6938 77782 7174
rect 77866 6938 78102 7174
rect 77546 6618 77782 6854
rect 77866 6618 78102 6854
rect 77546 -2502 77782 -2266
rect 77866 -2502 78102 -2266
rect 77546 -2822 77782 -2586
rect 77866 -2822 78102 -2586
rect 81266 82658 81502 82894
rect 81586 82658 81822 82894
rect 81266 82338 81502 82574
rect 81586 82338 81822 82574
rect 81266 46658 81502 46894
rect 81586 46658 81822 46894
rect 81266 46338 81502 46574
rect 81586 46338 81822 46574
rect 81266 10658 81502 10894
rect 81586 10658 81822 10894
rect 81266 10338 81502 10574
rect 81586 10338 81822 10574
rect 81266 -4422 81502 -4186
rect 81586 -4422 81822 -4186
rect 81266 -4742 81502 -4506
rect 81586 -4742 81822 -4506
rect 84986 86378 85222 86614
rect 85306 86378 85542 86614
rect 84986 86058 85222 86294
rect 85306 86058 85542 86294
rect 84986 50378 85222 50614
rect 85306 50378 85542 50614
rect 84986 50058 85222 50294
rect 85306 50058 85542 50294
rect 84986 14378 85222 14614
rect 85306 14378 85542 14614
rect 84986 14058 85222 14294
rect 85306 14058 85542 14294
rect 66986 -7302 67222 -7066
rect 67306 -7302 67542 -7066
rect 66986 -7622 67222 -7386
rect 67306 -7622 67542 -7386
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -1542 92062 -1306
rect 92146 -1542 92382 -1306
rect 91826 -1862 92062 -1626
rect 92146 -1862 92382 -1626
rect 95546 60938 95782 61174
rect 95866 60938 96102 61174
rect 95546 60618 95782 60854
rect 95866 60618 96102 60854
rect 95546 24938 95782 25174
rect 95866 24938 96102 25174
rect 95546 24618 95782 24854
rect 95866 24618 96102 24854
rect 95546 -3462 95782 -3226
rect 95866 -3462 96102 -3226
rect 95546 -3782 95782 -3546
rect 95866 -3782 96102 -3546
rect 99266 64658 99502 64894
rect 99586 64658 99822 64894
rect 99266 64338 99502 64574
rect 99586 64338 99822 64574
rect 99266 28658 99502 28894
rect 99586 28658 99822 28894
rect 99266 28338 99502 28574
rect 99586 28338 99822 28574
rect 99266 -5382 99502 -5146
rect 99586 -5382 99822 -5146
rect 99266 -5702 99502 -5466
rect 99586 -5702 99822 -5466
rect 102986 68378 103222 68614
rect 103306 68378 103542 68614
rect 102986 68058 103222 68294
rect 103306 68058 103542 68294
rect 102986 32378 103222 32614
rect 103306 32378 103542 32614
rect 102986 32058 103222 32294
rect 103306 32058 103542 32294
rect 84986 -6342 85222 -6106
rect 85306 -6342 85542 -6106
rect 84986 -6662 85222 -6426
rect 85306 -6662 85542 -6426
rect 109826 75218 110062 75454
rect 110146 75218 110382 75454
rect 109826 74898 110062 75134
rect 110146 74898 110382 75134
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 113546 78938 113782 79174
rect 113866 78938 114102 79174
rect 113546 78618 113782 78854
rect 113866 78618 114102 78854
rect 113546 42938 113782 43174
rect 113866 42938 114102 43174
rect 113546 42618 113782 42854
rect 113866 42618 114102 42854
rect 113546 6938 113782 7174
rect 113866 6938 114102 7174
rect 113546 6618 113782 6854
rect 113866 6618 114102 6854
rect 113546 -2502 113782 -2266
rect 113866 -2502 114102 -2266
rect 113546 -2822 113782 -2586
rect 113866 -2822 114102 -2586
rect 117266 82658 117502 82894
rect 117586 82658 117822 82894
rect 117266 82338 117502 82574
rect 117586 82338 117822 82574
rect 117266 46658 117502 46894
rect 117586 46658 117822 46894
rect 117266 46338 117502 46574
rect 117586 46338 117822 46574
rect 117266 10658 117502 10894
rect 117586 10658 117822 10894
rect 117266 10338 117502 10574
rect 117586 10338 117822 10574
rect 117266 -4422 117502 -4186
rect 117586 -4422 117822 -4186
rect 117266 -4742 117502 -4506
rect 117586 -4742 117822 -4506
rect 120986 86378 121222 86614
rect 121306 86378 121542 86614
rect 120986 86058 121222 86294
rect 121306 86058 121542 86294
rect 120986 50378 121222 50614
rect 121306 50378 121542 50614
rect 120986 50058 121222 50294
rect 121306 50058 121542 50294
rect 120986 14378 121222 14614
rect 121306 14378 121542 14614
rect 120986 14058 121222 14294
rect 121306 14058 121542 14294
rect 102986 -7302 103222 -7066
rect 103306 -7302 103542 -7066
rect 102986 -7622 103222 -7386
rect 103306 -7622 103542 -7386
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -1542 128062 -1306
rect 128146 -1542 128382 -1306
rect 127826 -1862 128062 -1626
rect 128146 -1862 128382 -1626
rect 131546 60938 131782 61174
rect 131866 60938 132102 61174
rect 131546 60618 131782 60854
rect 131866 60618 132102 60854
rect 131546 24938 131782 25174
rect 131866 24938 132102 25174
rect 131546 24618 131782 24854
rect 131866 24618 132102 24854
rect 131546 -3462 131782 -3226
rect 131866 -3462 132102 -3226
rect 131546 -3782 131782 -3546
rect 131866 -3782 132102 -3546
rect 135266 64658 135502 64894
rect 135586 64658 135822 64894
rect 135266 64338 135502 64574
rect 135586 64338 135822 64574
rect 135266 28658 135502 28894
rect 135586 28658 135822 28894
rect 135266 28338 135502 28574
rect 135586 28338 135822 28574
rect 135266 -5382 135502 -5146
rect 135586 -5382 135822 -5146
rect 135266 -5702 135502 -5466
rect 135586 -5702 135822 -5466
rect 138986 68378 139222 68614
rect 139306 68378 139542 68614
rect 138986 68058 139222 68294
rect 139306 68058 139542 68294
rect 138986 32378 139222 32614
rect 139306 32378 139542 32614
rect 138986 32058 139222 32294
rect 139306 32058 139542 32294
rect 120986 -6342 121222 -6106
rect 121306 -6342 121542 -6106
rect 120986 -6662 121222 -6426
rect 121306 -6662 121542 -6426
rect 145826 75218 146062 75454
rect 146146 75218 146382 75454
rect 145826 74898 146062 75134
rect 146146 74898 146382 75134
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 149546 78938 149782 79174
rect 149866 78938 150102 79174
rect 149546 78618 149782 78854
rect 149866 78618 150102 78854
rect 149546 42938 149782 43174
rect 149866 42938 150102 43174
rect 149546 42618 149782 42854
rect 149866 42618 150102 42854
rect 149546 6938 149782 7174
rect 149866 6938 150102 7174
rect 149546 6618 149782 6854
rect 149866 6618 150102 6854
rect 149546 -2502 149782 -2266
rect 149866 -2502 150102 -2266
rect 149546 -2822 149782 -2586
rect 149866 -2822 150102 -2586
rect 153266 82658 153502 82894
rect 153586 82658 153822 82894
rect 153266 82338 153502 82574
rect 153586 82338 153822 82574
rect 153266 46658 153502 46894
rect 153586 46658 153822 46894
rect 153266 46338 153502 46574
rect 153586 46338 153822 46574
rect 153266 10658 153502 10894
rect 153586 10658 153822 10894
rect 153266 10338 153502 10574
rect 153586 10338 153822 10574
rect 153266 -4422 153502 -4186
rect 153586 -4422 153822 -4186
rect 153266 -4742 153502 -4506
rect 153586 -4742 153822 -4506
rect 156986 86378 157222 86614
rect 157306 86378 157542 86614
rect 156986 86058 157222 86294
rect 157306 86058 157542 86294
rect 156986 50378 157222 50614
rect 157306 50378 157542 50614
rect 156986 50058 157222 50294
rect 157306 50058 157542 50294
rect 156986 14378 157222 14614
rect 157306 14378 157542 14614
rect 156986 14058 157222 14294
rect 157306 14058 157542 14294
rect 138986 -7302 139222 -7066
rect 139306 -7302 139542 -7066
rect 138986 -7622 139222 -7386
rect 139306 -7622 139542 -7386
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 167546 312938 167782 313174
rect 167866 312938 168102 313174
rect 167546 312618 167782 312854
rect 167866 312618 168102 312854
rect 167546 276938 167782 277174
rect 167866 276938 168102 277174
rect 167546 276618 167782 276854
rect 167866 276618 168102 276854
rect 167546 240938 167782 241174
rect 167866 240938 168102 241174
rect 167546 240618 167782 240854
rect 167866 240618 168102 240854
rect 171266 532658 171502 532894
rect 171586 532658 171822 532894
rect 171266 532338 171502 532574
rect 171586 532338 171822 532574
rect 171266 496658 171502 496894
rect 171586 496658 171822 496894
rect 171266 496338 171502 496574
rect 171586 496338 171822 496574
rect 171266 460658 171502 460894
rect 171586 460658 171822 460894
rect 171266 460338 171502 460574
rect 171586 460338 171822 460574
rect 171266 424658 171502 424894
rect 171586 424658 171822 424894
rect 171266 424338 171502 424574
rect 171586 424338 171822 424574
rect 171266 388658 171502 388894
rect 171586 388658 171822 388894
rect 171266 388338 171502 388574
rect 171586 388338 171822 388574
rect 171266 352658 171502 352894
rect 171586 352658 171822 352894
rect 171266 352338 171502 352574
rect 171586 352338 171822 352574
rect 192986 710362 193222 710598
rect 193306 710362 193542 710598
rect 192986 710042 193222 710278
rect 193306 710042 193542 710278
rect 189266 708442 189502 708678
rect 189586 708442 189822 708678
rect 189266 708122 189502 708358
rect 189586 708122 189822 708358
rect 185546 706522 185782 706758
rect 185866 706522 186102 706758
rect 185546 706202 185782 706438
rect 185866 706202 186102 706438
rect 174986 680378 175222 680614
rect 175306 680378 175542 680614
rect 174986 680058 175222 680294
rect 175306 680058 175542 680294
rect 174986 644378 175222 644614
rect 175306 644378 175542 644614
rect 174986 644058 175222 644294
rect 175306 644058 175542 644294
rect 174986 608378 175222 608614
rect 175306 608378 175542 608614
rect 174986 608058 175222 608294
rect 175306 608058 175542 608294
rect 174986 572378 175222 572614
rect 175306 572378 175542 572614
rect 174986 572058 175222 572294
rect 175306 572058 175542 572294
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 174986 536378 175222 536614
rect 175306 536378 175542 536614
rect 174986 536058 175222 536294
rect 175306 536058 175542 536294
rect 174986 500378 175222 500614
rect 175306 500378 175542 500614
rect 174986 500058 175222 500294
rect 175306 500058 175542 500294
rect 174986 464378 175222 464614
rect 175306 464378 175542 464614
rect 174986 464058 175222 464294
rect 175306 464058 175542 464294
rect 174986 428378 175222 428614
rect 175306 428378 175542 428614
rect 174986 428058 175222 428294
rect 175306 428058 175542 428294
rect 174986 392378 175222 392614
rect 175306 392378 175542 392614
rect 174986 392058 175222 392294
rect 175306 392058 175542 392294
rect 174986 356378 175222 356614
rect 175306 356378 175542 356614
rect 174986 356058 175222 356294
rect 175306 356058 175542 356294
rect 174986 320378 175222 320614
rect 175306 320378 175542 320614
rect 174986 320058 175222 320294
rect 175306 320058 175542 320294
rect 171266 316658 171502 316894
rect 171586 316658 171822 316894
rect 171266 316338 171502 316574
rect 171586 316338 171822 316574
rect 171266 280658 171502 280894
rect 171586 280658 171822 280894
rect 171266 280338 171502 280574
rect 171586 280338 171822 280574
rect 171266 244658 171502 244894
rect 171586 244658 171822 244894
rect 171266 244338 171502 244574
rect 171586 244338 171822 244574
rect 167546 204938 167782 205174
rect 167866 204938 168102 205174
rect 167546 204618 167782 204854
rect 167866 204618 168102 204854
rect 167546 168938 167782 169174
rect 167866 168938 168102 169174
rect 167546 168618 167782 168854
rect 167866 168618 168102 168854
rect 167546 132938 167782 133174
rect 167866 132938 168102 133174
rect 167546 132618 167782 132854
rect 167866 132618 168102 132854
rect 167546 96938 167782 97174
rect 167866 96938 168102 97174
rect 167546 96618 167782 96854
rect 167866 96618 168102 96854
rect 167546 60938 167782 61174
rect 167866 60938 168102 61174
rect 167546 60618 167782 60854
rect 167866 60618 168102 60854
rect 171266 208658 171502 208894
rect 171586 208658 171822 208894
rect 171266 208338 171502 208574
rect 171586 208338 171822 208574
rect 171266 172658 171502 172894
rect 171586 172658 171822 172894
rect 171266 172338 171502 172574
rect 171586 172338 171822 172574
rect 171266 136658 171502 136894
rect 171586 136658 171822 136894
rect 171266 136338 171502 136574
rect 171586 136338 171822 136574
rect 171266 100658 171502 100894
rect 171586 100658 171822 100894
rect 171266 100338 171502 100574
rect 171586 100338 171822 100574
rect 171266 64658 171502 64894
rect 171586 64658 171822 64894
rect 171266 64338 171502 64574
rect 171586 64338 171822 64574
rect 171266 28658 171502 28894
rect 171586 28658 171822 28894
rect 171266 28338 171502 28574
rect 171586 28338 171822 28574
rect 167546 24938 167782 25174
rect 167866 24938 168102 25174
rect 167546 24618 167782 24854
rect 167866 24618 168102 24854
rect 163826 -1542 164062 -1306
rect 164146 -1542 164382 -1306
rect 163826 -1862 164062 -1626
rect 164146 -1862 164382 -1626
rect 167546 -3462 167782 -3226
rect 167866 -3462 168102 -3226
rect 167546 -3782 167782 -3546
rect 167866 -3782 168102 -3546
rect 174986 284378 175222 284614
rect 175306 284378 175542 284614
rect 174986 284058 175222 284294
rect 175306 284058 175542 284294
rect 174986 248378 175222 248614
rect 175306 248378 175542 248614
rect 174986 248058 175222 248294
rect 175306 248058 175542 248294
rect 174986 212378 175222 212614
rect 175306 212378 175542 212614
rect 174986 212058 175222 212294
rect 175306 212058 175542 212294
rect 174986 176378 175222 176614
rect 175306 176378 175542 176614
rect 174986 176058 175222 176294
rect 175306 176058 175542 176294
rect 174986 140378 175222 140614
rect 175306 140378 175542 140614
rect 174986 140058 175222 140294
rect 175306 140058 175542 140294
rect 174986 104378 175222 104614
rect 175306 104378 175542 104614
rect 174986 104058 175222 104294
rect 175306 104058 175542 104294
rect 174986 68378 175222 68614
rect 175306 68378 175542 68614
rect 174986 68058 175222 68294
rect 175306 68058 175542 68294
rect 174986 32378 175222 32614
rect 175306 32378 175542 32614
rect 174986 32058 175222 32294
rect 175306 32058 175542 32294
rect 171266 -5382 171502 -5146
rect 171586 -5382 171822 -5146
rect 171266 -5702 171502 -5466
rect 171586 -5702 171822 -5466
rect 156986 -6342 157222 -6106
rect 157306 -6342 157542 -6106
rect 156986 -6662 157222 -6426
rect 157306 -6662 157542 -6426
rect 185546 690938 185782 691174
rect 185866 690938 186102 691174
rect 185546 690618 185782 690854
rect 185866 690618 186102 690854
rect 185546 654938 185782 655174
rect 185866 654938 186102 655174
rect 185546 654618 185782 654854
rect 185866 654618 186102 654854
rect 185546 618938 185782 619174
rect 185866 618938 186102 619174
rect 185546 618618 185782 618854
rect 185866 618618 186102 618854
rect 185546 582938 185782 583174
rect 185866 582938 186102 583174
rect 185546 582618 185782 582854
rect 185866 582618 186102 582854
rect 181826 543218 182062 543454
rect 182146 543218 182382 543454
rect 181826 542898 182062 543134
rect 182146 542898 182382 543134
rect 181826 507218 182062 507454
rect 182146 507218 182382 507454
rect 181826 506898 182062 507134
rect 182146 506898 182382 507134
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 181826 435218 182062 435454
rect 182146 435218 182382 435454
rect 181826 434898 182062 435134
rect 182146 434898 182382 435134
rect 181826 399218 182062 399454
rect 182146 399218 182382 399454
rect 181826 398898 182062 399134
rect 182146 398898 182382 399134
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 181826 327218 182062 327454
rect 182146 327218 182382 327454
rect 181826 326898 182062 327134
rect 182146 326898 182382 327134
rect 181826 291218 182062 291454
rect 182146 291218 182382 291454
rect 181826 290898 182062 291134
rect 182146 290898 182382 291134
rect 181826 255218 182062 255454
rect 182146 255218 182382 255454
rect 181826 254898 182062 255134
rect 182146 254898 182382 255134
rect 181826 219218 182062 219454
rect 182146 219218 182382 219454
rect 181826 218898 182062 219134
rect 182146 218898 182382 219134
rect 181826 183218 182062 183454
rect 182146 183218 182382 183454
rect 181826 182898 182062 183134
rect 182146 182898 182382 183134
rect 181826 147218 182062 147454
rect 182146 147218 182382 147454
rect 181826 146898 182062 147134
rect 182146 146898 182382 147134
rect 181826 111218 182062 111454
rect 182146 111218 182382 111454
rect 181826 110898 182062 111134
rect 182146 110898 182382 111134
rect 181826 75218 182062 75454
rect 182146 75218 182382 75454
rect 181826 74898 182062 75134
rect 182146 74898 182382 75134
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 185546 546938 185782 547174
rect 185866 546938 186102 547174
rect 185546 546618 185782 546854
rect 185866 546618 186102 546854
rect 185546 510938 185782 511174
rect 185866 510938 186102 511174
rect 185546 510618 185782 510854
rect 185866 510618 186102 510854
rect 189266 694658 189502 694894
rect 189586 694658 189822 694894
rect 189266 694338 189502 694574
rect 189586 694338 189822 694574
rect 189266 658658 189502 658894
rect 189586 658658 189822 658894
rect 189266 658338 189502 658574
rect 189586 658338 189822 658574
rect 189266 622658 189502 622894
rect 189586 622658 189822 622894
rect 189266 622338 189502 622574
rect 189586 622338 189822 622574
rect 189266 586658 189502 586894
rect 189586 586658 189822 586894
rect 189266 586338 189502 586574
rect 189586 586338 189822 586574
rect 189266 550658 189502 550894
rect 189586 550658 189822 550894
rect 189266 550338 189502 550574
rect 189586 550338 189822 550574
rect 210986 711322 211222 711558
rect 211306 711322 211542 711558
rect 210986 711002 211222 711238
rect 211306 711002 211542 711238
rect 207266 709402 207502 709638
rect 207586 709402 207822 709638
rect 207266 709082 207502 709318
rect 207586 709082 207822 709318
rect 203546 707482 203782 707718
rect 203866 707482 204102 707718
rect 203546 707162 203782 707398
rect 203866 707162 204102 707398
rect 192986 698378 193222 698614
rect 193306 698378 193542 698614
rect 192986 698058 193222 698294
rect 193306 698058 193542 698294
rect 192986 662378 193222 662614
rect 193306 662378 193542 662614
rect 192986 662058 193222 662294
rect 193306 662058 193542 662294
rect 192986 626378 193222 626614
rect 193306 626378 193542 626614
rect 192986 626058 193222 626294
rect 193306 626058 193542 626294
rect 192986 590378 193222 590614
rect 193306 590378 193542 590614
rect 192986 590058 193222 590294
rect 193306 590058 193542 590294
rect 192986 554378 193222 554614
rect 193306 554378 193542 554614
rect 192986 554058 193222 554294
rect 193306 554058 193542 554294
rect 199826 705562 200062 705798
rect 200146 705562 200382 705798
rect 199826 705242 200062 705478
rect 200146 705242 200382 705478
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 199826 633218 200062 633454
rect 200146 633218 200382 633454
rect 199826 632898 200062 633134
rect 200146 632898 200382 633134
rect 199826 597218 200062 597454
rect 200146 597218 200382 597454
rect 199826 596898 200062 597134
rect 200146 596898 200382 597134
rect 199826 561218 200062 561454
rect 200146 561218 200382 561454
rect 199826 560898 200062 561134
rect 200146 560898 200382 561134
rect 192986 518378 193222 518614
rect 193306 518378 193542 518614
rect 189266 514658 189502 514894
rect 189586 514658 189822 514894
rect 189266 514338 189502 514574
rect 189586 514338 189822 514574
rect 185546 474938 185782 475174
rect 185866 474938 186102 475174
rect 185546 474618 185782 474854
rect 185866 474618 186102 474854
rect 185546 438938 185782 439174
rect 185866 438938 186102 439174
rect 185546 438618 185782 438854
rect 185866 438618 186102 438854
rect 185546 402938 185782 403174
rect 185866 402938 186102 403174
rect 185546 402618 185782 402854
rect 185866 402618 186102 402854
rect 185546 366938 185782 367174
rect 185866 366938 186102 367174
rect 185546 366618 185782 366854
rect 185866 366618 186102 366854
rect 185546 330938 185782 331174
rect 185866 330938 186102 331174
rect 185546 330618 185782 330854
rect 185866 330618 186102 330854
rect 185546 294938 185782 295174
rect 185866 294938 186102 295174
rect 185546 294618 185782 294854
rect 185866 294618 186102 294854
rect 185546 258938 185782 259174
rect 185866 258938 186102 259174
rect 185546 258618 185782 258854
rect 185866 258618 186102 258854
rect 185546 222938 185782 223174
rect 185866 222938 186102 223174
rect 185546 222618 185782 222854
rect 185866 222618 186102 222854
rect 185546 186938 185782 187174
rect 185866 186938 186102 187174
rect 185546 186618 185782 186854
rect 185866 186618 186102 186854
rect 185546 150938 185782 151174
rect 185866 150938 186102 151174
rect 185546 150618 185782 150854
rect 185866 150618 186102 150854
rect 185546 114938 185782 115174
rect 185866 114938 186102 115174
rect 185546 114618 185782 114854
rect 185866 114618 186102 114854
rect 185546 78938 185782 79174
rect 185866 78938 186102 79174
rect 185546 78618 185782 78854
rect 185866 78618 186102 78854
rect 185546 42938 185782 43174
rect 185866 42938 186102 43174
rect 185546 42618 185782 42854
rect 185866 42618 186102 42854
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 189266 478658 189502 478894
rect 189586 478658 189822 478894
rect 189266 478338 189502 478574
rect 189586 478338 189822 478574
rect 189266 442658 189502 442894
rect 189586 442658 189822 442894
rect 189266 442338 189502 442574
rect 189586 442338 189822 442574
rect 189266 406658 189502 406894
rect 189586 406658 189822 406894
rect 189266 406338 189502 406574
rect 189586 406338 189822 406574
rect 189266 370658 189502 370894
rect 189586 370658 189822 370894
rect 189266 370338 189502 370574
rect 189586 370338 189822 370574
rect 189266 334658 189502 334894
rect 189586 334658 189822 334894
rect 189266 334338 189502 334574
rect 189586 334338 189822 334574
rect 189266 298658 189502 298894
rect 189586 298658 189822 298894
rect 189266 298338 189502 298574
rect 189586 298338 189822 298574
rect 189266 262658 189502 262894
rect 189586 262658 189822 262894
rect 189266 262338 189502 262574
rect 189586 262338 189822 262574
rect 189266 226658 189502 226894
rect 189586 226658 189822 226894
rect 189266 226338 189502 226574
rect 189586 226338 189822 226574
rect 189266 190658 189502 190894
rect 189586 190658 189822 190894
rect 189266 190338 189502 190574
rect 189586 190338 189822 190574
rect 189266 154658 189502 154894
rect 189586 154658 189822 154894
rect 189266 154338 189502 154574
rect 189586 154338 189822 154574
rect 189266 118658 189502 118894
rect 189586 118658 189822 118894
rect 189266 118338 189502 118574
rect 189586 118338 189822 118574
rect 192986 518058 193222 518294
rect 193306 518058 193542 518294
rect 192986 482378 193222 482614
rect 193306 482378 193542 482614
rect 192986 482058 193222 482294
rect 193306 482058 193542 482294
rect 192986 446378 193222 446614
rect 193306 446378 193542 446614
rect 192986 446058 193222 446294
rect 193306 446058 193542 446294
rect 192986 410378 193222 410614
rect 193306 410378 193542 410614
rect 192986 410058 193222 410294
rect 193306 410058 193542 410294
rect 192986 374378 193222 374614
rect 193306 374378 193542 374614
rect 192986 374058 193222 374294
rect 193306 374058 193542 374294
rect 192986 338378 193222 338614
rect 193306 338378 193542 338614
rect 192986 338058 193222 338294
rect 193306 338058 193542 338294
rect 192986 302378 193222 302614
rect 193306 302378 193542 302614
rect 192986 302058 193222 302294
rect 193306 302058 193542 302294
rect 192986 266378 193222 266614
rect 193306 266378 193542 266614
rect 192986 266058 193222 266294
rect 193306 266058 193542 266294
rect 203546 672938 203782 673174
rect 203866 672938 204102 673174
rect 203546 672618 203782 672854
rect 203866 672618 204102 672854
rect 203546 636938 203782 637174
rect 203866 636938 204102 637174
rect 203546 636618 203782 636854
rect 203866 636618 204102 636854
rect 203546 600938 203782 601174
rect 203866 600938 204102 601174
rect 203546 600618 203782 600854
rect 203866 600618 204102 600854
rect 203546 564938 203782 565174
rect 203866 564938 204102 565174
rect 203546 564618 203782 564854
rect 203866 564618 204102 564854
rect 207266 676658 207502 676894
rect 207586 676658 207822 676894
rect 207266 676338 207502 676574
rect 207586 676338 207822 676574
rect 207266 640658 207502 640894
rect 207586 640658 207822 640894
rect 207266 640338 207502 640574
rect 207586 640338 207822 640574
rect 207266 604658 207502 604894
rect 207586 604658 207822 604894
rect 207266 604338 207502 604574
rect 207586 604338 207822 604574
rect 207266 568658 207502 568894
rect 207586 568658 207822 568894
rect 207266 568338 207502 568574
rect 207586 568338 207822 568574
rect 228986 710362 229222 710598
rect 229306 710362 229542 710598
rect 228986 710042 229222 710278
rect 229306 710042 229542 710278
rect 225266 708442 225502 708678
rect 225586 708442 225822 708678
rect 225266 708122 225502 708358
rect 225586 708122 225822 708358
rect 221546 706522 221782 706758
rect 221866 706522 222102 706758
rect 221546 706202 221782 706438
rect 221866 706202 222102 706438
rect 210986 680378 211222 680614
rect 211306 680378 211542 680614
rect 210986 680058 211222 680294
rect 211306 680058 211542 680294
rect 210986 644378 211222 644614
rect 211306 644378 211542 644614
rect 210986 644058 211222 644294
rect 211306 644058 211542 644294
rect 210986 608378 211222 608614
rect 211306 608378 211542 608614
rect 210986 608058 211222 608294
rect 211306 608058 211542 608294
rect 210986 572378 211222 572614
rect 211306 572378 211542 572614
rect 210986 572058 211222 572294
rect 211306 572058 211542 572294
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 217826 543218 218062 543454
rect 218146 543218 218382 543454
rect 217826 542898 218062 543134
rect 218146 542898 218382 543134
rect 221546 690938 221782 691174
rect 221866 690938 222102 691174
rect 221546 690618 221782 690854
rect 221866 690618 222102 690854
rect 221546 654938 221782 655174
rect 221866 654938 222102 655174
rect 221546 654618 221782 654854
rect 221866 654618 222102 654854
rect 221546 618938 221782 619174
rect 221866 618938 222102 619174
rect 221546 618618 221782 618854
rect 221866 618618 222102 618854
rect 221546 582938 221782 583174
rect 221866 582938 222102 583174
rect 221546 582618 221782 582854
rect 221866 582618 222102 582854
rect 221546 546938 221782 547174
rect 221866 546938 222102 547174
rect 221546 546618 221782 546854
rect 221866 546618 222102 546854
rect 225266 694658 225502 694894
rect 225586 694658 225822 694894
rect 225266 694338 225502 694574
rect 225586 694338 225822 694574
rect 225266 658658 225502 658894
rect 225586 658658 225822 658894
rect 225266 658338 225502 658574
rect 225586 658338 225822 658574
rect 225266 622658 225502 622894
rect 225586 622658 225822 622894
rect 225266 622338 225502 622574
rect 225586 622338 225822 622574
rect 225266 586658 225502 586894
rect 225586 586658 225822 586894
rect 225266 586338 225502 586574
rect 225586 586338 225822 586574
rect 225266 550658 225502 550894
rect 225586 550658 225822 550894
rect 225266 550338 225502 550574
rect 225586 550338 225822 550574
rect 246986 711322 247222 711558
rect 247306 711322 247542 711558
rect 246986 711002 247222 711238
rect 247306 711002 247542 711238
rect 243266 709402 243502 709638
rect 243586 709402 243822 709638
rect 243266 709082 243502 709318
rect 243586 709082 243822 709318
rect 239546 707482 239782 707718
rect 239866 707482 240102 707718
rect 239546 707162 239782 707398
rect 239866 707162 240102 707398
rect 228986 698378 229222 698614
rect 229306 698378 229542 698614
rect 228986 698058 229222 698294
rect 229306 698058 229542 698294
rect 228986 662378 229222 662614
rect 229306 662378 229542 662614
rect 228986 662058 229222 662294
rect 229306 662058 229542 662294
rect 228986 626378 229222 626614
rect 229306 626378 229542 626614
rect 228986 626058 229222 626294
rect 229306 626058 229542 626294
rect 228986 590378 229222 590614
rect 229306 590378 229542 590614
rect 228986 590058 229222 590294
rect 229306 590058 229542 590294
rect 228986 554378 229222 554614
rect 229306 554378 229542 554614
rect 228986 554058 229222 554294
rect 229306 554058 229542 554294
rect 235826 705562 236062 705798
rect 236146 705562 236382 705798
rect 235826 705242 236062 705478
rect 236146 705242 236382 705478
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 235826 633218 236062 633454
rect 236146 633218 236382 633454
rect 235826 632898 236062 633134
rect 236146 632898 236382 633134
rect 235826 597218 236062 597454
rect 236146 597218 236382 597454
rect 235826 596898 236062 597134
rect 236146 596898 236382 597134
rect 235826 561218 236062 561454
rect 236146 561218 236382 561454
rect 235826 560898 236062 561134
rect 236146 560898 236382 561134
rect 239546 672938 239782 673174
rect 239866 672938 240102 673174
rect 239546 672618 239782 672854
rect 239866 672618 240102 672854
rect 239546 636938 239782 637174
rect 239866 636938 240102 637174
rect 239546 636618 239782 636854
rect 239866 636618 240102 636854
rect 239546 600938 239782 601174
rect 239866 600938 240102 601174
rect 239546 600618 239782 600854
rect 239866 600618 240102 600854
rect 239546 564938 239782 565174
rect 239866 564938 240102 565174
rect 239546 564618 239782 564854
rect 239866 564618 240102 564854
rect 243266 676658 243502 676894
rect 243586 676658 243822 676894
rect 243266 676338 243502 676574
rect 243586 676338 243822 676574
rect 243266 640658 243502 640894
rect 243586 640658 243822 640894
rect 243266 640338 243502 640574
rect 243586 640338 243822 640574
rect 243266 604658 243502 604894
rect 243586 604658 243822 604894
rect 243266 604338 243502 604574
rect 243586 604338 243822 604574
rect 243266 568658 243502 568894
rect 243586 568658 243822 568894
rect 243266 568338 243502 568574
rect 243586 568338 243822 568574
rect 264986 710362 265222 710598
rect 265306 710362 265542 710598
rect 264986 710042 265222 710278
rect 265306 710042 265542 710278
rect 261266 708442 261502 708678
rect 261586 708442 261822 708678
rect 261266 708122 261502 708358
rect 261586 708122 261822 708358
rect 257546 706522 257782 706758
rect 257866 706522 258102 706758
rect 257546 706202 257782 706438
rect 257866 706202 258102 706438
rect 246986 680378 247222 680614
rect 247306 680378 247542 680614
rect 246986 680058 247222 680294
rect 247306 680058 247542 680294
rect 246986 644378 247222 644614
rect 247306 644378 247542 644614
rect 246986 644058 247222 644294
rect 247306 644058 247542 644294
rect 246986 608378 247222 608614
rect 247306 608378 247542 608614
rect 246986 608058 247222 608294
rect 247306 608058 247542 608294
rect 246986 572378 247222 572614
rect 247306 572378 247542 572614
rect 246986 572058 247222 572294
rect 247306 572058 247542 572294
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 253826 615218 254062 615454
rect 254146 615218 254382 615454
rect 253826 614898 254062 615134
rect 254146 614898 254382 615134
rect 253826 579218 254062 579454
rect 254146 579218 254382 579454
rect 253826 578898 254062 579134
rect 254146 578898 254382 579134
rect 253826 543218 254062 543454
rect 254146 543218 254382 543454
rect 253826 542898 254062 543134
rect 254146 542898 254382 543134
rect 257546 690938 257782 691174
rect 257866 690938 258102 691174
rect 257546 690618 257782 690854
rect 257866 690618 258102 690854
rect 257546 654938 257782 655174
rect 257866 654938 258102 655174
rect 257546 654618 257782 654854
rect 257866 654618 258102 654854
rect 257546 618938 257782 619174
rect 257866 618938 258102 619174
rect 257546 618618 257782 618854
rect 257866 618618 258102 618854
rect 257546 582938 257782 583174
rect 257866 582938 258102 583174
rect 257546 582618 257782 582854
rect 257866 582618 258102 582854
rect 257546 546938 257782 547174
rect 257866 546938 258102 547174
rect 257546 546618 257782 546854
rect 257866 546618 258102 546854
rect 261266 694658 261502 694894
rect 261586 694658 261822 694894
rect 261266 694338 261502 694574
rect 261586 694338 261822 694574
rect 261266 658658 261502 658894
rect 261586 658658 261822 658894
rect 261266 658338 261502 658574
rect 261586 658338 261822 658574
rect 261266 622658 261502 622894
rect 261586 622658 261822 622894
rect 261266 622338 261502 622574
rect 261586 622338 261822 622574
rect 261266 586658 261502 586894
rect 261586 586658 261822 586894
rect 261266 586338 261502 586574
rect 261586 586338 261822 586574
rect 261266 550658 261502 550894
rect 261586 550658 261822 550894
rect 261266 550338 261502 550574
rect 261586 550338 261822 550574
rect 282986 711322 283222 711558
rect 283306 711322 283542 711558
rect 282986 711002 283222 711238
rect 283306 711002 283542 711238
rect 279266 709402 279502 709638
rect 279586 709402 279822 709638
rect 279266 709082 279502 709318
rect 279586 709082 279822 709318
rect 275546 707482 275782 707718
rect 275866 707482 276102 707718
rect 275546 707162 275782 707398
rect 275866 707162 276102 707398
rect 264986 698378 265222 698614
rect 265306 698378 265542 698614
rect 264986 698058 265222 698294
rect 265306 698058 265542 698294
rect 264986 662378 265222 662614
rect 265306 662378 265542 662614
rect 264986 662058 265222 662294
rect 265306 662058 265542 662294
rect 264986 626378 265222 626614
rect 265306 626378 265542 626614
rect 264986 626058 265222 626294
rect 265306 626058 265542 626294
rect 264986 590378 265222 590614
rect 265306 590378 265542 590614
rect 264986 590058 265222 590294
rect 265306 590058 265542 590294
rect 264986 554378 265222 554614
rect 265306 554378 265542 554614
rect 264986 554058 265222 554294
rect 265306 554058 265542 554294
rect 271826 705562 272062 705798
rect 272146 705562 272382 705798
rect 271826 705242 272062 705478
rect 272146 705242 272382 705478
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 271826 633218 272062 633454
rect 272146 633218 272382 633454
rect 271826 632898 272062 633134
rect 272146 632898 272382 633134
rect 271826 597218 272062 597454
rect 272146 597218 272382 597454
rect 271826 596898 272062 597134
rect 272146 596898 272382 597134
rect 271826 561218 272062 561454
rect 272146 561218 272382 561454
rect 271826 560898 272062 561134
rect 272146 560898 272382 561134
rect 275546 672938 275782 673174
rect 275866 672938 276102 673174
rect 275546 672618 275782 672854
rect 275866 672618 276102 672854
rect 275546 636938 275782 637174
rect 275866 636938 276102 637174
rect 275546 636618 275782 636854
rect 275866 636618 276102 636854
rect 275546 600938 275782 601174
rect 275866 600938 276102 601174
rect 275546 600618 275782 600854
rect 275866 600618 276102 600854
rect 275546 564938 275782 565174
rect 275866 564938 276102 565174
rect 275546 564618 275782 564854
rect 275866 564618 276102 564854
rect 279266 676658 279502 676894
rect 279586 676658 279822 676894
rect 279266 676338 279502 676574
rect 279586 676338 279822 676574
rect 279266 640658 279502 640894
rect 279586 640658 279822 640894
rect 279266 640338 279502 640574
rect 279586 640338 279822 640574
rect 279266 604658 279502 604894
rect 279586 604658 279822 604894
rect 279266 604338 279502 604574
rect 279586 604338 279822 604574
rect 279266 568658 279502 568894
rect 279586 568658 279822 568894
rect 279266 568338 279502 568574
rect 279586 568338 279822 568574
rect 300986 710362 301222 710598
rect 301306 710362 301542 710598
rect 300986 710042 301222 710278
rect 301306 710042 301542 710278
rect 297266 708442 297502 708678
rect 297586 708442 297822 708678
rect 297266 708122 297502 708358
rect 297586 708122 297822 708358
rect 293546 706522 293782 706758
rect 293866 706522 294102 706758
rect 293546 706202 293782 706438
rect 293866 706202 294102 706438
rect 282986 680378 283222 680614
rect 283306 680378 283542 680614
rect 282986 680058 283222 680294
rect 283306 680058 283542 680294
rect 282986 644378 283222 644614
rect 283306 644378 283542 644614
rect 282986 644058 283222 644294
rect 283306 644058 283542 644294
rect 282986 608378 283222 608614
rect 283306 608378 283542 608614
rect 282986 608058 283222 608294
rect 283306 608058 283542 608294
rect 282986 572378 283222 572614
rect 283306 572378 283542 572614
rect 282986 572058 283222 572294
rect 283306 572058 283542 572294
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 289826 543218 290062 543454
rect 290146 543218 290382 543454
rect 289826 542898 290062 543134
rect 290146 542898 290382 543134
rect 293546 690938 293782 691174
rect 293866 690938 294102 691174
rect 293546 690618 293782 690854
rect 293866 690618 294102 690854
rect 293546 654938 293782 655174
rect 293866 654938 294102 655174
rect 293546 654618 293782 654854
rect 293866 654618 294102 654854
rect 293546 618938 293782 619174
rect 293866 618938 294102 619174
rect 293546 618618 293782 618854
rect 293866 618618 294102 618854
rect 293546 582938 293782 583174
rect 293866 582938 294102 583174
rect 293546 582618 293782 582854
rect 293866 582618 294102 582854
rect 293546 546938 293782 547174
rect 293866 546938 294102 547174
rect 293546 546618 293782 546854
rect 293866 546618 294102 546854
rect 297266 694658 297502 694894
rect 297586 694658 297822 694894
rect 297266 694338 297502 694574
rect 297586 694338 297822 694574
rect 297266 658658 297502 658894
rect 297586 658658 297822 658894
rect 297266 658338 297502 658574
rect 297586 658338 297822 658574
rect 297266 622658 297502 622894
rect 297586 622658 297822 622894
rect 297266 622338 297502 622574
rect 297586 622338 297822 622574
rect 297266 586658 297502 586894
rect 297586 586658 297822 586894
rect 297266 586338 297502 586574
rect 297586 586338 297822 586574
rect 297266 550658 297502 550894
rect 297586 550658 297822 550894
rect 297266 550338 297502 550574
rect 297586 550338 297822 550574
rect 318986 711322 319222 711558
rect 319306 711322 319542 711558
rect 318986 711002 319222 711238
rect 319306 711002 319542 711238
rect 315266 709402 315502 709638
rect 315586 709402 315822 709638
rect 315266 709082 315502 709318
rect 315586 709082 315822 709318
rect 311546 707482 311782 707718
rect 311866 707482 312102 707718
rect 311546 707162 311782 707398
rect 311866 707162 312102 707398
rect 300986 698378 301222 698614
rect 301306 698378 301542 698614
rect 300986 698058 301222 698294
rect 301306 698058 301542 698294
rect 300986 662378 301222 662614
rect 301306 662378 301542 662614
rect 300986 662058 301222 662294
rect 301306 662058 301542 662294
rect 300986 626378 301222 626614
rect 301306 626378 301542 626614
rect 300986 626058 301222 626294
rect 301306 626058 301542 626294
rect 300986 590378 301222 590614
rect 301306 590378 301542 590614
rect 300986 590058 301222 590294
rect 301306 590058 301542 590294
rect 300986 554378 301222 554614
rect 301306 554378 301542 554614
rect 300986 554058 301222 554294
rect 301306 554058 301542 554294
rect 307826 705562 308062 705798
rect 308146 705562 308382 705798
rect 307826 705242 308062 705478
rect 308146 705242 308382 705478
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 307826 561218 308062 561454
rect 308146 561218 308382 561454
rect 307826 560898 308062 561134
rect 308146 560898 308382 561134
rect 311546 672938 311782 673174
rect 311866 672938 312102 673174
rect 311546 672618 311782 672854
rect 311866 672618 312102 672854
rect 311546 636938 311782 637174
rect 311866 636938 312102 637174
rect 311546 636618 311782 636854
rect 311866 636618 312102 636854
rect 311546 600938 311782 601174
rect 311866 600938 312102 601174
rect 311546 600618 311782 600854
rect 311866 600618 312102 600854
rect 311546 564938 311782 565174
rect 311866 564938 312102 565174
rect 311546 564618 311782 564854
rect 311866 564618 312102 564854
rect 315266 676658 315502 676894
rect 315586 676658 315822 676894
rect 315266 676338 315502 676574
rect 315586 676338 315822 676574
rect 315266 640658 315502 640894
rect 315586 640658 315822 640894
rect 315266 640338 315502 640574
rect 315586 640338 315822 640574
rect 315266 604658 315502 604894
rect 315586 604658 315822 604894
rect 315266 604338 315502 604574
rect 315586 604338 315822 604574
rect 315266 568658 315502 568894
rect 315586 568658 315822 568894
rect 315266 568338 315502 568574
rect 315586 568338 315822 568574
rect 336986 710362 337222 710598
rect 337306 710362 337542 710598
rect 336986 710042 337222 710278
rect 337306 710042 337542 710278
rect 333266 708442 333502 708678
rect 333586 708442 333822 708678
rect 333266 708122 333502 708358
rect 333586 708122 333822 708358
rect 329546 706522 329782 706758
rect 329866 706522 330102 706758
rect 329546 706202 329782 706438
rect 329866 706202 330102 706438
rect 318986 680378 319222 680614
rect 319306 680378 319542 680614
rect 318986 680058 319222 680294
rect 319306 680058 319542 680294
rect 318986 644378 319222 644614
rect 319306 644378 319542 644614
rect 318986 644058 319222 644294
rect 319306 644058 319542 644294
rect 318986 608378 319222 608614
rect 319306 608378 319542 608614
rect 318986 608058 319222 608294
rect 319306 608058 319542 608294
rect 318986 572378 319222 572614
rect 319306 572378 319542 572614
rect 318986 572058 319222 572294
rect 319306 572058 319542 572294
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 325826 543218 326062 543454
rect 326146 543218 326382 543454
rect 325826 542898 326062 543134
rect 326146 542898 326382 543134
rect 329546 690938 329782 691174
rect 329866 690938 330102 691174
rect 329546 690618 329782 690854
rect 329866 690618 330102 690854
rect 329546 654938 329782 655174
rect 329866 654938 330102 655174
rect 329546 654618 329782 654854
rect 329866 654618 330102 654854
rect 329546 618938 329782 619174
rect 329866 618938 330102 619174
rect 329546 618618 329782 618854
rect 329866 618618 330102 618854
rect 329546 582938 329782 583174
rect 329866 582938 330102 583174
rect 329546 582618 329782 582854
rect 329866 582618 330102 582854
rect 329546 546938 329782 547174
rect 329866 546938 330102 547174
rect 329546 546618 329782 546854
rect 329866 546618 330102 546854
rect 333266 694658 333502 694894
rect 333586 694658 333822 694894
rect 333266 694338 333502 694574
rect 333586 694338 333822 694574
rect 333266 658658 333502 658894
rect 333586 658658 333822 658894
rect 333266 658338 333502 658574
rect 333586 658338 333822 658574
rect 333266 622658 333502 622894
rect 333586 622658 333822 622894
rect 333266 622338 333502 622574
rect 333586 622338 333822 622574
rect 333266 586658 333502 586894
rect 333586 586658 333822 586894
rect 333266 586338 333502 586574
rect 333586 586338 333822 586574
rect 333266 550658 333502 550894
rect 333586 550658 333822 550894
rect 333266 550338 333502 550574
rect 333586 550338 333822 550574
rect 354986 711322 355222 711558
rect 355306 711322 355542 711558
rect 354986 711002 355222 711238
rect 355306 711002 355542 711238
rect 351266 709402 351502 709638
rect 351586 709402 351822 709638
rect 351266 709082 351502 709318
rect 351586 709082 351822 709318
rect 347546 707482 347782 707718
rect 347866 707482 348102 707718
rect 347546 707162 347782 707398
rect 347866 707162 348102 707398
rect 336986 698378 337222 698614
rect 337306 698378 337542 698614
rect 336986 698058 337222 698294
rect 337306 698058 337542 698294
rect 336986 662378 337222 662614
rect 337306 662378 337542 662614
rect 336986 662058 337222 662294
rect 337306 662058 337542 662294
rect 336986 626378 337222 626614
rect 337306 626378 337542 626614
rect 336986 626058 337222 626294
rect 337306 626058 337542 626294
rect 336986 590378 337222 590614
rect 337306 590378 337542 590614
rect 336986 590058 337222 590294
rect 337306 590058 337542 590294
rect 336986 554378 337222 554614
rect 337306 554378 337542 554614
rect 336986 554058 337222 554294
rect 337306 554058 337542 554294
rect 343826 705562 344062 705798
rect 344146 705562 344382 705798
rect 343826 705242 344062 705478
rect 344146 705242 344382 705478
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 343826 633218 344062 633454
rect 344146 633218 344382 633454
rect 343826 632898 344062 633134
rect 344146 632898 344382 633134
rect 343826 597218 344062 597454
rect 344146 597218 344382 597454
rect 343826 596898 344062 597134
rect 344146 596898 344382 597134
rect 343826 561218 344062 561454
rect 344146 561218 344382 561454
rect 343826 560898 344062 561134
rect 344146 560898 344382 561134
rect 347546 672938 347782 673174
rect 347866 672938 348102 673174
rect 347546 672618 347782 672854
rect 347866 672618 348102 672854
rect 347546 636938 347782 637174
rect 347866 636938 348102 637174
rect 347546 636618 347782 636854
rect 347866 636618 348102 636854
rect 347546 600938 347782 601174
rect 347866 600938 348102 601174
rect 347546 600618 347782 600854
rect 347866 600618 348102 600854
rect 347546 564938 347782 565174
rect 347866 564938 348102 565174
rect 347546 564618 347782 564854
rect 347866 564618 348102 564854
rect 351266 676658 351502 676894
rect 351586 676658 351822 676894
rect 351266 676338 351502 676574
rect 351586 676338 351822 676574
rect 351266 640658 351502 640894
rect 351586 640658 351822 640894
rect 351266 640338 351502 640574
rect 351586 640338 351822 640574
rect 351266 604658 351502 604894
rect 351586 604658 351822 604894
rect 351266 604338 351502 604574
rect 351586 604338 351822 604574
rect 351266 568658 351502 568894
rect 351586 568658 351822 568894
rect 351266 568338 351502 568574
rect 351586 568338 351822 568574
rect 372986 710362 373222 710598
rect 373306 710362 373542 710598
rect 372986 710042 373222 710278
rect 373306 710042 373542 710278
rect 369266 708442 369502 708678
rect 369586 708442 369822 708678
rect 369266 708122 369502 708358
rect 369586 708122 369822 708358
rect 365546 706522 365782 706758
rect 365866 706522 366102 706758
rect 365546 706202 365782 706438
rect 365866 706202 366102 706438
rect 354986 680378 355222 680614
rect 355306 680378 355542 680614
rect 354986 680058 355222 680294
rect 355306 680058 355542 680294
rect 354986 644378 355222 644614
rect 355306 644378 355542 644614
rect 354986 644058 355222 644294
rect 355306 644058 355542 644294
rect 354986 608378 355222 608614
rect 355306 608378 355542 608614
rect 354986 608058 355222 608294
rect 355306 608058 355542 608294
rect 354986 572378 355222 572614
rect 355306 572378 355542 572614
rect 354986 572058 355222 572294
rect 355306 572058 355542 572294
rect 219610 525218 219846 525454
rect 219610 524898 219846 525134
rect 250330 525218 250566 525454
rect 250330 524898 250566 525134
rect 281050 525218 281286 525454
rect 281050 524898 281286 525134
rect 311770 525218 312006 525454
rect 311770 524898 312006 525134
rect 342490 525218 342726 525454
rect 342490 524898 342726 525134
rect 204250 507218 204486 507454
rect 204250 506898 204486 507134
rect 234970 507218 235206 507454
rect 234970 506898 235206 507134
rect 265690 507218 265926 507454
rect 265690 506898 265926 507134
rect 296410 507218 296646 507454
rect 296410 506898 296646 507134
rect 327130 507218 327366 507454
rect 327130 506898 327366 507134
rect 219610 489218 219846 489454
rect 219610 488898 219846 489134
rect 250330 489218 250566 489454
rect 250330 488898 250566 489134
rect 281050 489218 281286 489454
rect 281050 488898 281286 489134
rect 311770 489218 312006 489454
rect 311770 488898 312006 489134
rect 342490 489218 342726 489454
rect 342490 488898 342726 489134
rect 204250 471218 204486 471454
rect 204250 470898 204486 471134
rect 234970 471218 235206 471454
rect 234970 470898 235206 471134
rect 265690 471218 265926 471454
rect 265690 470898 265926 471134
rect 296410 471218 296646 471454
rect 296410 470898 296646 471134
rect 327130 471218 327366 471454
rect 327130 470898 327366 471134
rect 192986 230378 193222 230614
rect 193306 230378 193542 230614
rect 192986 230058 193222 230294
rect 193306 230058 193542 230294
rect 219610 453218 219846 453454
rect 219610 452898 219846 453134
rect 250330 453218 250566 453454
rect 250330 452898 250566 453134
rect 281050 453218 281286 453454
rect 281050 452898 281286 453134
rect 311770 453218 312006 453454
rect 311770 452898 312006 453134
rect 342490 453218 342726 453454
rect 342490 452898 342726 453134
rect 204250 435218 204486 435454
rect 204250 434898 204486 435134
rect 234970 435218 235206 435454
rect 234970 434898 235206 435134
rect 265690 435218 265926 435454
rect 265690 434898 265926 435134
rect 296410 435218 296646 435454
rect 296410 434898 296646 435134
rect 327130 435218 327366 435454
rect 327130 434898 327366 435134
rect 219610 417218 219846 417454
rect 219610 416898 219846 417134
rect 250330 417218 250566 417454
rect 250330 416898 250566 417134
rect 281050 417218 281286 417454
rect 281050 416898 281286 417134
rect 311770 417218 312006 417454
rect 311770 416898 312006 417134
rect 342490 417218 342726 417454
rect 342490 416898 342726 417134
rect 204250 399218 204486 399454
rect 204250 398898 204486 399134
rect 234970 399218 235206 399454
rect 234970 398898 235206 399134
rect 265690 399218 265926 399454
rect 265690 398898 265926 399134
rect 296410 399218 296646 399454
rect 296410 398898 296646 399134
rect 327130 399218 327366 399454
rect 327130 398898 327366 399134
rect 219610 381218 219846 381454
rect 219610 380898 219846 381134
rect 250330 381218 250566 381454
rect 250330 380898 250566 381134
rect 281050 381218 281286 381454
rect 281050 380898 281286 381134
rect 311770 381218 312006 381454
rect 311770 380898 312006 381134
rect 342490 381218 342726 381454
rect 342490 380898 342726 381134
rect 199826 345218 200062 345454
rect 200146 345218 200382 345454
rect 199826 344898 200062 345134
rect 200146 344898 200382 345134
rect 199826 309218 200062 309454
rect 200146 309218 200382 309454
rect 199826 308898 200062 309134
rect 200146 308898 200382 309134
rect 203546 348938 203782 349174
rect 203866 348938 204102 349174
rect 203546 348618 203782 348854
rect 203866 348618 204102 348854
rect 207266 352658 207502 352894
rect 207586 352658 207822 352894
rect 207266 352338 207502 352574
rect 207586 352338 207822 352574
rect 210986 356378 211222 356614
rect 211306 356378 211542 356614
rect 210986 356058 211222 356294
rect 211306 356058 211542 356294
rect 207266 316658 207502 316894
rect 207586 316658 207822 316894
rect 207266 316338 207502 316574
rect 207586 316338 207822 316574
rect 203546 312938 203782 313174
rect 203866 312938 204102 313174
rect 203546 312618 203782 312854
rect 203866 312618 204102 312854
rect 204450 255218 204686 255454
rect 204450 254898 204686 255134
rect 217826 363218 218062 363454
rect 218146 363218 218382 363454
rect 217826 362898 218062 363134
rect 218146 362898 218382 363134
rect 210986 320378 211222 320614
rect 211306 320378 211542 320614
rect 210986 320058 211222 320294
rect 211306 320058 211542 320294
rect 199826 237218 200062 237454
rect 200146 237218 200382 237454
rect 199826 236898 200062 237134
rect 200146 236898 200382 237134
rect 192986 194378 193222 194614
rect 193306 194378 193542 194614
rect 192986 194058 193222 194294
rect 193306 194058 193542 194294
rect 199826 201218 200062 201454
rect 200146 201218 200382 201454
rect 199826 200898 200062 201134
rect 200146 200898 200382 201134
rect 192986 158378 193222 158614
rect 193306 158378 193542 158614
rect 192986 158058 193222 158294
rect 193306 158058 193542 158294
rect 192986 122378 193222 122614
rect 193306 122378 193542 122614
rect 192986 122058 193222 122294
rect 193306 122058 193542 122294
rect 199826 165218 200062 165454
rect 200146 165218 200382 165454
rect 199826 164898 200062 165134
rect 200146 164898 200382 165134
rect 199826 129218 200062 129454
rect 200146 129218 200382 129454
rect 199826 128898 200062 129134
rect 200146 128898 200382 129134
rect 192986 86378 193222 86614
rect 193306 86378 193542 86614
rect 192986 86058 193222 86294
rect 193306 86058 193542 86294
rect 189266 82658 189502 82894
rect 189586 82658 189822 82894
rect 189266 82338 189502 82574
rect 189586 82338 189822 82574
rect 189266 46658 189502 46894
rect 189586 46658 189822 46894
rect 189266 46338 189502 46574
rect 189586 46338 189822 46574
rect 185546 6938 185782 7174
rect 185866 6938 186102 7174
rect 185546 6618 185782 6854
rect 185866 6618 186102 6854
rect 185546 -2502 185782 -2266
rect 185866 -2502 186102 -2266
rect 185546 -2822 185782 -2586
rect 185866 -2822 186102 -2586
rect 189266 10658 189502 10894
rect 189586 10658 189822 10894
rect 189266 10338 189502 10574
rect 189586 10338 189822 10574
rect 189266 -4422 189502 -4186
rect 189586 -4422 189822 -4186
rect 189266 -4742 189502 -4506
rect 189586 -4742 189822 -4506
rect 192986 50378 193222 50614
rect 193306 50378 193542 50614
rect 192986 50058 193222 50294
rect 193306 50058 193542 50294
rect 192986 14378 193222 14614
rect 193306 14378 193542 14614
rect 192986 14058 193222 14294
rect 193306 14058 193542 14294
rect 174986 -7302 175222 -7066
rect 175306 -7302 175542 -7066
rect 174986 -7622 175222 -7386
rect 175306 -7622 175542 -7386
rect 199826 93218 200062 93454
rect 200146 93218 200382 93454
rect 199826 92898 200062 93134
rect 200146 92898 200382 93134
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -1542 200062 -1306
rect 200146 -1542 200382 -1306
rect 199826 -1862 200062 -1626
rect 200146 -1862 200382 -1626
rect 203546 204938 203782 205174
rect 203866 204938 204102 205174
rect 203546 204618 203782 204854
rect 203866 204618 204102 204854
rect 207266 208658 207502 208894
rect 207586 208658 207822 208894
rect 207266 208338 207502 208574
rect 207586 208338 207822 208574
rect 203546 168938 203782 169174
rect 203866 168938 204102 169174
rect 203546 168618 203782 168854
rect 203866 168618 204102 168854
rect 203546 132938 203782 133174
rect 203866 132938 204102 133174
rect 203546 132618 203782 132854
rect 203866 132618 204102 132854
rect 203546 96938 203782 97174
rect 203866 96938 204102 97174
rect 203546 96618 203782 96854
rect 203866 96618 204102 96854
rect 203546 60938 203782 61174
rect 203866 60938 204102 61174
rect 203546 60618 203782 60854
rect 203866 60618 204102 60854
rect 203546 24938 203782 25174
rect 203866 24938 204102 25174
rect 203546 24618 203782 24854
rect 203866 24618 204102 24854
rect 203546 -3462 203782 -3226
rect 203866 -3462 204102 -3226
rect 203546 -3782 203782 -3546
rect 203866 -3782 204102 -3546
rect 207266 172658 207502 172894
rect 207586 172658 207822 172894
rect 207266 172338 207502 172574
rect 207586 172338 207822 172574
rect 207266 136658 207502 136894
rect 207586 136658 207822 136894
rect 207266 136338 207502 136574
rect 207586 136338 207822 136574
rect 207266 100658 207502 100894
rect 207586 100658 207822 100894
rect 207266 100338 207502 100574
rect 207586 100338 207822 100574
rect 207266 64658 207502 64894
rect 207586 64658 207822 64894
rect 207266 64338 207502 64574
rect 207586 64338 207822 64574
rect 207266 28658 207502 28894
rect 207586 28658 207822 28894
rect 207266 28338 207502 28574
rect 207586 28338 207822 28574
rect 207266 -5382 207502 -5146
rect 207586 -5382 207822 -5146
rect 207266 -5702 207502 -5466
rect 207586 -5702 207822 -5466
rect 221546 366938 221782 367174
rect 221866 366938 222102 367174
rect 221546 366618 221782 366854
rect 221866 366618 222102 366854
rect 217826 327218 218062 327454
rect 218146 327218 218382 327454
rect 217826 326898 218062 327134
rect 218146 326898 218382 327134
rect 210986 212378 211222 212614
rect 211306 212378 211542 212614
rect 210986 212058 211222 212294
rect 211306 212058 211542 212294
rect 217826 291218 218062 291454
rect 218146 291218 218382 291454
rect 217826 290898 218062 291134
rect 218146 290898 218382 291134
rect 221546 330938 221782 331174
rect 221866 330938 222102 331174
rect 221546 330618 221782 330854
rect 221866 330618 222102 330854
rect 219810 273218 220046 273454
rect 219810 272898 220046 273134
rect 221546 294938 221782 295174
rect 221866 294938 222102 295174
rect 221546 294618 221782 294854
rect 221866 294618 222102 294854
rect 225266 370658 225502 370894
rect 225586 370658 225822 370894
rect 225266 370338 225502 370574
rect 225586 370338 225822 370574
rect 225266 334658 225502 334894
rect 225586 334658 225822 334894
rect 225266 334338 225502 334574
rect 225586 334338 225822 334574
rect 228986 374378 229222 374614
rect 229306 374378 229542 374614
rect 228986 374058 229222 374294
rect 229306 374058 229542 374294
rect 235826 345218 236062 345454
rect 236146 345218 236382 345454
rect 235826 344898 236062 345134
rect 236146 344898 236382 345134
rect 228986 338378 229222 338614
rect 229306 338378 229542 338614
rect 228986 338058 229222 338294
rect 229306 338058 229542 338294
rect 225266 298658 225502 298894
rect 225586 298658 225822 298894
rect 225266 298338 225502 298574
rect 225586 298338 225822 298574
rect 217826 219218 218062 219454
rect 218146 219218 218382 219454
rect 217826 218898 218062 219134
rect 218146 218898 218382 219134
rect 217826 183218 218062 183454
rect 218146 183218 218382 183454
rect 217826 182898 218062 183134
rect 218146 182898 218382 183134
rect 228986 302378 229222 302614
rect 229306 302378 229542 302614
rect 228986 302058 229222 302294
rect 229306 302058 229542 302294
rect 221546 222938 221782 223174
rect 221866 222938 222102 223174
rect 221546 222618 221782 222854
rect 221866 222618 222102 222854
rect 221546 186938 221782 187174
rect 221866 186938 222102 187174
rect 221546 186618 221782 186854
rect 221866 186618 222102 186854
rect 210986 176378 211222 176614
rect 211306 176378 211542 176614
rect 210986 176058 211222 176294
rect 211306 176058 211542 176294
rect 225266 226658 225502 226894
rect 225586 226658 225822 226894
rect 225266 226338 225502 226574
rect 225586 226338 225822 226574
rect 225266 190658 225502 190894
rect 225586 190658 225822 190894
rect 225266 190338 225502 190574
rect 225586 190338 225822 190574
rect 228986 230378 229222 230614
rect 229306 230378 229542 230614
rect 228986 230058 229222 230294
rect 229306 230058 229542 230294
rect 228986 194378 229222 194614
rect 229306 194378 229542 194614
rect 228986 194058 229222 194294
rect 229306 194058 229542 194294
rect 221249 165218 221485 165454
rect 221249 164898 221485 165134
rect 224513 165218 224749 165454
rect 224513 164898 224749 165134
rect 210986 140378 211222 140614
rect 211306 140378 211542 140614
rect 210986 140058 211222 140294
rect 211306 140058 211542 140294
rect 210986 104378 211222 104614
rect 211306 104378 211542 104614
rect 210986 104058 211222 104294
rect 211306 104058 211542 104294
rect 219617 147218 219853 147454
rect 219617 146898 219853 147134
rect 222881 147218 223117 147454
rect 222881 146898 223117 147134
rect 226145 147218 226381 147454
rect 226145 146898 226381 147134
rect 239546 348938 239782 349174
rect 239866 348938 240102 349174
rect 239546 348618 239782 348854
rect 239866 348618 240102 348854
rect 235826 309218 236062 309454
rect 236146 309218 236382 309454
rect 235826 308898 236062 309134
rect 236146 308898 236382 309134
rect 235170 255218 235406 255454
rect 235170 254898 235406 255134
rect 235826 237218 236062 237454
rect 236146 237218 236382 237454
rect 235826 236898 236062 237134
rect 236146 236898 236382 237134
rect 221249 129218 221485 129454
rect 221249 128898 221485 129134
rect 224513 129218 224749 129454
rect 224513 128898 224749 129134
rect 219617 111218 219853 111454
rect 219617 110898 219853 111134
rect 222881 111218 223117 111454
rect 222881 110898 223117 111134
rect 226145 111218 226381 111454
rect 226145 110898 226381 111134
rect 210986 68378 211222 68614
rect 211306 68378 211542 68614
rect 210986 68058 211222 68294
rect 211306 68058 211542 68294
rect 210986 32378 211222 32614
rect 211306 32378 211542 32614
rect 210986 32058 211222 32294
rect 211306 32058 211542 32294
rect 192986 -6342 193222 -6106
rect 193306 -6342 193542 -6106
rect 192986 -6662 193222 -6426
rect 193306 -6662 193542 -6426
rect 217826 75218 218062 75454
rect 218146 75218 218382 75454
rect 217826 74898 218062 75134
rect 218146 74898 218382 75134
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 221546 78938 221782 79174
rect 221866 78938 222102 79174
rect 221546 78618 221782 78854
rect 221866 78618 222102 78854
rect 221546 42938 221782 43174
rect 221866 42938 222102 43174
rect 221546 42618 221782 42854
rect 221866 42618 222102 42854
rect 221546 6938 221782 7174
rect 221866 6938 222102 7174
rect 221546 6618 221782 6854
rect 221866 6618 222102 6854
rect 221546 -2502 221782 -2266
rect 221866 -2502 222102 -2266
rect 221546 -2822 221782 -2586
rect 221866 -2822 222102 -2586
rect 225266 82658 225502 82894
rect 225586 82658 225822 82894
rect 225266 82338 225502 82574
rect 225586 82338 225822 82574
rect 225266 46658 225502 46894
rect 225586 46658 225822 46894
rect 225266 46338 225502 46574
rect 225586 46338 225822 46574
rect 225266 10658 225502 10894
rect 225586 10658 225822 10894
rect 225266 10338 225502 10574
rect 225586 10338 225822 10574
rect 228986 86378 229222 86614
rect 229306 86378 229542 86614
rect 228986 86058 229222 86294
rect 229306 86058 229542 86294
rect 228986 50378 229222 50614
rect 229306 50378 229542 50614
rect 228986 50058 229222 50294
rect 229306 50058 229542 50294
rect 235826 201218 236062 201454
rect 236146 201218 236382 201454
rect 235826 200898 236062 201134
rect 236146 200898 236382 201134
rect 239546 312938 239782 313174
rect 239866 312938 240102 313174
rect 239546 312618 239782 312854
rect 239866 312618 240102 312854
rect 235826 165218 236062 165454
rect 236146 165218 236382 165454
rect 235826 164898 236062 165134
rect 236146 164898 236382 165134
rect 243266 352658 243502 352894
rect 243586 352658 243822 352894
rect 243266 352338 243502 352574
rect 243586 352338 243822 352574
rect 246986 356378 247222 356614
rect 247306 356378 247542 356614
rect 246986 356058 247222 356294
rect 247306 356058 247542 356294
rect 243266 316658 243502 316894
rect 243586 316658 243822 316894
rect 243266 316338 243502 316574
rect 243586 316338 243822 316574
rect 246986 320378 247222 320614
rect 247306 320378 247542 320614
rect 246986 320058 247222 320294
rect 247306 320058 247542 320294
rect 246986 284378 247222 284614
rect 247306 284378 247542 284614
rect 246986 284058 247222 284294
rect 247306 284058 247542 284294
rect 239546 204938 239782 205174
rect 239866 204938 240102 205174
rect 239546 204618 239782 204854
rect 239866 204618 240102 204854
rect 239546 168938 239782 169174
rect 239866 168938 240102 169174
rect 239546 168618 239782 168854
rect 239866 168618 240102 168854
rect 235826 129218 236062 129454
rect 236146 129218 236382 129454
rect 235826 128898 236062 129134
rect 236146 128898 236382 129134
rect 235826 93218 236062 93454
rect 236146 93218 236382 93454
rect 235826 92898 236062 93134
rect 236146 92898 236382 93134
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 228986 14378 229222 14614
rect 229306 14378 229542 14614
rect 228986 14058 229222 14294
rect 229306 14058 229542 14294
rect 225266 -4422 225502 -4186
rect 225586 -4422 225822 -4186
rect 225266 -4742 225502 -4506
rect 225586 -4742 225822 -4506
rect 210986 -7302 211222 -7066
rect 211306 -7302 211542 -7066
rect 210986 -7622 211222 -7386
rect 211306 -7622 211542 -7386
rect 239546 132938 239782 133174
rect 239866 132938 240102 133174
rect 239546 132618 239782 132854
rect 239866 132618 240102 132854
rect 243266 208658 243502 208894
rect 243586 208658 243822 208894
rect 243266 208338 243502 208574
rect 243586 208338 243822 208574
rect 243266 172658 243502 172894
rect 243586 172658 243822 172894
rect 243266 172338 243502 172574
rect 243586 172338 243822 172574
rect 243266 136658 243502 136894
rect 243586 136658 243822 136894
rect 243266 136338 243502 136574
rect 243586 136338 243822 136574
rect 239546 96938 239782 97174
rect 239866 96938 240102 97174
rect 239546 96618 239782 96854
rect 239866 96618 240102 96854
rect 243266 100658 243502 100894
rect 243586 100658 243822 100894
rect 243266 100338 243502 100574
rect 243586 100338 243822 100574
rect 239546 60938 239782 61174
rect 239866 60938 240102 61174
rect 239546 60618 239782 60854
rect 239866 60618 240102 60854
rect 239546 24938 239782 25174
rect 239866 24938 240102 25174
rect 239546 24618 239782 24854
rect 239866 24618 240102 24854
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -1542 236062 -1306
rect 236146 -1542 236382 -1306
rect 235826 -1862 236062 -1626
rect 236146 -1862 236382 -1626
rect 239546 -3462 239782 -3226
rect 239866 -3462 240102 -3226
rect 239546 -3782 239782 -3546
rect 239866 -3782 240102 -3546
rect 243266 64658 243502 64894
rect 243586 64658 243822 64894
rect 243266 64338 243502 64574
rect 243586 64338 243822 64574
rect 243266 28658 243502 28894
rect 243586 28658 243822 28894
rect 243266 28338 243502 28574
rect 243586 28338 243822 28574
rect 246986 248378 247222 248614
rect 247306 248378 247542 248614
rect 246986 248058 247222 248294
rect 247306 248058 247542 248294
rect 246986 212378 247222 212614
rect 247306 212378 247542 212614
rect 246986 212058 247222 212294
rect 247306 212058 247542 212294
rect 246986 176378 247222 176614
rect 247306 176378 247542 176614
rect 246986 176058 247222 176294
rect 247306 176058 247542 176294
rect 246986 140378 247222 140614
rect 247306 140378 247542 140614
rect 246986 140058 247222 140294
rect 247306 140058 247542 140294
rect 246986 104378 247222 104614
rect 247306 104378 247542 104614
rect 246986 104058 247222 104294
rect 247306 104058 247542 104294
rect 246986 68378 247222 68614
rect 247306 68378 247542 68614
rect 246986 68058 247222 68294
rect 247306 68058 247542 68294
rect 253826 363218 254062 363454
rect 254146 363218 254382 363454
rect 253826 362898 254062 363134
rect 254146 362898 254382 363134
rect 253826 327218 254062 327454
rect 254146 327218 254382 327454
rect 253826 326898 254062 327134
rect 254146 326898 254382 327134
rect 257546 366938 257782 367174
rect 257866 366938 258102 367174
rect 257546 366618 257782 366854
rect 257866 366618 258102 366854
rect 257546 330938 257782 331174
rect 257866 330938 258102 331174
rect 257546 330618 257782 330854
rect 257866 330618 258102 330854
rect 253826 291218 254062 291454
rect 254146 291218 254382 291454
rect 253826 290898 254062 291134
rect 254146 290898 254382 291134
rect 253826 255218 254062 255454
rect 254146 255218 254382 255454
rect 253826 254898 254062 255134
rect 254146 254898 254382 255134
rect 253826 219218 254062 219454
rect 254146 219218 254382 219454
rect 253826 218898 254062 219134
rect 254146 218898 254382 219134
rect 261266 370658 261502 370894
rect 261586 370658 261822 370894
rect 261266 370338 261502 370574
rect 261586 370338 261822 370574
rect 261266 334658 261502 334894
rect 261586 334658 261822 334894
rect 261266 334338 261502 334574
rect 261586 334338 261822 334574
rect 257546 294938 257782 295174
rect 257866 294938 258102 295174
rect 257546 294618 257782 294854
rect 257866 294618 258102 294854
rect 257546 258938 257782 259174
rect 257866 258938 258102 259174
rect 257546 258618 257782 258854
rect 257866 258618 258102 258854
rect 261266 298658 261502 298894
rect 261586 298658 261822 298894
rect 261266 298338 261502 298574
rect 261586 298338 261822 298574
rect 261266 262658 261502 262894
rect 261586 262658 261822 262894
rect 261266 262338 261502 262574
rect 261586 262338 261822 262574
rect 257546 222938 257782 223174
rect 257866 222938 258102 223174
rect 257546 222618 257782 222854
rect 257866 222618 258102 222854
rect 253826 183218 254062 183454
rect 254146 183218 254382 183454
rect 253826 182898 254062 183134
rect 254146 182898 254382 183134
rect 253826 147218 254062 147454
rect 254146 147218 254382 147454
rect 253826 146898 254062 147134
rect 254146 146898 254382 147134
rect 253826 111218 254062 111454
rect 254146 111218 254382 111454
rect 253826 110898 254062 111134
rect 254146 110898 254382 111134
rect 253826 75218 254062 75454
rect 254146 75218 254382 75454
rect 253826 74898 254062 75134
rect 254146 74898 254382 75134
rect 246986 32378 247222 32614
rect 247306 32378 247542 32614
rect 246986 32058 247222 32294
rect 247306 32058 247542 32294
rect 243266 -5382 243502 -5146
rect 243586 -5382 243822 -5146
rect 243266 -5702 243502 -5466
rect 243586 -5702 243822 -5466
rect 228986 -6342 229222 -6106
rect 229306 -6342 229542 -6106
rect 228986 -6662 229222 -6426
rect 229306 -6662 229542 -6426
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 257546 186938 257782 187174
rect 257866 186938 258102 187174
rect 257546 186618 257782 186854
rect 257866 186618 258102 186854
rect 257546 150938 257782 151174
rect 257866 150938 258102 151174
rect 257546 150618 257782 150854
rect 257866 150618 258102 150854
rect 261266 226658 261502 226894
rect 261586 226658 261822 226894
rect 261266 226338 261502 226574
rect 261586 226338 261822 226574
rect 261266 190658 261502 190894
rect 261586 190658 261822 190894
rect 261266 190338 261502 190574
rect 261586 190338 261822 190574
rect 261266 154658 261502 154894
rect 261586 154658 261822 154894
rect 261266 154338 261502 154574
rect 261586 154338 261822 154574
rect 257546 114938 257782 115174
rect 257866 114938 258102 115174
rect 257546 114618 257782 114854
rect 257866 114618 258102 114854
rect 257546 78938 257782 79174
rect 257866 78938 258102 79174
rect 257546 78618 257782 78854
rect 257866 78618 258102 78854
rect 264986 374378 265222 374614
rect 265306 374378 265542 374614
rect 264986 374058 265222 374294
rect 265306 374058 265542 374294
rect 264986 338378 265222 338614
rect 265306 338378 265542 338614
rect 264986 338058 265222 338294
rect 265306 338058 265542 338294
rect 264986 302378 265222 302614
rect 265306 302378 265542 302614
rect 264986 302058 265222 302294
rect 265306 302058 265542 302294
rect 264986 266378 265222 266614
rect 265306 266378 265542 266614
rect 264986 266058 265222 266294
rect 265306 266058 265542 266294
rect 264986 230378 265222 230614
rect 265306 230378 265542 230614
rect 264986 230058 265222 230294
rect 265306 230058 265542 230294
rect 264986 194378 265222 194614
rect 265306 194378 265542 194614
rect 264986 194058 265222 194294
rect 265306 194058 265542 194294
rect 264986 158378 265222 158614
rect 265306 158378 265542 158614
rect 264986 158058 265222 158294
rect 265306 158058 265542 158294
rect 261266 118658 261502 118894
rect 261586 118658 261822 118894
rect 261266 118338 261502 118574
rect 261586 118338 261822 118574
rect 261266 82658 261502 82894
rect 261586 82658 261822 82894
rect 261266 82338 261502 82574
rect 261586 82338 261822 82574
rect 257546 42938 257782 43174
rect 257866 42938 258102 43174
rect 257546 42618 257782 42854
rect 257866 42618 258102 42854
rect 257546 6938 257782 7174
rect 257866 6938 258102 7174
rect 257546 6618 257782 6854
rect 257866 6618 258102 6854
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 257546 -2502 257782 -2266
rect 257866 -2502 258102 -2266
rect 257546 -2822 257782 -2586
rect 257866 -2822 258102 -2586
rect 264986 122378 265222 122614
rect 265306 122378 265542 122614
rect 264986 122058 265222 122294
rect 265306 122058 265542 122294
rect 264986 86378 265222 86614
rect 265306 86378 265542 86614
rect 264986 86058 265222 86294
rect 265306 86058 265542 86294
rect 261266 46658 261502 46894
rect 261586 46658 261822 46894
rect 261266 46338 261502 46574
rect 261586 46338 261822 46574
rect 261266 10658 261502 10894
rect 261586 10658 261822 10894
rect 261266 10338 261502 10574
rect 261586 10338 261822 10574
rect 261266 -4422 261502 -4186
rect 261586 -4422 261822 -4186
rect 261266 -4742 261502 -4506
rect 261586 -4742 261822 -4506
rect 264986 50378 265222 50614
rect 265306 50378 265542 50614
rect 264986 50058 265222 50294
rect 265306 50058 265542 50294
rect 271826 345218 272062 345454
rect 272146 345218 272382 345454
rect 271826 344898 272062 345134
rect 272146 344898 272382 345134
rect 271826 309218 272062 309454
rect 272146 309218 272382 309454
rect 271826 308898 272062 309134
rect 272146 308898 272382 309134
rect 271826 273218 272062 273454
rect 272146 273218 272382 273454
rect 271826 272898 272062 273134
rect 272146 272898 272382 273134
rect 271826 237218 272062 237454
rect 272146 237218 272382 237454
rect 271826 236898 272062 237134
rect 272146 236898 272382 237134
rect 271826 201218 272062 201454
rect 272146 201218 272382 201454
rect 271826 200898 272062 201134
rect 272146 200898 272382 201134
rect 275546 348938 275782 349174
rect 275866 348938 276102 349174
rect 275546 348618 275782 348854
rect 275866 348618 276102 348854
rect 275546 312938 275782 313174
rect 275866 312938 276102 313174
rect 275546 312618 275782 312854
rect 275866 312618 276102 312854
rect 275546 276938 275782 277174
rect 275866 276938 276102 277174
rect 275546 276618 275782 276854
rect 275866 276618 276102 276854
rect 275546 240938 275782 241174
rect 275866 240938 276102 241174
rect 275546 240618 275782 240854
rect 275866 240618 276102 240854
rect 275546 204938 275782 205174
rect 275866 204938 276102 205174
rect 275546 204618 275782 204854
rect 275866 204618 276102 204854
rect 279266 352658 279502 352894
rect 279586 352658 279822 352894
rect 279266 352338 279502 352574
rect 279586 352338 279822 352574
rect 279266 316658 279502 316894
rect 279586 316658 279822 316894
rect 279266 316338 279502 316574
rect 279586 316338 279822 316574
rect 279266 280658 279502 280894
rect 279586 280658 279822 280894
rect 279266 280338 279502 280574
rect 279586 280338 279822 280574
rect 282986 356378 283222 356614
rect 283306 356378 283542 356614
rect 282986 356058 283222 356294
rect 283306 356058 283542 356294
rect 282986 320378 283222 320614
rect 283306 320378 283542 320614
rect 282986 320058 283222 320294
rect 283306 320058 283542 320294
rect 282986 284378 283222 284614
rect 283306 284378 283542 284614
rect 282986 284058 283222 284294
rect 283306 284058 283542 284294
rect 279266 244658 279502 244894
rect 279586 244658 279822 244894
rect 279266 244338 279502 244574
rect 279586 244338 279822 244574
rect 279266 208658 279502 208894
rect 279586 208658 279822 208894
rect 279266 208338 279502 208574
rect 279586 208338 279822 208574
rect 272249 165218 272485 165454
rect 272249 164898 272485 165134
rect 275513 165218 275749 165454
rect 275513 164898 275749 165134
rect 270617 147218 270853 147454
rect 270617 146898 270853 147134
rect 273881 147218 274117 147454
rect 273881 146898 274117 147134
rect 277145 147218 277381 147454
rect 277145 146898 277381 147134
rect 272249 129218 272485 129454
rect 272249 128898 272485 129134
rect 275513 129218 275749 129454
rect 275513 128898 275749 129134
rect 270617 111218 270853 111454
rect 270617 110898 270853 111134
rect 273881 111218 274117 111454
rect 273881 110898 274117 111134
rect 277145 111218 277381 111454
rect 277145 110898 277381 111134
rect 282986 248378 283222 248614
rect 283306 248378 283542 248614
rect 282986 248058 283222 248294
rect 283306 248058 283542 248294
rect 282986 212378 283222 212614
rect 283306 212378 283542 212614
rect 282986 212058 283222 212294
rect 283306 212058 283542 212294
rect 282986 176378 283222 176614
rect 283306 176378 283542 176614
rect 282986 176058 283222 176294
rect 283306 176058 283542 176294
rect 282986 140378 283222 140614
rect 283306 140378 283542 140614
rect 282986 140058 283222 140294
rect 283306 140058 283542 140294
rect 282986 104378 283222 104614
rect 283306 104378 283542 104614
rect 282986 104058 283222 104294
rect 283306 104058 283542 104294
rect 271826 93218 272062 93454
rect 272146 93218 272382 93454
rect 271826 92898 272062 93134
rect 272146 92898 272382 93134
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 264986 14378 265222 14614
rect 265306 14378 265542 14614
rect 264986 14058 265222 14294
rect 265306 14058 265542 14294
rect 246986 -7302 247222 -7066
rect 247306 -7302 247542 -7066
rect 246986 -7622 247222 -7386
rect 247306 -7622 247542 -7386
rect 271826 -1542 272062 -1306
rect 272146 -1542 272382 -1306
rect 271826 -1862 272062 -1626
rect 272146 -1862 272382 -1626
rect 275546 60938 275782 61174
rect 275866 60938 276102 61174
rect 275546 60618 275782 60854
rect 275866 60618 276102 60854
rect 275546 24938 275782 25174
rect 275866 24938 276102 25174
rect 275546 24618 275782 24854
rect 275866 24618 276102 24854
rect 275546 -3462 275782 -3226
rect 275866 -3462 276102 -3226
rect 275546 -3782 275782 -3546
rect 275866 -3782 276102 -3546
rect 279266 64658 279502 64894
rect 279586 64658 279822 64894
rect 279266 64338 279502 64574
rect 279586 64338 279822 64574
rect 279266 28658 279502 28894
rect 279586 28658 279822 28894
rect 279266 28338 279502 28574
rect 279586 28338 279822 28574
rect 279266 -5382 279502 -5146
rect 279586 -5382 279822 -5146
rect 279266 -5702 279502 -5466
rect 279586 -5702 279822 -5466
rect 282986 68378 283222 68614
rect 283306 68378 283542 68614
rect 282986 68058 283222 68294
rect 283306 68058 283542 68294
rect 289826 363218 290062 363454
rect 290146 363218 290382 363454
rect 289826 362898 290062 363134
rect 290146 362898 290382 363134
rect 289826 327218 290062 327454
rect 290146 327218 290382 327454
rect 289826 326898 290062 327134
rect 290146 326898 290382 327134
rect 289826 291218 290062 291454
rect 290146 291218 290382 291454
rect 289826 290898 290062 291134
rect 290146 290898 290382 291134
rect 289826 255218 290062 255454
rect 290146 255218 290382 255454
rect 289826 254898 290062 255134
rect 290146 254898 290382 255134
rect 289826 219218 290062 219454
rect 290146 219218 290382 219454
rect 289826 218898 290062 219134
rect 290146 218898 290382 219134
rect 293546 366938 293782 367174
rect 293866 366938 294102 367174
rect 293546 366618 293782 366854
rect 293866 366618 294102 366854
rect 297266 370658 297502 370894
rect 297586 370658 297822 370894
rect 297266 370338 297502 370574
rect 297586 370338 297822 370574
rect 293546 330938 293782 331174
rect 293866 330938 294102 331174
rect 293546 330618 293782 330854
rect 293866 330618 294102 330854
rect 293546 294938 293782 295174
rect 293866 294938 294102 295174
rect 293546 294618 293782 294854
rect 293866 294618 294102 294854
rect 293546 258938 293782 259174
rect 293866 258938 294102 259174
rect 293546 258618 293782 258854
rect 293866 258618 294102 258854
rect 293546 222938 293782 223174
rect 293866 222938 294102 223174
rect 293546 222618 293782 222854
rect 293866 222618 294102 222854
rect 289826 183218 290062 183454
rect 290146 183218 290382 183454
rect 289826 182898 290062 183134
rect 290146 182898 290382 183134
rect 289826 147218 290062 147454
rect 290146 147218 290382 147454
rect 289826 146898 290062 147134
rect 290146 146898 290382 147134
rect 289826 111218 290062 111454
rect 290146 111218 290382 111454
rect 289826 110898 290062 111134
rect 290146 110898 290382 111134
rect 289826 75218 290062 75454
rect 290146 75218 290382 75454
rect 289826 74898 290062 75134
rect 290146 74898 290382 75134
rect 282986 32378 283222 32614
rect 283306 32378 283542 32614
rect 282986 32058 283222 32294
rect 283306 32058 283542 32294
rect 264986 -6342 265222 -6106
rect 265306 -6342 265542 -6106
rect 264986 -6662 265222 -6426
rect 265306 -6662 265542 -6426
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 293546 186938 293782 187174
rect 293866 186938 294102 187174
rect 293546 186618 293782 186854
rect 293866 186618 294102 186854
rect 293546 150938 293782 151174
rect 293866 150938 294102 151174
rect 293546 150618 293782 150854
rect 293866 150618 294102 150854
rect 293546 114938 293782 115174
rect 293866 114938 294102 115174
rect 293546 114618 293782 114854
rect 293866 114618 294102 114854
rect 293546 78938 293782 79174
rect 293866 78938 294102 79174
rect 293546 78618 293782 78854
rect 293866 78618 294102 78854
rect 293546 42938 293782 43174
rect 293866 42938 294102 43174
rect 293546 42618 293782 42854
rect 293866 42618 294102 42854
rect 297266 334658 297502 334894
rect 297586 334658 297822 334894
rect 297266 334338 297502 334574
rect 297586 334338 297822 334574
rect 297266 298658 297502 298894
rect 297586 298658 297822 298894
rect 297266 298338 297502 298574
rect 297586 298338 297822 298574
rect 297266 262658 297502 262894
rect 297586 262658 297822 262894
rect 297266 262338 297502 262574
rect 297586 262338 297822 262574
rect 297266 226658 297502 226894
rect 297586 226658 297822 226894
rect 297266 226338 297502 226574
rect 297586 226338 297822 226574
rect 300986 374378 301222 374614
rect 301306 374378 301542 374614
rect 300986 374058 301222 374294
rect 301306 374058 301542 374294
rect 300986 338378 301222 338614
rect 301306 338378 301542 338614
rect 300986 338058 301222 338294
rect 301306 338058 301542 338294
rect 300986 302378 301222 302614
rect 301306 302378 301542 302614
rect 300986 302058 301222 302294
rect 301306 302058 301542 302294
rect 300986 266378 301222 266614
rect 301306 266378 301542 266614
rect 300986 266058 301222 266294
rect 301306 266058 301542 266294
rect 300986 230378 301222 230614
rect 301306 230378 301542 230614
rect 300986 230058 301222 230294
rect 301306 230058 301542 230294
rect 297266 190658 297502 190894
rect 297586 190658 297822 190894
rect 297266 190338 297502 190574
rect 297586 190338 297822 190574
rect 297266 154658 297502 154894
rect 297586 154658 297822 154894
rect 297266 154338 297502 154574
rect 297586 154338 297822 154574
rect 300986 194378 301222 194614
rect 301306 194378 301542 194614
rect 300986 194058 301222 194294
rect 301306 194058 301542 194294
rect 297266 118658 297502 118894
rect 297586 118658 297822 118894
rect 297266 118338 297502 118574
rect 297586 118338 297822 118574
rect 297266 82658 297502 82894
rect 297586 82658 297822 82894
rect 297266 82338 297502 82574
rect 297586 82338 297822 82574
rect 297266 46658 297502 46894
rect 297586 46658 297822 46894
rect 297266 46338 297502 46574
rect 297586 46338 297822 46574
rect 293546 6938 293782 7174
rect 293866 6938 294102 7174
rect 293546 6618 293782 6854
rect 293866 6618 294102 6854
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 293546 -2502 293782 -2266
rect 293866 -2502 294102 -2266
rect 293546 -2822 293782 -2586
rect 293866 -2822 294102 -2586
rect 307826 345218 308062 345454
rect 308146 345218 308382 345454
rect 307826 344898 308062 345134
rect 308146 344898 308382 345134
rect 307826 309218 308062 309454
rect 308146 309218 308382 309454
rect 307826 308898 308062 309134
rect 308146 308898 308382 309134
rect 307826 273218 308062 273454
rect 308146 273218 308382 273454
rect 307826 272898 308062 273134
rect 308146 272898 308382 273134
rect 307826 237218 308062 237454
rect 308146 237218 308382 237454
rect 307826 236898 308062 237134
rect 308146 236898 308382 237134
rect 307826 201218 308062 201454
rect 308146 201218 308382 201454
rect 307826 200898 308062 201134
rect 308146 200898 308382 201134
rect 300986 158378 301222 158614
rect 301306 158378 301542 158614
rect 300986 158058 301222 158294
rect 301306 158058 301542 158294
rect 307826 165218 308062 165454
rect 308146 165218 308382 165454
rect 307826 164898 308062 165134
rect 308146 164898 308382 165134
rect 300986 122378 301222 122614
rect 301306 122378 301542 122614
rect 300986 122058 301222 122294
rect 301306 122058 301542 122294
rect 300986 86378 301222 86614
rect 301306 86378 301542 86614
rect 300986 86058 301222 86294
rect 301306 86058 301542 86294
rect 300986 50378 301222 50614
rect 301306 50378 301542 50614
rect 300986 50058 301222 50294
rect 301306 50058 301542 50294
rect 300986 14378 301222 14614
rect 301306 14378 301542 14614
rect 300986 14058 301222 14294
rect 301306 14058 301542 14294
rect 297266 10658 297502 10894
rect 297586 10658 297822 10894
rect 297266 10338 297502 10574
rect 297586 10338 297822 10574
rect 297266 -4422 297502 -4186
rect 297586 -4422 297822 -4186
rect 297266 -4742 297502 -4506
rect 297586 -4742 297822 -4506
rect 282986 -7302 283222 -7066
rect 283306 -7302 283542 -7066
rect 282986 -7622 283222 -7386
rect 283306 -7622 283542 -7386
rect 307826 129218 308062 129454
rect 308146 129218 308382 129454
rect 307826 128898 308062 129134
rect 308146 128898 308382 129134
rect 307826 93218 308062 93454
rect 308146 93218 308382 93454
rect 307826 92898 308062 93134
rect 308146 92898 308382 93134
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -1542 308062 -1306
rect 308146 -1542 308382 -1306
rect 307826 -1862 308062 -1626
rect 308146 -1862 308382 -1626
rect 311546 348938 311782 349174
rect 311866 348938 312102 349174
rect 311546 348618 311782 348854
rect 311866 348618 312102 348854
rect 311546 312938 311782 313174
rect 311866 312938 312102 313174
rect 311546 312618 311782 312854
rect 311866 312618 312102 312854
rect 311546 276938 311782 277174
rect 311866 276938 312102 277174
rect 311546 276618 311782 276854
rect 311866 276618 312102 276854
rect 311546 240938 311782 241174
rect 311866 240938 312102 241174
rect 311546 240618 311782 240854
rect 311866 240618 312102 240854
rect 311546 204938 311782 205174
rect 311866 204938 312102 205174
rect 311546 204618 311782 204854
rect 311866 204618 312102 204854
rect 311546 168938 311782 169174
rect 311866 168938 312102 169174
rect 311546 168618 311782 168854
rect 311866 168618 312102 168854
rect 311546 132938 311782 133174
rect 311866 132938 312102 133174
rect 311546 132618 311782 132854
rect 311866 132618 312102 132854
rect 311546 96938 311782 97174
rect 311866 96938 312102 97174
rect 311546 96618 311782 96854
rect 311866 96618 312102 96854
rect 311546 60938 311782 61174
rect 311866 60938 312102 61174
rect 311546 60618 311782 60854
rect 311866 60618 312102 60854
rect 311546 24938 311782 25174
rect 311866 24938 312102 25174
rect 311546 24618 311782 24854
rect 311866 24618 312102 24854
rect 311546 -3462 311782 -3226
rect 311866 -3462 312102 -3226
rect 311546 -3782 311782 -3546
rect 311866 -3782 312102 -3546
rect 315266 352658 315502 352894
rect 315586 352658 315822 352894
rect 315266 352338 315502 352574
rect 315586 352338 315822 352574
rect 315266 316658 315502 316894
rect 315586 316658 315822 316894
rect 315266 316338 315502 316574
rect 315586 316338 315822 316574
rect 315266 280658 315502 280894
rect 315586 280658 315822 280894
rect 315266 280338 315502 280574
rect 315586 280338 315822 280574
rect 315266 244658 315502 244894
rect 315586 244658 315822 244894
rect 315266 244338 315502 244574
rect 315586 244338 315822 244574
rect 315266 208658 315502 208894
rect 315586 208658 315822 208894
rect 315266 208338 315502 208574
rect 315586 208338 315822 208574
rect 315266 172658 315502 172894
rect 315586 172658 315822 172894
rect 315266 172338 315502 172574
rect 315586 172338 315822 172574
rect 315266 136658 315502 136894
rect 315586 136658 315822 136894
rect 315266 136338 315502 136574
rect 315586 136338 315822 136574
rect 315266 100658 315502 100894
rect 315586 100658 315822 100894
rect 315266 100338 315502 100574
rect 315586 100338 315822 100574
rect 315266 64658 315502 64894
rect 315586 64658 315822 64894
rect 315266 64338 315502 64574
rect 315586 64338 315822 64574
rect 315266 28658 315502 28894
rect 315586 28658 315822 28894
rect 315266 28338 315502 28574
rect 315586 28338 315822 28574
rect 315266 -5382 315502 -5146
rect 315586 -5382 315822 -5146
rect 315266 -5702 315502 -5466
rect 315586 -5702 315822 -5466
rect 318986 356378 319222 356614
rect 319306 356378 319542 356614
rect 318986 356058 319222 356294
rect 319306 356058 319542 356294
rect 318986 320378 319222 320614
rect 319306 320378 319542 320614
rect 318986 320058 319222 320294
rect 319306 320058 319542 320294
rect 318986 284378 319222 284614
rect 319306 284378 319542 284614
rect 318986 284058 319222 284294
rect 319306 284058 319542 284294
rect 318986 248378 319222 248614
rect 319306 248378 319542 248614
rect 318986 248058 319222 248294
rect 319306 248058 319542 248294
rect 318986 212378 319222 212614
rect 319306 212378 319542 212614
rect 318986 212058 319222 212294
rect 319306 212058 319542 212294
rect 318986 176378 319222 176614
rect 319306 176378 319542 176614
rect 318986 176058 319222 176294
rect 319306 176058 319542 176294
rect 318986 140378 319222 140614
rect 319306 140378 319542 140614
rect 318986 140058 319222 140294
rect 319306 140058 319542 140294
rect 318986 104378 319222 104614
rect 319306 104378 319542 104614
rect 318986 104058 319222 104294
rect 319306 104058 319542 104294
rect 318986 68378 319222 68614
rect 319306 68378 319542 68614
rect 318986 68058 319222 68294
rect 319306 68058 319542 68294
rect 318986 32378 319222 32614
rect 319306 32378 319542 32614
rect 318986 32058 319222 32294
rect 319306 32058 319542 32294
rect 300986 -6342 301222 -6106
rect 301306 -6342 301542 -6106
rect 300986 -6662 301222 -6426
rect 301306 -6662 301542 -6426
rect 325826 363218 326062 363454
rect 326146 363218 326382 363454
rect 325826 362898 326062 363134
rect 326146 362898 326382 363134
rect 325826 327218 326062 327454
rect 326146 327218 326382 327454
rect 325826 326898 326062 327134
rect 326146 326898 326382 327134
rect 325826 291218 326062 291454
rect 326146 291218 326382 291454
rect 325826 290898 326062 291134
rect 326146 290898 326382 291134
rect 325826 255218 326062 255454
rect 326146 255218 326382 255454
rect 325826 254898 326062 255134
rect 326146 254898 326382 255134
rect 325826 219218 326062 219454
rect 326146 219218 326382 219454
rect 325826 218898 326062 219134
rect 326146 218898 326382 219134
rect 325826 183218 326062 183454
rect 326146 183218 326382 183454
rect 325826 182898 326062 183134
rect 326146 182898 326382 183134
rect 325826 147218 326062 147454
rect 326146 147218 326382 147454
rect 325826 146898 326062 147134
rect 326146 146898 326382 147134
rect 325826 111218 326062 111454
rect 326146 111218 326382 111454
rect 325826 110898 326062 111134
rect 326146 110898 326382 111134
rect 325826 75218 326062 75454
rect 326146 75218 326382 75454
rect 325826 74898 326062 75134
rect 326146 74898 326382 75134
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 329546 366938 329782 367174
rect 329866 366938 330102 367174
rect 329546 366618 329782 366854
rect 329866 366618 330102 366854
rect 329546 330938 329782 331174
rect 329866 330938 330102 331174
rect 329546 330618 329782 330854
rect 329866 330618 330102 330854
rect 329546 294938 329782 295174
rect 329866 294938 330102 295174
rect 329546 294618 329782 294854
rect 329866 294618 330102 294854
rect 329546 258938 329782 259174
rect 329866 258938 330102 259174
rect 329546 258618 329782 258854
rect 329866 258618 330102 258854
rect 329546 222938 329782 223174
rect 329866 222938 330102 223174
rect 329546 222618 329782 222854
rect 329866 222618 330102 222854
rect 329546 186938 329782 187174
rect 329866 186938 330102 187174
rect 329546 186618 329782 186854
rect 329866 186618 330102 186854
rect 329546 150938 329782 151174
rect 329866 150938 330102 151174
rect 329546 150618 329782 150854
rect 329866 150618 330102 150854
rect 329546 114938 329782 115174
rect 329866 114938 330102 115174
rect 329546 114618 329782 114854
rect 329866 114618 330102 114854
rect 329546 78938 329782 79174
rect 329866 78938 330102 79174
rect 329546 78618 329782 78854
rect 329866 78618 330102 78854
rect 329546 42938 329782 43174
rect 329866 42938 330102 43174
rect 329546 42618 329782 42854
rect 329866 42618 330102 42854
rect 329546 6938 329782 7174
rect 329866 6938 330102 7174
rect 329546 6618 329782 6854
rect 329866 6618 330102 6854
rect 329546 -2502 329782 -2266
rect 329866 -2502 330102 -2266
rect 329546 -2822 329782 -2586
rect 329866 -2822 330102 -2586
rect 333266 370658 333502 370894
rect 333586 370658 333822 370894
rect 333266 370338 333502 370574
rect 333586 370338 333822 370574
rect 333266 334658 333502 334894
rect 333586 334658 333822 334894
rect 333266 334338 333502 334574
rect 333586 334338 333822 334574
rect 333266 298658 333502 298894
rect 333586 298658 333822 298894
rect 333266 298338 333502 298574
rect 333586 298338 333822 298574
rect 333266 262658 333502 262894
rect 333586 262658 333822 262894
rect 333266 262338 333502 262574
rect 333586 262338 333822 262574
rect 333266 226658 333502 226894
rect 333586 226658 333822 226894
rect 333266 226338 333502 226574
rect 333586 226338 333822 226574
rect 333266 190658 333502 190894
rect 333586 190658 333822 190894
rect 333266 190338 333502 190574
rect 333586 190338 333822 190574
rect 333266 154658 333502 154894
rect 333586 154658 333822 154894
rect 333266 154338 333502 154574
rect 333586 154338 333822 154574
rect 333266 118658 333502 118894
rect 333586 118658 333822 118894
rect 333266 118338 333502 118574
rect 333586 118338 333822 118574
rect 333266 82658 333502 82894
rect 333586 82658 333822 82894
rect 333266 82338 333502 82574
rect 333586 82338 333822 82574
rect 333266 46658 333502 46894
rect 333586 46658 333822 46894
rect 333266 46338 333502 46574
rect 333586 46338 333822 46574
rect 333266 10658 333502 10894
rect 333586 10658 333822 10894
rect 333266 10338 333502 10574
rect 333586 10338 333822 10574
rect 333266 -4422 333502 -4186
rect 333586 -4422 333822 -4186
rect 333266 -4742 333502 -4506
rect 333586 -4742 333822 -4506
rect 336986 374378 337222 374614
rect 337306 374378 337542 374614
rect 336986 374058 337222 374294
rect 337306 374058 337542 374294
rect 336986 338378 337222 338614
rect 337306 338378 337542 338614
rect 336986 338058 337222 338294
rect 337306 338058 337542 338294
rect 336986 302378 337222 302614
rect 337306 302378 337542 302614
rect 336986 302058 337222 302294
rect 337306 302058 337542 302294
rect 336986 266378 337222 266614
rect 337306 266378 337542 266614
rect 336986 266058 337222 266294
rect 337306 266058 337542 266294
rect 336986 230378 337222 230614
rect 337306 230378 337542 230614
rect 336986 230058 337222 230294
rect 337306 230058 337542 230294
rect 336986 194378 337222 194614
rect 337306 194378 337542 194614
rect 336986 194058 337222 194294
rect 337306 194058 337542 194294
rect 336986 158378 337222 158614
rect 337306 158378 337542 158614
rect 336986 158058 337222 158294
rect 337306 158058 337542 158294
rect 336986 122378 337222 122614
rect 337306 122378 337542 122614
rect 336986 122058 337222 122294
rect 337306 122058 337542 122294
rect 336986 86378 337222 86614
rect 337306 86378 337542 86614
rect 336986 86058 337222 86294
rect 337306 86058 337542 86294
rect 336986 50378 337222 50614
rect 337306 50378 337542 50614
rect 336986 50058 337222 50294
rect 337306 50058 337542 50294
rect 336986 14378 337222 14614
rect 337306 14378 337542 14614
rect 336986 14058 337222 14294
rect 337306 14058 337542 14294
rect 318986 -7302 319222 -7066
rect 319306 -7302 319542 -7066
rect 318986 -7622 319222 -7386
rect 319306 -7622 319542 -7386
rect 343826 345218 344062 345454
rect 344146 345218 344382 345454
rect 343826 344898 344062 345134
rect 344146 344898 344382 345134
rect 343826 309218 344062 309454
rect 344146 309218 344382 309454
rect 343826 308898 344062 309134
rect 344146 308898 344382 309134
rect 343826 273218 344062 273454
rect 344146 273218 344382 273454
rect 343826 272898 344062 273134
rect 344146 272898 344382 273134
rect 343826 237218 344062 237454
rect 344146 237218 344382 237454
rect 343826 236898 344062 237134
rect 344146 236898 344382 237134
rect 343826 201218 344062 201454
rect 344146 201218 344382 201454
rect 343826 200898 344062 201134
rect 344146 200898 344382 201134
rect 343826 165218 344062 165454
rect 344146 165218 344382 165454
rect 343826 164898 344062 165134
rect 344146 164898 344382 165134
rect 343826 129218 344062 129454
rect 344146 129218 344382 129454
rect 343826 128898 344062 129134
rect 344146 128898 344382 129134
rect 343826 93218 344062 93454
rect 344146 93218 344382 93454
rect 343826 92898 344062 93134
rect 344146 92898 344382 93134
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -1542 344062 -1306
rect 344146 -1542 344382 -1306
rect 343826 -1862 344062 -1626
rect 344146 -1862 344382 -1626
rect 347546 348938 347782 349174
rect 347866 348938 348102 349174
rect 347546 348618 347782 348854
rect 347866 348618 348102 348854
rect 347546 312938 347782 313174
rect 347866 312938 348102 313174
rect 347546 312618 347782 312854
rect 347866 312618 348102 312854
rect 347546 276938 347782 277174
rect 347866 276938 348102 277174
rect 347546 276618 347782 276854
rect 347866 276618 348102 276854
rect 347546 240938 347782 241174
rect 347866 240938 348102 241174
rect 347546 240618 347782 240854
rect 347866 240618 348102 240854
rect 347546 204938 347782 205174
rect 347866 204938 348102 205174
rect 347546 204618 347782 204854
rect 347866 204618 348102 204854
rect 347546 168938 347782 169174
rect 347866 168938 348102 169174
rect 347546 168618 347782 168854
rect 347866 168618 348102 168854
rect 347546 132938 347782 133174
rect 347866 132938 348102 133174
rect 347546 132618 347782 132854
rect 347866 132618 348102 132854
rect 347546 96938 347782 97174
rect 347866 96938 348102 97174
rect 347546 96618 347782 96854
rect 347866 96618 348102 96854
rect 347546 60938 347782 61174
rect 347866 60938 348102 61174
rect 347546 60618 347782 60854
rect 347866 60618 348102 60854
rect 347546 24938 347782 25174
rect 347866 24938 348102 25174
rect 347546 24618 347782 24854
rect 347866 24618 348102 24854
rect 347546 -3462 347782 -3226
rect 347866 -3462 348102 -3226
rect 347546 -3782 347782 -3546
rect 347866 -3782 348102 -3546
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 351266 352658 351502 352894
rect 351586 352658 351822 352894
rect 351266 352338 351502 352574
rect 351586 352338 351822 352574
rect 351266 316658 351502 316894
rect 351586 316658 351822 316894
rect 351266 316338 351502 316574
rect 351586 316338 351822 316574
rect 351266 280658 351502 280894
rect 351586 280658 351822 280894
rect 351266 280338 351502 280574
rect 351586 280338 351822 280574
rect 351266 244658 351502 244894
rect 351586 244658 351822 244894
rect 351266 244338 351502 244574
rect 351586 244338 351822 244574
rect 351266 208658 351502 208894
rect 351586 208658 351822 208894
rect 351266 208338 351502 208574
rect 351586 208338 351822 208574
rect 351266 172658 351502 172894
rect 351586 172658 351822 172894
rect 351266 172338 351502 172574
rect 351586 172338 351822 172574
rect 351266 136658 351502 136894
rect 351586 136658 351822 136894
rect 351266 136338 351502 136574
rect 351586 136338 351822 136574
rect 351266 100658 351502 100894
rect 351586 100658 351822 100894
rect 351266 100338 351502 100574
rect 351586 100338 351822 100574
rect 351266 64658 351502 64894
rect 351586 64658 351822 64894
rect 351266 64338 351502 64574
rect 351586 64338 351822 64574
rect 351266 28658 351502 28894
rect 351586 28658 351822 28894
rect 351266 28338 351502 28574
rect 351586 28338 351822 28574
rect 351266 -5382 351502 -5146
rect 351586 -5382 351822 -5146
rect 351266 -5702 351502 -5466
rect 351586 -5702 351822 -5466
rect 361826 543218 362062 543454
rect 362146 543218 362382 543454
rect 361826 542898 362062 543134
rect 362146 542898 362382 543134
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 354986 356378 355222 356614
rect 355306 356378 355542 356614
rect 354986 356058 355222 356294
rect 355306 356058 355542 356294
rect 354986 320378 355222 320614
rect 355306 320378 355542 320614
rect 354986 320058 355222 320294
rect 355306 320058 355542 320294
rect 354986 284378 355222 284614
rect 355306 284378 355542 284614
rect 354986 284058 355222 284294
rect 355306 284058 355542 284294
rect 354986 248378 355222 248614
rect 355306 248378 355542 248614
rect 354986 248058 355222 248294
rect 355306 248058 355542 248294
rect 354986 212378 355222 212614
rect 355306 212378 355542 212614
rect 354986 212058 355222 212294
rect 355306 212058 355542 212294
rect 354986 176378 355222 176614
rect 355306 176378 355542 176614
rect 354986 176058 355222 176294
rect 355306 176058 355542 176294
rect 354986 140378 355222 140614
rect 355306 140378 355542 140614
rect 354986 140058 355222 140294
rect 355306 140058 355542 140294
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 361826 435218 362062 435454
rect 362146 435218 362382 435454
rect 361826 434898 362062 435134
rect 362146 434898 362382 435134
rect 361826 399218 362062 399454
rect 362146 399218 362382 399454
rect 361826 398898 362062 399134
rect 362146 398898 362382 399134
rect 361826 363218 362062 363454
rect 362146 363218 362382 363454
rect 361826 362898 362062 363134
rect 362146 362898 362382 363134
rect 361826 327218 362062 327454
rect 362146 327218 362382 327454
rect 361826 326898 362062 327134
rect 362146 326898 362382 327134
rect 361826 291218 362062 291454
rect 362146 291218 362382 291454
rect 361826 290898 362062 291134
rect 362146 290898 362382 291134
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 361826 219218 362062 219454
rect 362146 219218 362382 219454
rect 361826 218898 362062 219134
rect 362146 218898 362382 219134
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 354986 104378 355222 104614
rect 355306 104378 355542 104614
rect 354986 104058 355222 104294
rect 355306 104058 355542 104294
rect 354986 68378 355222 68614
rect 355306 68378 355542 68614
rect 354986 68058 355222 68294
rect 355306 68058 355542 68294
rect 354986 32378 355222 32614
rect 355306 32378 355542 32614
rect 354986 32058 355222 32294
rect 355306 32058 355542 32294
rect 336986 -6342 337222 -6106
rect 337306 -6342 337542 -6106
rect 336986 -6662 337222 -6426
rect 337306 -6662 337542 -6426
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 365546 690938 365782 691174
rect 365866 690938 366102 691174
rect 365546 690618 365782 690854
rect 365866 690618 366102 690854
rect 365546 654938 365782 655174
rect 365866 654938 366102 655174
rect 365546 654618 365782 654854
rect 365866 654618 366102 654854
rect 365546 618938 365782 619174
rect 365866 618938 366102 619174
rect 365546 618618 365782 618854
rect 365866 618618 366102 618854
rect 365546 582938 365782 583174
rect 365866 582938 366102 583174
rect 365546 582618 365782 582854
rect 365866 582618 366102 582854
rect 365546 546938 365782 547174
rect 365866 546938 366102 547174
rect 365546 546618 365782 546854
rect 365866 546618 366102 546854
rect 365546 510938 365782 511174
rect 365866 510938 366102 511174
rect 365546 510618 365782 510854
rect 365866 510618 366102 510854
rect 365546 474938 365782 475174
rect 365866 474938 366102 475174
rect 365546 474618 365782 474854
rect 365866 474618 366102 474854
rect 365546 438938 365782 439174
rect 365866 438938 366102 439174
rect 365546 438618 365782 438854
rect 365866 438618 366102 438854
rect 365546 402938 365782 403174
rect 365866 402938 366102 403174
rect 365546 402618 365782 402854
rect 365866 402618 366102 402854
rect 365546 366938 365782 367174
rect 365866 366938 366102 367174
rect 365546 366618 365782 366854
rect 365866 366618 366102 366854
rect 365546 330938 365782 331174
rect 365866 330938 366102 331174
rect 365546 330618 365782 330854
rect 365866 330618 366102 330854
rect 365546 294938 365782 295174
rect 365866 294938 366102 295174
rect 365546 294618 365782 294854
rect 365866 294618 366102 294854
rect 365546 258938 365782 259174
rect 365866 258938 366102 259174
rect 365546 258618 365782 258854
rect 365866 258618 366102 258854
rect 365546 222938 365782 223174
rect 365866 222938 366102 223174
rect 365546 222618 365782 222854
rect 365866 222618 366102 222854
rect 365546 186938 365782 187174
rect 365866 186938 366102 187174
rect 365546 186618 365782 186854
rect 365866 186618 366102 186854
rect 365546 150938 365782 151174
rect 365866 150938 366102 151174
rect 365546 150618 365782 150854
rect 365866 150618 366102 150854
rect 365546 114938 365782 115174
rect 365866 114938 366102 115174
rect 365546 114618 365782 114854
rect 365866 114618 366102 114854
rect 365546 78938 365782 79174
rect 365866 78938 366102 79174
rect 365546 78618 365782 78854
rect 365866 78618 366102 78854
rect 365546 42938 365782 43174
rect 365866 42938 366102 43174
rect 365546 42618 365782 42854
rect 365866 42618 366102 42854
rect 365546 6938 365782 7174
rect 365866 6938 366102 7174
rect 365546 6618 365782 6854
rect 365866 6618 366102 6854
rect 365546 -2502 365782 -2266
rect 365866 -2502 366102 -2266
rect 365546 -2822 365782 -2586
rect 365866 -2822 366102 -2586
rect 369266 694658 369502 694894
rect 369586 694658 369822 694894
rect 369266 694338 369502 694574
rect 369586 694338 369822 694574
rect 369266 658658 369502 658894
rect 369586 658658 369822 658894
rect 369266 658338 369502 658574
rect 369586 658338 369822 658574
rect 369266 622658 369502 622894
rect 369586 622658 369822 622894
rect 369266 622338 369502 622574
rect 369586 622338 369822 622574
rect 369266 586658 369502 586894
rect 369586 586658 369822 586894
rect 369266 586338 369502 586574
rect 369586 586338 369822 586574
rect 369266 550658 369502 550894
rect 369586 550658 369822 550894
rect 369266 550338 369502 550574
rect 369586 550338 369822 550574
rect 369266 514658 369502 514894
rect 369586 514658 369822 514894
rect 369266 514338 369502 514574
rect 369586 514338 369822 514574
rect 369266 478658 369502 478894
rect 369586 478658 369822 478894
rect 369266 478338 369502 478574
rect 369586 478338 369822 478574
rect 369266 442658 369502 442894
rect 369586 442658 369822 442894
rect 369266 442338 369502 442574
rect 369586 442338 369822 442574
rect 369266 406658 369502 406894
rect 369586 406658 369822 406894
rect 369266 406338 369502 406574
rect 369586 406338 369822 406574
rect 369266 370658 369502 370894
rect 369586 370658 369822 370894
rect 369266 370338 369502 370574
rect 369586 370338 369822 370574
rect 369266 334658 369502 334894
rect 369586 334658 369822 334894
rect 369266 334338 369502 334574
rect 369586 334338 369822 334574
rect 369266 298658 369502 298894
rect 369586 298658 369822 298894
rect 369266 298338 369502 298574
rect 369586 298338 369822 298574
rect 369266 262658 369502 262894
rect 369586 262658 369822 262894
rect 369266 262338 369502 262574
rect 369586 262338 369822 262574
rect 369266 226658 369502 226894
rect 369586 226658 369822 226894
rect 369266 226338 369502 226574
rect 369586 226338 369822 226574
rect 369266 190658 369502 190894
rect 369586 190658 369822 190894
rect 369266 190338 369502 190574
rect 369586 190338 369822 190574
rect 369266 154658 369502 154894
rect 369586 154658 369822 154894
rect 369266 154338 369502 154574
rect 369586 154338 369822 154574
rect 369266 118658 369502 118894
rect 369586 118658 369822 118894
rect 369266 118338 369502 118574
rect 369586 118338 369822 118574
rect 369266 82658 369502 82894
rect 369586 82658 369822 82894
rect 369266 82338 369502 82574
rect 369586 82338 369822 82574
rect 369266 46658 369502 46894
rect 369586 46658 369822 46894
rect 369266 46338 369502 46574
rect 369586 46338 369822 46574
rect 369266 10658 369502 10894
rect 369586 10658 369822 10894
rect 369266 10338 369502 10574
rect 369586 10338 369822 10574
rect 369266 -4422 369502 -4186
rect 369586 -4422 369822 -4186
rect 369266 -4742 369502 -4506
rect 369586 -4742 369822 -4506
rect 390986 711322 391222 711558
rect 391306 711322 391542 711558
rect 390986 711002 391222 711238
rect 391306 711002 391542 711238
rect 387266 709402 387502 709638
rect 387586 709402 387822 709638
rect 387266 709082 387502 709318
rect 387586 709082 387822 709318
rect 383546 707482 383782 707718
rect 383866 707482 384102 707718
rect 383546 707162 383782 707398
rect 383866 707162 384102 707398
rect 372986 698378 373222 698614
rect 373306 698378 373542 698614
rect 372986 698058 373222 698294
rect 373306 698058 373542 698294
rect 372986 662378 373222 662614
rect 373306 662378 373542 662614
rect 372986 662058 373222 662294
rect 373306 662058 373542 662294
rect 372986 626378 373222 626614
rect 373306 626378 373542 626614
rect 372986 626058 373222 626294
rect 373306 626058 373542 626294
rect 372986 590378 373222 590614
rect 373306 590378 373542 590614
rect 372986 590058 373222 590294
rect 373306 590058 373542 590294
rect 372986 554378 373222 554614
rect 373306 554378 373542 554614
rect 372986 554058 373222 554294
rect 373306 554058 373542 554294
rect 372986 518378 373222 518614
rect 373306 518378 373542 518614
rect 372986 518058 373222 518294
rect 373306 518058 373542 518294
rect 372986 482378 373222 482614
rect 373306 482378 373542 482614
rect 372986 482058 373222 482294
rect 373306 482058 373542 482294
rect 372986 446378 373222 446614
rect 373306 446378 373542 446614
rect 372986 446058 373222 446294
rect 373306 446058 373542 446294
rect 372986 410378 373222 410614
rect 373306 410378 373542 410614
rect 372986 410058 373222 410294
rect 373306 410058 373542 410294
rect 372986 374378 373222 374614
rect 373306 374378 373542 374614
rect 372986 374058 373222 374294
rect 373306 374058 373542 374294
rect 372986 338378 373222 338614
rect 373306 338378 373542 338614
rect 372986 338058 373222 338294
rect 373306 338058 373542 338294
rect 372986 302378 373222 302614
rect 373306 302378 373542 302614
rect 372986 302058 373222 302294
rect 373306 302058 373542 302294
rect 372986 266378 373222 266614
rect 373306 266378 373542 266614
rect 372986 266058 373222 266294
rect 373306 266058 373542 266294
rect 372986 230378 373222 230614
rect 373306 230378 373542 230614
rect 372986 230058 373222 230294
rect 373306 230058 373542 230294
rect 372986 194378 373222 194614
rect 373306 194378 373542 194614
rect 372986 194058 373222 194294
rect 373306 194058 373542 194294
rect 372986 158378 373222 158614
rect 373306 158378 373542 158614
rect 372986 158058 373222 158294
rect 373306 158058 373542 158294
rect 372986 122378 373222 122614
rect 373306 122378 373542 122614
rect 372986 122058 373222 122294
rect 373306 122058 373542 122294
rect 372986 86378 373222 86614
rect 373306 86378 373542 86614
rect 372986 86058 373222 86294
rect 373306 86058 373542 86294
rect 372986 50378 373222 50614
rect 373306 50378 373542 50614
rect 372986 50058 373222 50294
rect 373306 50058 373542 50294
rect 372986 14378 373222 14614
rect 373306 14378 373542 14614
rect 372986 14058 373222 14294
rect 373306 14058 373542 14294
rect 354986 -7302 355222 -7066
rect 355306 -7302 355542 -7066
rect 354986 -7622 355222 -7386
rect 355306 -7622 355542 -7386
rect 379826 705562 380062 705798
rect 380146 705562 380382 705798
rect 379826 705242 380062 705478
rect 380146 705242 380382 705478
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 379826 633218 380062 633454
rect 380146 633218 380382 633454
rect 379826 632898 380062 633134
rect 380146 632898 380382 633134
rect 379826 597218 380062 597454
rect 380146 597218 380382 597454
rect 379826 596898 380062 597134
rect 380146 596898 380382 597134
rect 379826 561218 380062 561454
rect 380146 561218 380382 561454
rect 379826 560898 380062 561134
rect 380146 560898 380382 561134
rect 379826 525218 380062 525454
rect 380146 525218 380382 525454
rect 379826 524898 380062 525134
rect 380146 524898 380382 525134
rect 379826 489218 380062 489454
rect 380146 489218 380382 489454
rect 379826 488898 380062 489134
rect 380146 488898 380382 489134
rect 379826 453218 380062 453454
rect 380146 453218 380382 453454
rect 379826 452898 380062 453134
rect 380146 452898 380382 453134
rect 379826 417218 380062 417454
rect 380146 417218 380382 417454
rect 379826 416898 380062 417134
rect 380146 416898 380382 417134
rect 379826 381218 380062 381454
rect 380146 381218 380382 381454
rect 379826 380898 380062 381134
rect 380146 380898 380382 381134
rect 379826 345218 380062 345454
rect 380146 345218 380382 345454
rect 379826 344898 380062 345134
rect 380146 344898 380382 345134
rect 379826 309218 380062 309454
rect 380146 309218 380382 309454
rect 379826 308898 380062 309134
rect 380146 308898 380382 309134
rect 379826 273218 380062 273454
rect 380146 273218 380382 273454
rect 379826 272898 380062 273134
rect 380146 272898 380382 273134
rect 379826 237218 380062 237454
rect 380146 237218 380382 237454
rect 379826 236898 380062 237134
rect 380146 236898 380382 237134
rect 379826 201218 380062 201454
rect 380146 201218 380382 201454
rect 379826 200898 380062 201134
rect 380146 200898 380382 201134
rect 379826 165218 380062 165454
rect 380146 165218 380382 165454
rect 379826 164898 380062 165134
rect 380146 164898 380382 165134
rect 379826 129218 380062 129454
rect 380146 129218 380382 129454
rect 379826 128898 380062 129134
rect 380146 128898 380382 129134
rect 379826 93218 380062 93454
rect 380146 93218 380382 93454
rect 379826 92898 380062 93134
rect 380146 92898 380382 93134
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -1542 380062 -1306
rect 380146 -1542 380382 -1306
rect 379826 -1862 380062 -1626
rect 380146 -1862 380382 -1626
rect 383546 672938 383782 673174
rect 383866 672938 384102 673174
rect 383546 672618 383782 672854
rect 383866 672618 384102 672854
rect 383546 636938 383782 637174
rect 383866 636938 384102 637174
rect 383546 636618 383782 636854
rect 383866 636618 384102 636854
rect 383546 600938 383782 601174
rect 383866 600938 384102 601174
rect 383546 600618 383782 600854
rect 383866 600618 384102 600854
rect 383546 564938 383782 565174
rect 383866 564938 384102 565174
rect 383546 564618 383782 564854
rect 383866 564618 384102 564854
rect 383546 528938 383782 529174
rect 383866 528938 384102 529174
rect 383546 528618 383782 528854
rect 383866 528618 384102 528854
rect 383546 492938 383782 493174
rect 383866 492938 384102 493174
rect 383546 492618 383782 492854
rect 383866 492618 384102 492854
rect 383546 456938 383782 457174
rect 383866 456938 384102 457174
rect 383546 456618 383782 456854
rect 383866 456618 384102 456854
rect 383546 420938 383782 421174
rect 383866 420938 384102 421174
rect 383546 420618 383782 420854
rect 383866 420618 384102 420854
rect 383546 384938 383782 385174
rect 383866 384938 384102 385174
rect 383546 384618 383782 384854
rect 383866 384618 384102 384854
rect 383546 348938 383782 349174
rect 383866 348938 384102 349174
rect 383546 348618 383782 348854
rect 383866 348618 384102 348854
rect 383546 312938 383782 313174
rect 383866 312938 384102 313174
rect 383546 312618 383782 312854
rect 383866 312618 384102 312854
rect 383546 276938 383782 277174
rect 383866 276938 384102 277174
rect 383546 276618 383782 276854
rect 383866 276618 384102 276854
rect 383546 240938 383782 241174
rect 383866 240938 384102 241174
rect 383546 240618 383782 240854
rect 383866 240618 384102 240854
rect 383546 204938 383782 205174
rect 383866 204938 384102 205174
rect 383546 204618 383782 204854
rect 383866 204618 384102 204854
rect 383546 168938 383782 169174
rect 383866 168938 384102 169174
rect 383546 168618 383782 168854
rect 383866 168618 384102 168854
rect 383546 132938 383782 133174
rect 383866 132938 384102 133174
rect 383546 132618 383782 132854
rect 383866 132618 384102 132854
rect 383546 96938 383782 97174
rect 383866 96938 384102 97174
rect 383546 96618 383782 96854
rect 383866 96618 384102 96854
rect 383546 60938 383782 61174
rect 383866 60938 384102 61174
rect 383546 60618 383782 60854
rect 383866 60618 384102 60854
rect 383546 24938 383782 25174
rect 383866 24938 384102 25174
rect 383546 24618 383782 24854
rect 383866 24618 384102 24854
rect 383546 -3462 383782 -3226
rect 383866 -3462 384102 -3226
rect 383546 -3782 383782 -3546
rect 383866 -3782 384102 -3546
rect 387266 676658 387502 676894
rect 387586 676658 387822 676894
rect 387266 676338 387502 676574
rect 387586 676338 387822 676574
rect 387266 640658 387502 640894
rect 387586 640658 387822 640894
rect 387266 640338 387502 640574
rect 387586 640338 387822 640574
rect 387266 604658 387502 604894
rect 387586 604658 387822 604894
rect 387266 604338 387502 604574
rect 387586 604338 387822 604574
rect 387266 568658 387502 568894
rect 387586 568658 387822 568894
rect 387266 568338 387502 568574
rect 387586 568338 387822 568574
rect 387266 532658 387502 532894
rect 387586 532658 387822 532894
rect 387266 532338 387502 532574
rect 387586 532338 387822 532574
rect 387266 496658 387502 496894
rect 387586 496658 387822 496894
rect 387266 496338 387502 496574
rect 387586 496338 387822 496574
rect 387266 460658 387502 460894
rect 387586 460658 387822 460894
rect 387266 460338 387502 460574
rect 387586 460338 387822 460574
rect 387266 424658 387502 424894
rect 387586 424658 387822 424894
rect 387266 424338 387502 424574
rect 387586 424338 387822 424574
rect 387266 388658 387502 388894
rect 387586 388658 387822 388894
rect 387266 388338 387502 388574
rect 387586 388338 387822 388574
rect 387266 352658 387502 352894
rect 387586 352658 387822 352894
rect 387266 352338 387502 352574
rect 387586 352338 387822 352574
rect 387266 316658 387502 316894
rect 387586 316658 387822 316894
rect 387266 316338 387502 316574
rect 387586 316338 387822 316574
rect 387266 280658 387502 280894
rect 387586 280658 387822 280894
rect 387266 280338 387502 280574
rect 387586 280338 387822 280574
rect 387266 244658 387502 244894
rect 387586 244658 387822 244894
rect 387266 244338 387502 244574
rect 387586 244338 387822 244574
rect 387266 208658 387502 208894
rect 387586 208658 387822 208894
rect 387266 208338 387502 208574
rect 387586 208338 387822 208574
rect 387266 172658 387502 172894
rect 387586 172658 387822 172894
rect 387266 172338 387502 172574
rect 387586 172338 387822 172574
rect 387266 136658 387502 136894
rect 387586 136658 387822 136894
rect 387266 136338 387502 136574
rect 387586 136338 387822 136574
rect 387266 100658 387502 100894
rect 387586 100658 387822 100894
rect 387266 100338 387502 100574
rect 387586 100338 387822 100574
rect 387266 64658 387502 64894
rect 387586 64658 387822 64894
rect 387266 64338 387502 64574
rect 387586 64338 387822 64574
rect 387266 28658 387502 28894
rect 387586 28658 387822 28894
rect 387266 28338 387502 28574
rect 387586 28338 387822 28574
rect 387266 -5382 387502 -5146
rect 387586 -5382 387822 -5146
rect 387266 -5702 387502 -5466
rect 387586 -5702 387822 -5466
rect 408986 710362 409222 710598
rect 409306 710362 409542 710598
rect 408986 710042 409222 710278
rect 409306 710042 409542 710278
rect 405266 708442 405502 708678
rect 405586 708442 405822 708678
rect 405266 708122 405502 708358
rect 405586 708122 405822 708358
rect 401546 706522 401782 706758
rect 401866 706522 402102 706758
rect 401546 706202 401782 706438
rect 401866 706202 402102 706438
rect 390986 680378 391222 680614
rect 391306 680378 391542 680614
rect 390986 680058 391222 680294
rect 391306 680058 391542 680294
rect 390986 644378 391222 644614
rect 391306 644378 391542 644614
rect 390986 644058 391222 644294
rect 391306 644058 391542 644294
rect 390986 608378 391222 608614
rect 391306 608378 391542 608614
rect 390986 608058 391222 608294
rect 391306 608058 391542 608294
rect 390986 572378 391222 572614
rect 391306 572378 391542 572614
rect 390986 572058 391222 572294
rect 391306 572058 391542 572294
rect 390986 536378 391222 536614
rect 391306 536378 391542 536614
rect 390986 536058 391222 536294
rect 391306 536058 391542 536294
rect 390986 500378 391222 500614
rect 391306 500378 391542 500614
rect 390986 500058 391222 500294
rect 391306 500058 391542 500294
rect 390986 464378 391222 464614
rect 391306 464378 391542 464614
rect 390986 464058 391222 464294
rect 391306 464058 391542 464294
rect 390986 428378 391222 428614
rect 391306 428378 391542 428614
rect 390986 428058 391222 428294
rect 391306 428058 391542 428294
rect 390986 392378 391222 392614
rect 391306 392378 391542 392614
rect 390986 392058 391222 392294
rect 391306 392058 391542 392294
rect 390986 356378 391222 356614
rect 391306 356378 391542 356614
rect 390986 356058 391222 356294
rect 391306 356058 391542 356294
rect 390986 320378 391222 320614
rect 391306 320378 391542 320614
rect 390986 320058 391222 320294
rect 391306 320058 391542 320294
rect 390986 284378 391222 284614
rect 391306 284378 391542 284614
rect 390986 284058 391222 284294
rect 391306 284058 391542 284294
rect 390986 248378 391222 248614
rect 391306 248378 391542 248614
rect 390986 248058 391222 248294
rect 391306 248058 391542 248294
rect 390986 212378 391222 212614
rect 391306 212378 391542 212614
rect 390986 212058 391222 212294
rect 391306 212058 391542 212294
rect 390986 176378 391222 176614
rect 391306 176378 391542 176614
rect 390986 176058 391222 176294
rect 391306 176058 391542 176294
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 397826 543218 398062 543454
rect 398146 543218 398382 543454
rect 397826 542898 398062 543134
rect 398146 542898 398382 543134
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 397826 435218 398062 435454
rect 398146 435218 398382 435454
rect 397826 434898 398062 435134
rect 398146 434898 398382 435134
rect 397826 399218 398062 399454
rect 398146 399218 398382 399454
rect 397826 398898 398062 399134
rect 398146 398898 398382 399134
rect 401546 690938 401782 691174
rect 401866 690938 402102 691174
rect 401546 690618 401782 690854
rect 401866 690618 402102 690854
rect 401546 654938 401782 655174
rect 401866 654938 402102 655174
rect 401546 654618 401782 654854
rect 401866 654618 402102 654854
rect 401546 618938 401782 619174
rect 401866 618938 402102 619174
rect 401546 618618 401782 618854
rect 401866 618618 402102 618854
rect 401546 582938 401782 583174
rect 401866 582938 402102 583174
rect 401546 582618 401782 582854
rect 401866 582618 402102 582854
rect 401546 546938 401782 547174
rect 401866 546938 402102 547174
rect 401546 546618 401782 546854
rect 401866 546618 402102 546854
rect 401546 510938 401782 511174
rect 401866 510938 402102 511174
rect 401546 510618 401782 510854
rect 401866 510618 402102 510854
rect 401546 474938 401782 475174
rect 401866 474938 402102 475174
rect 401546 474618 401782 474854
rect 401866 474618 402102 474854
rect 401546 438938 401782 439174
rect 401866 438938 402102 439174
rect 401546 438618 401782 438854
rect 401866 438618 402102 438854
rect 401546 402938 401782 403174
rect 401866 402938 402102 403174
rect 401546 402618 401782 402854
rect 401866 402618 402102 402854
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 397826 327218 398062 327454
rect 398146 327218 398382 327454
rect 397826 326898 398062 327134
rect 398146 326898 398382 327134
rect 397826 291218 398062 291454
rect 398146 291218 398382 291454
rect 397826 290898 398062 291134
rect 398146 290898 398382 291134
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 397826 219218 398062 219454
rect 398146 219218 398382 219454
rect 397826 218898 398062 219134
rect 398146 218898 398382 219134
rect 397826 183218 398062 183454
rect 398146 183218 398382 183454
rect 397826 182898 398062 183134
rect 398146 182898 398382 183134
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 390986 140378 391222 140614
rect 391306 140378 391542 140614
rect 390986 140058 391222 140294
rect 391306 140058 391542 140294
rect 401546 366938 401782 367174
rect 401866 366938 402102 367174
rect 401546 366618 401782 366854
rect 401866 366618 402102 366854
rect 401546 330938 401782 331174
rect 401866 330938 402102 331174
rect 401546 330618 401782 330854
rect 401866 330618 402102 330854
rect 401546 294938 401782 295174
rect 401866 294938 402102 295174
rect 401546 294618 401782 294854
rect 401866 294618 402102 294854
rect 401546 258938 401782 259174
rect 401866 258938 402102 259174
rect 401546 258618 401782 258854
rect 401866 258618 402102 258854
rect 401546 222938 401782 223174
rect 401866 222938 402102 223174
rect 401546 222618 401782 222854
rect 401866 222618 402102 222854
rect 401546 186938 401782 187174
rect 401866 186938 402102 187174
rect 401546 186618 401782 186854
rect 401866 186618 402102 186854
rect 401546 150938 401782 151174
rect 401866 150938 402102 151174
rect 401546 150618 401782 150854
rect 401866 150618 402102 150854
rect 405266 694658 405502 694894
rect 405586 694658 405822 694894
rect 405266 694338 405502 694574
rect 405586 694338 405822 694574
rect 405266 658658 405502 658894
rect 405586 658658 405822 658894
rect 405266 658338 405502 658574
rect 405586 658338 405822 658574
rect 405266 622658 405502 622894
rect 405586 622658 405822 622894
rect 405266 622338 405502 622574
rect 405586 622338 405822 622574
rect 405266 586658 405502 586894
rect 405586 586658 405822 586894
rect 405266 586338 405502 586574
rect 405586 586338 405822 586574
rect 405266 550658 405502 550894
rect 405586 550658 405822 550894
rect 405266 550338 405502 550574
rect 405586 550338 405822 550574
rect 405266 514658 405502 514894
rect 405586 514658 405822 514894
rect 405266 514338 405502 514574
rect 405586 514338 405822 514574
rect 405266 478658 405502 478894
rect 405586 478658 405822 478894
rect 405266 478338 405502 478574
rect 405586 478338 405822 478574
rect 405266 442658 405502 442894
rect 405586 442658 405822 442894
rect 405266 442338 405502 442574
rect 405586 442338 405822 442574
rect 405266 406658 405502 406894
rect 405586 406658 405822 406894
rect 405266 406338 405502 406574
rect 405586 406338 405822 406574
rect 405266 370658 405502 370894
rect 405586 370658 405822 370894
rect 405266 370338 405502 370574
rect 405586 370338 405822 370574
rect 405266 334658 405502 334894
rect 405586 334658 405822 334894
rect 405266 334338 405502 334574
rect 405586 334338 405822 334574
rect 405266 298658 405502 298894
rect 405586 298658 405822 298894
rect 405266 298338 405502 298574
rect 405586 298338 405822 298574
rect 405266 262658 405502 262894
rect 405586 262658 405822 262894
rect 405266 262338 405502 262574
rect 405586 262338 405822 262574
rect 405266 226658 405502 226894
rect 405586 226658 405822 226894
rect 405266 226338 405502 226574
rect 405586 226338 405822 226574
rect 405266 190658 405502 190894
rect 405586 190658 405822 190894
rect 405266 190338 405502 190574
rect 405586 190338 405822 190574
rect 405266 154658 405502 154894
rect 405586 154658 405822 154894
rect 405266 154338 405502 154574
rect 405586 154338 405822 154574
rect 426986 711322 427222 711558
rect 427306 711322 427542 711558
rect 426986 711002 427222 711238
rect 427306 711002 427542 711238
rect 423266 709402 423502 709638
rect 423586 709402 423822 709638
rect 423266 709082 423502 709318
rect 423586 709082 423822 709318
rect 419546 707482 419782 707718
rect 419866 707482 420102 707718
rect 419546 707162 419782 707398
rect 419866 707162 420102 707398
rect 408986 698378 409222 698614
rect 409306 698378 409542 698614
rect 408986 698058 409222 698294
rect 409306 698058 409542 698294
rect 408986 662378 409222 662614
rect 409306 662378 409542 662614
rect 408986 662058 409222 662294
rect 409306 662058 409542 662294
rect 408986 626378 409222 626614
rect 409306 626378 409542 626614
rect 408986 626058 409222 626294
rect 409306 626058 409542 626294
rect 408986 590378 409222 590614
rect 409306 590378 409542 590614
rect 408986 590058 409222 590294
rect 409306 590058 409542 590294
rect 408986 554378 409222 554614
rect 409306 554378 409542 554614
rect 408986 554058 409222 554294
rect 409306 554058 409542 554294
rect 408986 518378 409222 518614
rect 409306 518378 409542 518614
rect 408986 518058 409222 518294
rect 409306 518058 409542 518294
rect 408986 482378 409222 482614
rect 409306 482378 409542 482614
rect 408986 482058 409222 482294
rect 409306 482058 409542 482294
rect 408986 446378 409222 446614
rect 409306 446378 409542 446614
rect 408986 446058 409222 446294
rect 409306 446058 409542 446294
rect 408986 410378 409222 410614
rect 409306 410378 409542 410614
rect 408986 410058 409222 410294
rect 409306 410058 409542 410294
rect 408986 374378 409222 374614
rect 409306 374378 409542 374614
rect 408986 374058 409222 374294
rect 409306 374058 409542 374294
rect 408986 338378 409222 338614
rect 409306 338378 409542 338614
rect 408986 338058 409222 338294
rect 409306 338058 409542 338294
rect 408986 302378 409222 302614
rect 409306 302378 409542 302614
rect 408986 302058 409222 302294
rect 409306 302058 409542 302294
rect 408986 266378 409222 266614
rect 409306 266378 409542 266614
rect 408986 266058 409222 266294
rect 409306 266058 409542 266294
rect 408986 230378 409222 230614
rect 409306 230378 409542 230614
rect 408986 230058 409222 230294
rect 409306 230058 409542 230294
rect 408986 194378 409222 194614
rect 409306 194378 409542 194614
rect 408986 194058 409222 194294
rect 409306 194058 409542 194294
rect 408986 158378 409222 158614
rect 409306 158378 409542 158614
rect 408986 158058 409222 158294
rect 409306 158058 409542 158294
rect 415826 705562 416062 705798
rect 416146 705562 416382 705798
rect 415826 705242 416062 705478
rect 416146 705242 416382 705478
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 415826 633218 416062 633454
rect 416146 633218 416382 633454
rect 415826 632898 416062 633134
rect 416146 632898 416382 633134
rect 415826 597218 416062 597454
rect 416146 597218 416382 597454
rect 415826 596898 416062 597134
rect 416146 596898 416382 597134
rect 415826 561218 416062 561454
rect 416146 561218 416382 561454
rect 415826 560898 416062 561134
rect 416146 560898 416382 561134
rect 415826 525218 416062 525454
rect 416146 525218 416382 525454
rect 415826 524898 416062 525134
rect 416146 524898 416382 525134
rect 415826 489218 416062 489454
rect 416146 489218 416382 489454
rect 415826 488898 416062 489134
rect 416146 488898 416382 489134
rect 415826 453218 416062 453454
rect 416146 453218 416382 453454
rect 415826 452898 416062 453134
rect 416146 452898 416382 453134
rect 415826 417218 416062 417454
rect 416146 417218 416382 417454
rect 415826 416898 416062 417134
rect 416146 416898 416382 417134
rect 415826 381218 416062 381454
rect 416146 381218 416382 381454
rect 415826 380898 416062 381134
rect 416146 380898 416382 381134
rect 415826 345218 416062 345454
rect 416146 345218 416382 345454
rect 415826 344898 416062 345134
rect 416146 344898 416382 345134
rect 415826 309218 416062 309454
rect 416146 309218 416382 309454
rect 415826 308898 416062 309134
rect 416146 308898 416382 309134
rect 415826 273218 416062 273454
rect 416146 273218 416382 273454
rect 415826 272898 416062 273134
rect 416146 272898 416382 273134
rect 415826 237218 416062 237454
rect 416146 237218 416382 237454
rect 415826 236898 416062 237134
rect 416146 236898 416382 237134
rect 415826 201218 416062 201454
rect 416146 201218 416382 201454
rect 415826 200898 416062 201134
rect 416146 200898 416382 201134
rect 415826 165218 416062 165454
rect 416146 165218 416382 165454
rect 415826 164898 416062 165134
rect 416146 164898 416382 165134
rect 402586 129218 402822 129454
rect 402586 128898 402822 129134
rect 405786 129218 406022 129454
rect 405786 128898 406022 129134
rect 408986 129218 409222 129454
rect 408986 128898 409222 129134
rect 404186 111218 404422 111454
rect 404186 110898 404422 111134
rect 407386 111218 407622 111454
rect 407386 110898 407622 111134
rect 390986 104378 391222 104614
rect 391306 104378 391542 104614
rect 390986 104058 391222 104294
rect 391306 104058 391542 104294
rect 390986 68378 391222 68614
rect 391306 68378 391542 68614
rect 390986 68058 391222 68294
rect 391306 68058 391542 68294
rect 390986 32378 391222 32614
rect 391306 32378 391542 32614
rect 390986 32058 391222 32294
rect 391306 32058 391542 32294
rect 372986 -6342 373222 -6106
rect 373306 -6342 373542 -6106
rect 372986 -6662 373222 -6426
rect 373306 -6662 373542 -6426
rect 397826 75218 398062 75454
rect 398146 75218 398382 75454
rect 397826 74898 398062 75134
rect 398146 74898 398382 75134
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 401546 78938 401782 79174
rect 401866 78938 402102 79174
rect 401546 78618 401782 78854
rect 401866 78618 402102 78854
rect 401546 42938 401782 43174
rect 401866 42938 402102 43174
rect 401546 42618 401782 42854
rect 401866 42618 402102 42854
rect 401546 6938 401782 7174
rect 401866 6938 402102 7174
rect 401546 6618 401782 6854
rect 401866 6618 402102 6854
rect 401546 -2502 401782 -2266
rect 401866 -2502 402102 -2266
rect 401546 -2822 401782 -2586
rect 401866 -2822 402102 -2586
rect 405266 82658 405502 82894
rect 405586 82658 405822 82894
rect 405266 82338 405502 82574
rect 405586 82338 405822 82574
rect 405266 46658 405502 46894
rect 405586 46658 405822 46894
rect 405266 46338 405502 46574
rect 405586 46338 405822 46574
rect 405266 10658 405502 10894
rect 405586 10658 405822 10894
rect 405266 10338 405502 10574
rect 405586 10338 405822 10574
rect 405266 -4422 405502 -4186
rect 405586 -4422 405822 -4186
rect 405266 -4742 405502 -4506
rect 405586 -4742 405822 -4506
rect 408986 86378 409222 86614
rect 409306 86378 409542 86614
rect 408986 86058 409222 86294
rect 409306 86058 409542 86294
rect 419546 672938 419782 673174
rect 419866 672938 420102 673174
rect 419546 672618 419782 672854
rect 419866 672618 420102 672854
rect 419546 636938 419782 637174
rect 419866 636938 420102 637174
rect 419546 636618 419782 636854
rect 419866 636618 420102 636854
rect 419546 600938 419782 601174
rect 419866 600938 420102 601174
rect 419546 600618 419782 600854
rect 419866 600618 420102 600854
rect 419546 564938 419782 565174
rect 419866 564938 420102 565174
rect 419546 564618 419782 564854
rect 419866 564618 420102 564854
rect 419546 528938 419782 529174
rect 419866 528938 420102 529174
rect 419546 528618 419782 528854
rect 419866 528618 420102 528854
rect 419546 492938 419782 493174
rect 419866 492938 420102 493174
rect 419546 492618 419782 492854
rect 419866 492618 420102 492854
rect 419546 456938 419782 457174
rect 419866 456938 420102 457174
rect 419546 456618 419782 456854
rect 419866 456618 420102 456854
rect 419546 420938 419782 421174
rect 419866 420938 420102 421174
rect 419546 420618 419782 420854
rect 419866 420618 420102 420854
rect 419546 384938 419782 385174
rect 419866 384938 420102 385174
rect 419546 384618 419782 384854
rect 419866 384618 420102 384854
rect 419546 348938 419782 349174
rect 419866 348938 420102 349174
rect 419546 348618 419782 348854
rect 419866 348618 420102 348854
rect 419546 312938 419782 313174
rect 419866 312938 420102 313174
rect 419546 312618 419782 312854
rect 419866 312618 420102 312854
rect 419546 276938 419782 277174
rect 419866 276938 420102 277174
rect 419546 276618 419782 276854
rect 419866 276618 420102 276854
rect 419546 240938 419782 241174
rect 419866 240938 420102 241174
rect 419546 240618 419782 240854
rect 419866 240618 420102 240854
rect 419546 204938 419782 205174
rect 419866 204938 420102 205174
rect 419546 204618 419782 204854
rect 419866 204618 420102 204854
rect 419546 168938 419782 169174
rect 419866 168938 420102 169174
rect 419546 168618 419782 168854
rect 419866 168618 420102 168854
rect 412186 129218 412422 129454
rect 412186 128898 412422 129134
rect 415386 129218 415622 129454
rect 415386 128898 415622 129134
rect 410586 111218 410822 111454
rect 410586 110898 410822 111134
rect 413786 111218 414022 111454
rect 413786 110898 414022 111134
rect 416986 111218 417222 111454
rect 416986 110898 417222 111134
rect 415826 93218 416062 93454
rect 416146 93218 416382 93454
rect 415826 92898 416062 93134
rect 416146 92898 416382 93134
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 408986 50378 409222 50614
rect 409306 50378 409542 50614
rect 408986 50058 409222 50294
rect 409306 50058 409542 50294
rect 408986 14378 409222 14614
rect 409306 14378 409542 14614
rect 408986 14058 409222 14294
rect 409306 14058 409542 14294
rect 390986 -7302 391222 -7066
rect 391306 -7302 391542 -7066
rect 390986 -7622 391222 -7386
rect 391306 -7622 391542 -7386
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 423266 676658 423502 676894
rect 423586 676658 423822 676894
rect 423266 676338 423502 676574
rect 423586 676338 423822 676574
rect 423266 640658 423502 640894
rect 423586 640658 423822 640894
rect 423266 640338 423502 640574
rect 423586 640338 423822 640574
rect 423266 604658 423502 604894
rect 423586 604658 423822 604894
rect 423266 604338 423502 604574
rect 423586 604338 423822 604574
rect 423266 568658 423502 568894
rect 423586 568658 423822 568894
rect 423266 568338 423502 568574
rect 423586 568338 423822 568574
rect 423266 532658 423502 532894
rect 423586 532658 423822 532894
rect 423266 532338 423502 532574
rect 423586 532338 423822 532574
rect 423266 496658 423502 496894
rect 423586 496658 423822 496894
rect 423266 496338 423502 496574
rect 423586 496338 423822 496574
rect 423266 460658 423502 460894
rect 423586 460658 423822 460894
rect 423266 460338 423502 460574
rect 423586 460338 423822 460574
rect 423266 424658 423502 424894
rect 423586 424658 423822 424894
rect 423266 424338 423502 424574
rect 423586 424338 423822 424574
rect 423266 388658 423502 388894
rect 423586 388658 423822 388894
rect 423266 388338 423502 388574
rect 423586 388338 423822 388574
rect 423266 352658 423502 352894
rect 423586 352658 423822 352894
rect 423266 352338 423502 352574
rect 423586 352338 423822 352574
rect 423266 316658 423502 316894
rect 423586 316658 423822 316894
rect 423266 316338 423502 316574
rect 423586 316338 423822 316574
rect 444986 710362 445222 710598
rect 445306 710362 445542 710598
rect 444986 710042 445222 710278
rect 445306 710042 445542 710278
rect 441266 708442 441502 708678
rect 441586 708442 441822 708678
rect 441266 708122 441502 708358
rect 441586 708122 441822 708358
rect 437546 706522 437782 706758
rect 437866 706522 438102 706758
rect 437546 706202 437782 706438
rect 437866 706202 438102 706438
rect 426986 680378 427222 680614
rect 427306 680378 427542 680614
rect 426986 680058 427222 680294
rect 427306 680058 427542 680294
rect 426986 644378 427222 644614
rect 427306 644378 427542 644614
rect 426986 644058 427222 644294
rect 427306 644058 427542 644294
rect 426986 608378 427222 608614
rect 427306 608378 427542 608614
rect 426986 608058 427222 608294
rect 427306 608058 427542 608294
rect 426986 572378 427222 572614
rect 427306 572378 427542 572614
rect 426986 572058 427222 572294
rect 427306 572058 427542 572294
rect 426986 536378 427222 536614
rect 427306 536378 427542 536614
rect 426986 536058 427222 536294
rect 427306 536058 427542 536294
rect 426986 500378 427222 500614
rect 427306 500378 427542 500614
rect 426986 500058 427222 500294
rect 427306 500058 427542 500294
rect 426986 464378 427222 464614
rect 427306 464378 427542 464614
rect 426986 464058 427222 464294
rect 427306 464058 427542 464294
rect 426986 428378 427222 428614
rect 427306 428378 427542 428614
rect 426986 428058 427222 428294
rect 427306 428058 427542 428294
rect 426986 392378 427222 392614
rect 427306 392378 427542 392614
rect 426986 392058 427222 392294
rect 427306 392058 427542 392294
rect 426986 356378 427222 356614
rect 427306 356378 427542 356614
rect 426986 356058 427222 356294
rect 427306 356058 427542 356294
rect 426986 320378 427222 320614
rect 427306 320378 427542 320614
rect 426986 320058 427222 320294
rect 427306 320058 427542 320294
rect 423266 280658 423502 280894
rect 423586 280658 423822 280894
rect 423266 280338 423502 280574
rect 423586 280338 423822 280574
rect 423266 244658 423502 244894
rect 423586 244658 423822 244894
rect 423266 244338 423502 244574
rect 423586 244338 423822 244574
rect 423266 208658 423502 208894
rect 423586 208658 423822 208894
rect 423266 208338 423502 208574
rect 423586 208338 423822 208574
rect 423266 172658 423502 172894
rect 423586 172658 423822 172894
rect 423266 172338 423502 172574
rect 423586 172338 423822 172574
rect 418586 129218 418822 129454
rect 418586 128898 418822 129134
rect 420186 111218 420422 111454
rect 420186 110898 420422 111134
rect 419546 96938 419782 97174
rect 419866 96938 420102 97174
rect 419546 96618 419782 96854
rect 419866 96618 420102 96854
rect 421786 129218 422022 129454
rect 421786 128898 422022 129134
rect 423386 111218 423622 111454
rect 423386 110898 423622 111134
rect 424986 129218 425222 129454
rect 424986 128898 425222 129134
rect 426986 284378 427222 284614
rect 427306 284378 427542 284614
rect 426986 284058 427222 284294
rect 427306 284058 427542 284294
rect 426986 248378 427222 248614
rect 427306 248378 427542 248614
rect 426986 248058 427222 248294
rect 427306 248058 427542 248294
rect 426986 212378 427222 212614
rect 427306 212378 427542 212614
rect 426986 212058 427222 212294
rect 427306 212058 427542 212294
rect 426986 176378 427222 176614
rect 427306 176378 427542 176614
rect 426986 176058 427222 176294
rect 427306 176058 427542 176294
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 433826 435218 434062 435454
rect 434146 435218 434382 435454
rect 433826 434898 434062 435134
rect 434146 434898 434382 435134
rect 433826 399218 434062 399454
rect 434146 399218 434382 399454
rect 433826 398898 434062 399134
rect 434146 398898 434382 399134
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 433826 291218 434062 291454
rect 434146 291218 434382 291454
rect 433826 290898 434062 291134
rect 434146 290898 434382 291134
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 433826 219218 434062 219454
rect 434146 219218 434382 219454
rect 433826 218898 434062 219134
rect 434146 218898 434382 219134
rect 433826 183218 434062 183454
rect 434146 183218 434382 183454
rect 433826 182898 434062 183134
rect 434146 182898 434382 183134
rect 433826 147218 434062 147454
rect 434146 147218 434382 147454
rect 433826 146898 434062 147134
rect 434146 146898 434382 147134
rect 419546 60938 419782 61174
rect 419866 60938 420102 61174
rect 419546 60618 419782 60854
rect 419866 60618 420102 60854
rect 419546 24938 419782 25174
rect 419866 24938 420102 25174
rect 419546 24618 419782 24854
rect 419866 24618 420102 24854
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -1542 416062 -1306
rect 416146 -1542 416382 -1306
rect 415826 -1862 416062 -1626
rect 416146 -1862 416382 -1626
rect 419546 -3462 419782 -3226
rect 419866 -3462 420102 -3226
rect 419546 -3782 419782 -3546
rect 419866 -3782 420102 -3546
rect 423266 64658 423502 64894
rect 423586 64658 423822 64894
rect 423266 64338 423502 64574
rect 423586 64338 423822 64574
rect 426586 111218 426822 111454
rect 426586 110898 426822 111134
rect 426986 68378 427222 68614
rect 427306 68378 427542 68614
rect 426986 68058 427222 68294
rect 427306 68058 427542 68294
rect 423266 28658 423502 28894
rect 423586 28658 423822 28894
rect 423266 28338 423502 28574
rect 423586 28338 423822 28574
rect 423266 -5382 423502 -5146
rect 423586 -5382 423822 -5146
rect 423266 -5702 423502 -5466
rect 423586 -5702 423822 -5466
rect 426986 32378 427222 32614
rect 427306 32378 427542 32614
rect 426986 32058 427222 32294
rect 427306 32058 427542 32294
rect 408986 -6342 409222 -6106
rect 409306 -6342 409542 -6106
rect 408986 -6662 409222 -6426
rect 409306 -6662 409542 -6426
rect 428186 129218 428422 129454
rect 428186 128898 428422 129134
rect 437546 690938 437782 691174
rect 437866 690938 438102 691174
rect 437546 690618 437782 690854
rect 437866 690618 438102 690854
rect 437546 654938 437782 655174
rect 437866 654938 438102 655174
rect 437546 654618 437782 654854
rect 437866 654618 438102 654854
rect 437546 618938 437782 619174
rect 437866 618938 438102 619174
rect 437546 618618 437782 618854
rect 437866 618618 438102 618854
rect 437546 582938 437782 583174
rect 437866 582938 438102 583174
rect 437546 582618 437782 582854
rect 437866 582618 438102 582854
rect 437546 546938 437782 547174
rect 437866 546938 438102 547174
rect 437546 546618 437782 546854
rect 437866 546618 438102 546854
rect 437546 510938 437782 511174
rect 437866 510938 438102 511174
rect 437546 510618 437782 510854
rect 437866 510618 438102 510854
rect 437546 474938 437782 475174
rect 437866 474938 438102 475174
rect 437546 474618 437782 474854
rect 437866 474618 438102 474854
rect 437546 438938 437782 439174
rect 437866 438938 438102 439174
rect 437546 438618 437782 438854
rect 437866 438618 438102 438854
rect 437546 402938 437782 403174
rect 437866 402938 438102 403174
rect 437546 402618 437782 402854
rect 437866 402618 438102 402854
rect 437546 366938 437782 367174
rect 437866 366938 438102 367174
rect 437546 366618 437782 366854
rect 437866 366618 438102 366854
rect 437546 330938 437782 331174
rect 437866 330938 438102 331174
rect 437546 330618 437782 330854
rect 437866 330618 438102 330854
rect 437546 294938 437782 295174
rect 437866 294938 438102 295174
rect 437546 294618 437782 294854
rect 437866 294618 438102 294854
rect 441266 694658 441502 694894
rect 441586 694658 441822 694894
rect 441266 694338 441502 694574
rect 441586 694338 441822 694574
rect 441266 658658 441502 658894
rect 441586 658658 441822 658894
rect 441266 658338 441502 658574
rect 441586 658338 441822 658574
rect 441266 622658 441502 622894
rect 441586 622658 441822 622894
rect 441266 622338 441502 622574
rect 441586 622338 441822 622574
rect 441266 586658 441502 586894
rect 441586 586658 441822 586894
rect 441266 586338 441502 586574
rect 441586 586338 441822 586574
rect 441266 550658 441502 550894
rect 441586 550658 441822 550894
rect 441266 550338 441502 550574
rect 441586 550338 441822 550574
rect 441266 514658 441502 514894
rect 441586 514658 441822 514894
rect 441266 514338 441502 514574
rect 441586 514338 441822 514574
rect 441266 478658 441502 478894
rect 441586 478658 441822 478894
rect 441266 478338 441502 478574
rect 441586 478338 441822 478574
rect 441266 442658 441502 442894
rect 441586 442658 441822 442894
rect 441266 442338 441502 442574
rect 441586 442338 441822 442574
rect 441266 406658 441502 406894
rect 441586 406658 441822 406894
rect 441266 406338 441502 406574
rect 441586 406338 441822 406574
rect 441266 370658 441502 370894
rect 441586 370658 441822 370894
rect 441266 370338 441502 370574
rect 441586 370338 441822 370574
rect 441266 334658 441502 334894
rect 441586 334658 441822 334894
rect 441266 334338 441502 334574
rect 441586 334338 441822 334574
rect 441266 298658 441502 298894
rect 441586 298658 441822 298894
rect 441266 298338 441502 298574
rect 441586 298338 441822 298574
rect 437546 258938 437782 259174
rect 437866 258938 438102 259174
rect 437546 258618 437782 258854
rect 437866 258618 438102 258854
rect 437546 222938 437782 223174
rect 437866 222938 438102 223174
rect 437546 222618 437782 222854
rect 437866 222618 438102 222854
rect 437546 186938 437782 187174
rect 437866 186938 438102 187174
rect 437546 186618 437782 186854
rect 437866 186618 438102 186854
rect 437546 150938 437782 151174
rect 437866 150938 438102 151174
rect 437546 150618 437782 150854
rect 437866 150618 438102 150854
rect 431386 129218 431622 129454
rect 431386 128898 431622 129134
rect 429786 111218 430022 111454
rect 429786 110898 430022 111134
rect 434586 129218 434822 129454
rect 434586 128898 434822 129134
rect 432986 111218 433222 111454
rect 432986 110898 433222 111134
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 437786 129218 438022 129454
rect 437786 128898 438022 129134
rect 441266 262658 441502 262894
rect 441586 262658 441822 262894
rect 441266 262338 441502 262574
rect 441586 262338 441822 262574
rect 441266 226658 441502 226894
rect 441586 226658 441822 226894
rect 441266 226338 441502 226574
rect 441586 226338 441822 226574
rect 462986 711322 463222 711558
rect 463306 711322 463542 711558
rect 462986 711002 463222 711238
rect 463306 711002 463542 711238
rect 459266 709402 459502 709638
rect 459586 709402 459822 709638
rect 459266 709082 459502 709318
rect 459586 709082 459822 709318
rect 455546 707482 455782 707718
rect 455866 707482 456102 707718
rect 455546 707162 455782 707398
rect 455866 707162 456102 707398
rect 444986 698378 445222 698614
rect 445306 698378 445542 698614
rect 444986 698058 445222 698294
rect 445306 698058 445542 698294
rect 444986 662378 445222 662614
rect 445306 662378 445542 662614
rect 444986 662058 445222 662294
rect 445306 662058 445542 662294
rect 444986 626378 445222 626614
rect 445306 626378 445542 626614
rect 444986 626058 445222 626294
rect 445306 626058 445542 626294
rect 444986 590378 445222 590614
rect 445306 590378 445542 590614
rect 444986 590058 445222 590294
rect 445306 590058 445542 590294
rect 444986 554378 445222 554614
rect 445306 554378 445542 554614
rect 444986 554058 445222 554294
rect 445306 554058 445542 554294
rect 444986 518378 445222 518614
rect 445306 518378 445542 518614
rect 444986 518058 445222 518294
rect 445306 518058 445542 518294
rect 444986 482378 445222 482614
rect 445306 482378 445542 482614
rect 444986 482058 445222 482294
rect 445306 482058 445542 482294
rect 444986 446378 445222 446614
rect 445306 446378 445542 446614
rect 444986 446058 445222 446294
rect 445306 446058 445542 446294
rect 444986 410378 445222 410614
rect 445306 410378 445542 410614
rect 444986 410058 445222 410294
rect 445306 410058 445542 410294
rect 444986 374378 445222 374614
rect 445306 374378 445542 374614
rect 444986 374058 445222 374294
rect 445306 374058 445542 374294
rect 444986 338378 445222 338614
rect 445306 338378 445542 338614
rect 444986 338058 445222 338294
rect 445306 338058 445542 338294
rect 444986 302378 445222 302614
rect 445306 302378 445542 302614
rect 444986 302058 445222 302294
rect 445306 302058 445542 302294
rect 444986 266378 445222 266614
rect 445306 266378 445542 266614
rect 444986 266058 445222 266294
rect 445306 266058 445542 266294
rect 444986 230378 445222 230614
rect 445306 230378 445542 230614
rect 444986 230058 445222 230294
rect 445306 230058 445542 230294
rect 441266 190658 441502 190894
rect 441586 190658 441822 190894
rect 441266 190338 441502 190574
rect 441586 190338 441822 190574
rect 441266 154658 441502 154894
rect 441586 154658 441822 154894
rect 441266 154338 441502 154574
rect 441586 154338 441822 154574
rect 436186 111218 436422 111454
rect 436186 110898 436422 111134
rect 437546 78938 437782 79174
rect 437866 78938 438102 79174
rect 437546 78618 437782 78854
rect 437866 78618 438102 78854
rect 437546 42938 437782 43174
rect 437866 42938 438102 43174
rect 437546 42618 437782 42854
rect 437866 42618 438102 42854
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 444986 194378 445222 194614
rect 445306 194378 445542 194614
rect 444986 194058 445222 194294
rect 445306 194058 445542 194294
rect 444986 158378 445222 158614
rect 445306 158378 445542 158614
rect 444986 158058 445222 158294
rect 445306 158058 445542 158294
rect 444986 122378 445222 122614
rect 445306 122378 445542 122614
rect 444986 122058 445222 122294
rect 445306 122058 445542 122294
rect 441266 82658 441502 82894
rect 441586 82658 441822 82894
rect 441266 82338 441502 82574
rect 441586 82338 441822 82574
rect 441266 46658 441502 46894
rect 441586 46658 441822 46894
rect 441266 46338 441502 46574
rect 441586 46338 441822 46574
rect 441266 10658 441502 10894
rect 441586 10658 441822 10894
rect 441266 10338 441502 10574
rect 441586 10338 441822 10574
rect 437546 6938 437782 7174
rect 437866 6938 438102 7174
rect 437546 6618 437782 6854
rect 437866 6618 438102 6854
rect 437546 -2502 437782 -2266
rect 437866 -2502 438102 -2266
rect 437546 -2822 437782 -2586
rect 437866 -2822 438102 -2586
rect 441266 -4422 441502 -4186
rect 441586 -4422 441822 -4186
rect 441266 -4742 441502 -4506
rect 441586 -4742 441822 -4506
rect 444986 86378 445222 86614
rect 445306 86378 445542 86614
rect 444986 86058 445222 86294
rect 445306 86058 445542 86294
rect 444986 50378 445222 50614
rect 445306 50378 445542 50614
rect 444986 50058 445222 50294
rect 445306 50058 445542 50294
rect 444986 14378 445222 14614
rect 445306 14378 445542 14614
rect 444986 14058 445222 14294
rect 445306 14058 445542 14294
rect 426986 -7302 427222 -7066
rect 427306 -7302 427542 -7066
rect 426986 -7622 427222 -7386
rect 427306 -7622 427542 -7386
rect 451826 705562 452062 705798
rect 452146 705562 452382 705798
rect 451826 705242 452062 705478
rect 452146 705242 452382 705478
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 451826 561218 452062 561454
rect 452146 561218 452382 561454
rect 451826 560898 452062 561134
rect 452146 560898 452382 561134
rect 451826 525218 452062 525454
rect 452146 525218 452382 525454
rect 451826 524898 452062 525134
rect 452146 524898 452382 525134
rect 451826 489218 452062 489454
rect 452146 489218 452382 489454
rect 451826 488898 452062 489134
rect 452146 488898 452382 489134
rect 451826 453218 452062 453454
rect 452146 453218 452382 453454
rect 451826 452898 452062 453134
rect 452146 452898 452382 453134
rect 451826 417218 452062 417454
rect 452146 417218 452382 417454
rect 451826 416898 452062 417134
rect 452146 416898 452382 417134
rect 451826 381218 452062 381454
rect 452146 381218 452382 381454
rect 451826 380898 452062 381134
rect 452146 380898 452382 381134
rect 451826 345218 452062 345454
rect 452146 345218 452382 345454
rect 451826 344898 452062 345134
rect 452146 344898 452382 345134
rect 451826 309218 452062 309454
rect 452146 309218 452382 309454
rect 451826 308898 452062 309134
rect 452146 308898 452382 309134
rect 451826 273218 452062 273454
rect 452146 273218 452382 273454
rect 451826 272898 452062 273134
rect 452146 272898 452382 273134
rect 451826 237218 452062 237454
rect 452146 237218 452382 237454
rect 451826 236898 452062 237134
rect 452146 236898 452382 237134
rect 451826 201218 452062 201454
rect 452146 201218 452382 201454
rect 451826 200898 452062 201134
rect 452146 200898 452382 201134
rect 451826 165218 452062 165454
rect 452146 165218 452382 165454
rect 451826 164898 452062 165134
rect 452146 164898 452382 165134
rect 451826 129218 452062 129454
rect 452146 129218 452382 129454
rect 451826 128898 452062 129134
rect 452146 128898 452382 129134
rect 451826 93218 452062 93454
rect 452146 93218 452382 93454
rect 451826 92898 452062 93134
rect 452146 92898 452382 93134
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -1542 452062 -1306
rect 452146 -1542 452382 -1306
rect 451826 -1862 452062 -1626
rect 452146 -1862 452382 -1626
rect 455546 672938 455782 673174
rect 455866 672938 456102 673174
rect 455546 672618 455782 672854
rect 455866 672618 456102 672854
rect 455546 636938 455782 637174
rect 455866 636938 456102 637174
rect 455546 636618 455782 636854
rect 455866 636618 456102 636854
rect 455546 600938 455782 601174
rect 455866 600938 456102 601174
rect 455546 600618 455782 600854
rect 455866 600618 456102 600854
rect 455546 564938 455782 565174
rect 455866 564938 456102 565174
rect 455546 564618 455782 564854
rect 455866 564618 456102 564854
rect 455546 528938 455782 529174
rect 455866 528938 456102 529174
rect 455546 528618 455782 528854
rect 455866 528618 456102 528854
rect 455546 492938 455782 493174
rect 455866 492938 456102 493174
rect 455546 492618 455782 492854
rect 455866 492618 456102 492854
rect 455546 456938 455782 457174
rect 455866 456938 456102 457174
rect 455546 456618 455782 456854
rect 455866 456618 456102 456854
rect 455546 420938 455782 421174
rect 455866 420938 456102 421174
rect 455546 420618 455782 420854
rect 455866 420618 456102 420854
rect 455546 384938 455782 385174
rect 455866 384938 456102 385174
rect 455546 384618 455782 384854
rect 455866 384618 456102 384854
rect 455546 348938 455782 349174
rect 455866 348938 456102 349174
rect 455546 348618 455782 348854
rect 455866 348618 456102 348854
rect 455546 312938 455782 313174
rect 455866 312938 456102 313174
rect 455546 312618 455782 312854
rect 455866 312618 456102 312854
rect 455546 276938 455782 277174
rect 455866 276938 456102 277174
rect 455546 276618 455782 276854
rect 455866 276618 456102 276854
rect 455546 240938 455782 241174
rect 455866 240938 456102 241174
rect 455546 240618 455782 240854
rect 455866 240618 456102 240854
rect 455546 204938 455782 205174
rect 455866 204938 456102 205174
rect 455546 204618 455782 204854
rect 455866 204618 456102 204854
rect 455546 168938 455782 169174
rect 455866 168938 456102 169174
rect 455546 168618 455782 168854
rect 455866 168618 456102 168854
rect 455546 132938 455782 133174
rect 455866 132938 456102 133174
rect 455546 132618 455782 132854
rect 455866 132618 456102 132854
rect 455546 96938 455782 97174
rect 455866 96938 456102 97174
rect 455546 96618 455782 96854
rect 455866 96618 456102 96854
rect 455546 60938 455782 61174
rect 455866 60938 456102 61174
rect 455546 60618 455782 60854
rect 455866 60618 456102 60854
rect 455546 24938 455782 25174
rect 455866 24938 456102 25174
rect 455546 24618 455782 24854
rect 455866 24618 456102 24854
rect 455546 -3462 455782 -3226
rect 455866 -3462 456102 -3226
rect 455546 -3782 455782 -3546
rect 455866 -3782 456102 -3546
rect 459266 676658 459502 676894
rect 459586 676658 459822 676894
rect 459266 676338 459502 676574
rect 459586 676338 459822 676574
rect 459266 640658 459502 640894
rect 459586 640658 459822 640894
rect 459266 640338 459502 640574
rect 459586 640338 459822 640574
rect 459266 604658 459502 604894
rect 459586 604658 459822 604894
rect 459266 604338 459502 604574
rect 459586 604338 459822 604574
rect 459266 568658 459502 568894
rect 459586 568658 459822 568894
rect 459266 568338 459502 568574
rect 459586 568338 459822 568574
rect 459266 532658 459502 532894
rect 459586 532658 459822 532894
rect 459266 532338 459502 532574
rect 459586 532338 459822 532574
rect 459266 496658 459502 496894
rect 459586 496658 459822 496894
rect 459266 496338 459502 496574
rect 459586 496338 459822 496574
rect 459266 460658 459502 460894
rect 459586 460658 459822 460894
rect 459266 460338 459502 460574
rect 459586 460338 459822 460574
rect 459266 424658 459502 424894
rect 459586 424658 459822 424894
rect 459266 424338 459502 424574
rect 459586 424338 459822 424574
rect 459266 388658 459502 388894
rect 459586 388658 459822 388894
rect 459266 388338 459502 388574
rect 459586 388338 459822 388574
rect 459266 352658 459502 352894
rect 459586 352658 459822 352894
rect 459266 352338 459502 352574
rect 459586 352338 459822 352574
rect 459266 316658 459502 316894
rect 459586 316658 459822 316894
rect 459266 316338 459502 316574
rect 459586 316338 459822 316574
rect 459266 280658 459502 280894
rect 459586 280658 459822 280894
rect 459266 280338 459502 280574
rect 459586 280338 459822 280574
rect 459266 244658 459502 244894
rect 459586 244658 459822 244894
rect 459266 244338 459502 244574
rect 459586 244338 459822 244574
rect 459266 208658 459502 208894
rect 459586 208658 459822 208894
rect 459266 208338 459502 208574
rect 459586 208338 459822 208574
rect 459266 172658 459502 172894
rect 459586 172658 459822 172894
rect 459266 172338 459502 172574
rect 459586 172338 459822 172574
rect 459266 136658 459502 136894
rect 459586 136658 459822 136894
rect 459266 136338 459502 136574
rect 459586 136338 459822 136574
rect 459266 100658 459502 100894
rect 459586 100658 459822 100894
rect 459266 100338 459502 100574
rect 459586 100338 459822 100574
rect 459266 64658 459502 64894
rect 459586 64658 459822 64894
rect 459266 64338 459502 64574
rect 459586 64338 459822 64574
rect 459266 28658 459502 28894
rect 459586 28658 459822 28894
rect 459266 28338 459502 28574
rect 459586 28338 459822 28574
rect 459266 -5382 459502 -5146
rect 459586 -5382 459822 -5146
rect 459266 -5702 459502 -5466
rect 459586 -5702 459822 -5466
rect 480986 710362 481222 710598
rect 481306 710362 481542 710598
rect 480986 710042 481222 710278
rect 481306 710042 481542 710278
rect 477266 708442 477502 708678
rect 477586 708442 477822 708678
rect 477266 708122 477502 708358
rect 477586 708122 477822 708358
rect 473546 706522 473782 706758
rect 473866 706522 474102 706758
rect 473546 706202 473782 706438
rect 473866 706202 474102 706438
rect 462986 680378 463222 680614
rect 463306 680378 463542 680614
rect 462986 680058 463222 680294
rect 463306 680058 463542 680294
rect 462986 644378 463222 644614
rect 463306 644378 463542 644614
rect 462986 644058 463222 644294
rect 463306 644058 463542 644294
rect 462986 608378 463222 608614
rect 463306 608378 463542 608614
rect 462986 608058 463222 608294
rect 463306 608058 463542 608294
rect 462986 572378 463222 572614
rect 463306 572378 463542 572614
rect 462986 572058 463222 572294
rect 463306 572058 463542 572294
rect 462986 536378 463222 536614
rect 463306 536378 463542 536614
rect 462986 536058 463222 536294
rect 463306 536058 463542 536294
rect 462986 500378 463222 500614
rect 463306 500378 463542 500614
rect 462986 500058 463222 500294
rect 463306 500058 463542 500294
rect 462986 464378 463222 464614
rect 463306 464378 463542 464614
rect 462986 464058 463222 464294
rect 463306 464058 463542 464294
rect 462986 428378 463222 428614
rect 463306 428378 463542 428614
rect 462986 428058 463222 428294
rect 463306 428058 463542 428294
rect 462986 392378 463222 392614
rect 463306 392378 463542 392614
rect 462986 392058 463222 392294
rect 463306 392058 463542 392294
rect 462986 356378 463222 356614
rect 463306 356378 463542 356614
rect 462986 356058 463222 356294
rect 463306 356058 463542 356294
rect 462986 320378 463222 320614
rect 463306 320378 463542 320614
rect 462986 320058 463222 320294
rect 463306 320058 463542 320294
rect 462986 284378 463222 284614
rect 463306 284378 463542 284614
rect 462986 284058 463222 284294
rect 463306 284058 463542 284294
rect 462986 248378 463222 248614
rect 463306 248378 463542 248614
rect 462986 248058 463222 248294
rect 463306 248058 463542 248294
rect 462986 212378 463222 212614
rect 463306 212378 463542 212614
rect 462986 212058 463222 212294
rect 463306 212058 463542 212294
rect 462986 176378 463222 176614
rect 463306 176378 463542 176614
rect 462986 176058 463222 176294
rect 463306 176058 463542 176294
rect 462986 140378 463222 140614
rect 463306 140378 463542 140614
rect 462986 140058 463222 140294
rect 463306 140058 463542 140294
rect 462986 104378 463222 104614
rect 463306 104378 463542 104614
rect 462986 104058 463222 104294
rect 463306 104058 463542 104294
rect 462986 68378 463222 68614
rect 463306 68378 463542 68614
rect 462986 68058 463222 68294
rect 463306 68058 463542 68294
rect 462986 32378 463222 32614
rect 463306 32378 463542 32614
rect 462986 32058 463222 32294
rect 463306 32058 463542 32294
rect 444986 -6342 445222 -6106
rect 445306 -6342 445542 -6106
rect 444986 -6662 445222 -6426
rect 445306 -6662 445542 -6426
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 469826 327218 470062 327454
rect 470146 327218 470382 327454
rect 469826 326898 470062 327134
rect 470146 326898 470382 327134
rect 469826 291218 470062 291454
rect 470146 291218 470382 291454
rect 469826 290898 470062 291134
rect 470146 290898 470382 291134
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 469826 219218 470062 219454
rect 470146 219218 470382 219454
rect 469826 218898 470062 219134
rect 470146 218898 470382 219134
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 473546 690938 473782 691174
rect 473866 690938 474102 691174
rect 473546 690618 473782 690854
rect 473866 690618 474102 690854
rect 473546 654938 473782 655174
rect 473866 654938 474102 655174
rect 473546 654618 473782 654854
rect 473866 654618 474102 654854
rect 473546 618938 473782 619174
rect 473866 618938 474102 619174
rect 473546 618618 473782 618854
rect 473866 618618 474102 618854
rect 473546 582938 473782 583174
rect 473866 582938 474102 583174
rect 473546 582618 473782 582854
rect 473866 582618 474102 582854
rect 473546 546938 473782 547174
rect 473866 546938 474102 547174
rect 473546 546618 473782 546854
rect 473866 546618 474102 546854
rect 473546 510938 473782 511174
rect 473866 510938 474102 511174
rect 473546 510618 473782 510854
rect 473866 510618 474102 510854
rect 473546 474938 473782 475174
rect 473866 474938 474102 475174
rect 473546 474618 473782 474854
rect 473866 474618 474102 474854
rect 473546 438938 473782 439174
rect 473866 438938 474102 439174
rect 473546 438618 473782 438854
rect 473866 438618 474102 438854
rect 473546 402938 473782 403174
rect 473866 402938 474102 403174
rect 473546 402618 473782 402854
rect 473866 402618 474102 402854
rect 473546 366938 473782 367174
rect 473866 366938 474102 367174
rect 473546 366618 473782 366854
rect 473866 366618 474102 366854
rect 473546 330938 473782 331174
rect 473866 330938 474102 331174
rect 473546 330618 473782 330854
rect 473866 330618 474102 330854
rect 473546 294938 473782 295174
rect 473866 294938 474102 295174
rect 473546 294618 473782 294854
rect 473866 294618 474102 294854
rect 473546 258938 473782 259174
rect 473866 258938 474102 259174
rect 473546 258618 473782 258854
rect 473866 258618 474102 258854
rect 473546 222938 473782 223174
rect 473866 222938 474102 223174
rect 473546 222618 473782 222854
rect 473866 222618 474102 222854
rect 473546 186938 473782 187174
rect 473866 186938 474102 187174
rect 473546 186618 473782 186854
rect 473866 186618 474102 186854
rect 473546 150938 473782 151174
rect 473866 150938 474102 151174
rect 473546 150618 473782 150854
rect 473866 150618 474102 150854
rect 473546 114938 473782 115174
rect 473866 114938 474102 115174
rect 473546 114618 473782 114854
rect 473866 114618 474102 114854
rect 473546 78938 473782 79174
rect 473866 78938 474102 79174
rect 473546 78618 473782 78854
rect 473866 78618 474102 78854
rect 473546 42938 473782 43174
rect 473866 42938 474102 43174
rect 473546 42618 473782 42854
rect 473866 42618 474102 42854
rect 473546 6938 473782 7174
rect 473866 6938 474102 7174
rect 473546 6618 473782 6854
rect 473866 6618 474102 6854
rect 473546 -2502 473782 -2266
rect 473866 -2502 474102 -2266
rect 473546 -2822 473782 -2586
rect 473866 -2822 474102 -2586
rect 477266 694658 477502 694894
rect 477586 694658 477822 694894
rect 477266 694338 477502 694574
rect 477586 694338 477822 694574
rect 477266 658658 477502 658894
rect 477586 658658 477822 658894
rect 477266 658338 477502 658574
rect 477586 658338 477822 658574
rect 477266 622658 477502 622894
rect 477586 622658 477822 622894
rect 477266 622338 477502 622574
rect 477586 622338 477822 622574
rect 477266 586658 477502 586894
rect 477586 586658 477822 586894
rect 477266 586338 477502 586574
rect 477586 586338 477822 586574
rect 477266 550658 477502 550894
rect 477586 550658 477822 550894
rect 477266 550338 477502 550574
rect 477586 550338 477822 550574
rect 477266 514658 477502 514894
rect 477586 514658 477822 514894
rect 477266 514338 477502 514574
rect 477586 514338 477822 514574
rect 477266 478658 477502 478894
rect 477586 478658 477822 478894
rect 477266 478338 477502 478574
rect 477586 478338 477822 478574
rect 477266 442658 477502 442894
rect 477586 442658 477822 442894
rect 477266 442338 477502 442574
rect 477586 442338 477822 442574
rect 477266 406658 477502 406894
rect 477586 406658 477822 406894
rect 477266 406338 477502 406574
rect 477586 406338 477822 406574
rect 477266 370658 477502 370894
rect 477586 370658 477822 370894
rect 477266 370338 477502 370574
rect 477586 370338 477822 370574
rect 477266 334658 477502 334894
rect 477586 334658 477822 334894
rect 477266 334338 477502 334574
rect 477586 334338 477822 334574
rect 477266 298658 477502 298894
rect 477586 298658 477822 298894
rect 477266 298338 477502 298574
rect 477586 298338 477822 298574
rect 477266 262658 477502 262894
rect 477586 262658 477822 262894
rect 477266 262338 477502 262574
rect 477586 262338 477822 262574
rect 477266 226658 477502 226894
rect 477586 226658 477822 226894
rect 477266 226338 477502 226574
rect 477586 226338 477822 226574
rect 477266 190658 477502 190894
rect 477586 190658 477822 190894
rect 477266 190338 477502 190574
rect 477586 190338 477822 190574
rect 477266 154658 477502 154894
rect 477586 154658 477822 154894
rect 477266 154338 477502 154574
rect 477586 154338 477822 154574
rect 477266 118658 477502 118894
rect 477586 118658 477822 118894
rect 477266 118338 477502 118574
rect 477586 118338 477822 118574
rect 477266 82658 477502 82894
rect 477586 82658 477822 82894
rect 477266 82338 477502 82574
rect 477586 82338 477822 82574
rect 477266 46658 477502 46894
rect 477586 46658 477822 46894
rect 477266 46338 477502 46574
rect 477586 46338 477822 46574
rect 477266 10658 477502 10894
rect 477586 10658 477822 10894
rect 477266 10338 477502 10574
rect 477586 10338 477822 10574
rect 477266 -4422 477502 -4186
rect 477586 -4422 477822 -4186
rect 477266 -4742 477502 -4506
rect 477586 -4742 477822 -4506
rect 498986 711322 499222 711558
rect 499306 711322 499542 711558
rect 498986 711002 499222 711238
rect 499306 711002 499542 711238
rect 495266 709402 495502 709638
rect 495586 709402 495822 709638
rect 495266 709082 495502 709318
rect 495586 709082 495822 709318
rect 491546 707482 491782 707718
rect 491866 707482 492102 707718
rect 491546 707162 491782 707398
rect 491866 707162 492102 707398
rect 480986 698378 481222 698614
rect 481306 698378 481542 698614
rect 480986 698058 481222 698294
rect 481306 698058 481542 698294
rect 480986 662378 481222 662614
rect 481306 662378 481542 662614
rect 480986 662058 481222 662294
rect 481306 662058 481542 662294
rect 480986 626378 481222 626614
rect 481306 626378 481542 626614
rect 480986 626058 481222 626294
rect 481306 626058 481542 626294
rect 480986 590378 481222 590614
rect 481306 590378 481542 590614
rect 480986 590058 481222 590294
rect 481306 590058 481542 590294
rect 480986 554378 481222 554614
rect 481306 554378 481542 554614
rect 480986 554058 481222 554294
rect 481306 554058 481542 554294
rect 480986 518378 481222 518614
rect 481306 518378 481542 518614
rect 480986 518058 481222 518294
rect 481306 518058 481542 518294
rect 480986 482378 481222 482614
rect 481306 482378 481542 482614
rect 480986 482058 481222 482294
rect 481306 482058 481542 482294
rect 480986 446378 481222 446614
rect 481306 446378 481542 446614
rect 480986 446058 481222 446294
rect 481306 446058 481542 446294
rect 480986 410378 481222 410614
rect 481306 410378 481542 410614
rect 480986 410058 481222 410294
rect 481306 410058 481542 410294
rect 480986 374378 481222 374614
rect 481306 374378 481542 374614
rect 480986 374058 481222 374294
rect 481306 374058 481542 374294
rect 480986 338378 481222 338614
rect 481306 338378 481542 338614
rect 480986 338058 481222 338294
rect 481306 338058 481542 338294
rect 480986 302378 481222 302614
rect 481306 302378 481542 302614
rect 480986 302058 481222 302294
rect 481306 302058 481542 302294
rect 480986 266378 481222 266614
rect 481306 266378 481542 266614
rect 480986 266058 481222 266294
rect 481306 266058 481542 266294
rect 480986 230378 481222 230614
rect 481306 230378 481542 230614
rect 480986 230058 481222 230294
rect 481306 230058 481542 230294
rect 480986 194378 481222 194614
rect 481306 194378 481542 194614
rect 480986 194058 481222 194294
rect 481306 194058 481542 194294
rect 480986 158378 481222 158614
rect 481306 158378 481542 158614
rect 480986 158058 481222 158294
rect 481306 158058 481542 158294
rect 480986 122378 481222 122614
rect 481306 122378 481542 122614
rect 480986 122058 481222 122294
rect 481306 122058 481542 122294
rect 480986 86378 481222 86614
rect 481306 86378 481542 86614
rect 480986 86058 481222 86294
rect 481306 86058 481542 86294
rect 480986 50378 481222 50614
rect 481306 50378 481542 50614
rect 480986 50058 481222 50294
rect 481306 50058 481542 50294
rect 480986 14378 481222 14614
rect 481306 14378 481542 14614
rect 480986 14058 481222 14294
rect 481306 14058 481542 14294
rect 462986 -7302 463222 -7066
rect 463306 -7302 463542 -7066
rect 462986 -7622 463222 -7386
rect 463306 -7622 463542 -7386
rect 487826 705562 488062 705798
rect 488146 705562 488382 705798
rect 487826 705242 488062 705478
rect 488146 705242 488382 705478
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 487826 633218 488062 633454
rect 488146 633218 488382 633454
rect 487826 632898 488062 633134
rect 488146 632898 488382 633134
rect 487826 597218 488062 597454
rect 488146 597218 488382 597454
rect 487826 596898 488062 597134
rect 488146 596898 488382 597134
rect 487826 561218 488062 561454
rect 488146 561218 488382 561454
rect 487826 560898 488062 561134
rect 488146 560898 488382 561134
rect 487826 525218 488062 525454
rect 488146 525218 488382 525454
rect 487826 524898 488062 525134
rect 488146 524898 488382 525134
rect 487826 489218 488062 489454
rect 488146 489218 488382 489454
rect 487826 488898 488062 489134
rect 488146 488898 488382 489134
rect 487826 453218 488062 453454
rect 488146 453218 488382 453454
rect 487826 452898 488062 453134
rect 488146 452898 488382 453134
rect 487826 417218 488062 417454
rect 488146 417218 488382 417454
rect 487826 416898 488062 417134
rect 488146 416898 488382 417134
rect 487826 381218 488062 381454
rect 488146 381218 488382 381454
rect 487826 380898 488062 381134
rect 488146 380898 488382 381134
rect 487826 345218 488062 345454
rect 488146 345218 488382 345454
rect 487826 344898 488062 345134
rect 488146 344898 488382 345134
rect 487826 309218 488062 309454
rect 488146 309218 488382 309454
rect 487826 308898 488062 309134
rect 488146 308898 488382 309134
rect 487826 273218 488062 273454
rect 488146 273218 488382 273454
rect 487826 272898 488062 273134
rect 488146 272898 488382 273134
rect 487826 237218 488062 237454
rect 488146 237218 488382 237454
rect 487826 236898 488062 237134
rect 488146 236898 488382 237134
rect 487826 201218 488062 201454
rect 488146 201218 488382 201454
rect 487826 200898 488062 201134
rect 488146 200898 488382 201134
rect 487826 165218 488062 165454
rect 488146 165218 488382 165454
rect 487826 164898 488062 165134
rect 488146 164898 488382 165134
rect 487826 129218 488062 129454
rect 488146 129218 488382 129454
rect 487826 128898 488062 129134
rect 488146 128898 488382 129134
rect 487826 93218 488062 93454
rect 488146 93218 488382 93454
rect 487826 92898 488062 93134
rect 488146 92898 488382 93134
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -1542 488062 -1306
rect 488146 -1542 488382 -1306
rect 487826 -1862 488062 -1626
rect 488146 -1862 488382 -1626
rect 491546 672938 491782 673174
rect 491866 672938 492102 673174
rect 491546 672618 491782 672854
rect 491866 672618 492102 672854
rect 491546 636938 491782 637174
rect 491866 636938 492102 637174
rect 491546 636618 491782 636854
rect 491866 636618 492102 636854
rect 491546 600938 491782 601174
rect 491866 600938 492102 601174
rect 491546 600618 491782 600854
rect 491866 600618 492102 600854
rect 491546 564938 491782 565174
rect 491866 564938 492102 565174
rect 491546 564618 491782 564854
rect 491866 564618 492102 564854
rect 491546 528938 491782 529174
rect 491866 528938 492102 529174
rect 491546 528618 491782 528854
rect 491866 528618 492102 528854
rect 491546 492938 491782 493174
rect 491866 492938 492102 493174
rect 491546 492618 491782 492854
rect 491866 492618 492102 492854
rect 491546 456938 491782 457174
rect 491866 456938 492102 457174
rect 491546 456618 491782 456854
rect 491866 456618 492102 456854
rect 491546 420938 491782 421174
rect 491866 420938 492102 421174
rect 491546 420618 491782 420854
rect 491866 420618 492102 420854
rect 491546 384938 491782 385174
rect 491866 384938 492102 385174
rect 491546 384618 491782 384854
rect 491866 384618 492102 384854
rect 491546 348938 491782 349174
rect 491866 348938 492102 349174
rect 491546 348618 491782 348854
rect 491866 348618 492102 348854
rect 491546 312938 491782 313174
rect 491866 312938 492102 313174
rect 491546 312618 491782 312854
rect 491866 312618 492102 312854
rect 491546 276938 491782 277174
rect 491866 276938 492102 277174
rect 491546 276618 491782 276854
rect 491866 276618 492102 276854
rect 491546 240938 491782 241174
rect 491866 240938 492102 241174
rect 491546 240618 491782 240854
rect 491866 240618 492102 240854
rect 491546 204938 491782 205174
rect 491866 204938 492102 205174
rect 491546 204618 491782 204854
rect 491866 204618 492102 204854
rect 491546 168938 491782 169174
rect 491866 168938 492102 169174
rect 491546 168618 491782 168854
rect 491866 168618 492102 168854
rect 491546 132938 491782 133174
rect 491866 132938 492102 133174
rect 491546 132618 491782 132854
rect 491866 132618 492102 132854
rect 491546 96938 491782 97174
rect 491866 96938 492102 97174
rect 491546 96618 491782 96854
rect 491866 96618 492102 96854
rect 491546 60938 491782 61174
rect 491866 60938 492102 61174
rect 491546 60618 491782 60854
rect 491866 60618 492102 60854
rect 491546 24938 491782 25174
rect 491866 24938 492102 25174
rect 491546 24618 491782 24854
rect 491866 24618 492102 24854
rect 491546 -3462 491782 -3226
rect 491866 -3462 492102 -3226
rect 491546 -3782 491782 -3546
rect 491866 -3782 492102 -3546
rect 495266 676658 495502 676894
rect 495586 676658 495822 676894
rect 495266 676338 495502 676574
rect 495586 676338 495822 676574
rect 495266 640658 495502 640894
rect 495586 640658 495822 640894
rect 495266 640338 495502 640574
rect 495586 640338 495822 640574
rect 495266 604658 495502 604894
rect 495586 604658 495822 604894
rect 495266 604338 495502 604574
rect 495586 604338 495822 604574
rect 495266 568658 495502 568894
rect 495586 568658 495822 568894
rect 495266 568338 495502 568574
rect 495586 568338 495822 568574
rect 495266 532658 495502 532894
rect 495586 532658 495822 532894
rect 495266 532338 495502 532574
rect 495586 532338 495822 532574
rect 495266 496658 495502 496894
rect 495586 496658 495822 496894
rect 495266 496338 495502 496574
rect 495586 496338 495822 496574
rect 495266 460658 495502 460894
rect 495586 460658 495822 460894
rect 495266 460338 495502 460574
rect 495586 460338 495822 460574
rect 495266 424658 495502 424894
rect 495586 424658 495822 424894
rect 495266 424338 495502 424574
rect 495586 424338 495822 424574
rect 495266 388658 495502 388894
rect 495586 388658 495822 388894
rect 495266 388338 495502 388574
rect 495586 388338 495822 388574
rect 495266 352658 495502 352894
rect 495586 352658 495822 352894
rect 495266 352338 495502 352574
rect 495586 352338 495822 352574
rect 495266 316658 495502 316894
rect 495586 316658 495822 316894
rect 495266 316338 495502 316574
rect 495586 316338 495822 316574
rect 495266 280658 495502 280894
rect 495586 280658 495822 280894
rect 495266 280338 495502 280574
rect 495586 280338 495822 280574
rect 495266 244658 495502 244894
rect 495586 244658 495822 244894
rect 495266 244338 495502 244574
rect 495586 244338 495822 244574
rect 495266 208658 495502 208894
rect 495586 208658 495822 208894
rect 495266 208338 495502 208574
rect 495586 208338 495822 208574
rect 495266 172658 495502 172894
rect 495586 172658 495822 172894
rect 495266 172338 495502 172574
rect 495586 172338 495822 172574
rect 495266 136658 495502 136894
rect 495586 136658 495822 136894
rect 495266 136338 495502 136574
rect 495586 136338 495822 136574
rect 495266 100658 495502 100894
rect 495586 100658 495822 100894
rect 495266 100338 495502 100574
rect 495586 100338 495822 100574
rect 495266 64658 495502 64894
rect 495586 64658 495822 64894
rect 495266 64338 495502 64574
rect 495586 64338 495822 64574
rect 495266 28658 495502 28894
rect 495586 28658 495822 28894
rect 495266 28338 495502 28574
rect 495586 28338 495822 28574
rect 495266 -5382 495502 -5146
rect 495586 -5382 495822 -5146
rect 495266 -5702 495502 -5466
rect 495586 -5702 495822 -5466
rect 516986 710362 517222 710598
rect 517306 710362 517542 710598
rect 516986 710042 517222 710278
rect 517306 710042 517542 710278
rect 513266 708442 513502 708678
rect 513586 708442 513822 708678
rect 513266 708122 513502 708358
rect 513586 708122 513822 708358
rect 509546 706522 509782 706758
rect 509866 706522 510102 706758
rect 509546 706202 509782 706438
rect 509866 706202 510102 706438
rect 498986 680378 499222 680614
rect 499306 680378 499542 680614
rect 498986 680058 499222 680294
rect 499306 680058 499542 680294
rect 498986 644378 499222 644614
rect 499306 644378 499542 644614
rect 498986 644058 499222 644294
rect 499306 644058 499542 644294
rect 498986 608378 499222 608614
rect 499306 608378 499542 608614
rect 498986 608058 499222 608294
rect 499306 608058 499542 608294
rect 498986 572378 499222 572614
rect 499306 572378 499542 572614
rect 498986 572058 499222 572294
rect 499306 572058 499542 572294
rect 498986 536378 499222 536614
rect 499306 536378 499542 536614
rect 498986 536058 499222 536294
rect 499306 536058 499542 536294
rect 498986 500378 499222 500614
rect 499306 500378 499542 500614
rect 498986 500058 499222 500294
rect 499306 500058 499542 500294
rect 498986 464378 499222 464614
rect 499306 464378 499542 464614
rect 498986 464058 499222 464294
rect 499306 464058 499542 464294
rect 498986 428378 499222 428614
rect 499306 428378 499542 428614
rect 498986 428058 499222 428294
rect 499306 428058 499542 428294
rect 498986 392378 499222 392614
rect 499306 392378 499542 392614
rect 498986 392058 499222 392294
rect 499306 392058 499542 392294
rect 498986 356378 499222 356614
rect 499306 356378 499542 356614
rect 498986 356058 499222 356294
rect 499306 356058 499542 356294
rect 498986 320378 499222 320614
rect 499306 320378 499542 320614
rect 498986 320058 499222 320294
rect 499306 320058 499542 320294
rect 498986 284378 499222 284614
rect 499306 284378 499542 284614
rect 498986 284058 499222 284294
rect 499306 284058 499542 284294
rect 498986 248378 499222 248614
rect 499306 248378 499542 248614
rect 498986 248058 499222 248294
rect 499306 248058 499542 248294
rect 498986 212378 499222 212614
rect 499306 212378 499542 212614
rect 498986 212058 499222 212294
rect 499306 212058 499542 212294
rect 498986 176378 499222 176614
rect 499306 176378 499542 176614
rect 498986 176058 499222 176294
rect 499306 176058 499542 176294
rect 498986 140378 499222 140614
rect 499306 140378 499542 140614
rect 498986 140058 499222 140294
rect 499306 140058 499542 140294
rect 498986 104378 499222 104614
rect 499306 104378 499542 104614
rect 498986 104058 499222 104294
rect 499306 104058 499542 104294
rect 498986 68378 499222 68614
rect 499306 68378 499542 68614
rect 498986 68058 499222 68294
rect 499306 68058 499542 68294
rect 498986 32378 499222 32614
rect 499306 32378 499542 32614
rect 498986 32058 499222 32294
rect 499306 32058 499542 32294
rect 480986 -6342 481222 -6106
rect 481306 -6342 481542 -6106
rect 480986 -6662 481222 -6426
rect 481306 -6662 481542 -6426
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 509546 690938 509782 691174
rect 509866 690938 510102 691174
rect 509546 690618 509782 690854
rect 509866 690618 510102 690854
rect 509546 654938 509782 655174
rect 509866 654938 510102 655174
rect 509546 654618 509782 654854
rect 509866 654618 510102 654854
rect 509546 618938 509782 619174
rect 509866 618938 510102 619174
rect 509546 618618 509782 618854
rect 509866 618618 510102 618854
rect 509546 582938 509782 583174
rect 509866 582938 510102 583174
rect 509546 582618 509782 582854
rect 509866 582618 510102 582854
rect 509546 546938 509782 547174
rect 509866 546938 510102 547174
rect 509546 546618 509782 546854
rect 509866 546618 510102 546854
rect 509546 510938 509782 511174
rect 509866 510938 510102 511174
rect 509546 510618 509782 510854
rect 509866 510618 510102 510854
rect 509546 474938 509782 475174
rect 509866 474938 510102 475174
rect 509546 474618 509782 474854
rect 509866 474618 510102 474854
rect 509546 438938 509782 439174
rect 509866 438938 510102 439174
rect 509546 438618 509782 438854
rect 509866 438618 510102 438854
rect 509546 402938 509782 403174
rect 509866 402938 510102 403174
rect 509546 402618 509782 402854
rect 509866 402618 510102 402854
rect 509546 366938 509782 367174
rect 509866 366938 510102 367174
rect 509546 366618 509782 366854
rect 509866 366618 510102 366854
rect 509546 330938 509782 331174
rect 509866 330938 510102 331174
rect 509546 330618 509782 330854
rect 509866 330618 510102 330854
rect 509546 294938 509782 295174
rect 509866 294938 510102 295174
rect 509546 294618 509782 294854
rect 509866 294618 510102 294854
rect 509546 258938 509782 259174
rect 509866 258938 510102 259174
rect 509546 258618 509782 258854
rect 509866 258618 510102 258854
rect 509546 222938 509782 223174
rect 509866 222938 510102 223174
rect 509546 222618 509782 222854
rect 509866 222618 510102 222854
rect 509546 186938 509782 187174
rect 509866 186938 510102 187174
rect 509546 186618 509782 186854
rect 509866 186618 510102 186854
rect 509546 150938 509782 151174
rect 509866 150938 510102 151174
rect 509546 150618 509782 150854
rect 509866 150618 510102 150854
rect 509546 114938 509782 115174
rect 509866 114938 510102 115174
rect 509546 114618 509782 114854
rect 509866 114618 510102 114854
rect 509546 78938 509782 79174
rect 509866 78938 510102 79174
rect 509546 78618 509782 78854
rect 509866 78618 510102 78854
rect 509546 42938 509782 43174
rect 509866 42938 510102 43174
rect 509546 42618 509782 42854
rect 509866 42618 510102 42854
rect 509546 6938 509782 7174
rect 509866 6938 510102 7174
rect 509546 6618 509782 6854
rect 509866 6618 510102 6854
rect 509546 -2502 509782 -2266
rect 509866 -2502 510102 -2266
rect 509546 -2822 509782 -2586
rect 509866 -2822 510102 -2586
rect 513266 694658 513502 694894
rect 513586 694658 513822 694894
rect 513266 694338 513502 694574
rect 513586 694338 513822 694574
rect 513266 658658 513502 658894
rect 513586 658658 513822 658894
rect 513266 658338 513502 658574
rect 513586 658338 513822 658574
rect 513266 622658 513502 622894
rect 513586 622658 513822 622894
rect 513266 622338 513502 622574
rect 513586 622338 513822 622574
rect 513266 586658 513502 586894
rect 513586 586658 513822 586894
rect 513266 586338 513502 586574
rect 513586 586338 513822 586574
rect 513266 550658 513502 550894
rect 513586 550658 513822 550894
rect 513266 550338 513502 550574
rect 513586 550338 513822 550574
rect 513266 514658 513502 514894
rect 513586 514658 513822 514894
rect 513266 514338 513502 514574
rect 513586 514338 513822 514574
rect 513266 478658 513502 478894
rect 513586 478658 513822 478894
rect 513266 478338 513502 478574
rect 513586 478338 513822 478574
rect 513266 442658 513502 442894
rect 513586 442658 513822 442894
rect 513266 442338 513502 442574
rect 513586 442338 513822 442574
rect 513266 406658 513502 406894
rect 513586 406658 513822 406894
rect 513266 406338 513502 406574
rect 513586 406338 513822 406574
rect 513266 370658 513502 370894
rect 513586 370658 513822 370894
rect 513266 370338 513502 370574
rect 513586 370338 513822 370574
rect 513266 334658 513502 334894
rect 513586 334658 513822 334894
rect 513266 334338 513502 334574
rect 513586 334338 513822 334574
rect 513266 298658 513502 298894
rect 513586 298658 513822 298894
rect 513266 298338 513502 298574
rect 513586 298338 513822 298574
rect 513266 262658 513502 262894
rect 513586 262658 513822 262894
rect 513266 262338 513502 262574
rect 513586 262338 513822 262574
rect 513266 226658 513502 226894
rect 513586 226658 513822 226894
rect 513266 226338 513502 226574
rect 513586 226338 513822 226574
rect 513266 190658 513502 190894
rect 513586 190658 513822 190894
rect 513266 190338 513502 190574
rect 513586 190338 513822 190574
rect 513266 154658 513502 154894
rect 513586 154658 513822 154894
rect 513266 154338 513502 154574
rect 513586 154338 513822 154574
rect 513266 118658 513502 118894
rect 513586 118658 513822 118894
rect 513266 118338 513502 118574
rect 513586 118338 513822 118574
rect 513266 82658 513502 82894
rect 513586 82658 513822 82894
rect 513266 82338 513502 82574
rect 513586 82338 513822 82574
rect 513266 46658 513502 46894
rect 513586 46658 513822 46894
rect 513266 46338 513502 46574
rect 513586 46338 513822 46574
rect 513266 10658 513502 10894
rect 513586 10658 513822 10894
rect 513266 10338 513502 10574
rect 513586 10338 513822 10574
rect 513266 -4422 513502 -4186
rect 513586 -4422 513822 -4186
rect 513266 -4742 513502 -4506
rect 513586 -4742 513822 -4506
rect 534986 711322 535222 711558
rect 535306 711322 535542 711558
rect 534986 711002 535222 711238
rect 535306 711002 535542 711238
rect 531266 709402 531502 709638
rect 531586 709402 531822 709638
rect 531266 709082 531502 709318
rect 531586 709082 531822 709318
rect 527546 707482 527782 707718
rect 527866 707482 528102 707718
rect 527546 707162 527782 707398
rect 527866 707162 528102 707398
rect 516986 698378 517222 698614
rect 517306 698378 517542 698614
rect 516986 698058 517222 698294
rect 517306 698058 517542 698294
rect 516986 662378 517222 662614
rect 517306 662378 517542 662614
rect 516986 662058 517222 662294
rect 517306 662058 517542 662294
rect 516986 626378 517222 626614
rect 517306 626378 517542 626614
rect 516986 626058 517222 626294
rect 517306 626058 517542 626294
rect 516986 590378 517222 590614
rect 517306 590378 517542 590614
rect 516986 590058 517222 590294
rect 517306 590058 517542 590294
rect 516986 554378 517222 554614
rect 517306 554378 517542 554614
rect 516986 554058 517222 554294
rect 517306 554058 517542 554294
rect 516986 518378 517222 518614
rect 517306 518378 517542 518614
rect 516986 518058 517222 518294
rect 517306 518058 517542 518294
rect 516986 482378 517222 482614
rect 517306 482378 517542 482614
rect 516986 482058 517222 482294
rect 517306 482058 517542 482294
rect 516986 446378 517222 446614
rect 517306 446378 517542 446614
rect 516986 446058 517222 446294
rect 517306 446058 517542 446294
rect 516986 410378 517222 410614
rect 517306 410378 517542 410614
rect 516986 410058 517222 410294
rect 517306 410058 517542 410294
rect 516986 374378 517222 374614
rect 517306 374378 517542 374614
rect 516986 374058 517222 374294
rect 517306 374058 517542 374294
rect 516986 338378 517222 338614
rect 517306 338378 517542 338614
rect 516986 338058 517222 338294
rect 517306 338058 517542 338294
rect 516986 302378 517222 302614
rect 517306 302378 517542 302614
rect 516986 302058 517222 302294
rect 517306 302058 517542 302294
rect 516986 266378 517222 266614
rect 517306 266378 517542 266614
rect 516986 266058 517222 266294
rect 517306 266058 517542 266294
rect 516986 230378 517222 230614
rect 517306 230378 517542 230614
rect 516986 230058 517222 230294
rect 517306 230058 517542 230294
rect 516986 194378 517222 194614
rect 517306 194378 517542 194614
rect 516986 194058 517222 194294
rect 517306 194058 517542 194294
rect 516986 158378 517222 158614
rect 517306 158378 517542 158614
rect 516986 158058 517222 158294
rect 517306 158058 517542 158294
rect 516986 122378 517222 122614
rect 517306 122378 517542 122614
rect 516986 122058 517222 122294
rect 517306 122058 517542 122294
rect 516986 86378 517222 86614
rect 517306 86378 517542 86614
rect 516986 86058 517222 86294
rect 517306 86058 517542 86294
rect 516986 50378 517222 50614
rect 517306 50378 517542 50614
rect 516986 50058 517222 50294
rect 517306 50058 517542 50294
rect 516986 14378 517222 14614
rect 517306 14378 517542 14614
rect 516986 14058 517222 14294
rect 517306 14058 517542 14294
rect 498986 -7302 499222 -7066
rect 499306 -7302 499542 -7066
rect 498986 -7622 499222 -7386
rect 499306 -7622 499542 -7386
rect 523826 705562 524062 705798
rect 524146 705562 524382 705798
rect 523826 705242 524062 705478
rect 524146 705242 524382 705478
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -1542 524062 -1306
rect 524146 -1542 524382 -1306
rect 523826 -1862 524062 -1626
rect 524146 -1862 524382 -1626
rect 527546 672938 527782 673174
rect 527866 672938 528102 673174
rect 527546 672618 527782 672854
rect 527866 672618 528102 672854
rect 527546 636938 527782 637174
rect 527866 636938 528102 637174
rect 527546 636618 527782 636854
rect 527866 636618 528102 636854
rect 527546 600938 527782 601174
rect 527866 600938 528102 601174
rect 527546 600618 527782 600854
rect 527866 600618 528102 600854
rect 527546 564938 527782 565174
rect 527866 564938 528102 565174
rect 527546 564618 527782 564854
rect 527866 564618 528102 564854
rect 527546 528938 527782 529174
rect 527866 528938 528102 529174
rect 527546 528618 527782 528854
rect 527866 528618 528102 528854
rect 527546 492938 527782 493174
rect 527866 492938 528102 493174
rect 527546 492618 527782 492854
rect 527866 492618 528102 492854
rect 527546 456938 527782 457174
rect 527866 456938 528102 457174
rect 527546 456618 527782 456854
rect 527866 456618 528102 456854
rect 527546 420938 527782 421174
rect 527866 420938 528102 421174
rect 527546 420618 527782 420854
rect 527866 420618 528102 420854
rect 527546 384938 527782 385174
rect 527866 384938 528102 385174
rect 527546 384618 527782 384854
rect 527866 384618 528102 384854
rect 527546 348938 527782 349174
rect 527866 348938 528102 349174
rect 527546 348618 527782 348854
rect 527866 348618 528102 348854
rect 527546 312938 527782 313174
rect 527866 312938 528102 313174
rect 527546 312618 527782 312854
rect 527866 312618 528102 312854
rect 527546 276938 527782 277174
rect 527866 276938 528102 277174
rect 527546 276618 527782 276854
rect 527866 276618 528102 276854
rect 527546 240938 527782 241174
rect 527866 240938 528102 241174
rect 527546 240618 527782 240854
rect 527866 240618 528102 240854
rect 527546 204938 527782 205174
rect 527866 204938 528102 205174
rect 527546 204618 527782 204854
rect 527866 204618 528102 204854
rect 527546 168938 527782 169174
rect 527866 168938 528102 169174
rect 527546 168618 527782 168854
rect 527866 168618 528102 168854
rect 527546 132938 527782 133174
rect 527866 132938 528102 133174
rect 527546 132618 527782 132854
rect 527866 132618 528102 132854
rect 527546 96938 527782 97174
rect 527866 96938 528102 97174
rect 527546 96618 527782 96854
rect 527866 96618 528102 96854
rect 527546 60938 527782 61174
rect 527866 60938 528102 61174
rect 527546 60618 527782 60854
rect 527866 60618 528102 60854
rect 527546 24938 527782 25174
rect 527866 24938 528102 25174
rect 527546 24618 527782 24854
rect 527866 24618 528102 24854
rect 527546 -3462 527782 -3226
rect 527866 -3462 528102 -3226
rect 527546 -3782 527782 -3546
rect 527866 -3782 528102 -3546
rect 531266 676658 531502 676894
rect 531586 676658 531822 676894
rect 531266 676338 531502 676574
rect 531586 676338 531822 676574
rect 531266 640658 531502 640894
rect 531586 640658 531822 640894
rect 531266 640338 531502 640574
rect 531586 640338 531822 640574
rect 531266 604658 531502 604894
rect 531586 604658 531822 604894
rect 531266 604338 531502 604574
rect 531586 604338 531822 604574
rect 531266 568658 531502 568894
rect 531586 568658 531822 568894
rect 531266 568338 531502 568574
rect 531586 568338 531822 568574
rect 531266 532658 531502 532894
rect 531586 532658 531822 532894
rect 531266 532338 531502 532574
rect 531586 532338 531822 532574
rect 531266 496658 531502 496894
rect 531586 496658 531822 496894
rect 531266 496338 531502 496574
rect 531586 496338 531822 496574
rect 531266 460658 531502 460894
rect 531586 460658 531822 460894
rect 531266 460338 531502 460574
rect 531586 460338 531822 460574
rect 531266 424658 531502 424894
rect 531586 424658 531822 424894
rect 531266 424338 531502 424574
rect 531586 424338 531822 424574
rect 531266 388658 531502 388894
rect 531586 388658 531822 388894
rect 531266 388338 531502 388574
rect 531586 388338 531822 388574
rect 531266 352658 531502 352894
rect 531586 352658 531822 352894
rect 531266 352338 531502 352574
rect 531586 352338 531822 352574
rect 531266 316658 531502 316894
rect 531586 316658 531822 316894
rect 531266 316338 531502 316574
rect 531586 316338 531822 316574
rect 531266 280658 531502 280894
rect 531586 280658 531822 280894
rect 531266 280338 531502 280574
rect 531586 280338 531822 280574
rect 531266 244658 531502 244894
rect 531586 244658 531822 244894
rect 531266 244338 531502 244574
rect 531586 244338 531822 244574
rect 531266 208658 531502 208894
rect 531586 208658 531822 208894
rect 531266 208338 531502 208574
rect 531586 208338 531822 208574
rect 531266 172658 531502 172894
rect 531586 172658 531822 172894
rect 531266 172338 531502 172574
rect 531586 172338 531822 172574
rect 531266 136658 531502 136894
rect 531586 136658 531822 136894
rect 531266 136338 531502 136574
rect 531586 136338 531822 136574
rect 531266 100658 531502 100894
rect 531586 100658 531822 100894
rect 531266 100338 531502 100574
rect 531586 100338 531822 100574
rect 531266 64658 531502 64894
rect 531586 64658 531822 64894
rect 531266 64338 531502 64574
rect 531586 64338 531822 64574
rect 531266 28658 531502 28894
rect 531586 28658 531822 28894
rect 531266 28338 531502 28574
rect 531586 28338 531822 28574
rect 531266 -5382 531502 -5146
rect 531586 -5382 531822 -5146
rect 531266 -5702 531502 -5466
rect 531586 -5702 531822 -5466
rect 552986 710362 553222 710598
rect 553306 710362 553542 710598
rect 552986 710042 553222 710278
rect 553306 710042 553542 710278
rect 549266 708442 549502 708678
rect 549586 708442 549822 708678
rect 549266 708122 549502 708358
rect 549586 708122 549822 708358
rect 545546 706522 545782 706758
rect 545866 706522 546102 706758
rect 545546 706202 545782 706438
rect 545866 706202 546102 706438
rect 534986 680378 535222 680614
rect 535306 680378 535542 680614
rect 534986 680058 535222 680294
rect 535306 680058 535542 680294
rect 534986 644378 535222 644614
rect 535306 644378 535542 644614
rect 534986 644058 535222 644294
rect 535306 644058 535542 644294
rect 534986 608378 535222 608614
rect 535306 608378 535542 608614
rect 534986 608058 535222 608294
rect 535306 608058 535542 608294
rect 534986 572378 535222 572614
rect 535306 572378 535542 572614
rect 534986 572058 535222 572294
rect 535306 572058 535542 572294
rect 534986 536378 535222 536614
rect 535306 536378 535542 536614
rect 534986 536058 535222 536294
rect 535306 536058 535542 536294
rect 534986 500378 535222 500614
rect 535306 500378 535542 500614
rect 534986 500058 535222 500294
rect 535306 500058 535542 500294
rect 534986 464378 535222 464614
rect 535306 464378 535542 464614
rect 534986 464058 535222 464294
rect 535306 464058 535542 464294
rect 534986 428378 535222 428614
rect 535306 428378 535542 428614
rect 534986 428058 535222 428294
rect 535306 428058 535542 428294
rect 534986 392378 535222 392614
rect 535306 392378 535542 392614
rect 534986 392058 535222 392294
rect 535306 392058 535542 392294
rect 534986 356378 535222 356614
rect 535306 356378 535542 356614
rect 534986 356058 535222 356294
rect 535306 356058 535542 356294
rect 534986 320378 535222 320614
rect 535306 320378 535542 320614
rect 534986 320058 535222 320294
rect 535306 320058 535542 320294
rect 534986 284378 535222 284614
rect 535306 284378 535542 284614
rect 534986 284058 535222 284294
rect 535306 284058 535542 284294
rect 534986 248378 535222 248614
rect 535306 248378 535542 248614
rect 534986 248058 535222 248294
rect 535306 248058 535542 248294
rect 534986 212378 535222 212614
rect 535306 212378 535542 212614
rect 534986 212058 535222 212294
rect 535306 212058 535542 212294
rect 534986 176378 535222 176614
rect 535306 176378 535542 176614
rect 534986 176058 535222 176294
rect 535306 176058 535542 176294
rect 534986 140378 535222 140614
rect 535306 140378 535542 140614
rect 534986 140058 535222 140294
rect 535306 140058 535542 140294
rect 534986 104378 535222 104614
rect 535306 104378 535542 104614
rect 534986 104058 535222 104294
rect 535306 104058 535542 104294
rect 534986 68378 535222 68614
rect 535306 68378 535542 68614
rect 534986 68058 535222 68294
rect 535306 68058 535542 68294
rect 534986 32378 535222 32614
rect 535306 32378 535542 32614
rect 534986 32058 535222 32294
rect 535306 32058 535542 32294
rect 516986 -6342 517222 -6106
rect 517306 -6342 517542 -6106
rect 516986 -6662 517222 -6426
rect 517306 -6662 517542 -6426
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 545546 690938 545782 691174
rect 545866 690938 546102 691174
rect 545546 690618 545782 690854
rect 545866 690618 546102 690854
rect 545546 654938 545782 655174
rect 545866 654938 546102 655174
rect 545546 654618 545782 654854
rect 545866 654618 546102 654854
rect 545546 618938 545782 619174
rect 545866 618938 546102 619174
rect 545546 618618 545782 618854
rect 545866 618618 546102 618854
rect 545546 582938 545782 583174
rect 545866 582938 546102 583174
rect 545546 582618 545782 582854
rect 545866 582618 546102 582854
rect 545546 546938 545782 547174
rect 545866 546938 546102 547174
rect 545546 546618 545782 546854
rect 545866 546618 546102 546854
rect 545546 510938 545782 511174
rect 545866 510938 546102 511174
rect 545546 510618 545782 510854
rect 545866 510618 546102 510854
rect 545546 474938 545782 475174
rect 545866 474938 546102 475174
rect 545546 474618 545782 474854
rect 545866 474618 546102 474854
rect 545546 438938 545782 439174
rect 545866 438938 546102 439174
rect 545546 438618 545782 438854
rect 545866 438618 546102 438854
rect 545546 402938 545782 403174
rect 545866 402938 546102 403174
rect 545546 402618 545782 402854
rect 545866 402618 546102 402854
rect 545546 366938 545782 367174
rect 545866 366938 546102 367174
rect 545546 366618 545782 366854
rect 545866 366618 546102 366854
rect 545546 330938 545782 331174
rect 545866 330938 546102 331174
rect 545546 330618 545782 330854
rect 545866 330618 546102 330854
rect 545546 294938 545782 295174
rect 545866 294938 546102 295174
rect 545546 294618 545782 294854
rect 545866 294618 546102 294854
rect 545546 258938 545782 259174
rect 545866 258938 546102 259174
rect 545546 258618 545782 258854
rect 545866 258618 546102 258854
rect 545546 222938 545782 223174
rect 545866 222938 546102 223174
rect 545546 222618 545782 222854
rect 545866 222618 546102 222854
rect 545546 186938 545782 187174
rect 545866 186938 546102 187174
rect 545546 186618 545782 186854
rect 545866 186618 546102 186854
rect 545546 150938 545782 151174
rect 545866 150938 546102 151174
rect 545546 150618 545782 150854
rect 545866 150618 546102 150854
rect 545546 114938 545782 115174
rect 545866 114938 546102 115174
rect 545546 114618 545782 114854
rect 545866 114618 546102 114854
rect 545546 78938 545782 79174
rect 545866 78938 546102 79174
rect 545546 78618 545782 78854
rect 545866 78618 546102 78854
rect 545546 42938 545782 43174
rect 545866 42938 546102 43174
rect 545546 42618 545782 42854
rect 545866 42618 546102 42854
rect 545546 6938 545782 7174
rect 545866 6938 546102 7174
rect 545546 6618 545782 6854
rect 545866 6618 546102 6854
rect 545546 -2502 545782 -2266
rect 545866 -2502 546102 -2266
rect 545546 -2822 545782 -2586
rect 545866 -2822 546102 -2586
rect 549266 694658 549502 694894
rect 549586 694658 549822 694894
rect 549266 694338 549502 694574
rect 549586 694338 549822 694574
rect 549266 658658 549502 658894
rect 549586 658658 549822 658894
rect 549266 658338 549502 658574
rect 549586 658338 549822 658574
rect 549266 622658 549502 622894
rect 549586 622658 549822 622894
rect 549266 622338 549502 622574
rect 549586 622338 549822 622574
rect 549266 586658 549502 586894
rect 549586 586658 549822 586894
rect 549266 586338 549502 586574
rect 549586 586338 549822 586574
rect 549266 550658 549502 550894
rect 549586 550658 549822 550894
rect 549266 550338 549502 550574
rect 549586 550338 549822 550574
rect 549266 514658 549502 514894
rect 549586 514658 549822 514894
rect 549266 514338 549502 514574
rect 549586 514338 549822 514574
rect 549266 478658 549502 478894
rect 549586 478658 549822 478894
rect 549266 478338 549502 478574
rect 549586 478338 549822 478574
rect 549266 442658 549502 442894
rect 549586 442658 549822 442894
rect 549266 442338 549502 442574
rect 549586 442338 549822 442574
rect 549266 406658 549502 406894
rect 549586 406658 549822 406894
rect 549266 406338 549502 406574
rect 549586 406338 549822 406574
rect 549266 370658 549502 370894
rect 549586 370658 549822 370894
rect 549266 370338 549502 370574
rect 549586 370338 549822 370574
rect 549266 334658 549502 334894
rect 549586 334658 549822 334894
rect 549266 334338 549502 334574
rect 549586 334338 549822 334574
rect 549266 298658 549502 298894
rect 549586 298658 549822 298894
rect 549266 298338 549502 298574
rect 549586 298338 549822 298574
rect 549266 262658 549502 262894
rect 549586 262658 549822 262894
rect 549266 262338 549502 262574
rect 549586 262338 549822 262574
rect 549266 226658 549502 226894
rect 549586 226658 549822 226894
rect 549266 226338 549502 226574
rect 549586 226338 549822 226574
rect 549266 190658 549502 190894
rect 549586 190658 549822 190894
rect 549266 190338 549502 190574
rect 549586 190338 549822 190574
rect 549266 154658 549502 154894
rect 549586 154658 549822 154894
rect 549266 154338 549502 154574
rect 549586 154338 549822 154574
rect 549266 118658 549502 118894
rect 549586 118658 549822 118894
rect 549266 118338 549502 118574
rect 549586 118338 549822 118574
rect 549266 82658 549502 82894
rect 549586 82658 549822 82894
rect 549266 82338 549502 82574
rect 549586 82338 549822 82574
rect 549266 46658 549502 46894
rect 549586 46658 549822 46894
rect 549266 46338 549502 46574
rect 549586 46338 549822 46574
rect 549266 10658 549502 10894
rect 549586 10658 549822 10894
rect 549266 10338 549502 10574
rect 549586 10338 549822 10574
rect 549266 -4422 549502 -4186
rect 549586 -4422 549822 -4186
rect 549266 -4742 549502 -4506
rect 549586 -4742 549822 -4506
rect 570986 711322 571222 711558
rect 571306 711322 571542 711558
rect 570986 711002 571222 711238
rect 571306 711002 571542 711238
rect 567266 709402 567502 709638
rect 567586 709402 567822 709638
rect 567266 709082 567502 709318
rect 567586 709082 567822 709318
rect 563546 707482 563782 707718
rect 563866 707482 564102 707718
rect 563546 707162 563782 707398
rect 563866 707162 564102 707398
rect 552986 698378 553222 698614
rect 553306 698378 553542 698614
rect 552986 698058 553222 698294
rect 553306 698058 553542 698294
rect 552986 662378 553222 662614
rect 553306 662378 553542 662614
rect 552986 662058 553222 662294
rect 553306 662058 553542 662294
rect 552986 626378 553222 626614
rect 553306 626378 553542 626614
rect 552986 626058 553222 626294
rect 553306 626058 553542 626294
rect 552986 590378 553222 590614
rect 553306 590378 553542 590614
rect 552986 590058 553222 590294
rect 553306 590058 553542 590294
rect 552986 554378 553222 554614
rect 553306 554378 553542 554614
rect 552986 554058 553222 554294
rect 553306 554058 553542 554294
rect 552986 518378 553222 518614
rect 553306 518378 553542 518614
rect 552986 518058 553222 518294
rect 553306 518058 553542 518294
rect 552986 482378 553222 482614
rect 553306 482378 553542 482614
rect 552986 482058 553222 482294
rect 553306 482058 553542 482294
rect 552986 446378 553222 446614
rect 553306 446378 553542 446614
rect 552986 446058 553222 446294
rect 553306 446058 553542 446294
rect 552986 410378 553222 410614
rect 553306 410378 553542 410614
rect 552986 410058 553222 410294
rect 553306 410058 553542 410294
rect 552986 374378 553222 374614
rect 553306 374378 553542 374614
rect 552986 374058 553222 374294
rect 553306 374058 553542 374294
rect 552986 338378 553222 338614
rect 553306 338378 553542 338614
rect 552986 338058 553222 338294
rect 553306 338058 553542 338294
rect 552986 302378 553222 302614
rect 553306 302378 553542 302614
rect 552986 302058 553222 302294
rect 553306 302058 553542 302294
rect 552986 266378 553222 266614
rect 553306 266378 553542 266614
rect 552986 266058 553222 266294
rect 553306 266058 553542 266294
rect 552986 230378 553222 230614
rect 553306 230378 553542 230614
rect 552986 230058 553222 230294
rect 553306 230058 553542 230294
rect 552986 194378 553222 194614
rect 553306 194378 553542 194614
rect 552986 194058 553222 194294
rect 553306 194058 553542 194294
rect 552986 158378 553222 158614
rect 553306 158378 553542 158614
rect 552986 158058 553222 158294
rect 553306 158058 553542 158294
rect 552986 122378 553222 122614
rect 553306 122378 553542 122614
rect 552986 122058 553222 122294
rect 553306 122058 553542 122294
rect 552986 86378 553222 86614
rect 553306 86378 553542 86614
rect 552986 86058 553222 86294
rect 553306 86058 553542 86294
rect 552986 50378 553222 50614
rect 553306 50378 553542 50614
rect 552986 50058 553222 50294
rect 553306 50058 553542 50294
rect 552986 14378 553222 14614
rect 553306 14378 553542 14614
rect 552986 14058 553222 14294
rect 553306 14058 553542 14294
rect 534986 -7302 535222 -7066
rect 535306 -7302 535542 -7066
rect 534986 -7622 535222 -7386
rect 535306 -7622 535542 -7386
rect 559826 705562 560062 705798
rect 560146 705562 560382 705798
rect 559826 705242 560062 705478
rect 560146 705242 560382 705478
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -1542 560062 -1306
rect 560146 -1542 560382 -1306
rect 559826 -1862 560062 -1626
rect 560146 -1862 560382 -1626
rect 563546 672938 563782 673174
rect 563866 672938 564102 673174
rect 563546 672618 563782 672854
rect 563866 672618 564102 672854
rect 563546 636938 563782 637174
rect 563866 636938 564102 637174
rect 563546 636618 563782 636854
rect 563866 636618 564102 636854
rect 563546 600938 563782 601174
rect 563866 600938 564102 601174
rect 563546 600618 563782 600854
rect 563866 600618 564102 600854
rect 563546 564938 563782 565174
rect 563866 564938 564102 565174
rect 563546 564618 563782 564854
rect 563866 564618 564102 564854
rect 563546 528938 563782 529174
rect 563866 528938 564102 529174
rect 563546 528618 563782 528854
rect 563866 528618 564102 528854
rect 563546 492938 563782 493174
rect 563866 492938 564102 493174
rect 563546 492618 563782 492854
rect 563866 492618 564102 492854
rect 563546 456938 563782 457174
rect 563866 456938 564102 457174
rect 563546 456618 563782 456854
rect 563866 456618 564102 456854
rect 563546 420938 563782 421174
rect 563866 420938 564102 421174
rect 563546 420618 563782 420854
rect 563866 420618 564102 420854
rect 563546 384938 563782 385174
rect 563866 384938 564102 385174
rect 563546 384618 563782 384854
rect 563866 384618 564102 384854
rect 563546 348938 563782 349174
rect 563866 348938 564102 349174
rect 563546 348618 563782 348854
rect 563866 348618 564102 348854
rect 563546 312938 563782 313174
rect 563866 312938 564102 313174
rect 563546 312618 563782 312854
rect 563866 312618 564102 312854
rect 563546 276938 563782 277174
rect 563866 276938 564102 277174
rect 563546 276618 563782 276854
rect 563866 276618 564102 276854
rect 563546 240938 563782 241174
rect 563866 240938 564102 241174
rect 563546 240618 563782 240854
rect 563866 240618 564102 240854
rect 563546 204938 563782 205174
rect 563866 204938 564102 205174
rect 563546 204618 563782 204854
rect 563866 204618 564102 204854
rect 563546 168938 563782 169174
rect 563866 168938 564102 169174
rect 563546 168618 563782 168854
rect 563866 168618 564102 168854
rect 563546 132938 563782 133174
rect 563866 132938 564102 133174
rect 563546 132618 563782 132854
rect 563866 132618 564102 132854
rect 563546 96938 563782 97174
rect 563866 96938 564102 97174
rect 563546 96618 563782 96854
rect 563866 96618 564102 96854
rect 563546 60938 563782 61174
rect 563866 60938 564102 61174
rect 563546 60618 563782 60854
rect 563866 60618 564102 60854
rect 563546 24938 563782 25174
rect 563866 24938 564102 25174
rect 563546 24618 563782 24854
rect 563866 24618 564102 24854
rect 563546 -3462 563782 -3226
rect 563866 -3462 564102 -3226
rect 563546 -3782 563782 -3546
rect 563866 -3782 564102 -3546
rect 567266 676658 567502 676894
rect 567586 676658 567822 676894
rect 567266 676338 567502 676574
rect 567586 676338 567822 676574
rect 567266 640658 567502 640894
rect 567586 640658 567822 640894
rect 567266 640338 567502 640574
rect 567586 640338 567822 640574
rect 567266 604658 567502 604894
rect 567586 604658 567822 604894
rect 567266 604338 567502 604574
rect 567586 604338 567822 604574
rect 567266 568658 567502 568894
rect 567586 568658 567822 568894
rect 567266 568338 567502 568574
rect 567586 568338 567822 568574
rect 567266 532658 567502 532894
rect 567586 532658 567822 532894
rect 567266 532338 567502 532574
rect 567586 532338 567822 532574
rect 567266 496658 567502 496894
rect 567586 496658 567822 496894
rect 567266 496338 567502 496574
rect 567586 496338 567822 496574
rect 567266 460658 567502 460894
rect 567586 460658 567822 460894
rect 567266 460338 567502 460574
rect 567586 460338 567822 460574
rect 567266 424658 567502 424894
rect 567586 424658 567822 424894
rect 567266 424338 567502 424574
rect 567586 424338 567822 424574
rect 567266 388658 567502 388894
rect 567586 388658 567822 388894
rect 567266 388338 567502 388574
rect 567586 388338 567822 388574
rect 567266 352658 567502 352894
rect 567586 352658 567822 352894
rect 567266 352338 567502 352574
rect 567586 352338 567822 352574
rect 567266 316658 567502 316894
rect 567586 316658 567822 316894
rect 567266 316338 567502 316574
rect 567586 316338 567822 316574
rect 567266 280658 567502 280894
rect 567586 280658 567822 280894
rect 567266 280338 567502 280574
rect 567586 280338 567822 280574
rect 567266 244658 567502 244894
rect 567586 244658 567822 244894
rect 567266 244338 567502 244574
rect 567586 244338 567822 244574
rect 567266 208658 567502 208894
rect 567586 208658 567822 208894
rect 567266 208338 567502 208574
rect 567586 208338 567822 208574
rect 567266 172658 567502 172894
rect 567586 172658 567822 172894
rect 567266 172338 567502 172574
rect 567586 172338 567822 172574
rect 567266 136658 567502 136894
rect 567586 136658 567822 136894
rect 567266 136338 567502 136574
rect 567586 136338 567822 136574
rect 567266 100658 567502 100894
rect 567586 100658 567822 100894
rect 567266 100338 567502 100574
rect 567586 100338 567822 100574
rect 567266 64658 567502 64894
rect 567586 64658 567822 64894
rect 567266 64338 567502 64574
rect 567586 64338 567822 64574
rect 567266 28658 567502 28894
rect 567586 28658 567822 28894
rect 567266 28338 567502 28574
rect 567586 28338 567822 28574
rect 567266 -5382 567502 -5146
rect 567586 -5382 567822 -5146
rect 567266 -5702 567502 -5466
rect 567586 -5702 567822 -5466
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 581546 706522 581782 706758
rect 581866 706522 582102 706758
rect 581546 706202 581782 706438
rect 581866 706202 582102 706438
rect 570986 680378 571222 680614
rect 571306 680378 571542 680614
rect 570986 680058 571222 680294
rect 571306 680058 571542 680294
rect 570986 644378 571222 644614
rect 571306 644378 571542 644614
rect 570986 644058 571222 644294
rect 571306 644058 571542 644294
rect 570986 608378 571222 608614
rect 571306 608378 571542 608614
rect 570986 608058 571222 608294
rect 571306 608058 571542 608294
rect 570986 572378 571222 572614
rect 571306 572378 571542 572614
rect 570986 572058 571222 572294
rect 571306 572058 571542 572294
rect 570986 536378 571222 536614
rect 571306 536378 571542 536614
rect 570986 536058 571222 536294
rect 571306 536058 571542 536294
rect 570986 500378 571222 500614
rect 571306 500378 571542 500614
rect 570986 500058 571222 500294
rect 571306 500058 571542 500294
rect 570986 464378 571222 464614
rect 571306 464378 571542 464614
rect 570986 464058 571222 464294
rect 571306 464058 571542 464294
rect 570986 428378 571222 428614
rect 571306 428378 571542 428614
rect 570986 428058 571222 428294
rect 571306 428058 571542 428294
rect 570986 392378 571222 392614
rect 571306 392378 571542 392614
rect 570986 392058 571222 392294
rect 571306 392058 571542 392294
rect 570986 356378 571222 356614
rect 571306 356378 571542 356614
rect 570986 356058 571222 356294
rect 571306 356058 571542 356294
rect 570986 320378 571222 320614
rect 571306 320378 571542 320614
rect 570986 320058 571222 320294
rect 571306 320058 571542 320294
rect 570986 284378 571222 284614
rect 571306 284378 571542 284614
rect 570986 284058 571222 284294
rect 571306 284058 571542 284294
rect 570986 248378 571222 248614
rect 571306 248378 571542 248614
rect 570986 248058 571222 248294
rect 571306 248058 571542 248294
rect 570986 212378 571222 212614
rect 571306 212378 571542 212614
rect 570986 212058 571222 212294
rect 571306 212058 571542 212294
rect 570986 176378 571222 176614
rect 571306 176378 571542 176614
rect 570986 176058 571222 176294
rect 571306 176058 571542 176294
rect 570986 140378 571222 140614
rect 571306 140378 571542 140614
rect 570986 140058 571222 140294
rect 571306 140058 571542 140294
rect 570986 104378 571222 104614
rect 571306 104378 571542 104614
rect 570986 104058 571222 104294
rect 571306 104058 571542 104294
rect 570986 68378 571222 68614
rect 571306 68378 571542 68614
rect 570986 68058 571222 68294
rect 571306 68058 571542 68294
rect 570986 32378 571222 32614
rect 571306 32378 571542 32614
rect 570986 32058 571222 32294
rect 571306 32058 571542 32294
rect 552986 -6342 553222 -6106
rect 553306 -6342 553542 -6106
rect 552986 -6662 553222 -6426
rect 553306 -6662 553542 -6426
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581546 690938 581782 691174
rect 581866 690938 582102 691174
rect 581546 690618 581782 690854
rect 581866 690618 582102 690854
rect 581546 654938 581782 655174
rect 581866 654938 582102 655174
rect 581546 654618 581782 654854
rect 581866 654618 582102 654854
rect 581546 618938 581782 619174
rect 581866 618938 582102 619174
rect 581546 618618 581782 618854
rect 581866 618618 582102 618854
rect 581546 582938 581782 583174
rect 581866 582938 582102 583174
rect 581546 582618 581782 582854
rect 581866 582618 582102 582854
rect 581546 546938 581782 547174
rect 581866 546938 582102 547174
rect 581546 546618 581782 546854
rect 581866 546618 582102 546854
rect 581546 510938 581782 511174
rect 581866 510938 582102 511174
rect 581546 510618 581782 510854
rect 581866 510618 582102 510854
rect 581546 474938 581782 475174
rect 581866 474938 582102 475174
rect 581546 474618 581782 474854
rect 581866 474618 582102 474854
rect 581546 438938 581782 439174
rect 581866 438938 582102 439174
rect 581546 438618 581782 438854
rect 581866 438618 582102 438854
rect 581546 402938 581782 403174
rect 581866 402938 582102 403174
rect 581546 402618 581782 402854
rect 581866 402618 582102 402854
rect 581546 366938 581782 367174
rect 581866 366938 582102 367174
rect 581546 366618 581782 366854
rect 581866 366618 582102 366854
rect 581546 330938 581782 331174
rect 581866 330938 582102 331174
rect 581546 330618 581782 330854
rect 581866 330618 582102 330854
rect 581546 294938 581782 295174
rect 581866 294938 582102 295174
rect 581546 294618 581782 294854
rect 581866 294618 582102 294854
rect 581546 258938 581782 259174
rect 581866 258938 582102 259174
rect 581546 258618 581782 258854
rect 581866 258618 582102 258854
rect 581546 222938 581782 223174
rect 581866 222938 582102 223174
rect 581546 222618 581782 222854
rect 581866 222618 582102 222854
rect 581546 186938 581782 187174
rect 581866 186938 582102 187174
rect 581546 186618 581782 186854
rect 581866 186618 582102 186854
rect 581546 150938 581782 151174
rect 581866 150938 582102 151174
rect 581546 150618 581782 150854
rect 581866 150618 582102 150854
rect 581546 114938 581782 115174
rect 581866 114938 582102 115174
rect 581546 114618 581782 114854
rect 581866 114618 582102 114854
rect 581546 78938 581782 79174
rect 581866 78938 582102 79174
rect 581546 78618 581782 78854
rect 581866 78618 582102 78854
rect 581546 42938 581782 43174
rect 581866 42938 582102 43174
rect 581546 42618 581782 42854
rect 581866 42618 582102 42854
rect 581546 6938 581782 7174
rect 581866 6938 582102 7174
rect 581546 6618 581782 6854
rect 581866 6618 582102 6854
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 669218 586538 669454
rect 586622 669218 586858 669454
rect 586302 668898 586538 669134
rect 586622 668898 586858 669134
rect 586302 633218 586538 633454
rect 586622 633218 586858 633454
rect 586302 632898 586538 633134
rect 586622 632898 586858 633134
rect 586302 597218 586538 597454
rect 586622 597218 586858 597454
rect 586302 596898 586538 597134
rect 586622 596898 586858 597134
rect 586302 561218 586538 561454
rect 586622 561218 586858 561454
rect 586302 560898 586538 561134
rect 586622 560898 586858 561134
rect 586302 525218 586538 525454
rect 586622 525218 586858 525454
rect 586302 524898 586538 525134
rect 586622 524898 586858 525134
rect 586302 489218 586538 489454
rect 586622 489218 586858 489454
rect 586302 488898 586538 489134
rect 586622 488898 586858 489134
rect 586302 453218 586538 453454
rect 586622 453218 586858 453454
rect 586302 452898 586538 453134
rect 586622 452898 586858 453134
rect 586302 417218 586538 417454
rect 586622 417218 586858 417454
rect 586302 416898 586538 417134
rect 586622 416898 586858 417134
rect 586302 381218 586538 381454
rect 586622 381218 586858 381454
rect 586302 380898 586538 381134
rect 586622 380898 586858 381134
rect 586302 345218 586538 345454
rect 586622 345218 586858 345454
rect 586302 344898 586538 345134
rect 586622 344898 586858 345134
rect 586302 309218 586538 309454
rect 586622 309218 586858 309454
rect 586302 308898 586538 309134
rect 586622 308898 586858 309134
rect 586302 273218 586538 273454
rect 586622 273218 586858 273454
rect 586302 272898 586538 273134
rect 586622 272898 586858 273134
rect 586302 237218 586538 237454
rect 586622 237218 586858 237454
rect 586302 236898 586538 237134
rect 586622 236898 586858 237134
rect 586302 201218 586538 201454
rect 586622 201218 586858 201454
rect 586302 200898 586538 201134
rect 586622 200898 586858 201134
rect 586302 165218 586538 165454
rect 586622 165218 586858 165454
rect 586302 164898 586538 165134
rect 586622 164898 586858 165134
rect 586302 129218 586538 129454
rect 586622 129218 586858 129454
rect 586302 128898 586538 129134
rect 586622 128898 586858 129134
rect 586302 93218 586538 93454
rect 586622 93218 586858 93454
rect 586302 92898 586538 93134
rect 586622 92898 586858 93134
rect 586302 57218 586538 57454
rect 586622 57218 586858 57454
rect 586302 56898 586538 57134
rect 586622 56898 586858 57134
rect 586302 21218 586538 21454
rect 586622 21218 586858 21454
rect 586302 20898 586538 21134
rect 586622 20898 586858 21134
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 690938 587498 691174
rect 587582 690938 587818 691174
rect 587262 690618 587498 690854
rect 587582 690618 587818 690854
rect 587262 654938 587498 655174
rect 587582 654938 587818 655174
rect 587262 654618 587498 654854
rect 587582 654618 587818 654854
rect 587262 618938 587498 619174
rect 587582 618938 587818 619174
rect 587262 618618 587498 618854
rect 587582 618618 587818 618854
rect 587262 582938 587498 583174
rect 587582 582938 587818 583174
rect 587262 582618 587498 582854
rect 587582 582618 587818 582854
rect 587262 546938 587498 547174
rect 587582 546938 587818 547174
rect 587262 546618 587498 546854
rect 587582 546618 587818 546854
rect 587262 510938 587498 511174
rect 587582 510938 587818 511174
rect 587262 510618 587498 510854
rect 587582 510618 587818 510854
rect 587262 474938 587498 475174
rect 587582 474938 587818 475174
rect 587262 474618 587498 474854
rect 587582 474618 587818 474854
rect 587262 438938 587498 439174
rect 587582 438938 587818 439174
rect 587262 438618 587498 438854
rect 587582 438618 587818 438854
rect 587262 402938 587498 403174
rect 587582 402938 587818 403174
rect 587262 402618 587498 402854
rect 587582 402618 587818 402854
rect 587262 366938 587498 367174
rect 587582 366938 587818 367174
rect 587262 366618 587498 366854
rect 587582 366618 587818 366854
rect 587262 330938 587498 331174
rect 587582 330938 587818 331174
rect 587262 330618 587498 330854
rect 587582 330618 587818 330854
rect 587262 294938 587498 295174
rect 587582 294938 587818 295174
rect 587262 294618 587498 294854
rect 587582 294618 587818 294854
rect 587262 258938 587498 259174
rect 587582 258938 587818 259174
rect 587262 258618 587498 258854
rect 587582 258618 587818 258854
rect 587262 222938 587498 223174
rect 587582 222938 587818 223174
rect 587262 222618 587498 222854
rect 587582 222618 587818 222854
rect 587262 186938 587498 187174
rect 587582 186938 587818 187174
rect 587262 186618 587498 186854
rect 587582 186618 587818 186854
rect 587262 150938 587498 151174
rect 587582 150938 587818 151174
rect 587262 150618 587498 150854
rect 587582 150618 587818 150854
rect 587262 114938 587498 115174
rect 587582 114938 587818 115174
rect 587262 114618 587498 114854
rect 587582 114618 587818 114854
rect 587262 78938 587498 79174
rect 587582 78938 587818 79174
rect 587262 78618 587498 78854
rect 587582 78618 587818 78854
rect 587262 42938 587498 43174
rect 587582 42938 587818 43174
rect 587262 42618 587498 42854
rect 587582 42618 587818 42854
rect 587262 6938 587498 7174
rect 587582 6938 587818 7174
rect 587262 6618 587498 6854
rect 587582 6618 587818 6854
rect 581546 -2502 581782 -2266
rect 581866 -2502 582102 -2266
rect 581546 -2822 581782 -2586
rect 581866 -2822 582102 -2586
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 672938 588458 673174
rect 588542 672938 588778 673174
rect 588222 672618 588458 672854
rect 588542 672618 588778 672854
rect 588222 636938 588458 637174
rect 588542 636938 588778 637174
rect 588222 636618 588458 636854
rect 588542 636618 588778 636854
rect 588222 600938 588458 601174
rect 588542 600938 588778 601174
rect 588222 600618 588458 600854
rect 588542 600618 588778 600854
rect 588222 564938 588458 565174
rect 588542 564938 588778 565174
rect 588222 564618 588458 564854
rect 588542 564618 588778 564854
rect 588222 528938 588458 529174
rect 588542 528938 588778 529174
rect 588222 528618 588458 528854
rect 588542 528618 588778 528854
rect 588222 492938 588458 493174
rect 588542 492938 588778 493174
rect 588222 492618 588458 492854
rect 588542 492618 588778 492854
rect 588222 456938 588458 457174
rect 588542 456938 588778 457174
rect 588222 456618 588458 456854
rect 588542 456618 588778 456854
rect 588222 420938 588458 421174
rect 588542 420938 588778 421174
rect 588222 420618 588458 420854
rect 588542 420618 588778 420854
rect 588222 384938 588458 385174
rect 588542 384938 588778 385174
rect 588222 384618 588458 384854
rect 588542 384618 588778 384854
rect 588222 348938 588458 349174
rect 588542 348938 588778 349174
rect 588222 348618 588458 348854
rect 588542 348618 588778 348854
rect 588222 312938 588458 313174
rect 588542 312938 588778 313174
rect 588222 312618 588458 312854
rect 588542 312618 588778 312854
rect 588222 276938 588458 277174
rect 588542 276938 588778 277174
rect 588222 276618 588458 276854
rect 588542 276618 588778 276854
rect 588222 240938 588458 241174
rect 588542 240938 588778 241174
rect 588222 240618 588458 240854
rect 588542 240618 588778 240854
rect 588222 204938 588458 205174
rect 588542 204938 588778 205174
rect 588222 204618 588458 204854
rect 588542 204618 588778 204854
rect 588222 168938 588458 169174
rect 588542 168938 588778 169174
rect 588222 168618 588458 168854
rect 588542 168618 588778 168854
rect 588222 132938 588458 133174
rect 588542 132938 588778 133174
rect 588222 132618 588458 132854
rect 588542 132618 588778 132854
rect 588222 96938 588458 97174
rect 588542 96938 588778 97174
rect 588222 96618 588458 96854
rect 588542 96618 588778 96854
rect 588222 60938 588458 61174
rect 588542 60938 588778 61174
rect 588222 60618 588458 60854
rect 588542 60618 588778 60854
rect 588222 24938 588458 25174
rect 588542 24938 588778 25174
rect 588222 24618 588458 24854
rect 588542 24618 588778 24854
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 694658 589418 694894
rect 589502 694658 589738 694894
rect 589182 694338 589418 694574
rect 589502 694338 589738 694574
rect 589182 658658 589418 658894
rect 589502 658658 589738 658894
rect 589182 658338 589418 658574
rect 589502 658338 589738 658574
rect 589182 622658 589418 622894
rect 589502 622658 589738 622894
rect 589182 622338 589418 622574
rect 589502 622338 589738 622574
rect 589182 586658 589418 586894
rect 589502 586658 589738 586894
rect 589182 586338 589418 586574
rect 589502 586338 589738 586574
rect 589182 550658 589418 550894
rect 589502 550658 589738 550894
rect 589182 550338 589418 550574
rect 589502 550338 589738 550574
rect 589182 514658 589418 514894
rect 589502 514658 589738 514894
rect 589182 514338 589418 514574
rect 589502 514338 589738 514574
rect 589182 478658 589418 478894
rect 589502 478658 589738 478894
rect 589182 478338 589418 478574
rect 589502 478338 589738 478574
rect 589182 442658 589418 442894
rect 589502 442658 589738 442894
rect 589182 442338 589418 442574
rect 589502 442338 589738 442574
rect 589182 406658 589418 406894
rect 589502 406658 589738 406894
rect 589182 406338 589418 406574
rect 589502 406338 589738 406574
rect 589182 370658 589418 370894
rect 589502 370658 589738 370894
rect 589182 370338 589418 370574
rect 589502 370338 589738 370574
rect 589182 334658 589418 334894
rect 589502 334658 589738 334894
rect 589182 334338 589418 334574
rect 589502 334338 589738 334574
rect 589182 298658 589418 298894
rect 589502 298658 589738 298894
rect 589182 298338 589418 298574
rect 589502 298338 589738 298574
rect 589182 262658 589418 262894
rect 589502 262658 589738 262894
rect 589182 262338 589418 262574
rect 589502 262338 589738 262574
rect 589182 226658 589418 226894
rect 589502 226658 589738 226894
rect 589182 226338 589418 226574
rect 589502 226338 589738 226574
rect 589182 190658 589418 190894
rect 589502 190658 589738 190894
rect 589182 190338 589418 190574
rect 589502 190338 589738 190574
rect 589182 154658 589418 154894
rect 589502 154658 589738 154894
rect 589182 154338 589418 154574
rect 589502 154338 589738 154574
rect 589182 118658 589418 118894
rect 589502 118658 589738 118894
rect 589182 118338 589418 118574
rect 589502 118338 589738 118574
rect 589182 82658 589418 82894
rect 589502 82658 589738 82894
rect 589182 82338 589418 82574
rect 589502 82338 589738 82574
rect 589182 46658 589418 46894
rect 589502 46658 589738 46894
rect 589182 46338 589418 46574
rect 589502 46338 589738 46574
rect 589182 10658 589418 10894
rect 589502 10658 589738 10894
rect 589182 10338 589418 10574
rect 589502 10338 589738 10574
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 676658 590378 676894
rect 590462 676658 590698 676894
rect 590142 676338 590378 676574
rect 590462 676338 590698 676574
rect 590142 640658 590378 640894
rect 590462 640658 590698 640894
rect 590142 640338 590378 640574
rect 590462 640338 590698 640574
rect 590142 604658 590378 604894
rect 590462 604658 590698 604894
rect 590142 604338 590378 604574
rect 590462 604338 590698 604574
rect 590142 568658 590378 568894
rect 590462 568658 590698 568894
rect 590142 568338 590378 568574
rect 590462 568338 590698 568574
rect 590142 532658 590378 532894
rect 590462 532658 590698 532894
rect 590142 532338 590378 532574
rect 590462 532338 590698 532574
rect 590142 496658 590378 496894
rect 590462 496658 590698 496894
rect 590142 496338 590378 496574
rect 590462 496338 590698 496574
rect 590142 460658 590378 460894
rect 590462 460658 590698 460894
rect 590142 460338 590378 460574
rect 590462 460338 590698 460574
rect 590142 424658 590378 424894
rect 590462 424658 590698 424894
rect 590142 424338 590378 424574
rect 590462 424338 590698 424574
rect 590142 388658 590378 388894
rect 590462 388658 590698 388894
rect 590142 388338 590378 388574
rect 590462 388338 590698 388574
rect 590142 352658 590378 352894
rect 590462 352658 590698 352894
rect 590142 352338 590378 352574
rect 590462 352338 590698 352574
rect 590142 316658 590378 316894
rect 590462 316658 590698 316894
rect 590142 316338 590378 316574
rect 590462 316338 590698 316574
rect 590142 280658 590378 280894
rect 590462 280658 590698 280894
rect 590142 280338 590378 280574
rect 590462 280338 590698 280574
rect 590142 244658 590378 244894
rect 590462 244658 590698 244894
rect 590142 244338 590378 244574
rect 590462 244338 590698 244574
rect 590142 208658 590378 208894
rect 590462 208658 590698 208894
rect 590142 208338 590378 208574
rect 590462 208338 590698 208574
rect 590142 172658 590378 172894
rect 590462 172658 590698 172894
rect 590142 172338 590378 172574
rect 590462 172338 590698 172574
rect 590142 136658 590378 136894
rect 590462 136658 590698 136894
rect 590142 136338 590378 136574
rect 590462 136338 590698 136574
rect 590142 100658 590378 100894
rect 590462 100658 590698 100894
rect 590142 100338 590378 100574
rect 590462 100338 590698 100574
rect 590142 64658 590378 64894
rect 590462 64658 590698 64894
rect 590142 64338 590378 64574
rect 590462 64338 590698 64574
rect 590142 28658 590378 28894
rect 590462 28658 590698 28894
rect 590142 28338 590378 28574
rect 590462 28338 590698 28574
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 698378 591338 698614
rect 591422 698378 591658 698614
rect 591102 698058 591338 698294
rect 591422 698058 591658 698294
rect 591102 662378 591338 662614
rect 591422 662378 591658 662614
rect 591102 662058 591338 662294
rect 591422 662058 591658 662294
rect 591102 626378 591338 626614
rect 591422 626378 591658 626614
rect 591102 626058 591338 626294
rect 591422 626058 591658 626294
rect 591102 590378 591338 590614
rect 591422 590378 591658 590614
rect 591102 590058 591338 590294
rect 591422 590058 591658 590294
rect 591102 554378 591338 554614
rect 591422 554378 591658 554614
rect 591102 554058 591338 554294
rect 591422 554058 591658 554294
rect 591102 518378 591338 518614
rect 591422 518378 591658 518614
rect 591102 518058 591338 518294
rect 591422 518058 591658 518294
rect 591102 482378 591338 482614
rect 591422 482378 591658 482614
rect 591102 482058 591338 482294
rect 591422 482058 591658 482294
rect 591102 446378 591338 446614
rect 591422 446378 591658 446614
rect 591102 446058 591338 446294
rect 591422 446058 591658 446294
rect 591102 410378 591338 410614
rect 591422 410378 591658 410614
rect 591102 410058 591338 410294
rect 591422 410058 591658 410294
rect 591102 374378 591338 374614
rect 591422 374378 591658 374614
rect 591102 374058 591338 374294
rect 591422 374058 591658 374294
rect 591102 338378 591338 338614
rect 591422 338378 591658 338614
rect 591102 338058 591338 338294
rect 591422 338058 591658 338294
rect 591102 302378 591338 302614
rect 591422 302378 591658 302614
rect 591102 302058 591338 302294
rect 591422 302058 591658 302294
rect 591102 266378 591338 266614
rect 591422 266378 591658 266614
rect 591102 266058 591338 266294
rect 591422 266058 591658 266294
rect 591102 230378 591338 230614
rect 591422 230378 591658 230614
rect 591102 230058 591338 230294
rect 591422 230058 591658 230294
rect 591102 194378 591338 194614
rect 591422 194378 591658 194614
rect 591102 194058 591338 194294
rect 591422 194058 591658 194294
rect 591102 158378 591338 158614
rect 591422 158378 591658 158614
rect 591102 158058 591338 158294
rect 591422 158058 591658 158294
rect 591102 122378 591338 122614
rect 591422 122378 591658 122614
rect 591102 122058 591338 122294
rect 591422 122058 591658 122294
rect 591102 86378 591338 86614
rect 591422 86378 591658 86614
rect 591102 86058 591338 86294
rect 591422 86058 591658 86294
rect 591102 50378 591338 50614
rect 591422 50378 591658 50614
rect 591102 50058 591338 50294
rect 591422 50058 591658 50294
rect 591102 14378 591338 14614
rect 591422 14378 591658 14614
rect 591102 14058 591338 14294
rect 591422 14058 591658 14294
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 680378 592298 680614
rect 592382 680378 592618 680614
rect 592062 680058 592298 680294
rect 592382 680058 592618 680294
rect 592062 644378 592298 644614
rect 592382 644378 592618 644614
rect 592062 644058 592298 644294
rect 592382 644058 592618 644294
rect 592062 608378 592298 608614
rect 592382 608378 592618 608614
rect 592062 608058 592298 608294
rect 592382 608058 592618 608294
rect 592062 572378 592298 572614
rect 592382 572378 592618 572614
rect 592062 572058 592298 572294
rect 592382 572058 592618 572294
rect 592062 536378 592298 536614
rect 592382 536378 592618 536614
rect 592062 536058 592298 536294
rect 592382 536058 592618 536294
rect 592062 500378 592298 500614
rect 592382 500378 592618 500614
rect 592062 500058 592298 500294
rect 592382 500058 592618 500294
rect 592062 464378 592298 464614
rect 592382 464378 592618 464614
rect 592062 464058 592298 464294
rect 592382 464058 592618 464294
rect 592062 428378 592298 428614
rect 592382 428378 592618 428614
rect 592062 428058 592298 428294
rect 592382 428058 592618 428294
rect 592062 392378 592298 392614
rect 592382 392378 592618 392614
rect 592062 392058 592298 392294
rect 592382 392058 592618 392294
rect 592062 356378 592298 356614
rect 592382 356378 592618 356614
rect 592062 356058 592298 356294
rect 592382 356058 592618 356294
rect 592062 320378 592298 320614
rect 592382 320378 592618 320614
rect 592062 320058 592298 320294
rect 592382 320058 592618 320294
rect 592062 284378 592298 284614
rect 592382 284378 592618 284614
rect 592062 284058 592298 284294
rect 592382 284058 592618 284294
rect 592062 248378 592298 248614
rect 592382 248378 592618 248614
rect 592062 248058 592298 248294
rect 592382 248058 592618 248294
rect 592062 212378 592298 212614
rect 592382 212378 592618 212614
rect 592062 212058 592298 212294
rect 592382 212058 592618 212294
rect 592062 176378 592298 176614
rect 592382 176378 592618 176614
rect 592062 176058 592298 176294
rect 592382 176058 592618 176294
rect 592062 140378 592298 140614
rect 592382 140378 592618 140614
rect 592062 140058 592298 140294
rect 592382 140058 592618 140294
rect 592062 104378 592298 104614
rect 592382 104378 592618 104614
rect 592062 104058 592298 104294
rect 592382 104058 592618 104294
rect 592062 68378 592298 68614
rect 592382 68378 592618 68614
rect 592062 68058 592298 68294
rect 592382 68058 592618 68294
rect 592062 32378 592298 32614
rect 592382 32378 592618 32614
rect 592062 32058 592298 32294
rect 592382 32058 592618 32294
rect 570986 -7302 571222 -7066
rect 571306 -7302 571542 -7066
rect 570986 -7622 571222 -7386
rect 571306 -7622 571542 -7386
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 592650 698614
rect -8726 698294 592650 698378
rect -8726 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 592650 698294
rect -8726 698026 592650 698058
rect -6806 694894 590730 694926
rect -6806 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 590730 694894
rect -6806 694574 590730 694658
rect -6806 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 590730 694574
rect -6806 694306 590730 694338
rect -4886 691174 588810 691206
rect -4886 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 588810 691174
rect -4886 690854 588810 690938
rect -4886 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 588810 690854
rect -4886 690586 588810 690618
rect -2966 687454 586890 687486
rect -2966 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 586890 687454
rect -2966 687134 586890 687218
rect -2966 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 586890 687134
rect -2966 686866 586890 686898
rect -8726 680614 592650 680646
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect -8726 680294 592650 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect -8726 680026 592650 680058
rect -6806 676894 590730 676926
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect -6806 676574 590730 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect -6806 676306 590730 676338
rect -4886 673174 588810 673206
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect -4886 672854 588810 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect -4886 672586 588810 672618
rect -2966 669454 586890 669486
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect -2966 669134 586890 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect -2966 668866 586890 668898
rect -8726 662614 592650 662646
rect -8726 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 592650 662614
rect -8726 662294 592650 662378
rect -8726 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 592650 662294
rect -8726 662026 592650 662058
rect -6806 658894 590730 658926
rect -6806 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 590730 658894
rect -6806 658574 590730 658658
rect -6806 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 590730 658574
rect -6806 658306 590730 658338
rect -4886 655174 588810 655206
rect -4886 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 588810 655174
rect -4886 654854 588810 654938
rect -4886 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 588810 654854
rect -4886 654586 588810 654618
rect -2966 651454 586890 651486
rect -2966 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 586890 651454
rect -2966 651134 586890 651218
rect -2966 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 586890 651134
rect -2966 650866 586890 650898
rect -8726 644614 592650 644646
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect -8726 644294 592650 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect -8726 644026 592650 644058
rect -6806 640894 590730 640926
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect -6806 640574 590730 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect -6806 640306 590730 640338
rect -4886 637174 588810 637206
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect -4886 636854 588810 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect -4886 636586 588810 636618
rect -2966 633454 586890 633486
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect -2966 633134 586890 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect -2966 632866 586890 632898
rect -8726 626614 592650 626646
rect -8726 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 592650 626614
rect -8726 626294 592650 626378
rect -8726 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 592650 626294
rect -8726 626026 592650 626058
rect -6806 622894 590730 622926
rect -6806 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 590730 622894
rect -6806 622574 590730 622658
rect -6806 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 590730 622574
rect -6806 622306 590730 622338
rect -4886 619174 588810 619206
rect -4886 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 588810 619174
rect -4886 618854 588810 618938
rect -4886 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 588810 618854
rect -4886 618586 588810 618618
rect -2966 615454 586890 615486
rect -2966 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 586890 615454
rect -2966 615134 586890 615218
rect -2966 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 586890 615134
rect -2966 614866 586890 614898
rect -8726 608614 592650 608646
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect -8726 608294 592650 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect -8726 608026 592650 608058
rect -6806 604894 590730 604926
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect -6806 604574 590730 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect -6806 604306 590730 604338
rect -4886 601174 588810 601206
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect -4886 600854 588810 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect -4886 600586 588810 600618
rect -2966 597454 586890 597486
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect -2966 597134 586890 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect -2966 596866 586890 596898
rect -8726 590614 592650 590646
rect -8726 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 592650 590614
rect -8726 590294 592650 590378
rect -8726 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 592650 590294
rect -8726 590026 592650 590058
rect -6806 586894 590730 586926
rect -6806 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 590730 586894
rect -6806 586574 590730 586658
rect -6806 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 590730 586574
rect -6806 586306 590730 586338
rect -4886 583174 588810 583206
rect -4886 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 588810 583174
rect -4886 582854 588810 582938
rect -4886 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 588810 582854
rect -4886 582586 588810 582618
rect -2966 579454 586890 579486
rect -2966 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 72721 579454
rect 72957 579218 78651 579454
rect 78887 579218 84582 579454
rect 84818 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 586890 579454
rect -2966 579134 586890 579218
rect -2966 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 72721 579134
rect 72957 578898 78651 579134
rect 78887 578898 84582 579134
rect 84818 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 586890 579134
rect -2966 578866 586890 578898
rect -8726 572614 592650 572646
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect -8726 572294 592650 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect -8726 572026 592650 572058
rect -6806 568894 590730 568926
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect -6806 568574 590730 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect -6806 568306 590730 568338
rect -4886 565174 588810 565206
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 95546 565174
rect 95782 564938 95866 565174
rect 96102 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 419546 565174
rect 419782 564938 419866 565174
rect 420102 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect -4886 564854 588810 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 95546 564854
rect 95782 564618 95866 564854
rect 96102 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 419546 564854
rect 419782 564618 419866 564854
rect 420102 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect -4886 564586 588810 564618
rect -2966 561454 586890 561486
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 75686 561454
rect 75922 561218 81617 561454
rect 81853 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect -2966 561134 586890 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 75686 561134
rect 75922 560898 81617 561134
rect 81853 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect -2966 560866 586890 560898
rect -8726 554614 592650 554646
rect -8726 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 592650 554614
rect -8726 554294 592650 554378
rect -8726 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 592650 554294
rect -8726 554026 592650 554058
rect -6806 550894 590730 550926
rect -6806 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 590730 550894
rect -6806 550574 590730 550658
rect -6806 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 590730 550574
rect -6806 550306 590730 550338
rect -4886 547174 588810 547206
rect -4886 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 588810 547174
rect -4886 546854 588810 546938
rect -4886 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 588810 546854
rect -4886 546586 588810 546618
rect -2966 543454 586890 543486
rect -2966 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 72721 543454
rect 72957 543218 78651 543454
rect 78887 543218 84582 543454
rect 84818 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 586890 543454
rect -2966 543134 586890 543218
rect -2966 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 72721 543134
rect 72957 542898 78651 543134
rect 78887 542898 84582 543134
rect 84818 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 586890 543134
rect -2966 542866 586890 542898
rect -8726 536614 592650 536646
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 102986 536614
rect 103222 536378 103306 536614
rect 103542 536378 138986 536614
rect 139222 536378 139306 536614
rect 139542 536378 174986 536614
rect 175222 536378 175306 536614
rect 175542 536378 390986 536614
rect 391222 536378 391306 536614
rect 391542 536378 426986 536614
rect 427222 536378 427306 536614
rect 427542 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect -8726 536294 592650 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 102986 536294
rect 103222 536058 103306 536294
rect 103542 536058 138986 536294
rect 139222 536058 139306 536294
rect 139542 536058 174986 536294
rect 175222 536058 175306 536294
rect 175542 536058 390986 536294
rect 391222 536058 391306 536294
rect 391542 536058 426986 536294
rect 427222 536058 427306 536294
rect 427542 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect -8726 536026 592650 536058
rect -6806 532894 590730 532926
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 99266 532894
rect 99502 532658 99586 532894
rect 99822 532658 135266 532894
rect 135502 532658 135586 532894
rect 135822 532658 171266 532894
rect 171502 532658 171586 532894
rect 171822 532658 387266 532894
rect 387502 532658 387586 532894
rect 387822 532658 423266 532894
rect 423502 532658 423586 532894
rect 423822 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect -6806 532574 590730 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 99266 532574
rect 99502 532338 99586 532574
rect 99822 532338 135266 532574
rect 135502 532338 135586 532574
rect 135822 532338 171266 532574
rect 171502 532338 171586 532574
rect 171822 532338 387266 532574
rect 387502 532338 387586 532574
rect 387822 532338 423266 532574
rect 423502 532338 423586 532574
rect 423822 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect -6806 532306 590730 532338
rect -4886 529174 588810 529206
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 95546 529174
rect 95782 528938 95866 529174
rect 96102 528938 131546 529174
rect 131782 528938 131866 529174
rect 132102 528938 167546 529174
rect 167782 528938 167866 529174
rect 168102 528938 383546 529174
rect 383782 528938 383866 529174
rect 384102 528938 419546 529174
rect 419782 528938 419866 529174
rect 420102 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect -4886 528854 588810 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 95546 528854
rect 95782 528618 95866 528854
rect 96102 528618 131546 528854
rect 131782 528618 131866 528854
rect 132102 528618 167546 528854
rect 167782 528618 167866 528854
rect 168102 528618 383546 528854
rect 383782 528618 383866 528854
rect 384102 528618 419546 528854
rect 419782 528618 419866 528854
rect 420102 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect -4886 528586 588810 528618
rect -2966 525454 586890 525486
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 219610 525454
rect 219846 525218 250330 525454
rect 250566 525218 281050 525454
rect 281286 525218 311770 525454
rect 312006 525218 342490 525454
rect 342726 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect -2966 525134 586890 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 219610 525134
rect 219846 524898 250330 525134
rect 250566 524898 281050 525134
rect 281286 524898 311770 525134
rect 312006 524898 342490 525134
rect 342726 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect -2966 524866 586890 524898
rect -8726 518614 592650 518646
rect -8726 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 592650 518614
rect -8726 518294 592650 518378
rect -8726 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 592650 518294
rect -8726 518026 592650 518058
rect -6806 514894 590730 514926
rect -6806 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 590730 514894
rect -6806 514574 590730 514658
rect -6806 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 590730 514574
rect -6806 514306 590730 514338
rect -4886 511174 588810 511206
rect -4886 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 588810 511174
rect -4886 510854 588810 510938
rect -4886 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 588810 510854
rect -4886 510586 588810 510618
rect -2966 507454 586890 507486
rect -2966 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 204250 507454
rect 204486 507218 234970 507454
rect 235206 507218 265690 507454
rect 265926 507218 296410 507454
rect 296646 507218 327130 507454
rect 327366 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 586890 507454
rect -2966 507134 586890 507218
rect -2966 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 204250 507134
rect 204486 506898 234970 507134
rect 235206 506898 265690 507134
rect 265926 506898 296410 507134
rect 296646 506898 327130 507134
rect 327366 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 586890 507134
rect -2966 506866 586890 506898
rect -8726 500614 592650 500646
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 102986 500614
rect 103222 500378 103306 500614
rect 103542 500378 138986 500614
rect 139222 500378 139306 500614
rect 139542 500378 174986 500614
rect 175222 500378 175306 500614
rect 175542 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect -8726 500294 592650 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 102986 500294
rect 103222 500058 103306 500294
rect 103542 500058 138986 500294
rect 139222 500058 139306 500294
rect 139542 500058 174986 500294
rect 175222 500058 175306 500294
rect 175542 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect -8726 500026 592650 500058
rect -6806 496894 590730 496926
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 99266 496894
rect 99502 496658 99586 496894
rect 99822 496658 135266 496894
rect 135502 496658 135586 496894
rect 135822 496658 171266 496894
rect 171502 496658 171586 496894
rect 171822 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect -6806 496574 590730 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 99266 496574
rect 99502 496338 99586 496574
rect 99822 496338 135266 496574
rect 135502 496338 135586 496574
rect 135822 496338 171266 496574
rect 171502 496338 171586 496574
rect 171822 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect -6806 496306 590730 496338
rect -4886 493174 588810 493206
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 95546 493174
rect 95782 492938 95866 493174
rect 96102 492938 131546 493174
rect 131782 492938 131866 493174
rect 132102 492938 167546 493174
rect 167782 492938 167866 493174
rect 168102 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect -4886 492854 588810 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 95546 492854
rect 95782 492618 95866 492854
rect 96102 492618 131546 492854
rect 131782 492618 131866 492854
rect 132102 492618 167546 492854
rect 167782 492618 167866 492854
rect 168102 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect -4886 492586 588810 492618
rect -2966 489454 586890 489486
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 219610 489454
rect 219846 489218 250330 489454
rect 250566 489218 281050 489454
rect 281286 489218 311770 489454
rect 312006 489218 342490 489454
rect 342726 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect -2966 489134 586890 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 219610 489134
rect 219846 488898 250330 489134
rect 250566 488898 281050 489134
rect 281286 488898 311770 489134
rect 312006 488898 342490 489134
rect 342726 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect -2966 488866 586890 488898
rect -8726 482614 592650 482646
rect -8726 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 592650 482614
rect -8726 482294 592650 482378
rect -8726 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 592650 482294
rect -8726 482026 592650 482058
rect -6806 478894 590730 478926
rect -6806 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 590730 478894
rect -6806 478574 590730 478658
rect -6806 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 590730 478574
rect -6806 478306 590730 478338
rect -4886 475174 588810 475206
rect -4886 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 588810 475174
rect -4886 474854 588810 474938
rect -4886 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 588810 474854
rect -4886 474586 588810 474618
rect -2966 471454 586890 471486
rect -2966 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 204250 471454
rect 204486 471218 234970 471454
rect 235206 471218 265690 471454
rect 265926 471218 296410 471454
rect 296646 471218 327130 471454
rect 327366 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 586890 471454
rect -2966 471134 586890 471218
rect -2966 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 204250 471134
rect 204486 470898 234970 471134
rect 235206 470898 265690 471134
rect 265926 470898 296410 471134
rect 296646 470898 327130 471134
rect 327366 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 586890 471134
rect -2966 470866 586890 470898
rect -8726 464614 592650 464646
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 66986 464614
rect 67222 464378 67306 464614
rect 67542 464378 102986 464614
rect 103222 464378 103306 464614
rect 103542 464378 138986 464614
rect 139222 464378 139306 464614
rect 139542 464378 174986 464614
rect 175222 464378 175306 464614
rect 175542 464378 390986 464614
rect 391222 464378 391306 464614
rect 391542 464378 426986 464614
rect 427222 464378 427306 464614
rect 427542 464378 462986 464614
rect 463222 464378 463306 464614
rect 463542 464378 498986 464614
rect 499222 464378 499306 464614
rect 499542 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect -8726 464294 592650 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 66986 464294
rect 67222 464058 67306 464294
rect 67542 464058 102986 464294
rect 103222 464058 103306 464294
rect 103542 464058 138986 464294
rect 139222 464058 139306 464294
rect 139542 464058 174986 464294
rect 175222 464058 175306 464294
rect 175542 464058 390986 464294
rect 391222 464058 391306 464294
rect 391542 464058 426986 464294
rect 427222 464058 427306 464294
rect 427542 464058 462986 464294
rect 463222 464058 463306 464294
rect 463542 464058 498986 464294
rect 499222 464058 499306 464294
rect 499542 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect -8726 464026 592650 464058
rect -6806 460894 590730 460926
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 63266 460894
rect 63502 460658 63586 460894
rect 63822 460658 99266 460894
rect 99502 460658 99586 460894
rect 99822 460658 135266 460894
rect 135502 460658 135586 460894
rect 135822 460658 171266 460894
rect 171502 460658 171586 460894
rect 171822 460658 387266 460894
rect 387502 460658 387586 460894
rect 387822 460658 423266 460894
rect 423502 460658 423586 460894
rect 423822 460658 459266 460894
rect 459502 460658 459586 460894
rect 459822 460658 495266 460894
rect 495502 460658 495586 460894
rect 495822 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect -6806 460574 590730 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 63266 460574
rect 63502 460338 63586 460574
rect 63822 460338 99266 460574
rect 99502 460338 99586 460574
rect 99822 460338 135266 460574
rect 135502 460338 135586 460574
rect 135822 460338 171266 460574
rect 171502 460338 171586 460574
rect 171822 460338 387266 460574
rect 387502 460338 387586 460574
rect 387822 460338 423266 460574
rect 423502 460338 423586 460574
rect 423822 460338 459266 460574
rect 459502 460338 459586 460574
rect 459822 460338 495266 460574
rect 495502 460338 495586 460574
rect 495822 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect -6806 460306 590730 460338
rect -4886 457174 588810 457206
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 59546 457174
rect 59782 456938 59866 457174
rect 60102 456938 95546 457174
rect 95782 456938 95866 457174
rect 96102 456938 131546 457174
rect 131782 456938 131866 457174
rect 132102 456938 167546 457174
rect 167782 456938 167866 457174
rect 168102 456938 383546 457174
rect 383782 456938 383866 457174
rect 384102 456938 419546 457174
rect 419782 456938 419866 457174
rect 420102 456938 455546 457174
rect 455782 456938 455866 457174
rect 456102 456938 491546 457174
rect 491782 456938 491866 457174
rect 492102 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect -4886 456854 588810 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 59546 456854
rect 59782 456618 59866 456854
rect 60102 456618 95546 456854
rect 95782 456618 95866 456854
rect 96102 456618 131546 456854
rect 131782 456618 131866 456854
rect 132102 456618 167546 456854
rect 167782 456618 167866 456854
rect 168102 456618 383546 456854
rect 383782 456618 383866 456854
rect 384102 456618 419546 456854
rect 419782 456618 419866 456854
rect 420102 456618 455546 456854
rect 455782 456618 455866 456854
rect 456102 456618 491546 456854
rect 491782 456618 491866 456854
rect 492102 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect -4886 456586 588810 456618
rect -2966 453454 586890 453486
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 219610 453454
rect 219846 453218 250330 453454
rect 250566 453218 281050 453454
rect 281286 453218 311770 453454
rect 312006 453218 342490 453454
rect 342726 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect -2966 453134 586890 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 219610 453134
rect 219846 452898 250330 453134
rect 250566 452898 281050 453134
rect 281286 452898 311770 453134
rect 312006 452898 342490 453134
rect 342726 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect -2966 452866 586890 452898
rect -8726 446614 592650 446646
rect -8726 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 156986 446614
rect 157222 446378 157306 446614
rect 157542 446378 192986 446614
rect 193222 446378 193306 446614
rect 193542 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 592650 446614
rect -8726 446294 592650 446378
rect -8726 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 156986 446294
rect 157222 446058 157306 446294
rect 157542 446058 192986 446294
rect 193222 446058 193306 446294
rect 193542 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 592650 446294
rect -8726 446026 592650 446058
rect -6806 442894 590730 442926
rect -6806 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 153266 442894
rect 153502 442658 153586 442894
rect 153822 442658 189266 442894
rect 189502 442658 189586 442894
rect 189822 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 441266 442894
rect 441502 442658 441586 442894
rect 441822 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 590730 442894
rect -6806 442574 590730 442658
rect -6806 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 153266 442574
rect 153502 442338 153586 442574
rect 153822 442338 189266 442574
rect 189502 442338 189586 442574
rect 189822 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 441266 442574
rect 441502 442338 441586 442574
rect 441822 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 590730 442574
rect -6806 442306 590730 442338
rect -4886 439174 588810 439206
rect -4886 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 149546 439174
rect 149782 438938 149866 439174
rect 150102 438938 185546 439174
rect 185782 438938 185866 439174
rect 186102 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 437546 439174
rect 437782 438938 437866 439174
rect 438102 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 588810 439174
rect -4886 438854 588810 438938
rect -4886 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 149546 438854
rect 149782 438618 149866 438854
rect 150102 438618 185546 438854
rect 185782 438618 185866 438854
rect 186102 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 437546 438854
rect 437782 438618 437866 438854
rect 438102 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 588810 438854
rect -4886 438586 588810 438618
rect -2966 435454 586890 435486
rect -2966 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 73020 435454
rect 73256 435218 103740 435454
rect 103976 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 204250 435454
rect 204486 435218 234970 435454
rect 235206 435218 265690 435454
rect 265926 435218 296410 435454
rect 296646 435218 327130 435454
rect 327366 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 586890 435454
rect -2966 435134 586890 435218
rect -2966 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 73020 435134
rect 73256 434898 103740 435134
rect 103976 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 204250 435134
rect 204486 434898 234970 435134
rect 235206 434898 265690 435134
rect 265926 434898 296410 435134
rect 296646 434898 327130 435134
rect 327366 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 586890 435134
rect -2966 434866 586890 434898
rect -8726 428614 592650 428646
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 138986 428614
rect 139222 428378 139306 428614
rect 139542 428378 174986 428614
rect 175222 428378 175306 428614
rect 175542 428378 390986 428614
rect 391222 428378 391306 428614
rect 391542 428378 426986 428614
rect 427222 428378 427306 428614
rect 427542 428378 462986 428614
rect 463222 428378 463306 428614
rect 463542 428378 498986 428614
rect 499222 428378 499306 428614
rect 499542 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect -8726 428294 592650 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 138986 428294
rect 139222 428058 139306 428294
rect 139542 428058 174986 428294
rect 175222 428058 175306 428294
rect 175542 428058 390986 428294
rect 391222 428058 391306 428294
rect 391542 428058 426986 428294
rect 427222 428058 427306 428294
rect 427542 428058 462986 428294
rect 463222 428058 463306 428294
rect 463542 428058 498986 428294
rect 499222 428058 499306 428294
rect 499542 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect -8726 428026 592650 428058
rect -6806 424894 590730 424926
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 63266 424894
rect 63502 424658 63586 424894
rect 63822 424658 135266 424894
rect 135502 424658 135586 424894
rect 135822 424658 171266 424894
rect 171502 424658 171586 424894
rect 171822 424658 387266 424894
rect 387502 424658 387586 424894
rect 387822 424658 423266 424894
rect 423502 424658 423586 424894
rect 423822 424658 459266 424894
rect 459502 424658 459586 424894
rect 459822 424658 495266 424894
rect 495502 424658 495586 424894
rect 495822 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect -6806 424574 590730 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 63266 424574
rect 63502 424338 63586 424574
rect 63822 424338 135266 424574
rect 135502 424338 135586 424574
rect 135822 424338 171266 424574
rect 171502 424338 171586 424574
rect 171822 424338 387266 424574
rect 387502 424338 387586 424574
rect 387822 424338 423266 424574
rect 423502 424338 423586 424574
rect 423822 424338 459266 424574
rect 459502 424338 459586 424574
rect 459822 424338 495266 424574
rect 495502 424338 495586 424574
rect 495822 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect -6806 424306 590730 424338
rect -4886 421174 588810 421206
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 59546 421174
rect 59782 420938 59866 421174
rect 60102 420938 131546 421174
rect 131782 420938 131866 421174
rect 132102 420938 167546 421174
rect 167782 420938 167866 421174
rect 168102 420938 383546 421174
rect 383782 420938 383866 421174
rect 384102 420938 419546 421174
rect 419782 420938 419866 421174
rect 420102 420938 455546 421174
rect 455782 420938 455866 421174
rect 456102 420938 491546 421174
rect 491782 420938 491866 421174
rect 492102 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect -4886 420854 588810 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 59546 420854
rect 59782 420618 59866 420854
rect 60102 420618 131546 420854
rect 131782 420618 131866 420854
rect 132102 420618 167546 420854
rect 167782 420618 167866 420854
rect 168102 420618 383546 420854
rect 383782 420618 383866 420854
rect 384102 420618 419546 420854
rect 419782 420618 419866 420854
rect 420102 420618 455546 420854
rect 455782 420618 455866 420854
rect 456102 420618 491546 420854
rect 491782 420618 491866 420854
rect 492102 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect -4886 420586 588810 420618
rect -2966 417454 586890 417486
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 88380 417454
rect 88616 417218 119100 417454
rect 119336 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 219610 417454
rect 219846 417218 250330 417454
rect 250566 417218 281050 417454
rect 281286 417218 311770 417454
rect 312006 417218 342490 417454
rect 342726 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect -2966 417134 586890 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 88380 417134
rect 88616 416898 119100 417134
rect 119336 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 219610 417134
rect 219846 416898 250330 417134
rect 250566 416898 281050 417134
rect 281286 416898 311770 417134
rect 312006 416898 342490 417134
rect 342726 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect -2966 416866 586890 416898
rect -8726 410614 592650 410646
rect -8726 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 156986 410614
rect 157222 410378 157306 410614
rect 157542 410378 192986 410614
rect 193222 410378 193306 410614
rect 193542 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 408986 410614
rect 409222 410378 409306 410614
rect 409542 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 592650 410614
rect -8726 410294 592650 410378
rect -8726 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 156986 410294
rect 157222 410058 157306 410294
rect 157542 410058 192986 410294
rect 193222 410058 193306 410294
rect 193542 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 408986 410294
rect 409222 410058 409306 410294
rect 409542 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 592650 410294
rect -8726 410026 592650 410058
rect -6806 406894 590730 406926
rect -6806 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 153266 406894
rect 153502 406658 153586 406894
rect 153822 406658 189266 406894
rect 189502 406658 189586 406894
rect 189822 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 405266 406894
rect 405502 406658 405586 406894
rect 405822 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 590730 406894
rect -6806 406574 590730 406658
rect -6806 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 153266 406574
rect 153502 406338 153586 406574
rect 153822 406338 189266 406574
rect 189502 406338 189586 406574
rect 189822 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 405266 406574
rect 405502 406338 405586 406574
rect 405822 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 590730 406574
rect -6806 406306 590730 406338
rect -4886 403174 588810 403206
rect -4886 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 149546 403174
rect 149782 402938 149866 403174
rect 150102 402938 185546 403174
rect 185782 402938 185866 403174
rect 186102 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 588810 403174
rect -4886 402854 588810 402938
rect -4886 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 149546 402854
rect 149782 402618 149866 402854
rect 150102 402618 185546 402854
rect 185782 402618 185866 402854
rect 186102 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 588810 402854
rect -4886 402586 588810 402618
rect -2966 399454 586890 399486
rect -2966 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 73020 399454
rect 73256 399218 103740 399454
rect 103976 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 204250 399454
rect 204486 399218 234970 399454
rect 235206 399218 265690 399454
rect 265926 399218 296410 399454
rect 296646 399218 327130 399454
rect 327366 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 586890 399454
rect -2966 399134 586890 399218
rect -2966 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 73020 399134
rect 73256 398898 103740 399134
rect 103976 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 204250 399134
rect 204486 398898 234970 399134
rect 235206 398898 265690 399134
rect 265926 398898 296410 399134
rect 296646 398898 327130 399134
rect 327366 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 586890 399134
rect -2966 398866 586890 398898
rect -8726 392614 592650 392646
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 138986 392614
rect 139222 392378 139306 392614
rect 139542 392378 174986 392614
rect 175222 392378 175306 392614
rect 175542 392378 390986 392614
rect 391222 392378 391306 392614
rect 391542 392378 426986 392614
rect 427222 392378 427306 392614
rect 427542 392378 462986 392614
rect 463222 392378 463306 392614
rect 463542 392378 498986 392614
rect 499222 392378 499306 392614
rect 499542 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect -8726 392294 592650 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 138986 392294
rect 139222 392058 139306 392294
rect 139542 392058 174986 392294
rect 175222 392058 175306 392294
rect 175542 392058 390986 392294
rect 391222 392058 391306 392294
rect 391542 392058 426986 392294
rect 427222 392058 427306 392294
rect 427542 392058 462986 392294
rect 463222 392058 463306 392294
rect 463542 392058 498986 392294
rect 499222 392058 499306 392294
rect 499542 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect -8726 392026 592650 392058
rect -6806 388894 590730 388926
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 63266 388894
rect 63502 388658 63586 388894
rect 63822 388658 135266 388894
rect 135502 388658 135586 388894
rect 135822 388658 171266 388894
rect 171502 388658 171586 388894
rect 171822 388658 387266 388894
rect 387502 388658 387586 388894
rect 387822 388658 423266 388894
rect 423502 388658 423586 388894
rect 423822 388658 459266 388894
rect 459502 388658 459586 388894
rect 459822 388658 495266 388894
rect 495502 388658 495586 388894
rect 495822 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect -6806 388574 590730 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 63266 388574
rect 63502 388338 63586 388574
rect 63822 388338 135266 388574
rect 135502 388338 135586 388574
rect 135822 388338 171266 388574
rect 171502 388338 171586 388574
rect 171822 388338 387266 388574
rect 387502 388338 387586 388574
rect 387822 388338 423266 388574
rect 423502 388338 423586 388574
rect 423822 388338 459266 388574
rect 459502 388338 459586 388574
rect 459822 388338 495266 388574
rect 495502 388338 495586 388574
rect 495822 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect -6806 388306 590730 388338
rect -4886 385174 588810 385206
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 59546 385174
rect 59782 384938 59866 385174
rect 60102 384938 95546 385174
rect 95782 384938 95866 385174
rect 96102 384938 131546 385174
rect 131782 384938 131866 385174
rect 132102 384938 167546 385174
rect 167782 384938 167866 385174
rect 168102 384938 383546 385174
rect 383782 384938 383866 385174
rect 384102 384938 419546 385174
rect 419782 384938 419866 385174
rect 420102 384938 455546 385174
rect 455782 384938 455866 385174
rect 456102 384938 491546 385174
rect 491782 384938 491866 385174
rect 492102 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect -4886 384854 588810 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 59546 384854
rect 59782 384618 59866 384854
rect 60102 384618 95546 384854
rect 95782 384618 95866 384854
rect 96102 384618 131546 384854
rect 131782 384618 131866 384854
rect 132102 384618 167546 384854
rect 167782 384618 167866 384854
rect 168102 384618 383546 384854
rect 383782 384618 383866 384854
rect 384102 384618 419546 384854
rect 419782 384618 419866 384854
rect 420102 384618 455546 384854
rect 455782 384618 455866 384854
rect 456102 384618 491546 384854
rect 491782 384618 491866 384854
rect 492102 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect -4886 384586 588810 384618
rect -2966 381454 586890 381486
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 219610 381454
rect 219846 381218 250330 381454
rect 250566 381218 281050 381454
rect 281286 381218 311770 381454
rect 312006 381218 342490 381454
rect 342726 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect -2966 381134 586890 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 219610 381134
rect 219846 380898 250330 381134
rect 250566 380898 281050 381134
rect 281286 380898 311770 381134
rect 312006 380898 342490 381134
rect 342726 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect -2966 380866 586890 380898
rect -8726 374614 592650 374646
rect -8726 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 84986 374614
rect 85222 374378 85306 374614
rect 85542 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 228986 374614
rect 229222 374378 229306 374614
rect 229542 374378 264986 374614
rect 265222 374378 265306 374614
rect 265542 374378 300986 374614
rect 301222 374378 301306 374614
rect 301542 374378 336986 374614
rect 337222 374378 337306 374614
rect 337542 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 592650 374614
rect -8726 374294 592650 374378
rect -8726 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 84986 374294
rect 85222 374058 85306 374294
rect 85542 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 228986 374294
rect 229222 374058 229306 374294
rect 229542 374058 264986 374294
rect 265222 374058 265306 374294
rect 265542 374058 300986 374294
rect 301222 374058 301306 374294
rect 301542 374058 336986 374294
rect 337222 374058 337306 374294
rect 337542 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 592650 374294
rect -8726 374026 592650 374058
rect -6806 370894 590730 370926
rect -6806 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 81266 370894
rect 81502 370658 81586 370894
rect 81822 370658 117266 370894
rect 117502 370658 117586 370894
rect 117822 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 225266 370894
rect 225502 370658 225586 370894
rect 225822 370658 261266 370894
rect 261502 370658 261586 370894
rect 261822 370658 297266 370894
rect 297502 370658 297586 370894
rect 297822 370658 333266 370894
rect 333502 370658 333586 370894
rect 333822 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 590730 370894
rect -6806 370574 590730 370658
rect -6806 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 81266 370574
rect 81502 370338 81586 370574
rect 81822 370338 117266 370574
rect 117502 370338 117586 370574
rect 117822 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 225266 370574
rect 225502 370338 225586 370574
rect 225822 370338 261266 370574
rect 261502 370338 261586 370574
rect 261822 370338 297266 370574
rect 297502 370338 297586 370574
rect 297822 370338 333266 370574
rect 333502 370338 333586 370574
rect 333822 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 590730 370574
rect -6806 370306 590730 370338
rect -4886 367174 588810 367206
rect -4886 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 77546 367174
rect 77782 366938 77866 367174
rect 78102 366938 113546 367174
rect 113782 366938 113866 367174
rect 114102 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 257546 367174
rect 257782 366938 257866 367174
rect 258102 366938 293546 367174
rect 293782 366938 293866 367174
rect 294102 366938 329546 367174
rect 329782 366938 329866 367174
rect 330102 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 588810 367174
rect -4886 366854 588810 366938
rect -4886 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 77546 366854
rect 77782 366618 77866 366854
rect 78102 366618 113546 366854
rect 113782 366618 113866 366854
rect 114102 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 257546 366854
rect 257782 366618 257866 366854
rect 258102 366618 293546 366854
rect 293782 366618 293866 366854
rect 294102 366618 329546 366854
rect 329782 366618 329866 366854
rect 330102 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 588810 366854
rect -4886 366586 588810 366618
rect -2966 363454 586890 363486
rect -2966 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 586890 363454
rect -2966 363134 586890 363218
rect -2966 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 586890 363134
rect -2966 362866 586890 362898
rect -8726 356614 592650 356646
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 66986 356614
rect 67222 356378 67306 356614
rect 67542 356378 102986 356614
rect 103222 356378 103306 356614
rect 103542 356378 138986 356614
rect 139222 356378 139306 356614
rect 139542 356378 174986 356614
rect 175222 356378 175306 356614
rect 175542 356378 210986 356614
rect 211222 356378 211306 356614
rect 211542 356378 246986 356614
rect 247222 356378 247306 356614
rect 247542 356378 282986 356614
rect 283222 356378 283306 356614
rect 283542 356378 318986 356614
rect 319222 356378 319306 356614
rect 319542 356378 354986 356614
rect 355222 356378 355306 356614
rect 355542 356378 390986 356614
rect 391222 356378 391306 356614
rect 391542 356378 426986 356614
rect 427222 356378 427306 356614
rect 427542 356378 462986 356614
rect 463222 356378 463306 356614
rect 463542 356378 498986 356614
rect 499222 356378 499306 356614
rect 499542 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect -8726 356294 592650 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 66986 356294
rect 67222 356058 67306 356294
rect 67542 356058 102986 356294
rect 103222 356058 103306 356294
rect 103542 356058 138986 356294
rect 139222 356058 139306 356294
rect 139542 356058 174986 356294
rect 175222 356058 175306 356294
rect 175542 356058 210986 356294
rect 211222 356058 211306 356294
rect 211542 356058 246986 356294
rect 247222 356058 247306 356294
rect 247542 356058 282986 356294
rect 283222 356058 283306 356294
rect 283542 356058 318986 356294
rect 319222 356058 319306 356294
rect 319542 356058 354986 356294
rect 355222 356058 355306 356294
rect 355542 356058 390986 356294
rect 391222 356058 391306 356294
rect 391542 356058 426986 356294
rect 427222 356058 427306 356294
rect 427542 356058 462986 356294
rect 463222 356058 463306 356294
rect 463542 356058 498986 356294
rect 499222 356058 499306 356294
rect 499542 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect -8726 356026 592650 356058
rect -6806 352894 590730 352926
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 63266 352894
rect 63502 352658 63586 352894
rect 63822 352658 99266 352894
rect 99502 352658 99586 352894
rect 99822 352658 135266 352894
rect 135502 352658 135586 352894
rect 135822 352658 171266 352894
rect 171502 352658 171586 352894
rect 171822 352658 207266 352894
rect 207502 352658 207586 352894
rect 207822 352658 243266 352894
rect 243502 352658 243586 352894
rect 243822 352658 279266 352894
rect 279502 352658 279586 352894
rect 279822 352658 315266 352894
rect 315502 352658 315586 352894
rect 315822 352658 351266 352894
rect 351502 352658 351586 352894
rect 351822 352658 387266 352894
rect 387502 352658 387586 352894
rect 387822 352658 423266 352894
rect 423502 352658 423586 352894
rect 423822 352658 459266 352894
rect 459502 352658 459586 352894
rect 459822 352658 495266 352894
rect 495502 352658 495586 352894
rect 495822 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect -6806 352574 590730 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 63266 352574
rect 63502 352338 63586 352574
rect 63822 352338 99266 352574
rect 99502 352338 99586 352574
rect 99822 352338 135266 352574
rect 135502 352338 135586 352574
rect 135822 352338 171266 352574
rect 171502 352338 171586 352574
rect 171822 352338 207266 352574
rect 207502 352338 207586 352574
rect 207822 352338 243266 352574
rect 243502 352338 243586 352574
rect 243822 352338 279266 352574
rect 279502 352338 279586 352574
rect 279822 352338 315266 352574
rect 315502 352338 315586 352574
rect 315822 352338 351266 352574
rect 351502 352338 351586 352574
rect 351822 352338 387266 352574
rect 387502 352338 387586 352574
rect 387822 352338 423266 352574
rect 423502 352338 423586 352574
rect 423822 352338 459266 352574
rect 459502 352338 459586 352574
rect 459822 352338 495266 352574
rect 495502 352338 495586 352574
rect 495822 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect -6806 352306 590730 352338
rect -4886 349174 588810 349206
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 59546 349174
rect 59782 348938 59866 349174
rect 60102 348938 95546 349174
rect 95782 348938 95866 349174
rect 96102 348938 131546 349174
rect 131782 348938 131866 349174
rect 132102 348938 167546 349174
rect 167782 348938 167866 349174
rect 168102 348938 203546 349174
rect 203782 348938 203866 349174
rect 204102 348938 239546 349174
rect 239782 348938 239866 349174
rect 240102 348938 275546 349174
rect 275782 348938 275866 349174
rect 276102 348938 311546 349174
rect 311782 348938 311866 349174
rect 312102 348938 347546 349174
rect 347782 348938 347866 349174
rect 348102 348938 383546 349174
rect 383782 348938 383866 349174
rect 384102 348938 419546 349174
rect 419782 348938 419866 349174
rect 420102 348938 455546 349174
rect 455782 348938 455866 349174
rect 456102 348938 491546 349174
rect 491782 348938 491866 349174
rect 492102 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect -4886 348854 588810 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 59546 348854
rect 59782 348618 59866 348854
rect 60102 348618 95546 348854
rect 95782 348618 95866 348854
rect 96102 348618 131546 348854
rect 131782 348618 131866 348854
rect 132102 348618 167546 348854
rect 167782 348618 167866 348854
rect 168102 348618 203546 348854
rect 203782 348618 203866 348854
rect 204102 348618 239546 348854
rect 239782 348618 239866 348854
rect 240102 348618 275546 348854
rect 275782 348618 275866 348854
rect 276102 348618 311546 348854
rect 311782 348618 311866 348854
rect 312102 348618 347546 348854
rect 347782 348618 347866 348854
rect 348102 348618 383546 348854
rect 383782 348618 383866 348854
rect 384102 348618 419546 348854
rect 419782 348618 419866 348854
rect 420102 348618 455546 348854
rect 455782 348618 455866 348854
rect 456102 348618 491546 348854
rect 491782 348618 491866 348854
rect 492102 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect -4886 348586 588810 348618
rect -2966 345454 586890 345486
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect -2966 345134 586890 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect -2966 344866 586890 344898
rect -8726 338614 592650 338646
rect -8726 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 84986 338614
rect 85222 338378 85306 338614
rect 85542 338378 120986 338614
rect 121222 338378 121306 338614
rect 121542 338378 156986 338614
rect 157222 338378 157306 338614
rect 157542 338378 192986 338614
rect 193222 338378 193306 338614
rect 193542 338378 228986 338614
rect 229222 338378 229306 338614
rect 229542 338378 264986 338614
rect 265222 338378 265306 338614
rect 265542 338378 300986 338614
rect 301222 338378 301306 338614
rect 301542 338378 336986 338614
rect 337222 338378 337306 338614
rect 337542 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 480986 338614
rect 481222 338378 481306 338614
rect 481542 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 592650 338614
rect -8726 338294 592650 338378
rect -8726 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 84986 338294
rect 85222 338058 85306 338294
rect 85542 338058 120986 338294
rect 121222 338058 121306 338294
rect 121542 338058 156986 338294
rect 157222 338058 157306 338294
rect 157542 338058 192986 338294
rect 193222 338058 193306 338294
rect 193542 338058 228986 338294
rect 229222 338058 229306 338294
rect 229542 338058 264986 338294
rect 265222 338058 265306 338294
rect 265542 338058 300986 338294
rect 301222 338058 301306 338294
rect 301542 338058 336986 338294
rect 337222 338058 337306 338294
rect 337542 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 480986 338294
rect 481222 338058 481306 338294
rect 481542 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 592650 338294
rect -8726 338026 592650 338058
rect -6806 334894 590730 334926
rect -6806 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 81266 334894
rect 81502 334658 81586 334894
rect 81822 334658 117266 334894
rect 117502 334658 117586 334894
rect 117822 334658 153266 334894
rect 153502 334658 153586 334894
rect 153822 334658 189266 334894
rect 189502 334658 189586 334894
rect 189822 334658 225266 334894
rect 225502 334658 225586 334894
rect 225822 334658 261266 334894
rect 261502 334658 261586 334894
rect 261822 334658 297266 334894
rect 297502 334658 297586 334894
rect 297822 334658 333266 334894
rect 333502 334658 333586 334894
rect 333822 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 405266 334894
rect 405502 334658 405586 334894
rect 405822 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 477266 334894
rect 477502 334658 477586 334894
rect 477822 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 590730 334894
rect -6806 334574 590730 334658
rect -6806 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 81266 334574
rect 81502 334338 81586 334574
rect 81822 334338 117266 334574
rect 117502 334338 117586 334574
rect 117822 334338 153266 334574
rect 153502 334338 153586 334574
rect 153822 334338 189266 334574
rect 189502 334338 189586 334574
rect 189822 334338 225266 334574
rect 225502 334338 225586 334574
rect 225822 334338 261266 334574
rect 261502 334338 261586 334574
rect 261822 334338 297266 334574
rect 297502 334338 297586 334574
rect 297822 334338 333266 334574
rect 333502 334338 333586 334574
rect 333822 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 405266 334574
rect 405502 334338 405586 334574
rect 405822 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 477266 334574
rect 477502 334338 477586 334574
rect 477822 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 590730 334574
rect -6806 334306 590730 334338
rect -4886 331174 588810 331206
rect -4886 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 185546 331174
rect 185782 330938 185866 331174
rect 186102 330938 221546 331174
rect 221782 330938 221866 331174
rect 222102 330938 257546 331174
rect 257782 330938 257866 331174
rect 258102 330938 293546 331174
rect 293782 330938 293866 331174
rect 294102 330938 329546 331174
rect 329782 330938 329866 331174
rect 330102 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 588810 331174
rect -4886 330854 588810 330938
rect -4886 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 185546 330854
rect 185782 330618 185866 330854
rect 186102 330618 221546 330854
rect 221782 330618 221866 330854
rect 222102 330618 257546 330854
rect 257782 330618 257866 330854
rect 258102 330618 293546 330854
rect 293782 330618 293866 330854
rect 294102 330618 329546 330854
rect 329782 330618 329866 330854
rect 330102 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 588810 330854
rect -4886 330586 588810 330618
rect -2966 327454 586890 327486
rect -2966 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 586890 327454
rect -2966 327134 586890 327218
rect -2966 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 586890 327134
rect -2966 326866 586890 326898
rect -8726 320614 592650 320646
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 174986 320614
rect 175222 320378 175306 320614
rect 175542 320378 210986 320614
rect 211222 320378 211306 320614
rect 211542 320378 246986 320614
rect 247222 320378 247306 320614
rect 247542 320378 282986 320614
rect 283222 320378 283306 320614
rect 283542 320378 318986 320614
rect 319222 320378 319306 320614
rect 319542 320378 354986 320614
rect 355222 320378 355306 320614
rect 355542 320378 390986 320614
rect 391222 320378 391306 320614
rect 391542 320378 426986 320614
rect 427222 320378 427306 320614
rect 427542 320378 462986 320614
rect 463222 320378 463306 320614
rect 463542 320378 498986 320614
rect 499222 320378 499306 320614
rect 499542 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect -8726 320294 592650 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 174986 320294
rect 175222 320058 175306 320294
rect 175542 320058 210986 320294
rect 211222 320058 211306 320294
rect 211542 320058 246986 320294
rect 247222 320058 247306 320294
rect 247542 320058 282986 320294
rect 283222 320058 283306 320294
rect 283542 320058 318986 320294
rect 319222 320058 319306 320294
rect 319542 320058 354986 320294
rect 355222 320058 355306 320294
rect 355542 320058 390986 320294
rect 391222 320058 391306 320294
rect 391542 320058 426986 320294
rect 427222 320058 427306 320294
rect 427542 320058 462986 320294
rect 463222 320058 463306 320294
rect 463542 320058 498986 320294
rect 499222 320058 499306 320294
rect 499542 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect -8726 320026 592650 320058
rect -6806 316894 590730 316926
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 63266 316894
rect 63502 316658 63586 316894
rect 63822 316658 171266 316894
rect 171502 316658 171586 316894
rect 171822 316658 207266 316894
rect 207502 316658 207586 316894
rect 207822 316658 243266 316894
rect 243502 316658 243586 316894
rect 243822 316658 279266 316894
rect 279502 316658 279586 316894
rect 279822 316658 315266 316894
rect 315502 316658 315586 316894
rect 315822 316658 351266 316894
rect 351502 316658 351586 316894
rect 351822 316658 387266 316894
rect 387502 316658 387586 316894
rect 387822 316658 423266 316894
rect 423502 316658 423586 316894
rect 423822 316658 459266 316894
rect 459502 316658 459586 316894
rect 459822 316658 495266 316894
rect 495502 316658 495586 316894
rect 495822 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect -6806 316574 590730 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 63266 316574
rect 63502 316338 63586 316574
rect 63822 316338 171266 316574
rect 171502 316338 171586 316574
rect 171822 316338 207266 316574
rect 207502 316338 207586 316574
rect 207822 316338 243266 316574
rect 243502 316338 243586 316574
rect 243822 316338 279266 316574
rect 279502 316338 279586 316574
rect 279822 316338 315266 316574
rect 315502 316338 315586 316574
rect 315822 316338 351266 316574
rect 351502 316338 351586 316574
rect 351822 316338 387266 316574
rect 387502 316338 387586 316574
rect 387822 316338 423266 316574
rect 423502 316338 423586 316574
rect 423822 316338 459266 316574
rect 459502 316338 459586 316574
rect 459822 316338 495266 316574
rect 495502 316338 495586 316574
rect 495822 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect -6806 316306 590730 316338
rect -4886 313174 588810 313206
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 59546 313174
rect 59782 312938 59866 313174
rect 60102 312938 167546 313174
rect 167782 312938 167866 313174
rect 168102 312938 203546 313174
rect 203782 312938 203866 313174
rect 204102 312938 239546 313174
rect 239782 312938 239866 313174
rect 240102 312938 275546 313174
rect 275782 312938 275866 313174
rect 276102 312938 311546 313174
rect 311782 312938 311866 313174
rect 312102 312938 347546 313174
rect 347782 312938 347866 313174
rect 348102 312938 383546 313174
rect 383782 312938 383866 313174
rect 384102 312938 419546 313174
rect 419782 312938 419866 313174
rect 420102 312938 455546 313174
rect 455782 312938 455866 313174
rect 456102 312938 491546 313174
rect 491782 312938 491866 313174
rect 492102 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect -4886 312854 588810 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 59546 312854
rect 59782 312618 59866 312854
rect 60102 312618 167546 312854
rect 167782 312618 167866 312854
rect 168102 312618 203546 312854
rect 203782 312618 203866 312854
rect 204102 312618 239546 312854
rect 239782 312618 239866 312854
rect 240102 312618 275546 312854
rect 275782 312618 275866 312854
rect 276102 312618 311546 312854
rect 311782 312618 311866 312854
rect 312102 312618 347546 312854
rect 347782 312618 347866 312854
rect 348102 312618 383546 312854
rect 383782 312618 383866 312854
rect 384102 312618 419546 312854
rect 419782 312618 419866 312854
rect 420102 312618 455546 312854
rect 455782 312618 455866 312854
rect 456102 312618 491546 312854
rect 491782 312618 491866 312854
rect 492102 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect -4886 312586 588810 312618
rect -2966 309454 586890 309486
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 88380 309454
rect 88616 309218 119100 309454
rect 119336 309218 149820 309454
rect 150056 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect -2966 309134 586890 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 88380 309134
rect 88616 308898 119100 309134
rect 119336 308898 149820 309134
rect 150056 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect -2966 308866 586890 308898
rect -8726 302614 592650 302646
rect -8726 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 192986 302614
rect 193222 302378 193306 302614
rect 193542 302378 228986 302614
rect 229222 302378 229306 302614
rect 229542 302378 264986 302614
rect 265222 302378 265306 302614
rect 265542 302378 300986 302614
rect 301222 302378 301306 302614
rect 301542 302378 336986 302614
rect 337222 302378 337306 302614
rect 337542 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 408986 302614
rect 409222 302378 409306 302614
rect 409542 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 592650 302614
rect -8726 302294 592650 302378
rect -8726 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 192986 302294
rect 193222 302058 193306 302294
rect 193542 302058 228986 302294
rect 229222 302058 229306 302294
rect 229542 302058 264986 302294
rect 265222 302058 265306 302294
rect 265542 302058 300986 302294
rect 301222 302058 301306 302294
rect 301542 302058 336986 302294
rect 337222 302058 337306 302294
rect 337542 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 408986 302294
rect 409222 302058 409306 302294
rect 409542 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 592650 302294
rect -8726 302026 592650 302058
rect -6806 298894 590730 298926
rect -6806 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 189266 298894
rect 189502 298658 189586 298894
rect 189822 298658 225266 298894
rect 225502 298658 225586 298894
rect 225822 298658 261266 298894
rect 261502 298658 261586 298894
rect 261822 298658 297266 298894
rect 297502 298658 297586 298894
rect 297822 298658 333266 298894
rect 333502 298658 333586 298894
rect 333822 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 405266 298894
rect 405502 298658 405586 298894
rect 405822 298658 441266 298894
rect 441502 298658 441586 298894
rect 441822 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 590730 298894
rect -6806 298574 590730 298658
rect -6806 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 189266 298574
rect 189502 298338 189586 298574
rect 189822 298338 225266 298574
rect 225502 298338 225586 298574
rect 225822 298338 261266 298574
rect 261502 298338 261586 298574
rect 261822 298338 297266 298574
rect 297502 298338 297586 298574
rect 297822 298338 333266 298574
rect 333502 298338 333586 298574
rect 333822 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 405266 298574
rect 405502 298338 405586 298574
rect 405822 298338 441266 298574
rect 441502 298338 441586 298574
rect 441822 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 590730 298574
rect -6806 298306 590730 298338
rect -4886 295174 588810 295206
rect -4886 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 185546 295174
rect 185782 294938 185866 295174
rect 186102 294938 221546 295174
rect 221782 294938 221866 295174
rect 222102 294938 257546 295174
rect 257782 294938 257866 295174
rect 258102 294938 293546 295174
rect 293782 294938 293866 295174
rect 294102 294938 329546 295174
rect 329782 294938 329866 295174
rect 330102 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 588810 295174
rect -4886 294854 588810 294938
rect -4886 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 185546 294854
rect 185782 294618 185866 294854
rect 186102 294618 221546 294854
rect 221782 294618 221866 294854
rect 222102 294618 257546 294854
rect 257782 294618 257866 294854
rect 258102 294618 293546 294854
rect 293782 294618 293866 294854
rect 294102 294618 329546 294854
rect 329782 294618 329866 294854
rect 330102 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 588810 294854
rect -4886 294586 588810 294618
rect -2966 291454 586890 291486
rect -2966 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 73020 291454
rect 73256 291218 103740 291454
rect 103976 291218 134460 291454
rect 134696 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 586890 291454
rect -2966 291134 586890 291218
rect -2966 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 73020 291134
rect 73256 290898 103740 291134
rect 103976 290898 134460 291134
rect 134696 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 586890 291134
rect -2966 290866 586890 290898
rect -8726 284614 592650 284646
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 174986 284614
rect 175222 284378 175306 284614
rect 175542 284378 246986 284614
rect 247222 284378 247306 284614
rect 247542 284378 282986 284614
rect 283222 284378 283306 284614
rect 283542 284378 318986 284614
rect 319222 284378 319306 284614
rect 319542 284378 354986 284614
rect 355222 284378 355306 284614
rect 355542 284378 390986 284614
rect 391222 284378 391306 284614
rect 391542 284378 426986 284614
rect 427222 284378 427306 284614
rect 427542 284378 462986 284614
rect 463222 284378 463306 284614
rect 463542 284378 498986 284614
rect 499222 284378 499306 284614
rect 499542 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect -8726 284294 592650 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 174986 284294
rect 175222 284058 175306 284294
rect 175542 284058 246986 284294
rect 247222 284058 247306 284294
rect 247542 284058 282986 284294
rect 283222 284058 283306 284294
rect 283542 284058 318986 284294
rect 319222 284058 319306 284294
rect 319542 284058 354986 284294
rect 355222 284058 355306 284294
rect 355542 284058 390986 284294
rect 391222 284058 391306 284294
rect 391542 284058 426986 284294
rect 427222 284058 427306 284294
rect 427542 284058 462986 284294
rect 463222 284058 463306 284294
rect 463542 284058 498986 284294
rect 499222 284058 499306 284294
rect 499542 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect -8726 284026 592650 284058
rect -6806 280894 590730 280926
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 63266 280894
rect 63502 280658 63586 280894
rect 63822 280658 171266 280894
rect 171502 280658 171586 280894
rect 171822 280658 279266 280894
rect 279502 280658 279586 280894
rect 279822 280658 315266 280894
rect 315502 280658 315586 280894
rect 315822 280658 351266 280894
rect 351502 280658 351586 280894
rect 351822 280658 387266 280894
rect 387502 280658 387586 280894
rect 387822 280658 423266 280894
rect 423502 280658 423586 280894
rect 423822 280658 459266 280894
rect 459502 280658 459586 280894
rect 459822 280658 495266 280894
rect 495502 280658 495586 280894
rect 495822 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect -6806 280574 590730 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 63266 280574
rect 63502 280338 63586 280574
rect 63822 280338 171266 280574
rect 171502 280338 171586 280574
rect 171822 280338 279266 280574
rect 279502 280338 279586 280574
rect 279822 280338 315266 280574
rect 315502 280338 315586 280574
rect 315822 280338 351266 280574
rect 351502 280338 351586 280574
rect 351822 280338 387266 280574
rect 387502 280338 387586 280574
rect 387822 280338 423266 280574
rect 423502 280338 423586 280574
rect 423822 280338 459266 280574
rect 459502 280338 459586 280574
rect 459822 280338 495266 280574
rect 495502 280338 495586 280574
rect 495822 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect -6806 280306 590730 280338
rect -4886 277174 588810 277206
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 59546 277174
rect 59782 276938 59866 277174
rect 60102 276938 167546 277174
rect 167782 276938 167866 277174
rect 168102 276938 275546 277174
rect 275782 276938 275866 277174
rect 276102 276938 311546 277174
rect 311782 276938 311866 277174
rect 312102 276938 347546 277174
rect 347782 276938 347866 277174
rect 348102 276938 383546 277174
rect 383782 276938 383866 277174
rect 384102 276938 419546 277174
rect 419782 276938 419866 277174
rect 420102 276938 455546 277174
rect 455782 276938 455866 277174
rect 456102 276938 491546 277174
rect 491782 276938 491866 277174
rect 492102 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect -4886 276854 588810 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 59546 276854
rect 59782 276618 59866 276854
rect 60102 276618 167546 276854
rect 167782 276618 167866 276854
rect 168102 276618 275546 276854
rect 275782 276618 275866 276854
rect 276102 276618 311546 276854
rect 311782 276618 311866 276854
rect 312102 276618 347546 276854
rect 347782 276618 347866 276854
rect 348102 276618 383546 276854
rect 383782 276618 383866 276854
rect 384102 276618 419546 276854
rect 419782 276618 419866 276854
rect 420102 276618 455546 276854
rect 455782 276618 455866 276854
rect 456102 276618 491546 276854
rect 491782 276618 491866 276854
rect 492102 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect -4886 276586 588810 276618
rect -2966 273454 586890 273486
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 88380 273454
rect 88616 273218 119100 273454
rect 119336 273218 149820 273454
rect 150056 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 219810 273454
rect 220046 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect -2966 273134 586890 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 88380 273134
rect 88616 272898 119100 273134
rect 119336 272898 149820 273134
rect 150056 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 219810 273134
rect 220046 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect -2966 272866 586890 272898
rect -8726 266614 592650 266646
rect -8726 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 192986 266614
rect 193222 266378 193306 266614
rect 193542 266378 264986 266614
rect 265222 266378 265306 266614
rect 265542 266378 300986 266614
rect 301222 266378 301306 266614
rect 301542 266378 336986 266614
rect 337222 266378 337306 266614
rect 337542 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 592650 266614
rect -8726 266294 592650 266378
rect -8726 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 192986 266294
rect 193222 266058 193306 266294
rect 193542 266058 264986 266294
rect 265222 266058 265306 266294
rect 265542 266058 300986 266294
rect 301222 266058 301306 266294
rect 301542 266058 336986 266294
rect 337222 266058 337306 266294
rect 337542 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 592650 266294
rect -8726 266026 592650 266058
rect -6806 262894 590730 262926
rect -6806 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 261266 262894
rect 261502 262658 261586 262894
rect 261822 262658 297266 262894
rect 297502 262658 297586 262894
rect 297822 262658 333266 262894
rect 333502 262658 333586 262894
rect 333822 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 590730 262894
rect -6806 262574 590730 262658
rect -6806 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 261266 262574
rect 261502 262338 261586 262574
rect 261822 262338 297266 262574
rect 297502 262338 297586 262574
rect 297822 262338 333266 262574
rect 333502 262338 333586 262574
rect 333822 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 590730 262574
rect -6806 262306 590730 262338
rect -4886 259174 588810 259206
rect -4886 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 257546 259174
rect 257782 258938 257866 259174
rect 258102 258938 293546 259174
rect 293782 258938 293866 259174
rect 294102 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 588810 259174
rect -4886 258854 588810 258938
rect -4886 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 257546 258854
rect 257782 258618 257866 258854
rect 258102 258618 293546 258854
rect 293782 258618 293866 258854
rect 294102 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 588810 258854
rect -4886 258586 588810 258618
rect -2966 255454 586890 255486
rect -2966 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 73020 255454
rect 73256 255218 103740 255454
rect 103976 255218 134460 255454
rect 134696 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 204450 255454
rect 204686 255218 235170 255454
rect 235406 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 586890 255454
rect -2966 255134 586890 255218
rect -2966 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 73020 255134
rect 73256 254898 103740 255134
rect 103976 254898 134460 255134
rect 134696 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 204450 255134
rect 204686 254898 235170 255134
rect 235406 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 586890 255134
rect -2966 254866 586890 254898
rect -8726 248614 592650 248646
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 174986 248614
rect 175222 248378 175306 248614
rect 175542 248378 246986 248614
rect 247222 248378 247306 248614
rect 247542 248378 282986 248614
rect 283222 248378 283306 248614
rect 283542 248378 318986 248614
rect 319222 248378 319306 248614
rect 319542 248378 354986 248614
rect 355222 248378 355306 248614
rect 355542 248378 390986 248614
rect 391222 248378 391306 248614
rect 391542 248378 426986 248614
rect 427222 248378 427306 248614
rect 427542 248378 462986 248614
rect 463222 248378 463306 248614
rect 463542 248378 498986 248614
rect 499222 248378 499306 248614
rect 499542 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect -8726 248294 592650 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 174986 248294
rect 175222 248058 175306 248294
rect 175542 248058 246986 248294
rect 247222 248058 247306 248294
rect 247542 248058 282986 248294
rect 283222 248058 283306 248294
rect 283542 248058 318986 248294
rect 319222 248058 319306 248294
rect 319542 248058 354986 248294
rect 355222 248058 355306 248294
rect 355542 248058 390986 248294
rect 391222 248058 391306 248294
rect 391542 248058 426986 248294
rect 427222 248058 427306 248294
rect 427542 248058 462986 248294
rect 463222 248058 463306 248294
rect 463542 248058 498986 248294
rect 499222 248058 499306 248294
rect 499542 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect -8726 248026 592650 248058
rect -6806 244894 590730 244926
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 63266 244894
rect 63502 244658 63586 244894
rect 63822 244658 171266 244894
rect 171502 244658 171586 244894
rect 171822 244658 279266 244894
rect 279502 244658 279586 244894
rect 279822 244658 315266 244894
rect 315502 244658 315586 244894
rect 315822 244658 351266 244894
rect 351502 244658 351586 244894
rect 351822 244658 387266 244894
rect 387502 244658 387586 244894
rect 387822 244658 423266 244894
rect 423502 244658 423586 244894
rect 423822 244658 459266 244894
rect 459502 244658 459586 244894
rect 459822 244658 495266 244894
rect 495502 244658 495586 244894
rect 495822 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect -6806 244574 590730 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 63266 244574
rect 63502 244338 63586 244574
rect 63822 244338 171266 244574
rect 171502 244338 171586 244574
rect 171822 244338 279266 244574
rect 279502 244338 279586 244574
rect 279822 244338 315266 244574
rect 315502 244338 315586 244574
rect 315822 244338 351266 244574
rect 351502 244338 351586 244574
rect 351822 244338 387266 244574
rect 387502 244338 387586 244574
rect 387822 244338 423266 244574
rect 423502 244338 423586 244574
rect 423822 244338 459266 244574
rect 459502 244338 459586 244574
rect 459822 244338 495266 244574
rect 495502 244338 495586 244574
rect 495822 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect -6806 244306 590730 244338
rect -4886 241174 588810 241206
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 59546 241174
rect 59782 240938 59866 241174
rect 60102 240938 167546 241174
rect 167782 240938 167866 241174
rect 168102 240938 275546 241174
rect 275782 240938 275866 241174
rect 276102 240938 311546 241174
rect 311782 240938 311866 241174
rect 312102 240938 347546 241174
rect 347782 240938 347866 241174
rect 348102 240938 383546 241174
rect 383782 240938 383866 241174
rect 384102 240938 419546 241174
rect 419782 240938 419866 241174
rect 420102 240938 455546 241174
rect 455782 240938 455866 241174
rect 456102 240938 491546 241174
rect 491782 240938 491866 241174
rect 492102 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect -4886 240854 588810 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 59546 240854
rect 59782 240618 59866 240854
rect 60102 240618 167546 240854
rect 167782 240618 167866 240854
rect 168102 240618 275546 240854
rect 275782 240618 275866 240854
rect 276102 240618 311546 240854
rect 311782 240618 311866 240854
rect 312102 240618 347546 240854
rect 347782 240618 347866 240854
rect 348102 240618 383546 240854
rect 383782 240618 383866 240854
rect 384102 240618 419546 240854
rect 419782 240618 419866 240854
rect 420102 240618 455546 240854
rect 455782 240618 455866 240854
rect 456102 240618 491546 240854
rect 491782 240618 491866 240854
rect 492102 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect -4886 240586 588810 240618
rect -2966 237454 586890 237486
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect -2966 237134 586890 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect -2966 236866 586890 236898
rect -8726 230614 592650 230646
rect -8726 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 84986 230614
rect 85222 230378 85306 230614
rect 85542 230378 120986 230614
rect 121222 230378 121306 230614
rect 121542 230378 156986 230614
rect 157222 230378 157306 230614
rect 157542 230378 192986 230614
rect 193222 230378 193306 230614
rect 193542 230378 228986 230614
rect 229222 230378 229306 230614
rect 229542 230378 264986 230614
rect 265222 230378 265306 230614
rect 265542 230378 300986 230614
rect 301222 230378 301306 230614
rect 301542 230378 336986 230614
rect 337222 230378 337306 230614
rect 337542 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 592650 230614
rect -8726 230294 592650 230378
rect -8726 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 84986 230294
rect 85222 230058 85306 230294
rect 85542 230058 120986 230294
rect 121222 230058 121306 230294
rect 121542 230058 156986 230294
rect 157222 230058 157306 230294
rect 157542 230058 192986 230294
rect 193222 230058 193306 230294
rect 193542 230058 228986 230294
rect 229222 230058 229306 230294
rect 229542 230058 264986 230294
rect 265222 230058 265306 230294
rect 265542 230058 300986 230294
rect 301222 230058 301306 230294
rect 301542 230058 336986 230294
rect 337222 230058 337306 230294
rect 337542 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 592650 230294
rect -8726 230026 592650 230058
rect -6806 226894 590730 226926
rect -6806 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 81266 226894
rect 81502 226658 81586 226894
rect 81822 226658 117266 226894
rect 117502 226658 117586 226894
rect 117822 226658 153266 226894
rect 153502 226658 153586 226894
rect 153822 226658 189266 226894
rect 189502 226658 189586 226894
rect 189822 226658 225266 226894
rect 225502 226658 225586 226894
rect 225822 226658 261266 226894
rect 261502 226658 261586 226894
rect 261822 226658 297266 226894
rect 297502 226658 297586 226894
rect 297822 226658 333266 226894
rect 333502 226658 333586 226894
rect 333822 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 405266 226894
rect 405502 226658 405586 226894
rect 405822 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 590730 226894
rect -6806 226574 590730 226658
rect -6806 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 81266 226574
rect 81502 226338 81586 226574
rect 81822 226338 117266 226574
rect 117502 226338 117586 226574
rect 117822 226338 153266 226574
rect 153502 226338 153586 226574
rect 153822 226338 189266 226574
rect 189502 226338 189586 226574
rect 189822 226338 225266 226574
rect 225502 226338 225586 226574
rect 225822 226338 261266 226574
rect 261502 226338 261586 226574
rect 261822 226338 297266 226574
rect 297502 226338 297586 226574
rect 297822 226338 333266 226574
rect 333502 226338 333586 226574
rect 333822 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 405266 226574
rect 405502 226338 405586 226574
rect 405822 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 590730 226574
rect -6806 226306 590730 226338
rect -4886 223174 588810 223206
rect -4886 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 77546 223174
rect 77782 222938 77866 223174
rect 78102 222938 113546 223174
rect 113782 222938 113866 223174
rect 114102 222938 149546 223174
rect 149782 222938 149866 223174
rect 150102 222938 185546 223174
rect 185782 222938 185866 223174
rect 186102 222938 221546 223174
rect 221782 222938 221866 223174
rect 222102 222938 257546 223174
rect 257782 222938 257866 223174
rect 258102 222938 293546 223174
rect 293782 222938 293866 223174
rect 294102 222938 329546 223174
rect 329782 222938 329866 223174
rect 330102 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 588810 223174
rect -4886 222854 588810 222938
rect -4886 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 77546 222854
rect 77782 222618 77866 222854
rect 78102 222618 113546 222854
rect 113782 222618 113866 222854
rect 114102 222618 149546 222854
rect 149782 222618 149866 222854
rect 150102 222618 185546 222854
rect 185782 222618 185866 222854
rect 186102 222618 221546 222854
rect 221782 222618 221866 222854
rect 222102 222618 257546 222854
rect 257782 222618 257866 222854
rect 258102 222618 293546 222854
rect 293782 222618 293866 222854
rect 294102 222618 329546 222854
rect 329782 222618 329866 222854
rect 330102 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 588810 222854
rect -4886 222586 588810 222618
rect -2966 219454 586890 219486
rect -2966 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 586890 219454
rect -2966 219134 586890 219218
rect -2966 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 586890 219134
rect -2966 218866 586890 218898
rect -8726 212614 592650 212646
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 66986 212614
rect 67222 212378 67306 212614
rect 67542 212378 102986 212614
rect 103222 212378 103306 212614
rect 103542 212378 138986 212614
rect 139222 212378 139306 212614
rect 139542 212378 174986 212614
rect 175222 212378 175306 212614
rect 175542 212378 210986 212614
rect 211222 212378 211306 212614
rect 211542 212378 246986 212614
rect 247222 212378 247306 212614
rect 247542 212378 282986 212614
rect 283222 212378 283306 212614
rect 283542 212378 318986 212614
rect 319222 212378 319306 212614
rect 319542 212378 354986 212614
rect 355222 212378 355306 212614
rect 355542 212378 390986 212614
rect 391222 212378 391306 212614
rect 391542 212378 426986 212614
rect 427222 212378 427306 212614
rect 427542 212378 462986 212614
rect 463222 212378 463306 212614
rect 463542 212378 498986 212614
rect 499222 212378 499306 212614
rect 499542 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect -8726 212294 592650 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 66986 212294
rect 67222 212058 67306 212294
rect 67542 212058 102986 212294
rect 103222 212058 103306 212294
rect 103542 212058 138986 212294
rect 139222 212058 139306 212294
rect 139542 212058 174986 212294
rect 175222 212058 175306 212294
rect 175542 212058 210986 212294
rect 211222 212058 211306 212294
rect 211542 212058 246986 212294
rect 247222 212058 247306 212294
rect 247542 212058 282986 212294
rect 283222 212058 283306 212294
rect 283542 212058 318986 212294
rect 319222 212058 319306 212294
rect 319542 212058 354986 212294
rect 355222 212058 355306 212294
rect 355542 212058 390986 212294
rect 391222 212058 391306 212294
rect 391542 212058 426986 212294
rect 427222 212058 427306 212294
rect 427542 212058 462986 212294
rect 463222 212058 463306 212294
rect 463542 212058 498986 212294
rect 499222 212058 499306 212294
rect 499542 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect -8726 212026 592650 212058
rect -6806 208894 590730 208926
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 63266 208894
rect 63502 208658 63586 208894
rect 63822 208658 99266 208894
rect 99502 208658 99586 208894
rect 99822 208658 135266 208894
rect 135502 208658 135586 208894
rect 135822 208658 171266 208894
rect 171502 208658 171586 208894
rect 171822 208658 207266 208894
rect 207502 208658 207586 208894
rect 207822 208658 243266 208894
rect 243502 208658 243586 208894
rect 243822 208658 279266 208894
rect 279502 208658 279586 208894
rect 279822 208658 315266 208894
rect 315502 208658 315586 208894
rect 315822 208658 351266 208894
rect 351502 208658 351586 208894
rect 351822 208658 387266 208894
rect 387502 208658 387586 208894
rect 387822 208658 423266 208894
rect 423502 208658 423586 208894
rect 423822 208658 459266 208894
rect 459502 208658 459586 208894
rect 459822 208658 495266 208894
rect 495502 208658 495586 208894
rect 495822 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect -6806 208574 590730 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 63266 208574
rect 63502 208338 63586 208574
rect 63822 208338 99266 208574
rect 99502 208338 99586 208574
rect 99822 208338 135266 208574
rect 135502 208338 135586 208574
rect 135822 208338 171266 208574
rect 171502 208338 171586 208574
rect 171822 208338 207266 208574
rect 207502 208338 207586 208574
rect 207822 208338 243266 208574
rect 243502 208338 243586 208574
rect 243822 208338 279266 208574
rect 279502 208338 279586 208574
rect 279822 208338 315266 208574
rect 315502 208338 315586 208574
rect 315822 208338 351266 208574
rect 351502 208338 351586 208574
rect 351822 208338 387266 208574
rect 387502 208338 387586 208574
rect 387822 208338 423266 208574
rect 423502 208338 423586 208574
rect 423822 208338 459266 208574
rect 459502 208338 459586 208574
rect 459822 208338 495266 208574
rect 495502 208338 495586 208574
rect 495822 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect -6806 208306 590730 208338
rect -4886 205174 588810 205206
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 59546 205174
rect 59782 204938 59866 205174
rect 60102 204938 95546 205174
rect 95782 204938 95866 205174
rect 96102 204938 131546 205174
rect 131782 204938 131866 205174
rect 132102 204938 167546 205174
rect 167782 204938 167866 205174
rect 168102 204938 203546 205174
rect 203782 204938 203866 205174
rect 204102 204938 239546 205174
rect 239782 204938 239866 205174
rect 240102 204938 275546 205174
rect 275782 204938 275866 205174
rect 276102 204938 311546 205174
rect 311782 204938 311866 205174
rect 312102 204938 347546 205174
rect 347782 204938 347866 205174
rect 348102 204938 383546 205174
rect 383782 204938 383866 205174
rect 384102 204938 419546 205174
rect 419782 204938 419866 205174
rect 420102 204938 455546 205174
rect 455782 204938 455866 205174
rect 456102 204938 491546 205174
rect 491782 204938 491866 205174
rect 492102 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect -4886 204854 588810 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 59546 204854
rect 59782 204618 59866 204854
rect 60102 204618 95546 204854
rect 95782 204618 95866 204854
rect 96102 204618 131546 204854
rect 131782 204618 131866 204854
rect 132102 204618 167546 204854
rect 167782 204618 167866 204854
rect 168102 204618 203546 204854
rect 203782 204618 203866 204854
rect 204102 204618 239546 204854
rect 239782 204618 239866 204854
rect 240102 204618 275546 204854
rect 275782 204618 275866 204854
rect 276102 204618 311546 204854
rect 311782 204618 311866 204854
rect 312102 204618 347546 204854
rect 347782 204618 347866 204854
rect 348102 204618 383546 204854
rect 383782 204618 383866 204854
rect 384102 204618 419546 204854
rect 419782 204618 419866 204854
rect 420102 204618 455546 204854
rect 455782 204618 455866 204854
rect 456102 204618 491546 204854
rect 491782 204618 491866 204854
rect 492102 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect -4886 204586 588810 204618
rect -2966 201454 586890 201486
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect -2966 201134 586890 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect -2966 200866 586890 200898
rect -8726 194614 592650 194646
rect -8726 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 84986 194614
rect 85222 194378 85306 194614
rect 85542 194378 120986 194614
rect 121222 194378 121306 194614
rect 121542 194378 156986 194614
rect 157222 194378 157306 194614
rect 157542 194378 192986 194614
rect 193222 194378 193306 194614
rect 193542 194378 228986 194614
rect 229222 194378 229306 194614
rect 229542 194378 264986 194614
rect 265222 194378 265306 194614
rect 265542 194378 300986 194614
rect 301222 194378 301306 194614
rect 301542 194378 336986 194614
rect 337222 194378 337306 194614
rect 337542 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 592650 194614
rect -8726 194294 592650 194378
rect -8726 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 84986 194294
rect 85222 194058 85306 194294
rect 85542 194058 120986 194294
rect 121222 194058 121306 194294
rect 121542 194058 156986 194294
rect 157222 194058 157306 194294
rect 157542 194058 192986 194294
rect 193222 194058 193306 194294
rect 193542 194058 228986 194294
rect 229222 194058 229306 194294
rect 229542 194058 264986 194294
rect 265222 194058 265306 194294
rect 265542 194058 300986 194294
rect 301222 194058 301306 194294
rect 301542 194058 336986 194294
rect 337222 194058 337306 194294
rect 337542 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 592650 194294
rect -8726 194026 592650 194058
rect -6806 190894 590730 190926
rect -6806 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 81266 190894
rect 81502 190658 81586 190894
rect 81822 190658 117266 190894
rect 117502 190658 117586 190894
rect 117822 190658 153266 190894
rect 153502 190658 153586 190894
rect 153822 190658 189266 190894
rect 189502 190658 189586 190894
rect 189822 190658 225266 190894
rect 225502 190658 225586 190894
rect 225822 190658 261266 190894
rect 261502 190658 261586 190894
rect 261822 190658 297266 190894
rect 297502 190658 297586 190894
rect 297822 190658 333266 190894
rect 333502 190658 333586 190894
rect 333822 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 590730 190894
rect -6806 190574 590730 190658
rect -6806 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 81266 190574
rect 81502 190338 81586 190574
rect 81822 190338 117266 190574
rect 117502 190338 117586 190574
rect 117822 190338 153266 190574
rect 153502 190338 153586 190574
rect 153822 190338 189266 190574
rect 189502 190338 189586 190574
rect 189822 190338 225266 190574
rect 225502 190338 225586 190574
rect 225822 190338 261266 190574
rect 261502 190338 261586 190574
rect 261822 190338 297266 190574
rect 297502 190338 297586 190574
rect 297822 190338 333266 190574
rect 333502 190338 333586 190574
rect 333822 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 590730 190574
rect -6806 190306 590730 190338
rect -4886 187174 588810 187206
rect -4886 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 77546 187174
rect 77782 186938 77866 187174
rect 78102 186938 113546 187174
rect 113782 186938 113866 187174
rect 114102 186938 149546 187174
rect 149782 186938 149866 187174
rect 150102 186938 185546 187174
rect 185782 186938 185866 187174
rect 186102 186938 221546 187174
rect 221782 186938 221866 187174
rect 222102 186938 257546 187174
rect 257782 186938 257866 187174
rect 258102 186938 293546 187174
rect 293782 186938 293866 187174
rect 294102 186938 329546 187174
rect 329782 186938 329866 187174
rect 330102 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 588810 187174
rect -4886 186854 588810 186938
rect -4886 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 77546 186854
rect 77782 186618 77866 186854
rect 78102 186618 113546 186854
rect 113782 186618 113866 186854
rect 114102 186618 149546 186854
rect 149782 186618 149866 186854
rect 150102 186618 185546 186854
rect 185782 186618 185866 186854
rect 186102 186618 221546 186854
rect 221782 186618 221866 186854
rect 222102 186618 257546 186854
rect 257782 186618 257866 186854
rect 258102 186618 293546 186854
rect 293782 186618 293866 186854
rect 294102 186618 329546 186854
rect 329782 186618 329866 186854
rect 330102 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 588810 186854
rect -4886 186586 588810 186618
rect -2966 183454 586890 183486
rect -2966 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 586890 183454
rect -2966 183134 586890 183218
rect -2966 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 586890 183134
rect -2966 182866 586890 182898
rect -8726 176614 592650 176646
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 174986 176614
rect 175222 176378 175306 176614
rect 175542 176378 210986 176614
rect 211222 176378 211306 176614
rect 211542 176378 246986 176614
rect 247222 176378 247306 176614
rect 247542 176378 282986 176614
rect 283222 176378 283306 176614
rect 283542 176378 318986 176614
rect 319222 176378 319306 176614
rect 319542 176378 354986 176614
rect 355222 176378 355306 176614
rect 355542 176378 390986 176614
rect 391222 176378 391306 176614
rect 391542 176378 426986 176614
rect 427222 176378 427306 176614
rect 427542 176378 462986 176614
rect 463222 176378 463306 176614
rect 463542 176378 498986 176614
rect 499222 176378 499306 176614
rect 499542 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect -8726 176294 592650 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 174986 176294
rect 175222 176058 175306 176294
rect 175542 176058 210986 176294
rect 211222 176058 211306 176294
rect 211542 176058 246986 176294
rect 247222 176058 247306 176294
rect 247542 176058 282986 176294
rect 283222 176058 283306 176294
rect 283542 176058 318986 176294
rect 319222 176058 319306 176294
rect 319542 176058 354986 176294
rect 355222 176058 355306 176294
rect 355542 176058 390986 176294
rect 391222 176058 391306 176294
rect 391542 176058 426986 176294
rect 427222 176058 427306 176294
rect 427542 176058 462986 176294
rect 463222 176058 463306 176294
rect 463542 176058 498986 176294
rect 499222 176058 499306 176294
rect 499542 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect -8726 176026 592650 176058
rect -6806 172894 590730 172926
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 63266 172894
rect 63502 172658 63586 172894
rect 63822 172658 171266 172894
rect 171502 172658 171586 172894
rect 171822 172658 207266 172894
rect 207502 172658 207586 172894
rect 207822 172658 243266 172894
rect 243502 172658 243586 172894
rect 243822 172658 315266 172894
rect 315502 172658 315586 172894
rect 315822 172658 351266 172894
rect 351502 172658 351586 172894
rect 351822 172658 387266 172894
rect 387502 172658 387586 172894
rect 387822 172658 423266 172894
rect 423502 172658 423586 172894
rect 423822 172658 459266 172894
rect 459502 172658 459586 172894
rect 459822 172658 495266 172894
rect 495502 172658 495586 172894
rect 495822 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect -6806 172574 590730 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 63266 172574
rect 63502 172338 63586 172574
rect 63822 172338 171266 172574
rect 171502 172338 171586 172574
rect 171822 172338 207266 172574
rect 207502 172338 207586 172574
rect 207822 172338 243266 172574
rect 243502 172338 243586 172574
rect 243822 172338 315266 172574
rect 315502 172338 315586 172574
rect 315822 172338 351266 172574
rect 351502 172338 351586 172574
rect 351822 172338 387266 172574
rect 387502 172338 387586 172574
rect 387822 172338 423266 172574
rect 423502 172338 423586 172574
rect 423822 172338 459266 172574
rect 459502 172338 459586 172574
rect 459822 172338 495266 172574
rect 495502 172338 495586 172574
rect 495822 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect -6806 172306 590730 172338
rect -4886 169174 588810 169206
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 59546 169174
rect 59782 168938 59866 169174
rect 60102 168938 167546 169174
rect 167782 168938 167866 169174
rect 168102 168938 203546 169174
rect 203782 168938 203866 169174
rect 204102 168938 239546 169174
rect 239782 168938 239866 169174
rect 240102 168938 311546 169174
rect 311782 168938 311866 169174
rect 312102 168938 347546 169174
rect 347782 168938 347866 169174
rect 348102 168938 383546 169174
rect 383782 168938 383866 169174
rect 384102 168938 419546 169174
rect 419782 168938 419866 169174
rect 420102 168938 455546 169174
rect 455782 168938 455866 169174
rect 456102 168938 491546 169174
rect 491782 168938 491866 169174
rect 492102 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect -4886 168854 588810 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 59546 168854
rect 59782 168618 59866 168854
rect 60102 168618 167546 168854
rect 167782 168618 167866 168854
rect 168102 168618 203546 168854
rect 203782 168618 203866 168854
rect 204102 168618 239546 168854
rect 239782 168618 239866 168854
rect 240102 168618 311546 168854
rect 311782 168618 311866 168854
rect 312102 168618 347546 168854
rect 347782 168618 347866 168854
rect 348102 168618 383546 168854
rect 383782 168618 383866 168854
rect 384102 168618 419546 168854
rect 419782 168618 419866 168854
rect 420102 168618 455546 168854
rect 455782 168618 455866 168854
rect 456102 168618 491546 168854
rect 491782 168618 491866 168854
rect 492102 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect -4886 168586 588810 168618
rect -2966 165454 586890 165486
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 69128 165454
rect 69364 165218 164192 165454
rect 164428 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 221249 165454
rect 221485 165218 224513 165454
rect 224749 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 272249 165454
rect 272485 165218 275513 165454
rect 275749 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect -2966 165134 586890 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 69128 165134
rect 69364 164898 164192 165134
rect 164428 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 221249 165134
rect 221485 164898 224513 165134
rect 224749 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 272249 165134
rect 272485 164898 275513 165134
rect 275749 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect -2966 164866 586890 164898
rect -8726 158614 592650 158646
rect -8726 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 192986 158614
rect 193222 158378 193306 158614
rect 193542 158378 264986 158614
rect 265222 158378 265306 158614
rect 265542 158378 300986 158614
rect 301222 158378 301306 158614
rect 301542 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 592650 158614
rect -8726 158294 592650 158378
rect -8726 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 192986 158294
rect 193222 158058 193306 158294
rect 193542 158058 264986 158294
rect 265222 158058 265306 158294
rect 265542 158058 300986 158294
rect 301222 158058 301306 158294
rect 301542 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 592650 158294
rect -8726 158026 592650 158058
rect -6806 154894 590730 154926
rect -6806 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 189266 154894
rect 189502 154658 189586 154894
rect 189822 154658 261266 154894
rect 261502 154658 261586 154894
rect 261822 154658 297266 154894
rect 297502 154658 297586 154894
rect 297822 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 441266 154894
rect 441502 154658 441586 154894
rect 441822 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 590730 154894
rect -6806 154574 590730 154658
rect -6806 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 189266 154574
rect 189502 154338 189586 154574
rect 189822 154338 261266 154574
rect 261502 154338 261586 154574
rect 261822 154338 297266 154574
rect 297502 154338 297586 154574
rect 297822 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 441266 154574
rect 441502 154338 441586 154574
rect 441822 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 590730 154574
rect -6806 154306 590730 154338
rect -4886 151174 588810 151206
rect -4886 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 257546 151174
rect 257782 150938 257866 151174
rect 258102 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 588810 151174
rect -4886 150854 588810 150938
rect -4886 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 257546 150854
rect 257782 150618 257866 150854
rect 258102 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 588810 150854
rect -4886 150586 588810 150618
rect -2966 147454 586890 147486
rect -2966 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 69808 147454
rect 70044 147218 163512 147454
rect 163748 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 219617 147454
rect 219853 147218 222881 147454
rect 223117 147218 226145 147454
rect 226381 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 270617 147454
rect 270853 147218 273881 147454
rect 274117 147218 277145 147454
rect 277381 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 586890 147454
rect -2966 147134 586890 147218
rect -2966 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 69808 147134
rect 70044 146898 163512 147134
rect 163748 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 219617 147134
rect 219853 146898 222881 147134
rect 223117 146898 226145 147134
rect 226381 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 270617 147134
rect 270853 146898 273881 147134
rect 274117 146898 277145 147134
rect 277381 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 586890 147134
rect -2966 146866 586890 146898
rect -8726 140614 592650 140646
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 174986 140614
rect 175222 140378 175306 140614
rect 175542 140378 210986 140614
rect 211222 140378 211306 140614
rect 211542 140378 246986 140614
rect 247222 140378 247306 140614
rect 247542 140378 282986 140614
rect 283222 140378 283306 140614
rect 283542 140378 318986 140614
rect 319222 140378 319306 140614
rect 319542 140378 354986 140614
rect 355222 140378 355306 140614
rect 355542 140378 390986 140614
rect 391222 140378 391306 140614
rect 391542 140378 462986 140614
rect 463222 140378 463306 140614
rect 463542 140378 498986 140614
rect 499222 140378 499306 140614
rect 499542 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect -8726 140294 592650 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 174986 140294
rect 175222 140058 175306 140294
rect 175542 140058 210986 140294
rect 211222 140058 211306 140294
rect 211542 140058 246986 140294
rect 247222 140058 247306 140294
rect 247542 140058 282986 140294
rect 283222 140058 283306 140294
rect 283542 140058 318986 140294
rect 319222 140058 319306 140294
rect 319542 140058 354986 140294
rect 355222 140058 355306 140294
rect 355542 140058 390986 140294
rect 391222 140058 391306 140294
rect 391542 140058 462986 140294
rect 463222 140058 463306 140294
rect 463542 140058 498986 140294
rect 499222 140058 499306 140294
rect 499542 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect -8726 140026 592650 140058
rect -6806 136894 590730 136926
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 63266 136894
rect 63502 136658 63586 136894
rect 63822 136658 171266 136894
rect 171502 136658 171586 136894
rect 171822 136658 207266 136894
rect 207502 136658 207586 136894
rect 207822 136658 243266 136894
rect 243502 136658 243586 136894
rect 243822 136658 315266 136894
rect 315502 136658 315586 136894
rect 315822 136658 351266 136894
rect 351502 136658 351586 136894
rect 351822 136658 387266 136894
rect 387502 136658 387586 136894
rect 387822 136658 459266 136894
rect 459502 136658 459586 136894
rect 459822 136658 495266 136894
rect 495502 136658 495586 136894
rect 495822 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect -6806 136574 590730 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 63266 136574
rect 63502 136338 63586 136574
rect 63822 136338 171266 136574
rect 171502 136338 171586 136574
rect 171822 136338 207266 136574
rect 207502 136338 207586 136574
rect 207822 136338 243266 136574
rect 243502 136338 243586 136574
rect 243822 136338 315266 136574
rect 315502 136338 315586 136574
rect 315822 136338 351266 136574
rect 351502 136338 351586 136574
rect 351822 136338 387266 136574
rect 387502 136338 387586 136574
rect 387822 136338 459266 136574
rect 459502 136338 459586 136574
rect 459822 136338 495266 136574
rect 495502 136338 495586 136574
rect 495822 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect -6806 136306 590730 136338
rect -4886 133174 588810 133206
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 59546 133174
rect 59782 132938 59866 133174
rect 60102 132938 167546 133174
rect 167782 132938 167866 133174
rect 168102 132938 203546 133174
rect 203782 132938 203866 133174
rect 204102 132938 239546 133174
rect 239782 132938 239866 133174
rect 240102 132938 311546 133174
rect 311782 132938 311866 133174
rect 312102 132938 347546 133174
rect 347782 132938 347866 133174
rect 348102 132938 383546 133174
rect 383782 132938 383866 133174
rect 384102 132938 455546 133174
rect 455782 132938 455866 133174
rect 456102 132938 491546 133174
rect 491782 132938 491866 133174
rect 492102 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect -4886 132854 588810 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 59546 132854
rect 59782 132618 59866 132854
rect 60102 132618 167546 132854
rect 167782 132618 167866 132854
rect 168102 132618 203546 132854
rect 203782 132618 203866 132854
rect 204102 132618 239546 132854
rect 239782 132618 239866 132854
rect 240102 132618 311546 132854
rect 311782 132618 311866 132854
rect 312102 132618 347546 132854
rect 347782 132618 347866 132854
rect 348102 132618 383546 132854
rect 383782 132618 383866 132854
rect 384102 132618 455546 132854
rect 455782 132618 455866 132854
rect 456102 132618 491546 132854
rect 491782 132618 491866 132854
rect 492102 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect -4886 132586 588810 132618
rect -2966 129454 586890 129486
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 69128 129454
rect 69364 129218 164192 129454
rect 164428 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 221249 129454
rect 221485 129218 224513 129454
rect 224749 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 272249 129454
rect 272485 129218 275513 129454
rect 275749 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 402586 129454
rect 402822 129218 405786 129454
rect 406022 129218 408986 129454
rect 409222 129218 412186 129454
rect 412422 129218 415386 129454
rect 415622 129218 418586 129454
rect 418822 129218 421786 129454
rect 422022 129218 424986 129454
rect 425222 129218 428186 129454
rect 428422 129218 431386 129454
rect 431622 129218 434586 129454
rect 434822 129218 437786 129454
rect 438022 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect -2966 129134 586890 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 69128 129134
rect 69364 128898 164192 129134
rect 164428 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 221249 129134
rect 221485 128898 224513 129134
rect 224749 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 272249 129134
rect 272485 128898 275513 129134
rect 275749 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 402586 129134
rect 402822 128898 405786 129134
rect 406022 128898 408986 129134
rect 409222 128898 412186 129134
rect 412422 128898 415386 129134
rect 415622 128898 418586 129134
rect 418822 128898 421786 129134
rect 422022 128898 424986 129134
rect 425222 128898 428186 129134
rect 428422 128898 431386 129134
rect 431622 128898 434586 129134
rect 434822 128898 437786 129134
rect 438022 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect -2966 128866 586890 128898
rect -8726 122614 592650 122646
rect -8726 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 192986 122614
rect 193222 122378 193306 122614
rect 193542 122378 264986 122614
rect 265222 122378 265306 122614
rect 265542 122378 300986 122614
rect 301222 122378 301306 122614
rect 301542 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 444986 122614
rect 445222 122378 445306 122614
rect 445542 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 592650 122614
rect -8726 122294 592650 122378
rect -8726 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 192986 122294
rect 193222 122058 193306 122294
rect 193542 122058 264986 122294
rect 265222 122058 265306 122294
rect 265542 122058 300986 122294
rect 301222 122058 301306 122294
rect 301542 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 444986 122294
rect 445222 122058 445306 122294
rect 445542 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 592650 122294
rect -8726 122026 592650 122058
rect -6806 118894 590730 118926
rect -6806 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 189266 118894
rect 189502 118658 189586 118894
rect 189822 118658 261266 118894
rect 261502 118658 261586 118894
rect 261822 118658 297266 118894
rect 297502 118658 297586 118894
rect 297822 118658 333266 118894
rect 333502 118658 333586 118894
rect 333822 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 590730 118894
rect -6806 118574 590730 118658
rect -6806 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 189266 118574
rect 189502 118338 189586 118574
rect 189822 118338 261266 118574
rect 261502 118338 261586 118574
rect 261822 118338 297266 118574
rect 297502 118338 297586 118574
rect 297822 118338 333266 118574
rect 333502 118338 333586 118574
rect 333822 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 590730 118574
rect -6806 118306 590730 118338
rect -4886 115174 588810 115206
rect -4886 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 185546 115174
rect 185782 114938 185866 115174
rect 186102 114938 257546 115174
rect 257782 114938 257866 115174
rect 258102 114938 293546 115174
rect 293782 114938 293866 115174
rect 294102 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 588810 115174
rect -4886 114854 588810 114938
rect -4886 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 185546 114854
rect 185782 114618 185866 114854
rect 186102 114618 257546 114854
rect 257782 114618 257866 114854
rect 258102 114618 293546 114854
rect 293782 114618 293866 114854
rect 294102 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 588810 114854
rect -4886 114586 588810 114618
rect -2966 111454 586890 111486
rect -2966 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 69808 111454
rect 70044 111218 163512 111454
rect 163748 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 219617 111454
rect 219853 111218 222881 111454
rect 223117 111218 226145 111454
rect 226381 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 270617 111454
rect 270853 111218 273881 111454
rect 274117 111218 277145 111454
rect 277381 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 404186 111454
rect 404422 111218 407386 111454
rect 407622 111218 410586 111454
rect 410822 111218 413786 111454
rect 414022 111218 416986 111454
rect 417222 111218 420186 111454
rect 420422 111218 423386 111454
rect 423622 111218 426586 111454
rect 426822 111218 429786 111454
rect 430022 111218 432986 111454
rect 433222 111218 436186 111454
rect 436422 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 586890 111454
rect -2966 111134 586890 111218
rect -2966 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 69808 111134
rect 70044 110898 163512 111134
rect 163748 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 219617 111134
rect 219853 110898 222881 111134
rect 223117 110898 226145 111134
rect 226381 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 270617 111134
rect 270853 110898 273881 111134
rect 274117 110898 277145 111134
rect 277381 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 404186 111134
rect 404422 110898 407386 111134
rect 407622 110898 410586 111134
rect 410822 110898 413786 111134
rect 414022 110898 416986 111134
rect 417222 110898 420186 111134
rect 420422 110898 423386 111134
rect 423622 110898 426586 111134
rect 426822 110898 429786 111134
rect 430022 110898 432986 111134
rect 433222 110898 436186 111134
rect 436422 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 586890 111134
rect -2966 110866 586890 110898
rect -8726 104614 592650 104646
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 174986 104614
rect 175222 104378 175306 104614
rect 175542 104378 210986 104614
rect 211222 104378 211306 104614
rect 211542 104378 246986 104614
rect 247222 104378 247306 104614
rect 247542 104378 282986 104614
rect 283222 104378 283306 104614
rect 283542 104378 318986 104614
rect 319222 104378 319306 104614
rect 319542 104378 354986 104614
rect 355222 104378 355306 104614
rect 355542 104378 390986 104614
rect 391222 104378 391306 104614
rect 391542 104378 462986 104614
rect 463222 104378 463306 104614
rect 463542 104378 498986 104614
rect 499222 104378 499306 104614
rect 499542 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect -8726 104294 592650 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 174986 104294
rect 175222 104058 175306 104294
rect 175542 104058 210986 104294
rect 211222 104058 211306 104294
rect 211542 104058 246986 104294
rect 247222 104058 247306 104294
rect 247542 104058 282986 104294
rect 283222 104058 283306 104294
rect 283542 104058 318986 104294
rect 319222 104058 319306 104294
rect 319542 104058 354986 104294
rect 355222 104058 355306 104294
rect 355542 104058 390986 104294
rect 391222 104058 391306 104294
rect 391542 104058 462986 104294
rect 463222 104058 463306 104294
rect 463542 104058 498986 104294
rect 499222 104058 499306 104294
rect 499542 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect -8726 104026 592650 104058
rect -6806 100894 590730 100926
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 63266 100894
rect 63502 100658 63586 100894
rect 63822 100658 171266 100894
rect 171502 100658 171586 100894
rect 171822 100658 207266 100894
rect 207502 100658 207586 100894
rect 207822 100658 243266 100894
rect 243502 100658 243586 100894
rect 243822 100658 315266 100894
rect 315502 100658 315586 100894
rect 315822 100658 351266 100894
rect 351502 100658 351586 100894
rect 351822 100658 387266 100894
rect 387502 100658 387586 100894
rect 387822 100658 459266 100894
rect 459502 100658 459586 100894
rect 459822 100658 495266 100894
rect 495502 100658 495586 100894
rect 495822 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect -6806 100574 590730 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 63266 100574
rect 63502 100338 63586 100574
rect 63822 100338 171266 100574
rect 171502 100338 171586 100574
rect 171822 100338 207266 100574
rect 207502 100338 207586 100574
rect 207822 100338 243266 100574
rect 243502 100338 243586 100574
rect 243822 100338 315266 100574
rect 315502 100338 315586 100574
rect 315822 100338 351266 100574
rect 351502 100338 351586 100574
rect 351822 100338 387266 100574
rect 387502 100338 387586 100574
rect 387822 100338 459266 100574
rect 459502 100338 459586 100574
rect 459822 100338 495266 100574
rect 495502 100338 495586 100574
rect 495822 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect -6806 100306 590730 100338
rect -4886 97174 588810 97206
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 59546 97174
rect 59782 96938 59866 97174
rect 60102 96938 167546 97174
rect 167782 96938 167866 97174
rect 168102 96938 203546 97174
rect 203782 96938 203866 97174
rect 204102 96938 239546 97174
rect 239782 96938 239866 97174
rect 240102 96938 311546 97174
rect 311782 96938 311866 97174
rect 312102 96938 347546 97174
rect 347782 96938 347866 97174
rect 348102 96938 383546 97174
rect 383782 96938 383866 97174
rect 384102 96938 419546 97174
rect 419782 96938 419866 97174
rect 420102 96938 455546 97174
rect 455782 96938 455866 97174
rect 456102 96938 491546 97174
rect 491782 96938 491866 97174
rect 492102 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect -4886 96854 588810 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 59546 96854
rect 59782 96618 59866 96854
rect 60102 96618 167546 96854
rect 167782 96618 167866 96854
rect 168102 96618 203546 96854
rect 203782 96618 203866 96854
rect 204102 96618 239546 96854
rect 239782 96618 239866 96854
rect 240102 96618 311546 96854
rect 311782 96618 311866 96854
rect 312102 96618 347546 96854
rect 347782 96618 347866 96854
rect 348102 96618 383546 96854
rect 383782 96618 383866 96854
rect 384102 96618 419546 96854
rect 419782 96618 419866 96854
rect 420102 96618 455546 96854
rect 455782 96618 455866 96854
rect 456102 96618 491546 96854
rect 491782 96618 491866 96854
rect 492102 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect -4886 96586 588810 96618
rect -2966 93454 586890 93486
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect -2966 93134 586890 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect -2966 92866 586890 92898
rect -8726 86614 592650 86646
rect -8726 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 84986 86614
rect 85222 86378 85306 86614
rect 85542 86378 120986 86614
rect 121222 86378 121306 86614
rect 121542 86378 156986 86614
rect 157222 86378 157306 86614
rect 157542 86378 192986 86614
rect 193222 86378 193306 86614
rect 193542 86378 228986 86614
rect 229222 86378 229306 86614
rect 229542 86378 264986 86614
rect 265222 86378 265306 86614
rect 265542 86378 300986 86614
rect 301222 86378 301306 86614
rect 301542 86378 336986 86614
rect 337222 86378 337306 86614
rect 337542 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 592650 86614
rect -8726 86294 592650 86378
rect -8726 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 84986 86294
rect 85222 86058 85306 86294
rect 85542 86058 120986 86294
rect 121222 86058 121306 86294
rect 121542 86058 156986 86294
rect 157222 86058 157306 86294
rect 157542 86058 192986 86294
rect 193222 86058 193306 86294
rect 193542 86058 228986 86294
rect 229222 86058 229306 86294
rect 229542 86058 264986 86294
rect 265222 86058 265306 86294
rect 265542 86058 300986 86294
rect 301222 86058 301306 86294
rect 301542 86058 336986 86294
rect 337222 86058 337306 86294
rect 337542 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 592650 86294
rect -8726 86026 592650 86058
rect -6806 82894 590730 82926
rect -6806 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 81266 82894
rect 81502 82658 81586 82894
rect 81822 82658 117266 82894
rect 117502 82658 117586 82894
rect 117822 82658 153266 82894
rect 153502 82658 153586 82894
rect 153822 82658 189266 82894
rect 189502 82658 189586 82894
rect 189822 82658 225266 82894
rect 225502 82658 225586 82894
rect 225822 82658 261266 82894
rect 261502 82658 261586 82894
rect 261822 82658 297266 82894
rect 297502 82658 297586 82894
rect 297822 82658 333266 82894
rect 333502 82658 333586 82894
rect 333822 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 590730 82894
rect -6806 82574 590730 82658
rect -6806 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 81266 82574
rect 81502 82338 81586 82574
rect 81822 82338 117266 82574
rect 117502 82338 117586 82574
rect 117822 82338 153266 82574
rect 153502 82338 153586 82574
rect 153822 82338 189266 82574
rect 189502 82338 189586 82574
rect 189822 82338 225266 82574
rect 225502 82338 225586 82574
rect 225822 82338 261266 82574
rect 261502 82338 261586 82574
rect 261822 82338 297266 82574
rect 297502 82338 297586 82574
rect 297822 82338 333266 82574
rect 333502 82338 333586 82574
rect 333822 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 590730 82574
rect -6806 82306 590730 82338
rect -4886 79174 588810 79206
rect -4886 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 77546 79174
rect 77782 78938 77866 79174
rect 78102 78938 113546 79174
rect 113782 78938 113866 79174
rect 114102 78938 149546 79174
rect 149782 78938 149866 79174
rect 150102 78938 185546 79174
rect 185782 78938 185866 79174
rect 186102 78938 221546 79174
rect 221782 78938 221866 79174
rect 222102 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 588810 79174
rect -4886 78854 588810 78938
rect -4886 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 77546 78854
rect 77782 78618 77866 78854
rect 78102 78618 113546 78854
rect 113782 78618 113866 78854
rect 114102 78618 149546 78854
rect 149782 78618 149866 78854
rect 150102 78618 185546 78854
rect 185782 78618 185866 78854
rect 186102 78618 221546 78854
rect 221782 78618 221866 78854
rect 222102 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 588810 78854
rect -4886 78586 588810 78618
rect -2966 75454 586890 75486
rect -2966 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 586890 75454
rect -2966 75134 586890 75218
rect -2966 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 586890 75134
rect -2966 74866 586890 74898
rect -8726 68614 592650 68646
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 66986 68614
rect 67222 68378 67306 68614
rect 67542 68378 102986 68614
rect 103222 68378 103306 68614
rect 103542 68378 138986 68614
rect 139222 68378 139306 68614
rect 139542 68378 174986 68614
rect 175222 68378 175306 68614
rect 175542 68378 210986 68614
rect 211222 68378 211306 68614
rect 211542 68378 246986 68614
rect 247222 68378 247306 68614
rect 247542 68378 282986 68614
rect 283222 68378 283306 68614
rect 283542 68378 318986 68614
rect 319222 68378 319306 68614
rect 319542 68378 354986 68614
rect 355222 68378 355306 68614
rect 355542 68378 390986 68614
rect 391222 68378 391306 68614
rect 391542 68378 426986 68614
rect 427222 68378 427306 68614
rect 427542 68378 462986 68614
rect 463222 68378 463306 68614
rect 463542 68378 498986 68614
rect 499222 68378 499306 68614
rect 499542 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect -8726 68294 592650 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 66986 68294
rect 67222 68058 67306 68294
rect 67542 68058 102986 68294
rect 103222 68058 103306 68294
rect 103542 68058 138986 68294
rect 139222 68058 139306 68294
rect 139542 68058 174986 68294
rect 175222 68058 175306 68294
rect 175542 68058 210986 68294
rect 211222 68058 211306 68294
rect 211542 68058 246986 68294
rect 247222 68058 247306 68294
rect 247542 68058 282986 68294
rect 283222 68058 283306 68294
rect 283542 68058 318986 68294
rect 319222 68058 319306 68294
rect 319542 68058 354986 68294
rect 355222 68058 355306 68294
rect 355542 68058 390986 68294
rect 391222 68058 391306 68294
rect 391542 68058 426986 68294
rect 427222 68058 427306 68294
rect 427542 68058 462986 68294
rect 463222 68058 463306 68294
rect 463542 68058 498986 68294
rect 499222 68058 499306 68294
rect 499542 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect -8726 68026 592650 68058
rect -6806 64894 590730 64926
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 63266 64894
rect 63502 64658 63586 64894
rect 63822 64658 99266 64894
rect 99502 64658 99586 64894
rect 99822 64658 135266 64894
rect 135502 64658 135586 64894
rect 135822 64658 171266 64894
rect 171502 64658 171586 64894
rect 171822 64658 207266 64894
rect 207502 64658 207586 64894
rect 207822 64658 243266 64894
rect 243502 64658 243586 64894
rect 243822 64658 279266 64894
rect 279502 64658 279586 64894
rect 279822 64658 315266 64894
rect 315502 64658 315586 64894
rect 315822 64658 351266 64894
rect 351502 64658 351586 64894
rect 351822 64658 387266 64894
rect 387502 64658 387586 64894
rect 387822 64658 423266 64894
rect 423502 64658 423586 64894
rect 423822 64658 459266 64894
rect 459502 64658 459586 64894
rect 459822 64658 495266 64894
rect 495502 64658 495586 64894
rect 495822 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect -6806 64574 590730 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 63266 64574
rect 63502 64338 63586 64574
rect 63822 64338 99266 64574
rect 99502 64338 99586 64574
rect 99822 64338 135266 64574
rect 135502 64338 135586 64574
rect 135822 64338 171266 64574
rect 171502 64338 171586 64574
rect 171822 64338 207266 64574
rect 207502 64338 207586 64574
rect 207822 64338 243266 64574
rect 243502 64338 243586 64574
rect 243822 64338 279266 64574
rect 279502 64338 279586 64574
rect 279822 64338 315266 64574
rect 315502 64338 315586 64574
rect 315822 64338 351266 64574
rect 351502 64338 351586 64574
rect 351822 64338 387266 64574
rect 387502 64338 387586 64574
rect 387822 64338 423266 64574
rect 423502 64338 423586 64574
rect 423822 64338 459266 64574
rect 459502 64338 459586 64574
rect 459822 64338 495266 64574
rect 495502 64338 495586 64574
rect 495822 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect -6806 64306 590730 64338
rect -4886 61174 588810 61206
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 59546 61174
rect 59782 60938 59866 61174
rect 60102 60938 95546 61174
rect 95782 60938 95866 61174
rect 96102 60938 131546 61174
rect 131782 60938 131866 61174
rect 132102 60938 167546 61174
rect 167782 60938 167866 61174
rect 168102 60938 203546 61174
rect 203782 60938 203866 61174
rect 204102 60938 239546 61174
rect 239782 60938 239866 61174
rect 240102 60938 275546 61174
rect 275782 60938 275866 61174
rect 276102 60938 311546 61174
rect 311782 60938 311866 61174
rect 312102 60938 347546 61174
rect 347782 60938 347866 61174
rect 348102 60938 383546 61174
rect 383782 60938 383866 61174
rect 384102 60938 419546 61174
rect 419782 60938 419866 61174
rect 420102 60938 455546 61174
rect 455782 60938 455866 61174
rect 456102 60938 491546 61174
rect 491782 60938 491866 61174
rect 492102 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect -4886 60854 588810 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 59546 60854
rect 59782 60618 59866 60854
rect 60102 60618 95546 60854
rect 95782 60618 95866 60854
rect 96102 60618 131546 60854
rect 131782 60618 131866 60854
rect 132102 60618 167546 60854
rect 167782 60618 167866 60854
rect 168102 60618 203546 60854
rect 203782 60618 203866 60854
rect 204102 60618 239546 60854
rect 239782 60618 239866 60854
rect 240102 60618 275546 60854
rect 275782 60618 275866 60854
rect 276102 60618 311546 60854
rect 311782 60618 311866 60854
rect 312102 60618 347546 60854
rect 347782 60618 347866 60854
rect 348102 60618 383546 60854
rect 383782 60618 383866 60854
rect 384102 60618 419546 60854
rect 419782 60618 419866 60854
rect 420102 60618 455546 60854
rect 455782 60618 455866 60854
rect 456102 60618 491546 60854
rect 491782 60618 491866 60854
rect 492102 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect -4886 60586 588810 60618
rect -2966 57454 586890 57486
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect -2966 57134 586890 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect -2966 56866 586890 56898
rect -8726 50614 592650 50646
rect -8726 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 592650 50614
rect -8726 50294 592650 50378
rect -8726 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 592650 50294
rect -8726 50026 592650 50058
rect -6806 46894 590730 46926
rect -6806 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 590730 46894
rect -6806 46574 590730 46658
rect -6806 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 590730 46574
rect -6806 46306 590730 46338
rect -4886 43174 588810 43206
rect -4886 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 588810 43174
rect -4886 42854 588810 42938
rect -4886 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 588810 42854
rect -4886 42586 588810 42618
rect -2966 39454 586890 39486
rect -2966 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 586890 39454
rect -2966 39134 586890 39218
rect -2966 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 586890 39134
rect -2966 38866 586890 38898
rect -8726 32614 592650 32646
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect -8726 32294 592650 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect -8726 32026 592650 32058
rect -6806 28894 590730 28926
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect -6806 28574 590730 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect -6806 28306 590730 28338
rect -4886 25174 588810 25206
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect -4886 24854 588810 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect -4886 24586 588810 24618
rect -2966 21454 586890 21486
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect -2966 21134 586890 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect -2966 20866 586890 20898
rect -8726 14614 592650 14646
rect -8726 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 592650 14614
rect -8726 14294 592650 14378
rect -8726 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 592650 14294
rect -8726 14026 592650 14058
rect -6806 10894 590730 10926
rect -6806 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 590730 10894
rect -6806 10574 590730 10658
rect -6806 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 590730 10574
rect -6806 10306 590730 10338
rect -4886 7174 588810 7206
rect -4886 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 588810 7174
rect -4886 6854 588810 6938
rect -4886 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 588810 6854
rect -4886 6586 588810 6618
rect -2966 3454 586890 3486
rect -2966 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 586890 3454
rect -2966 3134 586890 3218
rect -2966 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 586890 3134
rect -2966 2866 586890 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use wrapped_spell  wrapped_spell_1
timestamp 1640693535
transform 1 0 68770 0 1 241592
box 0 0 88000 88000
use wrapped_skullfet  wrapped_skullfet_5
timestamp 1640693535
transform 1 0 400000 0 1 100000
box -10 0 40000 40000
use wrapped_silife  wrapped_silife_4
timestamp 1640693535
transform 1 0 200000 0 1 377600
box -10 0 156249 158393
use wrapped_ppm_decoder  wrapped_ppm_decoder_3
timestamp 1640693535
transform 1 0 68770 0 1 539166
box -10 0 20000 50000
use wrapped_ppm_coder  wrapped_ppm_coder_2
timestamp 1640693535
transform 1 0 68770 0 1 390356
box -10 0 51907 54051
use wrapped_function_generator  wrapped_function_generator_0
timestamp 1640693535
transform 1 0 200200 0 1 240182
box 0 0 44000 44000
use wb_openram_wrapper  wb_openram_wrapper
timestamp 1640693535
transform 1 0 217000 0 1 96000
box 0 144 12000 79688
use wb_bridge_2way  wb_bridge_2way
timestamp 1640693535
transform 1 0 268000 0 1 96000
box 0 0 12000 79688
use sky130_sram_1kbyte_1rw1r_32x256_8  openram_1kB
timestamp 1640693535
transform 1 0 68800 0 1 95100
box 0 0 95956 79500
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 30 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 31 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 32 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 33 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 37 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 38 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 39 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 41 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 42 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 44 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 45 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 46 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 47 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 48 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 49 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 50 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 51 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 52 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 53 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 54 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 55 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 56 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 57 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 58 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 59 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 61 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 62 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 63 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 64 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 65 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 66 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 67 nsew signal tristate
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 68 nsew signal tristate
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 69 nsew signal tristate
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 70 nsew signal tristate
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 71 nsew signal tristate
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 72 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 73 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 74 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 75 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 76 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 77 nsew signal tristate
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 78 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 79 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 80 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 81 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 82 nsew signal tristate
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 83 nsew signal tristate
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 84 nsew signal tristate
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 85 nsew signal tristate
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 86 nsew signal tristate
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 87 nsew signal tristate
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 88 nsew signal tristate
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 89 nsew signal tristate
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 90 nsew signal tristate
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 91 nsew signal tristate
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 92 nsew signal tristate
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 93 nsew signal tristate
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 94 nsew signal tristate
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 95 nsew signal tristate
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 96 nsew signal tristate
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 97 nsew signal tristate
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 98 nsew signal tristate
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 99 nsew signal tristate
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 100 nsew signal tristate
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 101 nsew signal tristate
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 102 nsew signal tristate
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 103 nsew signal tristate
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 104 nsew signal tristate
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 105 nsew signal tristate
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 106 nsew signal tristate
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 107 nsew signal tristate
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 108 nsew signal tristate
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 109 nsew signal tristate
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 110 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 111 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 112 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 113 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 114 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 115 nsew signal tristate
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 116 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 117 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 118 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 119 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 120 nsew signal tristate
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 121 nsew signal tristate
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 122 nsew signal tristate
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 123 nsew signal tristate
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 124 nsew signal tristate
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 125 nsew signal tristate
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 126 nsew signal tristate
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 127 nsew signal tristate
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 128 nsew signal tristate
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 129 nsew signal tristate
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 130 nsew signal tristate
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 131 nsew signal tristate
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 132 nsew signal tristate
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 133 nsew signal tristate
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 134 nsew signal tristate
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 135 nsew signal tristate
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 136 nsew signal tristate
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 137 nsew signal tristate
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 138 nsew signal tristate
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 139 nsew signal tristate
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 140 nsew signal tristate
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 141 nsew signal tristate
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 142 nsew signal tristate
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 271 nsew signal tristate
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 274 nsew signal tristate
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 276 nsew signal tristate
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 278 nsew signal tristate
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 279 nsew signal tristate
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 282 nsew signal tristate
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 283 nsew signal tristate
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 284 nsew signal tristate
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 287 nsew signal tristate
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 290 nsew signal tristate
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 292 nsew signal tristate
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 293 nsew signal tristate
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 295 nsew signal tristate
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 296 nsew signal tristate
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 304 nsew signal tristate
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 305 nsew signal tristate
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 306 nsew signal tristate
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 307 nsew signal tristate
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 311 nsew signal tristate
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 312 nsew signal tristate
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 313 nsew signal tristate
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 316 nsew signal tristate
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 322 nsew signal tristate
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 323 nsew signal tristate
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 326 nsew signal tristate
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 330 nsew signal tristate
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 332 nsew signal tristate
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 333 nsew signal tristate
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 335 nsew signal tristate
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 336 nsew signal tristate
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 343 nsew signal tristate
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 345 nsew signal tristate
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 347 nsew signal tristate
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 352 nsew signal tristate
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 356 nsew signal tristate
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 358 nsew signal tristate
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 361 nsew signal tristate
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 362 nsew signal tristate
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 374 nsew signal tristate
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 376 nsew signal tristate
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 378 nsew signal tristate
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 379 nsew signal tristate
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 380 nsew signal tristate
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 383 nsew signal tristate
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 384 nsew signal tristate
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 386 nsew signal tristate
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 387 nsew signal tristate
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 396 nsew signal tristate
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 397 nsew signal tristate
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 404 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 407 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 410 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 411 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 414 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 416 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 421 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 422 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 424 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 428 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 429 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 430 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 432 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 433 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 435 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 436 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 438 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 441 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 442 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 443 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 445 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 449 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 451 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 452 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 454 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 455 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 457 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 458 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 461 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 462 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 463 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 464 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 466 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 468 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 472 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 473 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 476 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 478 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 479 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 482 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 483 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 488 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 493 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 494 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 495 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 496 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 497 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 498 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 499 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 500 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 504 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 505 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 506 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 507 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 508 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 509 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 510 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 512 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 515 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 518 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 520 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 522 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 526 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 527 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 528 nsew signal tristate
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 529 nsew signal tristate
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 530 nsew signal tristate
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 531 nsew power input
rlabel metal5 s -2966 2866 586890 3486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 38866 586890 39486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 74866 586890 75486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 110866 586890 111486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 146866 586890 147486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 182866 586890 183486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 218866 586890 219486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 254866 586890 255486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 290866 586890 291486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 326866 586890 327486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 362866 586890 363486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 398866 586890 399486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 434866 586890 435486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 470866 586890 471486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 506866 586890 507486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 542866 586890 543486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 578866 586890 579486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 614866 586890 615486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 650866 586890 651486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 686866 586890 687486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 -1894 74414 93100 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 -1894 110414 93100 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 -1894 146414 93100 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 -1894 218414 94000 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 -1894 398414 98000 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 -1894 434414 98000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 178000 218414 238182 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 176600 74414 239592 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 176600 110414 239592 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 176600 146414 239592 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 286182 218414 375600 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 -1894 254414 375600 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 -1894 290414 375600 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 -1894 326414 375600 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 331592 74414 388356 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 331592 110414 388356 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 446407 74414 537166 6 vccd1
port 531 nsew power input
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 531 nsew power input
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 1794 -1894 2414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 -1894 38414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 591166 74414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 446407 110414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 331592 146414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 -1894 182414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 537993 218414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 537993 254414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 537993 290414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 537993 326414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 -1894 362414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 142000 398414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 142000 434414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 -1894 470414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 -1894 506414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 -1894 542414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 577794 -1894 578414 705830 6 vccd1
port 531 nsew power input
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 532 nsew power input
rlabel metal5 s -4886 6586 588810 7206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 42586 588810 43206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 78586 588810 79206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 114586 588810 115206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 150586 588810 151206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 186586 588810 187206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 222586 588810 223206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 258586 588810 259206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 294586 588810 295206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 330586 588810 331206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 366586 588810 367206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 402586 588810 403206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 438586 588810 439206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 474586 588810 475206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 510586 588810 511206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 546586 588810 547206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 582586 588810 583206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 618586 588810 619206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 654586 588810 655206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 690586 588810 691206 6 vccd2
port 532 nsew power input
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 -3814 78134 93100 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 -3814 114134 93100 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 -3814 150134 93100 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 -3814 222134 94000 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 -3814 402134 98000 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 -3814 438134 98000 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 178000 222134 238182 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 176600 78134 239592 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 176600 114134 239592 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 176600 150134 239592 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 286182 222134 375600 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 -3814 258134 375600 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 -3814 294134 375600 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 -3814 330134 375600 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 331592 78134 388356 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 331592 114134 388356 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 446407 78134 537166 6 vccd2
port 532 nsew power input
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 532 nsew power input
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 5514 -3814 6134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 41514 -3814 42134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 591166 78134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 446407 114134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 331592 150134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 -3814 186134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 537993 222134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 537993 258134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 537993 294134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 537993 330134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 -3814 366134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 142000 402134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 142000 438134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 -3814 474134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 -3814 510134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 545514 -3814 546134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 581514 -3814 582134 707750 6 vccd2
port 532 nsew power input
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 533 nsew power input
rlabel metal5 s -6806 10306 590730 10926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 46306 590730 46926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 82306 590730 82926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 118306 590730 118926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 154306 590730 154926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 190306 590730 190926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 226306 590730 226926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 262306 590730 262926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 298306 590730 298926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 334306 590730 334926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 370306 590730 370926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 406306 590730 406926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 442306 590730 442926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 478306 590730 478926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 514306 590730 514926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 550306 590730 550926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 586306 590730 586926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 622306 590730 622926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 658306 590730 658926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 694306 590730 694926 6 vdda1
port 533 nsew power input
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 -5734 81854 93100 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 -5734 117854 93100 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 -5734 153854 93100 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 -5734 225854 94000 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 -5734 405854 98000 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 -5734 441854 98000 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 178000 225854 238182 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 176600 81854 239592 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 176600 117854 239592 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 176600 153854 239592 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 286182 225854 375600 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 -5734 261854 375600 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 -5734 297854 375600 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 -5734 333854 375600 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 331592 81854 388356 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 331592 117854 388356 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 446407 81854 537166 6 vdda1
port 533 nsew power input
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 533 nsew power input
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 9234 -5734 9854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 45234 -5734 45854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 591166 81854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 446407 117854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 331592 153854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 -5734 189854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 537993 225854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 537993 261854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 537993 297854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 537993 333854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 -5734 369854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 142000 405854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 142000 441854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 -5734 477854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 -5734 513854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 549234 -5734 549854 709670 6 vdda1
port 533 nsew power input
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 534 nsew power input
rlabel metal5 s -8726 14026 592650 14646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 50026 592650 50646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 86026 592650 86646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 122026 592650 122646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 158026 592650 158646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 194026 592650 194646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 230026 592650 230646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 266026 592650 266646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 302026 592650 302646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 338026 592650 338646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 374026 592650 374646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 410026 592650 410646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 446026 592650 446646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 482026 592650 482646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 518026 592650 518646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 554026 592650 554646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 590026 592650 590646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 626026 592650 626646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 662026 592650 662646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 698026 592650 698646 6 vdda2
port 534 nsew power input
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 -7654 85574 93100 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 -7654 121574 93100 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 -7654 157574 93100 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 -7654 229574 94000 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 -7654 409574 98000 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 178000 229574 238182 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 176600 85574 239592 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 176600 121574 239592 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 176600 157574 239592 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 286182 229574 375600 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 -7654 265574 375600 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 -7654 301574 375600 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 -7654 337574 375600 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 331592 85574 388356 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 331592 121574 388356 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 446407 85574 537166 6 vdda2
port 534 nsew power input
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 534 nsew power input
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 12954 -7654 13574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 48954 -7654 49574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 591166 85574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 446407 121574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 331592 157574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 -7654 193574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 537993 229574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 537993 265574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 537993 301574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 537993 337574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 -7654 373574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 142000 409574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 -7654 445574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 -7654 481574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 -7654 517574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 552954 -7654 553574 711590 6 vdda2
port 534 nsew power input
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 28306 590730 28926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 64306 590730 64926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 100306 590730 100926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 136306 590730 136926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 172306 590730 172926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 208306 590730 208926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 244306 590730 244926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 280306 590730 280926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 316306 590730 316926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 352306 590730 352926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 388306 590730 388926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 424306 590730 424926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 460306 590730 460926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 496306 590730 496926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 532306 590730 532926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 568306 590730 568926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 604306 590730 604926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 640306 590730 640926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 676306 590730 676926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 -5734 99854 93100 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 -5734 135854 93100 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 -5734 279854 94000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 -5734 423854 98000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 -5734 207854 238182 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 -5734 243854 238182 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 176600 99854 239592 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 176600 135854 239592 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 286182 207854 375600 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 286182 243854 375600 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 178000 279854 375600 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 -5734 315854 375600 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 -5734 351854 375600 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 331592 99854 388356 6 vssa1
port 535 nsew ground input
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 535 nsew ground input
rlabel metal4 s 27234 -5734 27854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 -5734 63854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 446407 99854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 331592 135854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 -5734 171854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 537993 207854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 537993 243854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 537993 279854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 537993 315854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 537993 351854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 -5734 387854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 142000 423854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 -5734 459854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 -5734 495854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 -5734 531854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 567234 -5734 567854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 32026 592650 32646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 68026 592650 68646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 104026 592650 104646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 140026 592650 140646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 176026 592650 176646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 212026 592650 212646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 248026 592650 248646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 284026 592650 284646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 320026 592650 320646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 356026 592650 356646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 392026 592650 392646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 428026 592650 428646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 464026 592650 464646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 500026 592650 500646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 536026 592650 536646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 572026 592650 572646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 608026 592650 608646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 644026 592650 644646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 680026 592650 680646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 -7654 67574 93100 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 -7654 103574 93100 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 -7654 139574 93100 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 -7654 427574 98000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 -7654 211574 238182 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 176600 67574 239592 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 176600 103574 239592 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 176600 139574 239592 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 286182 211574 375600 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 -7654 247574 375600 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 -7654 283574 375600 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 -7654 319574 375600 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 -7654 355574 375600 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 331592 67574 388356 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 331592 103574 388356 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 446407 67574 537166 6 vssa2
port 536 nsew ground input
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 536 nsew ground input
rlabel metal4 s 30954 -7654 31574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 591166 67574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 446407 103574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 331592 139574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 -7654 175574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 537993 211574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 537993 247574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 537993 283574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 537993 319574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 537993 355574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 -7654 391574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 142000 427574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 -7654 463574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 -7654 499574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 -7654 535574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 570954 -7654 571574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 20866 586890 21486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 56866 586890 57486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 92866 586890 93486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 128866 586890 129486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 164866 586890 165486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 200866 586890 201486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 236866 586890 237486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 272866 586890 273486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 308866 586890 309486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 344866 586890 345486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 380866 586890 381486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 416866 586890 417486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 452866 586890 453486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 488866 586890 489486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 524866 586890 525486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 560866 586890 561486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 596866 586890 597486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 632866 586890 633486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 668866 586890 669486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 -1894 92414 93100 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 -1894 128414 93100 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 -1894 164414 93100 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 -1894 272414 94000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 -1894 416414 98000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 -1894 200414 238182 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 -1894 236414 238182 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 176600 92414 239592 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 176600 128414 239592 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 286182 200414 375600 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 286182 236414 375600 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 178000 272414 375600 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 -1894 308414 375600 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 -1894 344414 375600 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 331592 92414 388356 6 vssd1
port 537 nsew ground input
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 537 nsew ground input
rlabel metal4 s 19794 -1894 20414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 -1894 56414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 446407 92414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 331592 128414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 176600 164414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 537993 200414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 537993 236414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 537993 272414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 537993 308414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 537993 344414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 -1894 380414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 142000 416414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 -1894 452414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 -1894 488414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 523794 -1894 524414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 559794 -1894 560414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 24586 588810 25206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 60586 588810 61206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 96586 588810 97206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 132586 588810 133206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 168586 588810 169206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 204586 588810 205206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 240586 588810 241206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 276586 588810 277206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 312586 588810 313206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 348586 588810 349206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 384586 588810 385206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 420586 588810 421206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 456586 588810 457206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 492586 588810 493206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 528586 588810 529206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 564586 588810 565206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 600586 588810 601206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 636586 588810 637206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 672586 588810 673206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 -3814 96134 93100 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 -3814 132134 93100 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 -3814 276134 94000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 -3814 420134 98000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 -3814 204134 238182 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 -3814 240134 238182 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 176600 96134 239592 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 176600 132134 239592 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 286182 204134 375600 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 286182 240134 375600 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 178000 276134 375600 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 -3814 312134 375600 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 -3814 348134 375600 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 331592 96134 388356 6 vssd2
port 538 nsew ground input
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 538 nsew ground input
rlabel metal4 s 23514 -3814 24134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 -3814 60134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 446407 96134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 331592 132134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 -3814 168134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 537993 204134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 537993 240134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 537993 276134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 537993 312134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 537993 348134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 -3814 384134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 142000 420134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 -3814 456134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 -3814 492134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 -3814 528134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 563514 -3814 564134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 539 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 540 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 541 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 542 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 543 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 544 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 545 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 546 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 547 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 548 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 549 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 550 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 551 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 552 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 553 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 554 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 555 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 556 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 557 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 558 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 559 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 560 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 561 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 562 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 563 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 564 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 565 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 566 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 567 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 568 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 569 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 570 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 571 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 572 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 573 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 574 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 575 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 576 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 577 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 578 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 579 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 580 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 581 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 582 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 583 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 584 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 585 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 586 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 587 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 588 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 589 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 590 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 591 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 592 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 593 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 594 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 595 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 596 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 597 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 598 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 599 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 600 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 601 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 602 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 603 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 604 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 605 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 606 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 607 nsew signal tristate
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 608 nsew signal tristate
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 609 nsew signal tristate
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 610 nsew signal tristate
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 611 nsew signal tristate
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 612 nsew signal tristate
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 613 nsew signal tristate
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 614 nsew signal tristate
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 615 nsew signal tristate
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 616 nsew signal tristate
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 617 nsew signal tristate
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 618 nsew signal tristate
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 619 nsew signal tristate
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 620 nsew signal tristate
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 621 nsew signal tristate
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 622 nsew signal tristate
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 623 nsew signal tristate
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 624 nsew signal tristate
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 625 nsew signal tristate
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 626 nsew signal tristate
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 627 nsew signal tristate
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 628 nsew signal tristate
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 629 nsew signal tristate
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 630 nsew signal tristate
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 631 nsew signal tristate
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 632 nsew signal tristate
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 633 nsew signal tristate
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 634 nsew signal tristate
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 635 nsew signal tristate
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 636 nsew signal tristate
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 637 nsew signal tristate
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 638 nsew signal tristate
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 639 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 640 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 641 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 642 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 643 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
