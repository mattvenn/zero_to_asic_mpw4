VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wrapped_ppm_decoder
  CLASS BLOCK ;
  FOREIGN wrapped_ppm_decoder ;
  ORIGIN 0.000 0.000 ;
  SIZE 100.000 BY 250.000 ;
  PIN active
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 242.120 100.000 242.720 ;
    END
  END active
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 97.960 100.000 98.560 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 219.000 4.000 219.600 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.840 4.000 109.440 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.650 246.000 85.930 250.000 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.650 246.000 62.930 250.000 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.440 4.000 123.040 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.050 246.000 12.330 250.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.890 0.000 37.170 4.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 228.520 100.000 229.120 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 57.160 100.000 57.760 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.050 246.000 81.330 250.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 137.400 4.000 138.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 178.200 4.000 178.800 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 140.120 100.000 140.720 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 4.000 21.040 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 185.000 4.000 185.600 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.450 246.000 30.730 250.000 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 235.320 100.000 235.920 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 43.560 100.000 44.160 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 111.560 100.000 112.160 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 246.000 26.130 250.000 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.890 0.000 83.170 4.000 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 153.720 100.000 154.320 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 4.000 116.240 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 4.000 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.690 0.000 50.970 4.000 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 70.760 100.000 71.360 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 151.000 4.000 151.600 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.530 246.000 6.810 250.000 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 119.720 100.000 120.320 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 160.520 100.000 161.120 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.650 246.000 39.930 250.000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 133.320 100.000 133.920 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.250 246.000 44.530 250.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.450 246.000 53.730 250.000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.850 246.000 72.130 250.000 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.450 246.000 99.730 250.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 214.920 100.000 215.520 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.490 0.000 18.770 4.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 232.600 4.000 233.200 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.890 0.000 60.170 4.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.290 0.000 78.570 4.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 221.720 100.000 222.320 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 29.960 100.000 30.560 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 180.920 100.000 181.520 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.250 246.000 21.530 250.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 4.000 95.840 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 246.200 4.000 246.800 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.050 246.000 35.330 250.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 9.560 100.000 10.160 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.490 0.000 41.770 4.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 104.760 100.000 105.360 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.930 246.000 2.210 250.000 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 187.720 100.000 188.320 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.290 0.000 9.570 4.000 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 36.760 100.000 37.360 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 91.160 100.000 91.760 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.850 246.000 95.130 250.000 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 164.600 4.000 165.200 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 16.360 100.000 16.960 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.290 0.000 55.570 4.000 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 157.800 4.000 158.400 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 201.320 100.000 201.920 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 4.000 89.040 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 63.960 100.000 64.560 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 198.600 4.000 199.200 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 225.800 4.000 226.400 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 4.000 129.840 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.610 0.000 97.890 4.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.890 0.000 14.170 4.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 4.000 82.240 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 50.360 100.000 50.960 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 167.320 100.000 167.920 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 126.520 100.000 127.120 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 2.760 100.000 3.360 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 144.200 4.000 144.800 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 84.360 100.000 84.960 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.040 4.000 102.640 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 4.000 7.440 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 194.520 100.000 195.120 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 23.160 100.000 23.760 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 208.120 100.000 208.720 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.090 0.000 69.370 4.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 4.000 41.440 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.490 0.000 87.770 4.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 212.200 4.000 212.800 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.650 246.000 16.930 250.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 246.000 58.330 250.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 13.640 4.000 14.240 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.090 0.000 23.370 4.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.690 0.000 4.970 4.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.450 246.000 76.730 250.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.850 246.000 49.130 250.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 4.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 246.000 90.530 250.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 77.560 100.000 78.160 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 191.800 4.000 192.400 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.690 0.000 27.970 4.000 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.090 0.000 46.370 4.000 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 174.120 100.000 174.720 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.690 0.000 73.970 4.000 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.250 246.000 67.530 250.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 205.400 4.000 206.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 239.400 4.000 240.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.010 0.000 93.290 4.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 171.400 4.000 172.000 ;
    END
  END io_out[9]
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 19.545 10.640 21.145 236.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 49.195 10.640 50.795 236.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.850 10.640 80.450 236.880 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 34.370 10.640 35.970 236.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 64.025 10.640 65.625 236.880 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 146.920 100.000 147.520 ;
    END
  END wb_clk_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 95.075 236.725 ;
      LAYER met1 ;
        RECT 0.070 10.640 99.750 236.880 ;
      LAYER met2 ;
        RECT 0.100 245.720 1.650 246.005 ;
        RECT 2.490 245.720 6.250 246.005 ;
        RECT 7.090 245.720 11.770 246.005 ;
        RECT 12.610 245.720 16.370 246.005 ;
        RECT 17.210 245.720 20.970 246.005 ;
        RECT 21.810 245.720 25.570 246.005 ;
        RECT 26.410 245.720 30.170 246.005 ;
        RECT 31.010 245.720 34.770 246.005 ;
        RECT 35.610 245.720 39.370 246.005 ;
        RECT 40.210 245.720 43.970 246.005 ;
        RECT 44.810 245.720 48.570 246.005 ;
        RECT 49.410 245.720 53.170 246.005 ;
        RECT 54.010 245.720 57.770 246.005 ;
        RECT 58.610 245.720 62.370 246.005 ;
        RECT 63.210 245.720 66.970 246.005 ;
        RECT 67.810 245.720 71.570 246.005 ;
        RECT 72.410 245.720 76.170 246.005 ;
        RECT 77.010 245.720 80.770 246.005 ;
        RECT 81.610 245.720 85.370 246.005 ;
        RECT 86.210 245.720 89.970 246.005 ;
        RECT 90.810 245.720 94.570 246.005 ;
        RECT 95.410 245.720 99.170 246.005 ;
        RECT 0.100 4.280 99.720 245.720 ;
        RECT 0.650 2.875 4.410 4.280 ;
        RECT 5.250 2.875 9.010 4.280 ;
        RECT 9.850 2.875 13.610 4.280 ;
        RECT 14.450 2.875 18.210 4.280 ;
        RECT 19.050 2.875 22.810 4.280 ;
        RECT 23.650 2.875 27.410 4.280 ;
        RECT 28.250 2.875 32.010 4.280 ;
        RECT 32.850 2.875 36.610 4.280 ;
        RECT 37.450 2.875 41.210 4.280 ;
        RECT 42.050 2.875 45.810 4.280 ;
        RECT 46.650 2.875 50.410 4.280 ;
        RECT 51.250 2.875 55.010 4.280 ;
        RECT 55.850 2.875 59.610 4.280 ;
        RECT 60.450 2.875 64.210 4.280 ;
        RECT 65.050 2.875 68.810 4.280 ;
        RECT 69.650 2.875 73.410 4.280 ;
        RECT 74.250 2.875 78.010 4.280 ;
        RECT 78.850 2.875 82.610 4.280 ;
        RECT 83.450 2.875 87.210 4.280 ;
        RECT 88.050 2.875 92.730 4.280 ;
        RECT 93.570 2.875 97.330 4.280 ;
        RECT 98.170 2.875 99.720 4.280 ;
      LAYER met3 ;
        RECT 4.400 245.800 96.000 246.650 ;
        RECT 4.000 243.120 96.000 245.800 ;
        RECT 4.000 241.720 95.600 243.120 ;
        RECT 4.000 240.400 96.000 241.720 ;
        RECT 4.400 239.000 96.000 240.400 ;
        RECT 4.000 236.320 96.000 239.000 ;
        RECT 4.000 234.920 95.600 236.320 ;
        RECT 4.000 233.600 96.000 234.920 ;
        RECT 4.400 232.200 96.000 233.600 ;
        RECT 4.000 229.520 96.000 232.200 ;
        RECT 4.000 228.120 95.600 229.520 ;
        RECT 4.000 226.800 96.000 228.120 ;
        RECT 4.400 225.400 96.000 226.800 ;
        RECT 4.000 222.720 96.000 225.400 ;
        RECT 4.000 221.320 95.600 222.720 ;
        RECT 4.000 220.000 96.000 221.320 ;
        RECT 4.400 218.600 96.000 220.000 ;
        RECT 4.000 215.920 96.000 218.600 ;
        RECT 4.000 214.520 95.600 215.920 ;
        RECT 4.000 213.200 96.000 214.520 ;
        RECT 4.400 211.800 96.000 213.200 ;
        RECT 4.000 209.120 96.000 211.800 ;
        RECT 4.000 207.720 95.600 209.120 ;
        RECT 4.000 206.400 96.000 207.720 ;
        RECT 4.400 205.000 96.000 206.400 ;
        RECT 4.000 202.320 96.000 205.000 ;
        RECT 4.000 200.920 95.600 202.320 ;
        RECT 4.000 199.600 96.000 200.920 ;
        RECT 4.400 198.200 96.000 199.600 ;
        RECT 4.000 195.520 96.000 198.200 ;
        RECT 4.000 194.120 95.600 195.520 ;
        RECT 4.000 192.800 96.000 194.120 ;
        RECT 4.400 191.400 96.000 192.800 ;
        RECT 4.000 188.720 96.000 191.400 ;
        RECT 4.000 187.320 95.600 188.720 ;
        RECT 4.000 186.000 96.000 187.320 ;
        RECT 4.400 184.600 96.000 186.000 ;
        RECT 4.000 181.920 96.000 184.600 ;
        RECT 4.000 180.520 95.600 181.920 ;
        RECT 4.000 179.200 96.000 180.520 ;
        RECT 4.400 177.800 96.000 179.200 ;
        RECT 4.000 175.120 96.000 177.800 ;
        RECT 4.000 173.720 95.600 175.120 ;
        RECT 4.000 172.400 96.000 173.720 ;
        RECT 4.400 171.000 96.000 172.400 ;
        RECT 4.000 168.320 96.000 171.000 ;
        RECT 4.000 166.920 95.600 168.320 ;
        RECT 4.000 165.600 96.000 166.920 ;
        RECT 4.400 164.200 96.000 165.600 ;
        RECT 4.000 161.520 96.000 164.200 ;
        RECT 4.000 160.120 95.600 161.520 ;
        RECT 4.000 158.800 96.000 160.120 ;
        RECT 4.400 157.400 96.000 158.800 ;
        RECT 4.000 154.720 96.000 157.400 ;
        RECT 4.000 153.320 95.600 154.720 ;
        RECT 4.000 152.000 96.000 153.320 ;
        RECT 4.400 150.600 96.000 152.000 ;
        RECT 4.000 147.920 96.000 150.600 ;
        RECT 4.000 146.520 95.600 147.920 ;
        RECT 4.000 145.200 96.000 146.520 ;
        RECT 4.400 143.800 96.000 145.200 ;
        RECT 4.000 141.120 96.000 143.800 ;
        RECT 4.000 139.720 95.600 141.120 ;
        RECT 4.000 138.400 96.000 139.720 ;
        RECT 4.400 137.000 96.000 138.400 ;
        RECT 4.000 134.320 96.000 137.000 ;
        RECT 4.000 132.920 95.600 134.320 ;
        RECT 4.000 130.240 96.000 132.920 ;
        RECT 4.400 128.840 96.000 130.240 ;
        RECT 4.000 127.520 96.000 128.840 ;
        RECT 4.000 126.120 95.600 127.520 ;
        RECT 4.000 123.440 96.000 126.120 ;
        RECT 4.400 122.040 96.000 123.440 ;
        RECT 4.000 120.720 96.000 122.040 ;
        RECT 4.000 119.320 95.600 120.720 ;
        RECT 4.000 116.640 96.000 119.320 ;
        RECT 4.400 115.240 96.000 116.640 ;
        RECT 4.000 112.560 96.000 115.240 ;
        RECT 4.000 111.160 95.600 112.560 ;
        RECT 4.000 109.840 96.000 111.160 ;
        RECT 4.400 108.440 96.000 109.840 ;
        RECT 4.000 105.760 96.000 108.440 ;
        RECT 4.000 104.360 95.600 105.760 ;
        RECT 4.000 103.040 96.000 104.360 ;
        RECT 4.400 101.640 96.000 103.040 ;
        RECT 4.000 98.960 96.000 101.640 ;
        RECT 4.000 97.560 95.600 98.960 ;
        RECT 4.000 96.240 96.000 97.560 ;
        RECT 4.400 94.840 96.000 96.240 ;
        RECT 4.000 92.160 96.000 94.840 ;
        RECT 4.000 90.760 95.600 92.160 ;
        RECT 4.000 89.440 96.000 90.760 ;
        RECT 4.400 88.040 96.000 89.440 ;
        RECT 4.000 85.360 96.000 88.040 ;
        RECT 4.000 83.960 95.600 85.360 ;
        RECT 4.000 82.640 96.000 83.960 ;
        RECT 4.400 81.240 96.000 82.640 ;
        RECT 4.000 78.560 96.000 81.240 ;
        RECT 4.000 77.160 95.600 78.560 ;
        RECT 4.000 75.840 96.000 77.160 ;
        RECT 4.400 74.440 96.000 75.840 ;
        RECT 4.000 71.760 96.000 74.440 ;
        RECT 4.000 70.360 95.600 71.760 ;
        RECT 4.000 69.040 96.000 70.360 ;
        RECT 4.400 67.640 96.000 69.040 ;
        RECT 4.000 64.960 96.000 67.640 ;
        RECT 4.000 63.560 95.600 64.960 ;
        RECT 4.000 62.240 96.000 63.560 ;
        RECT 4.400 60.840 96.000 62.240 ;
        RECT 4.000 58.160 96.000 60.840 ;
        RECT 4.000 56.760 95.600 58.160 ;
        RECT 4.000 55.440 96.000 56.760 ;
        RECT 4.400 54.040 96.000 55.440 ;
        RECT 4.000 51.360 96.000 54.040 ;
        RECT 4.000 49.960 95.600 51.360 ;
        RECT 4.000 48.640 96.000 49.960 ;
        RECT 4.400 47.240 96.000 48.640 ;
        RECT 4.000 44.560 96.000 47.240 ;
        RECT 4.000 43.160 95.600 44.560 ;
        RECT 4.000 41.840 96.000 43.160 ;
        RECT 4.400 40.440 96.000 41.840 ;
        RECT 4.000 37.760 96.000 40.440 ;
        RECT 4.000 36.360 95.600 37.760 ;
        RECT 4.000 35.040 96.000 36.360 ;
        RECT 4.400 33.640 96.000 35.040 ;
        RECT 4.000 30.960 96.000 33.640 ;
        RECT 4.000 29.560 95.600 30.960 ;
        RECT 4.000 28.240 96.000 29.560 ;
        RECT 4.400 26.840 96.000 28.240 ;
        RECT 4.000 24.160 96.000 26.840 ;
        RECT 4.000 22.760 95.600 24.160 ;
        RECT 4.000 21.440 96.000 22.760 ;
        RECT 4.400 20.040 96.000 21.440 ;
        RECT 4.000 17.360 96.000 20.040 ;
        RECT 4.000 15.960 95.600 17.360 ;
        RECT 4.000 14.640 96.000 15.960 ;
        RECT 4.400 13.240 96.000 14.640 ;
        RECT 4.000 10.560 96.000 13.240 ;
        RECT 4.000 9.160 95.600 10.560 ;
        RECT 4.000 7.840 96.000 9.160 ;
        RECT 4.400 6.440 96.000 7.840 ;
        RECT 4.000 3.760 96.000 6.440 ;
        RECT 4.000 2.895 95.600 3.760 ;
  END
END wrapped_ppm_decoder
END LIBRARY

